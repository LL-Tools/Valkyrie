

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654;

  AND2_X1 U7512 ( .A1(n7664), .A2(n7663), .ZN(n14318) );
  INV_X1 U7513 ( .A(n8029), .ZN(n16040) );
  XNOR2_X1 U7514 ( .A(n13449), .B(n14012), .ZN(n13983) );
  INV_X1 U7515 ( .A(n11533), .ZN(n12771) );
  OR2_X1 U7516 ( .A1(n10958), .A2(n10969), .ZN(n11059) );
  AND2_X1 U7517 ( .A1(n7668), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15934) );
  CLKBUF_X1 U7518 ( .A(n11144), .Z(n7442) );
  CLKBUF_X2 U7519 ( .A(n9249), .Z(n9805) );
  AND2_X2 U7521 ( .A1(n9147), .A2(n9930), .ZN(n9820) );
  BUF_X1 U7522 ( .A(n9190), .Z(n7439) );
  NAND2_X1 U7523 ( .A1(n13212), .A2(n9963), .ZN(n10876) );
  NAND3_X1 U7524 ( .A1(n9569), .A2(n9577), .A3(n8009), .ZN(n9628) );
  INV_X2 U7525 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n10117) );
  NAND3_X1 U7526 ( .A1(n12471), .A2(n8115), .A3(n12781), .ZN(n7643) );
  NAND2_X1 U7527 ( .A1(n15958), .A2(n15957), .ZN(n7586) );
  OAI211_X1 U7528 ( .C1(n8039), .C2(n8032), .A(n7411), .B(n8034), .ZN(n8038)
         );
  NAND2_X1 U7529 ( .A1(n7588), .A2(n7589), .ZN(n7411) );
  NAND3_X1 U7530 ( .A1(n8433), .A2(n7962), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7961) );
  INV_X2 U7531 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8433) );
  INV_X4 U7532 ( .A(n10899), .ZN(n10919) );
  OR2_X1 U7533 ( .A1(n8978), .A2(n8977), .ZN(n13967) );
  INV_X2 U7534 ( .A(n11490), .ZN(n14244) );
  INV_X1 U7535 ( .A(n10714), .ZN(n10702) );
  INV_X1 U7536 ( .A(n10981), .ZN(n13313) );
  OR2_X1 U7537 ( .A1(n8757), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8784) );
  OR2_X1 U7539 ( .A1(n8801), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8818) );
  INV_X1 U7540 ( .A(n13983), .ZN(n13994) );
  CLKBUF_X3 U7541 ( .A(n8494), .Z(n13351) );
  CLKBUF_X3 U7542 ( .A(n8467), .Z(n8923) );
  INV_X1 U7543 ( .A(n12328), .ZN(n8970) );
  INV_X1 U7544 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8626) );
  INV_X1 U7545 ( .A(n10876), .ZN(n10682) );
  INV_X1 U7546 ( .A(n9820), .ZN(n9796) );
  INV_X1 U7547 ( .A(n11209), .ZN(n9930) );
  AND4_X1 U7548 ( .A1(n8540), .A2(n8539), .A3(n8538), .A4(n8537), .ZN(n12988)
         );
  AND4_X1 U7549 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n12850)
         );
  INV_X1 U7550 ( .A(n11771), .ZN(n11772) );
  NAND2_X1 U7551 ( .A1(n13909), .A2(n13463), .ZN(n13893) );
  NAND2_X1 U7552 ( .A1(n9002), .A2(n8409), .ZN(n9005) );
  NAND2_X1 U7553 ( .A1(n9379), .A2(n9378), .ZN(n12928) );
  CLKBUF_X3 U7554 ( .A(n9754), .Z(n7433) );
  AOI211_X1 U7555 ( .C1(n13802), .C2(n16262), .A(n13801), .B(n13800), .ZN(
        n13803) );
  NAND4_X1 U7556 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n14384) );
  INV_X1 U7557 ( .A(n10848), .ZN(n10329) );
  XNOR2_X1 U7558 ( .A(n9097), .B(n9096), .ZN(n13209) );
  AND4_X1 U7559 ( .A1(n10320), .A2(n7413), .A3(n9922), .A4(n9921), .ZN(n7412)
         );
  NAND2_X2 U7560 ( .A1(n13210), .A2(n9104), .ZN(n9249) );
  AND2_X2 U7561 ( .A1(n8086), .A2(n8406), .ZN(n9002) );
  NAND2_X1 U7562 ( .A1(n9103), .A2(n13209), .ZN(n9190) );
  INV_X1 U7563 ( .A(n9103), .ZN(n13210) );
  BUF_X1 U7564 ( .A(n10319), .Z(n7413) );
  INV_X1 U7565 ( .A(n9963), .ZN(n14776) );
  INV_X2 U7566 ( .A(n9874), .ZN(n13032) );
  NOR2_X2 U7567 ( .A1(n15103), .A2(n8240), .ZN(n8239) );
  OAI21_X2 U7568 ( .B1(n13893), .B2(n13467), .A(n13461), .ZN(n13880) );
  OR2_X1 U7569 ( .A1(n10646), .A2(n9824), .ZN(n11092) );
  NAND2_X1 U7570 ( .A1(n10646), .A2(n12846), .ZN(n10958) );
  XNOR2_X2 U7571 ( .A(n9887), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10646) );
  AND2_X1 U7572 ( .A1(n10867), .A2(n10866), .ZN(n7600) );
  XNOR2_X2 U7573 ( .A(n8219), .B(n14365), .ZN(n10867) );
  BUF_X4 U7574 ( .A(n13766), .Z(n7414) );
  XNOR2_X1 U7575 ( .A(n8431), .B(n7942), .ZN(n13766) );
  AOI21_X2 U7576 ( .B1(n12581), .B2(n16055), .A(n16054), .ZN(n16063) );
  NOR2_X2 U7577 ( .A1(n15930), .A2(n15929), .ZN(n16096) );
  AND2_X1 U7578 ( .A1(n7959), .A2(n7955), .ZN(n7954) );
  NOR2_X1 U7579 ( .A1(n14744), .A2(n14493), .ZN(n8281) );
  CLKBUF_X1 U7580 ( .A(n10493), .Z(n10494) );
  OAI21_X1 U7581 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(n9768) );
  NAND2_X1 U7582 ( .A1(n10201), .A2(n10200), .ZN(n14710) );
  NAND2_X1 U7583 ( .A1(n10557), .A2(n10623), .ZN(n12551) );
  NAND2_X1 U7584 ( .A1(n8754), .A2(n8753), .ZN(n13449) );
  NAND2_X1 U7585 ( .A1(n8972), .A2(n13388), .ZN(n12738) );
  NAND2_X1 U7586 ( .A1(n13378), .A2(n13376), .ZN(n13515) );
  NAND2_X1 U7587 ( .A1(n13715), .A2(n8448), .ZN(n13367) );
  INV_X4 U7588 ( .A(n9260), .ZN(n7415) );
  CLKBUF_X2 U7589 ( .A(n10714), .Z(n10899) );
  BUF_X1 U7590 ( .A(n12846), .Z(n7436) );
  BUF_X1 U7591 ( .A(n9191), .Z(n7450) );
  BUF_X1 U7592 ( .A(n9754), .Z(n7434) );
  CLKBUF_X2 U7593 ( .A(n9190), .Z(n7438) );
  INV_X1 U7594 ( .A(n13209), .ZN(n9104) );
  NAND2_X2 U7595 ( .A1(n14784), .A2(n11308), .ZN(n11300) );
  NAND4_X1 U7596 ( .A1(n10120), .A2(n10117), .A3(n9919), .A4(n9918), .ZN(
        n10172) );
  OAI21_X1 U7597 ( .B1(n7520), .B2(n16598), .A(n10692), .ZN(n10693) );
  OR2_X1 U7598 ( .A1(n10945), .A2(n8229), .ZN(n10951) );
  NAND2_X1 U7599 ( .A1(n14840), .A2(n13292), .ZN(n14895) );
  NAND2_X1 U7600 ( .A1(n10916), .A2(n11852), .ZN(n10930) );
  AOI211_X1 U7601 ( .C1(n16588), .C2(n14662), .A(n14661), .B(n14660), .ZN(
        n14737) );
  XNOR2_X1 U7602 ( .A(n7423), .B(n14460), .ZN(n14462) );
  OAI22_X1 U7603 ( .A1(n14489), .A2(n8279), .B1(n8278), .B2(n7485), .ZN(n10373) );
  NAND2_X1 U7604 ( .A1(n14491), .A2(n14490), .ZN(n14489) );
  INV_X1 U7605 ( .A(n8280), .ZN(n7422) );
  AOI21_X1 U7606 ( .B1(n8280), .B2(n7421), .A(n8281), .ZN(n7420) );
  NAND2_X1 U7607 ( .A1(n14541), .A2(n10366), .ZN(n14533) );
  NAND2_X1 U7608 ( .A1(n14542), .A2(n14549), .ZN(n14541) );
  INV_X1 U7609 ( .A(n14490), .ZN(n7421) );
  NAND2_X1 U7610 ( .A1(n14558), .A2(n10365), .ZN(n14542) );
  NAND2_X1 U7611 ( .A1(n14559), .A2(n14570), .ZN(n14558) );
  OAI21_X1 U7612 ( .B1(n14574), .B2(n10364), .A(n10847), .ZN(n14559) );
  NAND2_X1 U7613 ( .A1(n10298), .A2(n10297), .ZN(n14467) );
  AND2_X1 U7614 ( .A1(n10494), .A2(n10495), .ZN(n7955) );
  NAND2_X1 U7615 ( .A1(n9816), .A2(n9795), .ZN(n13213) );
  NAND2_X1 U7616 ( .A1(n14599), .A2(n10363), .ZN(n14574) );
  NAND2_X1 U7617 ( .A1(n14601), .A2(n14600), .ZN(n14599) );
  AOI21_X1 U7618 ( .B1(n13788), .B2(n16213), .A(n13787), .ZN(n16238) );
  NAND2_X1 U7619 ( .A1(n7418), .A2(n7417), .ZN(n14601) );
  NAND2_X1 U7620 ( .A1(n9660), .A2(n9659), .ZN(n15718) );
  XNOR2_X1 U7621 ( .A(n9788), .B(n9787), .ZN(n13208) );
  OAI21_X1 U7622 ( .B1(n13130), .B2(n8923), .A(n8903), .ZN(n8915) );
  OAI21_X1 U7623 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9788) );
  OAI21_X1 U7624 ( .B1(n10211), .B2(n8342), .A(n8341), .ZN(n14581) );
  NAND2_X1 U7625 ( .A1(n7746), .A2(n7744), .ZN(n14906) );
  AND2_X1 U7626 ( .A1(n11061), .A2(n8214), .ZN(n8213) );
  NAND2_X1 U7627 ( .A1(n14631), .A2(n7419), .ZN(n7418) );
  OAI21_X1 U7628 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(n9784) );
  NAND2_X1 U7629 ( .A1(n7480), .A2(n11060), .ZN(n11061) );
  NAND2_X1 U7630 ( .A1(n14631), .A2(n10360), .ZN(n14614) );
  NAND2_X1 U7631 ( .A1(n10361), .A2(n10362), .ZN(n7417) );
  AND2_X1 U7632 ( .A1(n10361), .A2(n10360), .ZN(n7419) );
  OR2_X1 U7633 ( .A1(n16232), .A2(n7827), .ZN(n7826) );
  NAND2_X1 U7634 ( .A1(n8268), .A2(n9680), .ZN(n9725) );
  XNOR2_X1 U7635 ( .A(n13729), .B(n16243), .ZN(n16232) );
  AND2_X1 U7636 ( .A1(n14710), .A2(n14603), .ZN(n10362) );
  OR2_X1 U7637 ( .A1(n14710), .A2(n14603), .ZN(n10361) );
  NAND2_X1 U7638 ( .A1(n9551), .A2(n9550), .ZN(n15753) );
  NAND2_X1 U7639 ( .A1(n10217), .A2(n10216), .ZN(n14594) );
  NAND2_X1 U7640 ( .A1(n7426), .A2(n7424), .ZN(n10356) );
  NAND2_X1 U7641 ( .A1(n7426), .A2(n10354), .ZN(n16580) );
  NAND2_X1 U7642 ( .A1(n12701), .A2(n12705), .ZN(n7426) );
  NOR2_X1 U7643 ( .A1(n7464), .A2(n7425), .ZN(n7424) );
  OR2_X1 U7644 ( .A1(n9544), .A2(n11694), .ZN(n9569) );
  AND2_X1 U7645 ( .A1(n7534), .A2(n7834), .ZN(n16178) );
  AND2_X1 U7646 ( .A1(n16600), .A2(n12931), .ZN(n7464) );
  INV_X1 U7647 ( .A(n10354), .ZN(n7425) );
  NAND2_X1 U7648 ( .A1(n10181), .A2(n10180), .ZN(n14720) );
  AND2_X1 U7649 ( .A1(n12374), .A2(n10351), .ZN(n12457) );
  NAND2_X1 U7650 ( .A1(n10140), .A2(n10139), .ZN(n12863) );
  NAND2_X1 U7651 ( .A1(n12373), .A2(n7427), .ZN(n12374) );
  NAND2_X1 U7652 ( .A1(n8973), .A2(n7503), .ZN(n13073) );
  AND2_X1 U7653 ( .A1(n12375), .A2(n12372), .ZN(n7427) );
  NOR2_X1 U7654 ( .A1(n16141), .A2(n13721), .ZN(n13722) );
  NAND2_X1 U7655 ( .A1(n10125), .A2(n10124), .ZN(n12770) );
  OAI21_X1 U7656 ( .B1(n16125), .B2(n8016), .A(n8015), .ZN(n16141) );
  NAND2_X1 U7657 ( .A1(n10109), .A2(n10108), .ZN(n12644) );
  AND2_X1 U7658 ( .A1(n10351), .A2(n10103), .ZN(n12375) );
  NAND2_X1 U7659 ( .A1(n9404), .A2(n9403), .ZN(n12614) );
  NAND2_X1 U7660 ( .A1(n12211), .A2(n12210), .ZN(n12373) );
  NAND2_X1 U7661 ( .A1(n12131), .A2(n10350), .ZN(n12211) );
  OAI21_X1 U7662 ( .B1(n8209), .B2(n8208), .A(n8206), .ZN(n12565) );
  XNOR2_X1 U7663 ( .A(n9420), .B(n9419), .ZN(n11344) );
  NOR2_X1 U7664 ( .A1(n16007), .A2(n16006), .ZN(n16014) );
  NAND2_X1 U7665 ( .A1(n10348), .A2(n10347), .ZN(n12130) );
  AND2_X1 U7666 ( .A1(n7573), .A2(n7754), .ZN(n11882) );
  NAND2_X2 U7667 ( .A1(n9399), .A2(n9398), .ZN(n9420) );
  OAI21_X1 U7668 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n16012), .A(n16011), .ZN(
        n16018) );
  NAND2_X1 U7669 ( .A1(n9369), .A2(n7775), .ZN(n11251) );
  NAND2_X1 U7670 ( .A1(n7428), .A2(n8287), .ZN(n12081) );
  AND2_X1 U7671 ( .A1(n8308), .A2(n10031), .ZN(n8307) );
  OR2_X1 U7672 ( .A1(n15998), .A2(n15999), .ZN(n8026) );
  NAND2_X1 U7673 ( .A1(n7429), .A2(n10344), .ZN(n11702) );
  AND2_X1 U7674 ( .A1(n9859), .A2(n12178), .ZN(n11994) );
  NOR2_X1 U7675 ( .A1(n15995), .A2(n15994), .ZN(n16003) );
  AND2_X1 U7676 ( .A1(n13390), .A2(n13387), .ZN(n13512) );
  AND2_X1 U7677 ( .A1(n13364), .A2(n13367), .ZN(n8388) );
  NAND2_X1 U7678 ( .A1(n10339), .A2(n10338), .ZN(n7430) );
  AND2_X1 U7679 ( .A1(n16109), .A2(n11939), .ZN(n12110) );
  XNOR2_X1 U7680 ( .A(n15977), .B(n7670), .ZN(n15979) );
  NAND2_X1 U7681 ( .A1(n10605), .A2(n10604), .ZN(n16342) );
  INV_X1 U7682 ( .A(n10438), .ZN(n13713) );
  INV_X2 U7683 ( .A(n16398), .ZN(n7416) );
  OR2_X1 U7684 ( .A1(n15967), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U7685 ( .A1(n10333), .A2(n10334), .ZN(n10336) );
  NAND2_X1 U7686 ( .A1(n15975), .A2(n15976), .ZN(n15977) );
  AND3_X1 U7687 ( .A1(n8514), .A2(n8513), .A3(n8512), .ZN(n12670) );
  NAND4_X1 U7688 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n13585)
         );
  AND2_X1 U7689 ( .A1(n7837), .A2(n8020), .ZN(n16112) );
  NAND2_X1 U7690 ( .A1(n9996), .A2(n9997), .ZN(n12045) );
  NAND2_X4 U7691 ( .A1(n16566), .A2(n13302), .ZN(n10968) );
  AND3_X1 U7692 ( .A1(n8460), .A2(n8459), .A3(n7542), .ZN(n11919) );
  CLKBUF_X2 U7693 ( .A(n10705), .Z(n7435) );
  INV_X4 U7694 ( .A(n11059), .ZN(n13316) );
  NAND2_X1 U7695 ( .A1(n9184), .A2(n9161), .ZN(n9232) );
  NAND2_X1 U7696 ( .A1(n9194), .A2(n7511), .ZN(n14941) );
  NAND4_X1 U7697 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n14386)
         );
  NAND2_X1 U7698 ( .A1(n11724), .A2(n11209), .ZN(n8494) );
  NAND2_X1 U7699 ( .A1(n9163), .A2(n9164), .ZN(n9184) );
  AND3_X2 U7700 ( .A1(n9150), .A2(n9149), .A3(n9148), .ZN(n16314) );
  NAND2_X1 U7701 ( .A1(n8950), .A2(n9034), .ZN(n12413) );
  INV_X1 U7702 ( .A(n10035), .ZN(n9998) );
  OR2_X1 U7703 ( .A1(n9999), .A2(n12053), .ZN(n9968) );
  INV_X1 U7704 ( .A(n11092), .ZN(n10647) );
  CLKBUF_X1 U7705 ( .A(n10035), .Z(n10878) );
  INV_X2 U7706 ( .A(n7449), .ZN(n9318) );
  CLKBUF_X1 U7707 ( .A(n9191), .Z(n7449) );
  OR2_X1 U7708 ( .A1(n8427), .A2(n8411), .ZN(n8428) );
  XNOR2_X1 U7709 ( .A(n9127), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U7710 ( .A1(n9209), .A2(n11222), .ZN(n9235) );
  XNOR2_X1 U7711 ( .A(n9951), .B(n14770), .ZN(n9942) );
  NAND2_X2 U7712 ( .A1(n11300), .A2(n9930), .ZN(n10873) );
  NAND2_X2 U7713 ( .A1(n11300), .A2(n11209), .ZN(n10845) );
  NAND2_X2 U7714 ( .A1(n14769), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9951) );
  NOR2_X1 U7715 ( .A1(n8944), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U7716 ( .A1(n15792), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9094) );
  XNOR2_X1 U7717 ( .A(n8270), .B(n9929), .ZN(n14784) );
  NAND2_X1 U7718 ( .A1(n7412), .A2(n9938), .ZN(n14769) );
  XNOR2_X1 U7719 ( .A(n8269), .B(n9922), .ZN(n11308) );
  NOR2_X1 U7720 ( .A1(n9548), .A2(n8265), .ZN(n9117) );
  OR2_X1 U7721 ( .A1(n7412), .A2(n9939), .ZN(n9940) );
  OR2_X1 U7722 ( .A1(n8737), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8944) );
  XNOR2_X1 U7723 ( .A(n7665), .B(P2_IR_REG_20__SCAN_IN), .ZN(n10848) );
  NAND2_X2 U7724 ( .A1(n11208), .A2(P1_U3086), .ZN(n15805) );
  XNOR2_X1 U7725 ( .A(n9113), .B(n9112), .ZN(n14954) );
  NAND2_X2 U7726 ( .A1(n11208), .A2(P2_U3088), .ZN(n14792) );
  OR2_X1 U7727 ( .A1(n9108), .A2(n7761), .ZN(n9110) );
  NAND2_X1 U7728 ( .A1(n8302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8269) );
  NOR2_X2 U7729 ( .A1(n8475), .A2(n8474), .ZN(n11838) );
  NOR2_X1 U7730 ( .A1(n8087), .A2(n8089), .ZN(n8086) );
  NAND2_X1 U7731 ( .A1(n15936), .A2(n7676), .ZN(n15943) );
  NOR2_X1 U7732 ( .A1(n9920), .A2(n10172), .ZN(n10319) );
  NAND3_X1 U7733 ( .A1(n10059), .A2(n9913), .A3(n9981), .ZN(n10091) );
  NAND2_X1 U7734 ( .A1(n7960), .A2(n16084), .ZN(n8435) );
  AND2_X1 U7735 ( .A1(n8023), .A2(n8022), .ZN(n11736) );
  AND2_X1 U7736 ( .A1(n8350), .A2(n8349), .ZN(n9913) );
  AND2_X1 U7737 ( .A1(n8407), .A2(n8091), .ZN(n8090) );
  AND4_X1 U7738 ( .A1(n8404), .A2(n8403), .A3(n8648), .A4(n8645), .ZN(n8405)
         );
  AND3_X2 U7739 ( .A1(n8023), .A2(n8022), .A3(n8399), .ZN(n8458) );
  CLKBUF_X1 U7740 ( .A(n9116), .Z(n9888) );
  AND2_X1 U7741 ( .A1(n8946), .A2(n8408), .ZN(n7904) );
  AND2_X1 U7742 ( .A1(n7432), .A2(n7431), .ZN(n10059) );
  AND3_X1 U7743 ( .A1(n8528), .A2(n8509), .A3(n8473), .ZN(n8005) );
  INV_X1 U7744 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10391) );
  INV_X1 U7745 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n16084) );
  INV_X1 U7746 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n15636) );
  INV_X1 U7747 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10388) );
  INV_X1 U7748 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9918) );
  INV_X1 U7749 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8509) );
  INV_X1 U7750 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9919) );
  INV_X1 U7751 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8528) );
  INV_X4 U7752 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7753 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8403) );
  INV_X4 U7754 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7755 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9981) );
  INV_X1 U7756 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8022) );
  INV_X1 U7757 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9890) );
  INV_X1 U7758 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8023) );
  NOR2_X1 U7759 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8398) );
  INV_X1 U7760 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8648) );
  INV_X1 U7761 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10398) );
  INV_X1 U7762 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n10326) );
  INV_X1 U7763 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8645) );
  INV_X1 U7764 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n10120) );
  INV_X1 U7765 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8399) );
  INV_X1 U7766 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7691) );
  INV_X2 U7767 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7690) );
  INV_X1 U7768 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8473) );
  INV_X1 U7769 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n15631) );
  NOR2_X1 U7770 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8350) );
  INV_X1 U7771 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8946) );
  NOR2_X1 U7772 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8349) );
  NOR2_X1 U7773 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7431) );
  NOR2_X1 U7774 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7432) );
  OAI21_X1 U7775 ( .B1(n14491), .B2(n7422), .A(n7420), .ZN(n7423) );
  INV_X1 U7776 ( .A(n12205), .ZN(n12210) );
  INV_X2 U7777 ( .A(n10091), .ZN(n10320) );
  NAND2_X1 U7778 ( .A1(n8289), .A2(n11702), .ZN(n7428) );
  NAND2_X1 U7779 ( .A1(n11613), .A2(n10343), .ZN(n7429) );
  NAND2_X1 U7780 ( .A1(n7430), .A2(n10852), .ZN(n10342) );
  XNOR2_X1 U7781 ( .A(n7430), .B(n11686), .ZN(n11688) );
  XNOR2_X2 U7782 ( .A(n10705), .B(n11668), .ZN(n10333) );
  NAND3_X1 U7783 ( .A1(n7483), .A2(n9970), .A3(n9971), .ZN(n10705) );
  OR2_X2 U7784 ( .A1(n10819), .A2(n7459), .ZN(n7884) );
  NOR3_X4 U7785 ( .A1(n15131), .A2(n15691), .A3(n7952), .ZN(n15083) );
  AOI21_X2 U7786 ( .B1(n12529), .B2(n12530), .A(n10449), .ZN(n12520) );
  NAND2_X1 U7787 ( .A1(n9104), .A2(n9103), .ZN(n9754) );
  INV_X2 U7788 ( .A(n16314), .ZN(n9154) );
  OR2_X1 U7789 ( .A1(n7438), .A2(n11150), .ZN(n8397) );
  XNOR2_X1 U7790 ( .A(n8201), .B(P1_IR_REG_20__SCAN_IN), .ZN(n12846) );
  AND3_X1 U7791 ( .A1(n9079), .A2(n9135), .A3(n8215), .ZN(n9243) );
  AOI21_X2 U7792 ( .B1(n13131), .B2(n10477), .A(n8387), .ZN(n13623) );
  OR2_X1 U7793 ( .A1(n9095), .A2(n7761), .ZN(n9097) );
  BUF_X4 U7794 ( .A(n8481), .Z(n7437) );
  AND3_X4 U7795 ( .A1(n10901), .A2(n10696), .A3(n10695), .ZN(n10714) );
  AND4_X2 U7796 ( .A1(n9089), .A2(n9088), .A3(n9087), .A4(n9086), .ZN(n9486)
         );
  NAND2_X1 U7797 ( .A1(n12330), .A2(n10429), .ZN(n13366) );
  NAND2_X1 U7798 ( .A1(n10637), .A2(n10636), .ZN(n15701) );
  NAND2_X2 U7799 ( .A1(n12218), .A2(n12221), .ZN(n12217) );
  AND2_X1 U7800 ( .A1(n9147), .A2(n9930), .ZN(n7440) );
  NAND2_X2 U7801 ( .A1(n7448), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9131) );
  AND2_X1 U7802 ( .A1(n9896), .A2(n9111), .ZN(n15803) );
  NAND4_X2 U7803 ( .A1(n9133), .A2(n9132), .A3(n8397), .A4(n9131), .ZN(n10603)
         );
  CLKBUF_X1 U7804 ( .A(n11144), .Z(n7441) );
  INV_X2 U7805 ( .A(n9147), .ZN(n11144) );
  AND2_X1 U7806 ( .A1(n9147), .A2(n11209), .ZN(n7444) );
  AND2_X1 U7807 ( .A1(n9147), .A2(n11209), .ZN(n7445) );
  INV_X1 U7808 ( .A(n7444), .ZN(n7446) );
  AND2_X1 U7809 ( .A1(n9147), .A2(n11209), .ZN(n9186) );
  INV_X1 U7810 ( .A(n9249), .ZN(n7447) );
  INV_X1 U7811 ( .A(n9249), .ZN(n7448) );
  NAND2_X1 U7812 ( .A1(n13210), .A2(n13209), .ZN(n9191) );
  OAI21_X2 U7813 ( .B1(n12954), .B2(n8168), .A(n8167), .ZN(n15258) );
  NAND2_X2 U7814 ( .A1(n10626), .A2(n10560), .ZN(n12954) );
  OAI22_X2 U7815 ( .A1(n12196), .A2(n12197), .B1(n14935), .B2(n12891), .ZN(
        n12367) );
  OR2_X1 U7816 ( .A1(n8985), .A2(n8984), .ZN(n8986) );
  XNOR2_X1 U7817 ( .A(n14676), .B(n14492), .ZN(n10866) );
  INV_X1 U7818 ( .A(n11072), .ZN(n8196) );
  INV_X1 U7819 ( .A(n10957), .ZN(n10969) );
  AND2_X1 U7820 ( .A1(n8663), .A2(n8662), .ZN(n8678) );
  CLKBUF_X3 U7821 ( .A(n9998), .Z(n10683) );
  NOR2_X1 U7822 ( .A1(n10799), .A2(n10802), .ZN(n8364) );
  NAND2_X1 U7823 ( .A1(n10798), .A2(n10797), .ZN(n10800) );
  NOR2_X1 U7824 ( .A1(n7451), .A2(n10813), .ZN(n7870) );
  NAND2_X1 U7825 ( .A1(n9141), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7766) );
  NOR2_X1 U7826 ( .A1(n16176), .A2(n7838), .ZN(n13726) );
  AND2_X1 U7827 ( .A1(n16185), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7838) );
  AND2_X1 U7828 ( .A1(n13828), .A2(n8916), .ZN(n9062) );
  NAND2_X1 U7829 ( .A1(n7922), .A2(n7927), .ZN(n13828) );
  NAND2_X1 U7830 ( .A1(n13912), .A2(n8823), .ZN(n7908) );
  NAND2_X1 U7831 ( .A1(n11724), .A2(n9930), .ZN(n8467) );
  INV_X2 U7832 ( .A(n13487), .ZN(n13466) );
  AND2_X1 U7833 ( .A1(n8398), .A2(n8402), .ZN(n8006) );
  XNOR2_X1 U7834 ( .A(n11490), .B(n12271), .ZN(n11486) );
  NAND2_X1 U7835 ( .A1(n7892), .A2(n10832), .ZN(n7891) );
  NOR2_X1 U7836 ( .A1(n10834), .A2(n10837), .ZN(n8369) );
  NAND2_X1 U7837 ( .A1(n10834), .A2(n10837), .ZN(n8368) );
  AND2_X1 U7838 ( .A1(n10868), .A2(n14463), .ZN(n7582) );
  AND2_X1 U7839 ( .A1(n7533), .A2(n10369), .ZN(n8280) );
  NOR2_X1 U7840 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n10385) );
  OR2_X1 U7841 ( .A1(n14859), .A2(n8196), .ZN(n8195) );
  NAND2_X1 U7842 ( .A1(n7753), .A2(n7752), .ZN(n8209) );
  INV_X1 U7843 ( .A(n11884), .ZN(n7752) );
  NAND2_X1 U7844 ( .A1(n11882), .A2(n11883), .ZN(n7753) );
  XNOR2_X1 U7845 ( .A(n15696), .B(n14922), .ZN(n8152) );
  NAND2_X1 U7846 ( .A1(n10645), .A2(n14925), .ZN(n9640) );
  NOR2_X1 U7847 ( .A1(n16625), .A2(n8176), .ZN(n8175) );
  INV_X1 U7848 ( .A(n10627), .ZN(n8176) );
  BUF_X1 U7849 ( .A(n9147), .Z(n9590) );
  AND2_X1 U7850 ( .A1(n9580), .A2(n9627), .ZN(n9581) );
  AOI21_X1 U7851 ( .B1(n7980), .B2(n7982), .A(n7978), .ZN(n7977) );
  OAI21_X1 U7852 ( .B1(n11209), .B2(n9207), .A(n9206), .ZN(n9208) );
  NAND2_X1 U7853 ( .A1(n11209), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U7854 ( .A1(n7964), .A2(n7965), .ZN(n13687) );
  INV_X1 U7855 ( .A(n7966), .ZN(n7965) );
  OAI21_X1 U7856 ( .B1(n7968), .B2(n7967), .A(n13689), .ZN(n7966) );
  NAND2_X1 U7857 ( .A1(n7970), .A2(n7968), .ZN(n13610) );
  CLKBUF_X1 U7858 ( .A(n8631), .Z(n8932) );
  NAND3_X1 U7859 ( .A1(n9039), .A2(n9038), .A3(n9037), .ZN(n10955) );
  XNOR2_X1 U7860 ( .A(n13726), .B(n16197), .ZN(n16206) );
  OR2_X1 U7861 ( .A1(n16206), .A2(n16207), .ZN(n8014) );
  OR2_X1 U7862 ( .A1(n12972), .A2(n13409), .ZN(n8973) );
  AND2_X1 U7863 ( .A1(n8986), .A2(n13931), .ZN(n8085) );
  INV_X1 U7864 ( .A(n13351), .ZN(n8780) );
  INV_X1 U7865 ( .A(n8923), .ZN(n13353) );
  AND2_X1 U7866 ( .A1(n10529), .A2(n13466), .ZN(n13987) );
  AND2_X1 U7867 ( .A1(n9013), .A2(n9039), .ZN(n11376) );
  AND2_X1 U7868 ( .A1(n8792), .A2(n8774), .ZN(n8775) );
  INV_X1 U7869 ( .A(n7818), .ZN(n7817) );
  OAI21_X1 U7870 ( .B1(n8064), .B2(n7819), .A(n8772), .ZN(n7818) );
  INV_X1 U7871 ( .A(n8734), .ZN(n7819) );
  AND2_X1 U7872 ( .A1(n7807), .A2(n7806), .ZN(n8677) );
  OR2_X1 U7873 ( .A1(n8547), .A2(n8546), .ZN(n8569) );
  NAND2_X1 U7874 ( .A1(n14318), .A2(n7655), .ZN(n7647) );
  OAI21_X1 U7875 ( .B1(n14318), .B2(n7650), .A(n7648), .ZN(n14349) );
  INV_X1 U7876 ( .A(n7653), .ZN(n7650) );
  AOI21_X1 U7877 ( .B1(n7653), .B2(n7658), .A(n7649), .ZN(n7648) );
  INV_X1 U7878 ( .A(n14351), .ZN(n7649) );
  AND2_X1 U7879 ( .A1(n10896), .A2(n10895), .ZN(n10933) );
  NOR2_X1 U7880 ( .A1(n7791), .A2(n7782), .ZN(n7788) );
  INV_X1 U7881 ( .A(n7789), .ZN(n7787) );
  AOI21_X1 U7882 ( .B1(n14477), .B2(n7790), .A(n14463), .ZN(n7789) );
  NAND2_X1 U7883 ( .A1(n8332), .A2(n8329), .ZN(n14478) );
  NAND2_X1 U7884 ( .A1(n10275), .A2(n8330), .ZN(n8332) );
  NAND2_X1 U7885 ( .A1(n8274), .A2(n7486), .ZN(n8272) );
  AND2_X1 U7886 ( .A1(n10273), .A2(n10272), .ZN(n14512) );
  NAND2_X1 U7887 ( .A1(n7856), .A2(n14370), .ZN(n10366) );
  NAND2_X1 U7888 ( .A1(n10356), .A2(n8293), .ZN(n8292) );
  AND2_X1 U7889 ( .A1(n7501), .A2(n10355), .ZN(n8293) );
  NAND2_X1 U7890 ( .A1(n10371), .A2(n10370), .ZN(n16584) );
  OAI211_X1 U7891 ( .C1(n11671), .C2(n8304), .A(n11686), .B(n8303), .ZN(n11681) );
  NAND2_X1 U7892 ( .A1(n10849), .A2(n9991), .ZN(n8303) );
  INV_X1 U7893 ( .A(n9991), .ZN(n8304) );
  NOR2_X1 U7894 ( .A1(n14443), .A2(n8297), .ZN(n14658) );
  INV_X1 U7895 ( .A(n8298), .ZN(n8297) );
  NAND2_X1 U7896 ( .A1(n10867), .A2(n7454), .ZN(n8316) );
  INV_X1 U7897 ( .A(n8210), .ZN(n8207) );
  AOI21_X1 U7898 ( .B1(n8211), .B2(n11114), .A(n11120), .ZN(n8210) );
  INV_X1 U7899 ( .A(n8212), .ZN(n8211) );
  NOR2_X1 U7900 ( .A1(n8204), .A2(n8203), .ZN(n8202) );
  INV_X1 U7901 ( .A(n13168), .ZN(n8204) );
  INV_X1 U7902 ( .A(n11037), .ZN(n8203) );
  XNOR2_X1 U7903 ( .A(n7727), .B(n10643), .ZN(n10967) );
  OAI21_X1 U7904 ( .B1(n16550), .B2(n7748), .A(n14907), .ZN(n7747) );
  NAND2_X1 U7905 ( .A1(n7749), .A2(n7751), .ZN(n7748) );
  INV_X1 U7906 ( .A(n7750), .ZN(n7749) );
  NAND2_X1 U7907 ( .A1(n10641), .A2(n10640), .ZN(n8161) );
  AND2_X1 U7908 ( .A1(n10640), .A2(n9853), .ZN(n15090) );
  NAND2_X1 U7909 ( .A1(n7708), .A2(n7476), .ZN(n15074) );
  INV_X1 U7910 ( .A(n8152), .ZN(n15103) );
  OAI21_X1 U7911 ( .B1(n15210), .B2(n7711), .A(n7709), .ZN(n15177) );
  AND2_X1 U7912 ( .A1(n9854), .A2(n7710), .ZN(n7709) );
  OR2_X1 U7913 ( .A1(n7712), .A2(n7711), .ZN(n7710) );
  INV_X1 U7914 ( .A(n15174), .ZN(n7711) );
  NAND2_X1 U7915 ( .A1(n10628), .A2(n8177), .ZN(n8168) );
  NAND2_X1 U7916 ( .A1(n8171), .A2(n10628), .ZN(n8167) );
  NAND2_X1 U7917 ( .A1(n12551), .A2(n8234), .ZN(n12835) );
  NOR2_X1 U7918 ( .A1(n8236), .A2(n8235), .ZN(n8234) );
  INV_X1 U7919 ( .A(n10558), .ZN(n8235) );
  INV_X1 U7920 ( .A(n7760), .ZN(n7759) );
  OAI21_X1 U7921 ( .B1(n7489), .B2(n7761), .A(P1_IR_REG_26__SCAN_IN), .ZN(
        n7760) );
  XNOR2_X1 U7922 ( .A(n9701), .B(n9700), .ZN(n14789) );
  NAND2_X1 U7923 ( .A1(n16010), .A2(n16009), .ZN(n16011) );
  NAND2_X1 U7924 ( .A1(n8956), .A2(P3_U3897), .ZN(n16190) );
  NAND2_X1 U7925 ( .A1(n10265), .A2(n10264), .ZN(n14527) );
  NAND2_X1 U7926 ( .A1(n10304), .A2(n10303), .ZN(n14367) );
  NAND2_X1 U7927 ( .A1(n10296), .A2(n10295), .ZN(n14493) );
  AND2_X1 U7928 ( .A1(n14613), .A2(n10675), .ZN(n14648) );
  AOI22_X1 U7929 ( .A1(n10701), .A2(n10700), .B1(n10699), .B2(n11492), .ZN(
        n10708) );
  MUX2_X1 U7930 ( .A(n10700), .B(n10702), .S(n14387), .Z(n10699) );
  NAND2_X1 U7931 ( .A1(n7878), .A2(n7877), .ZN(n10724) );
  NAND2_X1 U7932 ( .A1(n12045), .A2(n10919), .ZN(n7878) );
  NAND2_X1 U7933 ( .A1(n14384), .A2(n10899), .ZN(n7877) );
  NAND2_X1 U7934 ( .A1(n9260), .A2(n14938), .ZN(n7616) );
  AOI21_X1 U7935 ( .B1(n7894), .B2(n10737), .A(n7893), .ZN(n8371) );
  INV_X1 U7936 ( .A(n10736), .ZN(n7893) );
  INV_X1 U7937 ( .A(n10743), .ZN(n8372) );
  NAND2_X1 U7938 ( .A1(n7603), .A2(n7601), .ZN(n10762) );
  NAND2_X1 U7939 ( .A1(n10758), .A2(n7602), .ZN(n7601) );
  NAND2_X1 U7940 ( .A1(n9493), .A2(n7612), .ZN(n7613) );
  NAND2_X1 U7941 ( .A1(n9508), .A2(n8262), .ZN(n8261) );
  AND2_X1 U7942 ( .A1(n9644), .A2(n9636), .ZN(n9637) );
  OAI21_X1 U7943 ( .B1(n10800), .B2(n8364), .A(n7887), .ZN(n10807) );
  AND2_X1 U7944 ( .A1(n10806), .A2(n8363), .ZN(n7887) );
  NAND2_X1 U7945 ( .A1(n7875), .A2(n10813), .ZN(n7874) );
  NOR2_X1 U7946 ( .A1(n10822), .A2(n10825), .ZN(n8359) );
  NAND2_X1 U7947 ( .A1(n10822), .A2(n10825), .ZN(n8358) );
  NOR2_X1 U7948 ( .A1(n10817), .A2(n10814), .ZN(n8354) );
  INV_X1 U7949 ( .A(n10814), .ZN(n8353) );
  INV_X1 U7950 ( .A(n10818), .ZN(n7886) );
  NOR2_X1 U7951 ( .A1(n8359), .A2(n7883), .ZN(n7882) );
  INV_X1 U7952 ( .A(n7885), .ZN(n7883) );
  INV_X1 U7953 ( .A(n8358), .ZN(n7880) );
  AOI21_X1 U7954 ( .B1(n7490), .B2(n7634), .A(n7465), .ZN(n7631) );
  NOR2_X1 U7955 ( .A1(n7633), .A2(n9704), .ZN(n7634) );
  NAND2_X1 U7956 ( .A1(n13493), .A2(n13492), .ZN(n13494) );
  NAND2_X1 U7957 ( .A1(n13359), .A2(n13360), .ZN(n13486) );
  OR2_X1 U7958 ( .A1(n8915), .A2(n13839), .ZN(n13481) );
  NOR2_X1 U7959 ( .A1(n7599), .A2(n10870), .ZN(n7598) );
  OR2_X1 U7960 ( .A1(n8281), .A2(n8280), .ZN(n8277) );
  INV_X1 U7961 ( .A(n13042), .ZN(n7735) );
  NAND2_X1 U7962 ( .A1(n7529), .A2(n7460), .ZN(n7705) );
  NAND2_X1 U7963 ( .A1(n8182), .A2(n15213), .ZN(n8181) );
  INV_X1 U7964 ( .A(n10631), .ZN(n8182) );
  NOR2_X1 U7965 ( .A1(n9483), .A2(n7984), .ZN(n7983) );
  INV_X1 U7966 ( .A(n9461), .ZN(n7984) );
  NAND2_X1 U7967 ( .A1(n7961), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n8434) );
  INV_X1 U7968 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7962) );
  OAI21_X1 U7969 ( .B1(n15944), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n15945), .ZN(
        n15946) );
  AND2_X1 U7970 ( .A1(n7969), .A2(n13611), .ZN(n7968) );
  NAND2_X1 U7971 ( .A1(n13638), .A2(n10500), .ZN(n7969) );
  OAI21_X1 U7972 ( .B1(n9069), .B2(n8054), .A(n8052), .ZN(n8051) );
  INV_X1 U7973 ( .A(n8053), .ZN(n8052) );
  OAI21_X1 U7974 ( .B1(n9063), .B2(n8054), .A(n13498), .ZN(n8053) );
  INV_X1 U7975 ( .A(n13486), .ZN(n13533) );
  NAND2_X1 U7976 ( .A1(n11813), .A2(n11776), .ZN(n11778) );
  NAND2_X1 U7977 ( .A1(n11801), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U7978 ( .A1(n13738), .A2(n7638), .ZN(n13739) );
  NAND2_X1 U7979 ( .A1(n13717), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U7980 ( .A1(n16179), .A2(n7576), .ZN(n13748) );
  NAND2_X1 U7981 ( .A1(n16217), .A2(n13750), .ZN(n13751) );
  AND2_X1 U7982 ( .A1(n8993), .A2(n13485), .ZN(n8097) );
  NOR2_X1 U7983 ( .A1(n13360), .A2(n8389), .ZN(n7927) );
  INV_X1 U7984 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15524) );
  INV_X1 U7985 ( .A(n14067), .ZN(n8655) );
  NAND2_X1 U7986 ( .A1(n13851), .A2(n13850), .ZN(n13853) );
  OR2_X1 U7987 ( .A1(n13467), .A2(n13468), .ZN(n13531) );
  OR2_X1 U7988 ( .A1(n9051), .A2(n9000), .ZN(n9048) );
  AND2_X1 U7989 ( .A1(n8951), .A2(n8945), .ZN(n8948) );
  INV_X1 U7990 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8945) );
  AND2_X1 U7991 ( .A1(n7825), .A2(n8583), .ZN(n7824) );
  INV_X1 U7992 ( .A(n8586), .ZN(n7825) );
  INV_X1 U7993 ( .A(n8493), .ZN(n8075) );
  INV_X1 U7994 ( .A(n8074), .ZN(n8073) );
  OAI21_X1 U7995 ( .B1(n8491), .B2(n8075), .A(n8506), .ZN(n8074) );
  NOR2_X1 U7996 ( .A1(n10183), .A2(n15867), .ZN(n10182) );
  NOR2_X1 U7997 ( .A1(n8114), .A2(n8110), .ZN(n8109) );
  INV_X1 U7998 ( .A(n13059), .ZN(n8110) );
  INV_X1 U7999 ( .A(n13158), .ZN(n8114) );
  INV_X1 U8000 ( .A(n13184), .ZN(n8112) );
  AND2_X1 U8001 ( .A1(n7656), .A2(n7654), .ZN(n7653) );
  OR2_X1 U8002 ( .A1(n14311), .A2(n7657), .ZN(n7656) );
  NAND2_X1 U8003 ( .A1(n7655), .A2(n14319), .ZN(n7654) );
  INV_X1 U8004 ( .A(n7659), .ZN(n7657) );
  NAND2_X1 U8005 ( .A1(n8218), .A2(n8217), .ZN(n10913) );
  NOR2_X1 U8006 ( .A1(n14467), .A2(n7860), .ZN(n7858) );
  OR2_X1 U8007 ( .A1(n10866), .A2(n8338), .ZN(n8337) );
  INV_X1 U8008 ( .A(n10274), .ZN(n8338) );
  INV_X1 U8009 ( .A(n14514), .ZN(n8294) );
  OR2_X1 U8010 ( .A1(n14752), .A2(n14369), .ZN(n8383) );
  NOR2_X1 U8011 ( .A1(n14566), .A2(n14698), .ZN(n7857) );
  INV_X1 U8012 ( .A(n8324), .ZN(n8327) );
  OAI21_X1 U8013 ( .B1(n10855), .B2(n8328), .A(n12205), .ZN(n8324) );
  INV_X1 U8014 ( .A(n10078), .ZN(n8328) );
  AND2_X1 U8015 ( .A1(n10346), .A2(n10345), .ZN(n8288) );
  AND2_X1 U8016 ( .A1(n12245), .A2(n10346), .ZN(n8289) );
  AND2_X2 U8017 ( .A1(n10902), .A2(n10329), .ZN(n10901) );
  INV_X1 U8018 ( .A(n9920), .ZN(n8374) );
  NOR2_X1 U8019 ( .A1(n10172), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8375) );
  INV_X1 U8020 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8142) );
  INV_X1 U8021 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10178) );
  AND2_X1 U8022 ( .A1(n10178), .A2(n10189), .ZN(n8143) );
  INV_X1 U8023 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10189) );
  INV_X1 U8024 ( .A(n10175), .ZN(n8144) );
  OR2_X1 U8025 ( .A1(n10020), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n10046) );
  INV_X1 U8026 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9980) );
  NOR2_X1 U8027 ( .A1(n7735), .A2(n7738), .ZN(n7733) );
  NOR2_X1 U8028 ( .A1(n7735), .A2(n12920), .ZN(n7734) );
  NOR2_X1 U8029 ( .A1(n7735), .A2(n7731), .ZN(n7730) );
  INV_X1 U8030 ( .A(n7571), .ZN(n7731) );
  NOR2_X1 U8031 ( .A1(n9618), .A2(n11105), .ZN(n9600) );
  NAND2_X1 U8032 ( .A1(n7635), .A2(n8223), .ZN(n9830) );
  NAND2_X1 U8033 ( .A1(n8224), .A2(n9774), .ZN(n8223) );
  OR2_X1 U8034 ( .A1(n15696), .A2(n15123), .ZN(n7953) );
  INV_X1 U8035 ( .A(n10573), .ZN(n8240) );
  AND2_X1 U8036 ( .A1(n15192), .A2(n10568), .ZN(n7712) );
  NAND2_X1 U8037 ( .A1(n8173), .A2(n8177), .ZN(n8172) );
  INV_X1 U8038 ( .A(n8175), .ZN(n8173) );
  NAND2_X1 U8039 ( .A1(n9786), .A2(n9785), .ZN(n15679) );
  INV_X1 U8040 ( .A(n11235), .ZN(n10599) );
  NAND2_X1 U8041 ( .A1(n7993), .A2(n7997), .ZN(n8268) );
  NOR2_X1 U8042 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n9084) );
  AOI21_X1 U8043 ( .B1(n7974), .B2(n7976), .A(n7566), .ZN(n7972) );
  NAND2_X1 U8044 ( .A1(n8222), .A2(n8221), .ZN(n8009) );
  INV_X1 U8045 ( .A(n9546), .ZN(n8221) );
  NAND2_X1 U8046 ( .A1(n7715), .A2(n7718), .ZN(n9439) );
  INV_X1 U8047 ( .A(n9444), .ZN(n9443) );
  XNOR2_X1 U8048 ( .A(n15960), .B(n8048), .ZN(n15961) );
  INV_X1 U8049 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n8048) );
  INV_X1 U8050 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16005) );
  INV_X1 U8051 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8036) );
  INV_X1 U8052 ( .A(n7671), .ZN(n16057) );
  OAI21_X1 U8053 ( .B1(n16049), .B2(n16050), .A(n7672), .ZN(n7671) );
  NAND2_X1 U8054 ( .A1(n16051), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n7672) );
  XNOR2_X1 U8055 ( .A(n16071), .B(n7688), .ZN(n16072) );
  NOR2_X1 U8056 ( .A1(n7992), .A2(n12387), .ZN(n7991) );
  INV_X1 U8057 ( .A(n10443), .ZN(n7992) );
  NOR2_X1 U8058 ( .A1(n7990), .A2(n7987), .ZN(n7986) );
  INV_X1 U8059 ( .A(n13678), .ZN(n7987) );
  INV_X1 U8060 ( .A(n13573), .ZN(n7990) );
  INV_X1 U8061 ( .A(n10483), .ZN(n7989) );
  XNOR2_X1 U8062 ( .A(n10429), .B(n10507), .ZN(n10431) );
  NAND2_X1 U8063 ( .A1(n8741), .A2(n15541), .ZN(n8757) );
  OAI21_X1 U8064 ( .B1(n11771), .B2(n11766), .A(n7640), .ZN(n11819) );
  NAND2_X1 U8065 ( .A1(n11771), .A2(n11766), .ZN(n7640) );
  NAND2_X1 U8066 ( .A1(n8458), .A2(n8473), .ZN(n8487) );
  NAND2_X1 U8067 ( .A1(n8021), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8020) );
  OAI21_X1 U8068 ( .B1(n12109), .B2(n12744), .A(n7513), .ZN(n12114) );
  NAND2_X1 U8069 ( .A1(n12114), .A2(n12113), .ZN(n12289) );
  INV_X1 U8070 ( .A(n12115), .ZN(n12113) );
  OAI211_X1 U8071 ( .C1(n12289), .C2(n12688), .A(n7831), .B(n7832), .ZN(n12291) );
  OR2_X1 U8072 ( .A1(n12288), .A2(n12688), .ZN(n7832) );
  NAND2_X1 U8073 ( .A1(n12289), .A2(n7833), .ZN(n7831) );
  AND2_X1 U8074 ( .A1(n12288), .A2(n12688), .ZN(n7833) );
  NOR2_X1 U8075 ( .A1(n12291), .A2(n12290), .ZN(n12689) );
  XNOR2_X1 U8076 ( .A(n13739), .B(n13768), .ZN(n16128) );
  NAND2_X1 U8077 ( .A1(n16128), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n16127) );
  INV_X1 U8078 ( .A(n16134), .ZN(n13768) );
  NAND2_X1 U8079 ( .A1(n7605), .A2(n7604), .ZN(n16165) );
  INV_X1 U8080 ( .A(n16162), .ZN(n7604) );
  INV_X1 U8081 ( .A(n16163), .ZN(n7605) );
  XNOR2_X1 U8082 ( .A(n13722), .B(n16159), .ZN(n16169) );
  OR2_X1 U8083 ( .A1(n16169), .A2(n16170), .ZN(n7834) );
  NAND2_X1 U8084 ( .A1(n7488), .A2(n8014), .ZN(n8013) );
  NAND2_X1 U8085 ( .A1(n8013), .A2(n8012), .ZN(n16223) );
  INV_X1 U8086 ( .A(n16224), .ZN(n8012) );
  NAND2_X1 U8087 ( .A1(n16223), .A2(n13728), .ZN(n13729) );
  XNOR2_X1 U8088 ( .A(n13751), .B(n13756), .ZN(n16235) );
  NAND2_X1 U8089 ( .A1(n16235), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n16234) );
  INV_X1 U8090 ( .A(n13509), .ZN(n8994) );
  NAND2_X1 U8091 ( .A1(n9069), .A2(n9063), .ZN(n9071) );
  AOI21_X1 U8092 ( .B1(n7921), .B2(n13979), .A(n7928), .ZN(n7919) );
  NAND2_X1 U8093 ( .A1(n7930), .A2(n7929), .ZN(n7928) );
  INV_X1 U8094 ( .A(n7923), .ZN(n7921) );
  NAND2_X1 U8095 ( .A1(n13857), .A2(n13987), .ZN(n7929) );
  AND2_X1 U8096 ( .A1(n13873), .A2(n7937), .ZN(n7936) );
  INV_X1 U8097 ( .A(n8385), .ZN(n7937) );
  NAND2_X1 U8098 ( .A1(n8817), .A2(n15532), .ZN(n8834) );
  INV_X1 U8099 ( .A(n8818), .ZN(n8817) );
  NAND2_X1 U8100 ( .A1(n14030), .A2(n8691), .ZN(n14029) );
  NAND2_X1 U8101 ( .A1(n13073), .A2(n13412), .ZN(n14092) );
  NAND2_X1 U8102 ( .A1(n12984), .A2(n8573), .ZN(n12973) );
  AOI21_X1 U8103 ( .B1(n8082), .B2(n8084), .A(n8080), .ZN(n8079) );
  INV_X1 U8104 ( .A(n13405), .ZN(n8080) );
  OAI21_X1 U8105 ( .B1(n12492), .B2(n7917), .A(n7915), .ZN(n12739) );
  AND2_X1 U8106 ( .A1(n7916), .A2(n13514), .ZN(n7915) );
  OR2_X1 U8107 ( .A1(n7479), .A2(n7917), .ZN(n7916) );
  INV_X1 U8108 ( .A(n8533), .ZN(n7917) );
  NAND2_X1 U8109 ( .A1(n12492), .A2(n7479), .ZN(n12848) );
  INV_X1 U8110 ( .A(n12413), .ZN(n13363) );
  OAI211_X1 U8111 ( .C1(n14209), .C2(n12403), .A(n12402), .B(n12401), .ZN(
        n12440) );
  NAND2_X1 U8112 ( .A1(n8844), .A2(n8843), .ZN(n13563) );
  INV_X1 U8113 ( .A(n13531), .ZN(n13895) );
  NAND2_X1 U8114 ( .A1(n13927), .A2(n8989), .ZN(n13909) );
  NAND2_X1 U8115 ( .A1(n13929), .A2(n8807), .ZN(n13912) );
  NAND2_X1 U8116 ( .A1(n8782), .A2(n8781), .ZN(n13570) );
  INV_X1 U8117 ( .A(n12828), .ZN(n16462) );
  AND2_X1 U8118 ( .A1(n14210), .A2(n10955), .ZN(n11722) );
  NAND2_X1 U8119 ( .A1(n9019), .A2(n9018), .ZN(n9045) );
  XNOR2_X1 U8120 ( .A(n9012), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9039) );
  AND2_X1 U8121 ( .A1(n9009), .A2(n9011), .ZN(n9038) );
  OAI21_X1 U8122 ( .B1(n8862), .B2(n8076), .A(n8864), .ZN(n8880) );
  INV_X1 U8123 ( .A(n8405), .ZN(n8087) );
  NAND2_X1 U8124 ( .A1(n8948), .A2(n8946), .ZN(n9034) );
  AOI21_X1 U8125 ( .B1(n7817), .B2(n7819), .A(n7816), .ZN(n7815) );
  INV_X1 U8126 ( .A(n8775), .ZN(n7816) );
  AOI21_X1 U8127 ( .B1(n8067), .B2(n8069), .A(n8065), .ZN(n8064) );
  INV_X1 U8128 ( .A(n8732), .ZN(n8065) );
  INV_X1 U8129 ( .A(n8068), .ZN(n8067) );
  OAI21_X1 U8130 ( .B1(n8697), .B2(n8069), .A(n8748), .ZN(n8068) );
  INV_X1 U8131 ( .A(n8729), .ZN(n8069) );
  NAND2_X1 U8132 ( .A1(n8658), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8660) );
  INV_X1 U8133 ( .A(n8661), .ZN(n7812) );
  NAND2_X1 U8134 ( .A1(n8660), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7813) );
  AND2_X1 U8135 ( .A1(n8639), .A2(n8622), .ZN(n8623) );
  AOI21_X1 U8136 ( .B1(n8604), .B2(n8063), .A(n8062), .ZN(n8061) );
  INV_X1 U8137 ( .A(n8620), .ZN(n8062) );
  INV_X1 U8138 ( .A(n8599), .ZN(n8063) );
  OAI21_X1 U8139 ( .B1(n8584), .B2(n7823), .A(n7820), .ZN(n8640) );
  INV_X1 U8140 ( .A(n8061), .ZN(n7823) );
  AND2_X1 U8141 ( .A1(n8059), .A2(n7821), .ZN(n7820) );
  AOI21_X1 U8142 ( .B1(n8061), .B2(n8603), .A(n8060), .ZN(n8059) );
  NAND2_X1 U8143 ( .A1(n8600), .A2(n8599), .ZN(n8605) );
  NAND2_X1 U8144 ( .A1(n8584), .A2(n7824), .ZN(n8600) );
  NAND2_X1 U8145 ( .A1(n7793), .A2(n8544), .ZN(n8547) );
  NAND2_X1 U8146 ( .A1(n8543), .A2(n8542), .ZN(n7793) );
  XNOR2_X1 U8147 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8506) );
  XNOR2_X1 U8148 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8491) );
  XNOR2_X1 U8149 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8439) );
  NAND2_X1 U8150 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7841) );
  INV_X1 U8151 ( .A(n8107), .ZN(n8103) );
  OR2_X1 U8152 ( .A1(n14290), .A2(n14264), .ZN(n8123) );
  AOI21_X1 U8153 ( .B1(n8102), .B2(n11962), .A(n8101), .ZN(n8100) );
  INV_X1 U8154 ( .A(n11976), .ZN(n8101) );
  NOR2_X1 U8155 ( .A1(n8120), .A2(n8116), .ZN(n8115) );
  INV_X1 U8156 ( .A(n12472), .ZN(n8116) );
  INV_X1 U8157 ( .A(n12630), .ZN(n8120) );
  AOI21_X1 U8158 ( .B1(n12630), .B2(n8119), .A(n8118), .ZN(n8117) );
  INV_X1 U8159 ( .A(n12627), .ZN(n8119) );
  INV_X1 U8160 ( .A(n12778), .ZN(n8118) );
  OR2_X1 U8161 ( .A1(n10279), .A2(n10278), .ZN(n10289) );
  INV_X1 U8162 ( .A(n11528), .ZN(n8126) );
  NAND2_X1 U8163 ( .A1(n12471), .A2(n12472), .ZN(n12628) );
  NAND2_X1 U8164 ( .A1(n13058), .A2(n13059), .ZN(n13156) );
  AOI21_X1 U8165 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(n8366) );
  INV_X1 U8166 ( .A(n10841), .ZN(n8367) );
  NOR2_X1 U8167 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  NAND2_X1 U8168 ( .A1(n10910), .A2(n10909), .ZN(n10932) );
  AND4_X1 U8169 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        n11647) );
  AND2_X1 U8170 ( .A1(n11511), .A2(n10953), .ZN(n11302) );
  OR2_X1 U8171 ( .A1(n10064), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U8172 ( .A1(n8294), .A2(n7858), .ZN(n14465) );
  OR2_X1 U8173 ( .A1(n14490), .A2(n8335), .ZN(n8331) );
  INV_X1 U8174 ( .A(n8340), .ZN(n8335) );
  OR2_X1 U8175 ( .A1(n8337), .A2(n8339), .ZN(n8336) );
  INV_X1 U8176 ( .A(n10275), .ZN(n8339) );
  NAND2_X1 U8177 ( .A1(n14533), .A2(n8383), .ZN(n8276) );
  OR2_X1 U8178 ( .A1(n14527), .A2(n14512), .ZN(n10367) );
  INV_X1 U8179 ( .A(n8276), .ZN(n8275) );
  NAND2_X1 U8180 ( .A1(n10866), .A2(n10367), .ZN(n8274) );
  INV_X1 U8181 ( .A(n10866), .ZN(n14509) );
  OR2_X1 U8182 ( .A1(n14566), .A2(n14343), .ZN(n10365) );
  XNOR2_X1 U8183 ( .A(n14551), .B(n14370), .ZN(n14549) );
  OR2_X1 U8184 ( .A1(n14548), .A2(n14549), .ZN(n14546) );
  INV_X1 U8185 ( .A(n8343), .ZN(n8342) );
  AOI21_X1 U8186 ( .B1(n8343), .B2(n14626), .A(n7508), .ZN(n8341) );
  AND2_X1 U8187 ( .A1(n14592), .A2(n10212), .ZN(n8343) );
  NAND2_X1 U8188 ( .A1(n13085), .A2(n10187), .ZN(n7779) );
  INV_X1 U8189 ( .A(n10187), .ZN(n7780) );
  NAND2_X1 U8190 ( .A1(n8346), .A2(n8344), .ZN(n13090) );
  OR2_X1 U8191 ( .A1(n8348), .A2(n8345), .ZN(n8344) );
  INV_X1 U8192 ( .A(n10171), .ZN(n8345) );
  NAND2_X1 U8193 ( .A1(n13090), .A2(n13089), .ZN(n13088) );
  AND2_X1 U8194 ( .A1(n13085), .A2(n7495), .ZN(n8291) );
  AND2_X1 U8195 ( .A1(n12912), .A2(n10156), .ZN(n8348) );
  OR2_X1 U8196 ( .A1(n10142), .A2(n12876), .ZN(n10162) );
  NAND2_X1 U8197 ( .A1(n16572), .A2(n16581), .ZN(n16574) );
  NAND2_X1 U8198 ( .A1(n7771), .A2(n7769), .ZN(n8311) );
  NOR2_X1 U8199 ( .A1(n7516), .A2(n7770), .ZN(n7769) );
  INV_X1 U8200 ( .A(n10115), .ZN(n7770) );
  NAND2_X1 U8201 ( .A1(n8311), .A2(n8310), .ZN(n12708) );
  AND2_X1 U8202 ( .A1(n10858), .A2(n10135), .ZN(n8310) );
  NAND2_X1 U8203 ( .A1(n12448), .A2(n12449), .ZN(n7771) );
  NOR2_X1 U8204 ( .A1(n7850), .A2(n7849), .ZN(n7848) );
  NAND2_X1 U8205 ( .A1(n10077), .A2(n10855), .ZN(n12125) );
  NAND2_X1 U8206 ( .A1(n12130), .A2(n10349), .ZN(n12131) );
  NAND2_X1 U8207 ( .A1(n11703), .A2(n8309), .ZN(n8308) );
  NAND2_X1 U8208 ( .A1(n11308), .A2(n11501), .ZN(n14604) );
  XNOR2_X1 U8209 ( .A(n11612), .B(n11647), .ZN(n11614) );
  NAND2_X1 U8210 ( .A1(n11661), .A2(n9977), .ZN(n11671) );
  NAND2_X1 U8211 ( .A1(n11671), .A2(n11675), .ZN(n11670) );
  AOI21_X1 U8212 ( .B1(n14478), .B2(n7783), .A(n7524), .ZN(n10666) );
  NOR2_X1 U8213 ( .A1(n7785), .A2(n7474), .ZN(n7783) );
  INV_X1 U8214 ( .A(n7788), .ZN(n7785) );
  NAND2_X1 U8215 ( .A1(n10383), .A2(n14298), .ZN(n14449) );
  INV_X1 U8216 ( .A(n10413), .ZN(n15818) );
  INV_X1 U8217 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9948) );
  INV_X1 U8218 ( .A(n8200), .ZN(n8199) );
  OAI21_X1 U8219 ( .B1(n14896), .B2(n13301), .A(n14796), .ZN(n8200) );
  INV_X1 U8220 ( .A(n15076), .ZN(n14897) );
  INV_X1 U8221 ( .A(n15114), .ZN(n14843) );
  NAND2_X1 U8222 ( .A1(n8213), .A2(n14906), .ZN(n14849) );
  INV_X1 U8223 ( .A(n14851), .ZN(n8214) );
  NAND2_X1 U8224 ( .A1(n11841), .A2(n11842), .ZN(n7754) );
  AOI21_X1 U8225 ( .B1(n7455), .B2(n8196), .A(n7515), .ZN(n8194) );
  NAND2_X1 U8226 ( .A1(n14857), .A2(n7455), .ZN(n7765) );
  INV_X1 U8227 ( .A(n11445), .ZN(n7714) );
  AOI21_X1 U8228 ( .B1(n12883), .B2(n7737), .A(n7571), .ZN(n7736) );
  INV_X1 U8229 ( .A(n14941), .ZN(n11846) );
  NAND2_X1 U8230 ( .A1(n13291), .A2(n14838), .ZN(n14840) );
  NOR2_X1 U8231 ( .A1(n11054), .A2(n7751), .ZN(n7750) );
  NAND2_X1 U8232 ( .A1(n9522), .A2(n9081), .ZN(n9548) );
  NOR3_X1 U8233 ( .A1(n15131), .A2(n15691), .A3(n7953), .ZN(n15082) );
  AND2_X1 U8234 ( .A1(n15130), .A2(n7472), .ZN(n8165) );
  AND2_X1 U8235 ( .A1(n15159), .A2(n7555), .ZN(n8148) );
  NAND2_X1 U8236 ( .A1(n15811), .A2(n9590), .ZN(n10645) );
  NAND2_X1 U8237 ( .A1(n10571), .A2(n9640), .ZN(n15159) );
  NAND2_X1 U8238 ( .A1(n8150), .A2(n15175), .ZN(n15183) );
  INV_X1 U8239 ( .A(n10567), .ZN(n8225) );
  INV_X1 U8240 ( .A(n10629), .ZN(n8187) );
  NAND2_X1 U8241 ( .A1(n15231), .A2(n15230), .ZN(n15229) );
  OAI21_X1 U8242 ( .B1(n16620), .B2(n7697), .A(n7695), .ZN(n15248) );
  AOI21_X1 U8243 ( .B1(n7698), .B2(n7701), .A(n7696), .ZN(n7695) );
  INV_X1 U8244 ( .A(n7698), .ZN(n7697) );
  OR2_X1 U8245 ( .A1(n8226), .A2(n7699), .ZN(n7698) );
  INV_X1 U8246 ( .A(n10565), .ZN(n7699) );
  NAND2_X1 U8247 ( .A1(n12954), .A2(n8175), .ZN(n8169) );
  NOR2_X1 U8248 ( .A1(n8228), .A2(n8227), .ZN(n8226) );
  INV_X1 U8249 ( .A(n10562), .ZN(n8227) );
  NAND2_X1 U8250 ( .A1(n16620), .A2(n16625), .ZN(n16619) );
  NAND2_X1 U8251 ( .A1(n9492), .A2(n9491), .ZN(n11055) );
  OR2_X1 U8252 ( .A1(n11093), .A2(n14957), .ZN(n15218) );
  OR2_X1 U8253 ( .A1(n11093), .A2(n9908), .ZN(n15216) );
  NAND2_X2 U8254 ( .A1(n9855), .A2(n10541), .ZN(n16349) );
  NAND2_X1 U8255 ( .A1(n9634), .A2(n9633), .ZN(n15739) );
  NOR2_X1 U8256 ( .A1(n10560), .A2(n8233), .ZN(n8232) );
  INV_X1 U8257 ( .A(n10559), .ZN(n8233) );
  NAND2_X1 U8258 ( .A1(n16324), .A2(n12308), .ZN(n16568) );
  OR2_X1 U8259 ( .A1(n9794), .A2(n9793), .ZN(n9816) );
  INV_X1 U8260 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7763) );
  INV_X1 U8261 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U8262 ( .A1(n8000), .A2(SI_22_), .ZN(n9588) );
  NAND2_X1 U8263 ( .A1(n7996), .A2(n8830), .ZN(n9657) );
  AND2_X1 U8264 ( .A1(n9657), .A2(n9588), .ZN(n9656) );
  NAND2_X1 U8265 ( .A1(n7609), .A2(n7608), .ZN(n9126) );
  INV_X1 U8266 ( .A(n9548), .ZN(n7609) );
  NAND2_X1 U8267 ( .A1(n9544), .A2(n11694), .ZN(n8222) );
  INV_X1 U8268 ( .A(n8009), .ZN(n8008) );
  NAND2_X1 U8269 ( .A1(n9439), .A2(n7475), .ZN(n9462) );
  INV_X1 U8270 ( .A(n9438), .ZN(n7717) );
  INV_X1 U8271 ( .A(n9419), .ZN(n7721) );
  NAND2_X1 U8272 ( .A1(n9369), .A2(n9368), .ZN(n9373) );
  NAND2_X1 U8273 ( .A1(n9373), .A2(n9372), .ZN(n9399) );
  INV_X1 U8274 ( .A(n9208), .ZN(n9209) );
  XNOR2_X1 U8275 ( .A(n15961), .B(n15950), .ZN(n15956) );
  NAND2_X1 U8276 ( .A1(n8046), .A2(n8045), .ZN(n15981) );
  INV_X1 U8277 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U8278 ( .A1(n8027), .A2(n8026), .ZN(n16006) );
  NAND2_X1 U8279 ( .A1(n8028), .A2(n16001), .ZN(n8027) );
  NAND2_X1 U8280 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n16133), .ZN(n7686) );
  OAI21_X1 U8281 ( .B1(n16029), .B2(n16028), .A(n16027), .ZN(n16033) );
  AND2_X1 U8282 ( .A1(n7680), .A2(n7682), .ZN(n16036) );
  NAND2_X1 U8283 ( .A1(n7675), .A2(n7673), .ZN(n16049) );
  NAND2_X1 U8284 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n7674), .ZN(n7673) );
  NAND2_X1 U8285 ( .A1(n16045), .A2(n16046), .ZN(n7675) );
  INV_X1 U8286 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n7674) );
  XNOR2_X1 U8287 ( .A(n16072), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n16067) );
  AND3_X1 U8288 ( .A1(n8554), .A2(n8553), .A3(n8552), .ZN(n12663) );
  NOR2_X1 U8289 ( .A1(n12895), .A2(n8004), .ZN(n8003) );
  INV_X1 U8290 ( .A(n10462), .ZN(n8004) );
  NAND2_X1 U8291 ( .A1(n12822), .A2(n10462), .ZN(n12896) );
  NAND2_X1 U8292 ( .A1(n8925), .A2(n8924), .ZN(n13245) );
  AND2_X1 U8293 ( .A1(n8875), .A2(n8874), .ZN(n13838) );
  AND3_X1 U8294 ( .A1(n8849), .A2(n8848), .A3(n8847), .ZN(n13897) );
  INV_X1 U8295 ( .A(n13675), .ZN(n13690) );
  INV_X1 U8296 ( .A(n16610), .ZN(n13137) );
  AND2_X1 U8297 ( .A1(n7803), .A2(n7801), .ZN(n7800) );
  INV_X1 U8298 ( .A(n13838), .ZN(n13870) );
  AND2_X1 U8299 ( .A1(n11742), .A2(n11741), .ZN(n16265) );
  OR2_X1 U8300 ( .A1(n16125), .A2(n16126), .ZN(n8018) );
  AND2_X1 U8301 ( .A1(n9068), .A2(n9067), .ZN(n13827) );
  INV_X1 U8302 ( .A(n14182), .ZN(n13921) );
  NAND2_X1 U8303 ( .A1(n8684), .A2(n8683), .ZN(n16534) );
  AND2_X1 U8304 ( .A1(n8740), .A2(n8739), .ZN(n14199) );
  INV_X1 U8305 ( .A(n16618), .ZN(n9044) );
  INV_X1 U8306 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7941) );
  INV_X1 U8307 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14215) );
  NOR2_X1 U8308 ( .A1(n8425), .A2(n8424), .ZN(n8429) );
  NOR2_X1 U8309 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8424) );
  NAND2_X1 U8310 ( .A1(n10277), .A2(n10276), .ZN(n14498) );
  NAND2_X1 U8311 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  OR2_X1 U8312 ( .A1(n12341), .A2(n10845), .ZN(n10201) );
  OAI21_X2 U8313 ( .B1(n11506), .B2(n11505), .A(n14640), .ZN(n14324) );
  INV_X1 U8314 ( .A(n14332), .ZN(n14355) );
  AND4_X1 U8315 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n12772) );
  OR2_X1 U8316 ( .A1(n11321), .A2(n14784), .ZN(n15897) );
  AOI21_X1 U8317 ( .B1(n14658), .B2(n14645), .A(n10691), .ZN(n10692) );
  NAND2_X1 U8318 ( .A1(n9932), .A2(n9931), .ZN(n14676) );
  NAND2_X2 U8319 ( .A1(n10672), .A2(n15823), .ZN(n14640) );
  OR2_X1 U8320 ( .A1(n16598), .A2(n10674), .ZN(n14613) );
  NAND2_X1 U8321 ( .A1(n7591), .A2(n16588), .ZN(n7590) );
  INV_X1 U8322 ( .A(n14659), .ZN(n7591) );
  NOR2_X1 U8323 ( .A1(n14736), .A2(n14708), .ZN(n10418) );
  NOR2_X1 U8324 ( .A1(n14740), .A2(n14708), .ZN(n7596) );
  AND2_X1 U8325 ( .A1(n8323), .A2(n7540), .ZN(n8319) );
  INV_X1 U8326 ( .A(n14658), .ZN(n8296) );
  NAND2_X1 U8327 ( .A1(n8313), .A2(n10867), .ZN(n8312) );
  INV_X1 U8328 ( .A(n10666), .ZN(n8313) );
  NAND2_X1 U8329 ( .A1(n10666), .A2(n8315), .ZN(n8314) );
  NOR2_X1 U8330 ( .A1(n10867), .A2(n7454), .ZN(n8315) );
  AND2_X1 U8331 ( .A1(n16595), .A2(n16588), .ZN(n8318) );
  NOR2_X1 U8332 ( .A1(n14449), .A2(n7583), .ZN(n14733) );
  NAND2_X1 U8333 ( .A1(n7585), .A2(n7584), .ZN(n7583) );
  INV_X1 U8334 ( .A(n14455), .ZN(n7584) );
  NAND2_X1 U8335 ( .A1(n14454), .A2(n16588), .ZN(n7585) );
  OAI21_X1 U8336 ( .B1(n10413), .B2(P2_D_REG_0__SCAN_IN), .A(n10412), .ZN(
        n15822) );
  INV_X1 U8337 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U8338 ( .A1(n15803), .A2(n9905), .ZN(n10957) );
  XNOR2_X1 U8339 ( .A(n9891), .B(n9890), .ZN(n11146) );
  NOR2_X1 U8340 ( .A1(n11113), .A2(n8212), .ZN(n11121) );
  AND2_X1 U8341 ( .A1(n16545), .A2(n16546), .ZN(n11050) );
  OR2_X1 U8342 ( .A1(n10975), .A2(n10974), .ZN(n10976) );
  NAND2_X1 U8343 ( .A1(n9572), .A2(n9571), .ZN(n15748) );
  NAND2_X1 U8344 ( .A1(n7724), .A2(n10643), .ZN(n7725) );
  NAND2_X1 U8345 ( .A1(n11461), .A2(n11462), .ZN(n7723) );
  INV_X1 U8346 ( .A(n11462), .ZN(n7724) );
  NAND2_X1 U8347 ( .A1(n9614), .A2(n9613), .ZN(n15729) );
  NAND2_X1 U8348 ( .A1(n9507), .A2(n9506), .ZN(n15762) );
  INV_X1 U8349 ( .A(n15235), .ZN(n14888) );
  NAND2_X1 U8350 ( .A1(n9654), .A2(n9653), .ZN(n14924) );
  NAND2_X1 U8351 ( .A1(n9609), .A2(n9608), .ZN(n15194) );
  NAND2_X1 U8352 ( .A1(n10583), .A2(n16631), .ZN(n15682) );
  INV_X1 U8353 ( .A(n8158), .ZN(n8157) );
  OAI21_X1 U8354 ( .B1(n8162), .B2(n8161), .A(n8159), .ZN(n8158) );
  AOI21_X1 U8355 ( .B1(n13220), .B2(n16631), .A(n13219), .ZN(n15693) );
  NAND2_X1 U8356 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  OAI21_X1 U8357 ( .B1(n10637), .B2(n8154), .A(n8151), .ZN(n15106) );
  NAND2_X1 U8358 ( .A1(n15701), .A2(n10638), .ZN(n15104) );
  NAND2_X1 U8359 ( .A1(n7416), .A2(n16327), .ZN(n16493) );
  AND2_X1 U8360 ( .A1(n12233), .A2(n12035), .ZN(n15247) );
  AND2_X1 U8361 ( .A1(n7436), .A2(n9874), .ZN(n16295) );
  NAND2_X1 U8362 ( .A1(n15771), .A2(n16635), .ZN(n15268) );
  NOR2_X1 U8363 ( .A1(n15803), .A2(n10586), .ZN(n11242) );
  INV_X1 U8364 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12340) );
  AND2_X1 U8365 ( .A1(n8047), .A2(n7462), .ZN(n16092) );
  AND2_X1 U8366 ( .A1(n16006), .A2(n16007), .ZN(n16015) );
  OR2_X1 U8367 ( .A1(n16014), .A2(n8037), .ZN(n8030) );
  INV_X1 U8368 ( .A(n16015), .ZN(n8039) );
  OR2_X1 U8369 ( .A1(n16014), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U8370 ( .A(n16033), .B(n16034), .ZN(n16035) );
  XNOR2_X1 U8371 ( .A(n16067), .B(n7687), .ZN(n16069) );
  NAND2_X1 U8372 ( .A1(n8043), .A2(n8044), .ZN(n8042) );
  NAND2_X1 U8373 ( .A1(n16065), .A2(n16066), .ZN(n8043) );
  OR2_X1 U8374 ( .A1(n10724), .A2(n8380), .ZN(n8379) );
  NAND2_X1 U8375 ( .A1(n8351), .A2(n10733), .ZN(n10741) );
  OR2_X1 U8376 ( .A1(n8259), .A2(n9288), .ZN(n8258) );
  NAND2_X1 U8377 ( .A1(n9288), .A2(n8259), .ZN(n7615) );
  INV_X1 U8378 ( .A(n10746), .ZN(n7895) );
  NOR2_X1 U8379 ( .A1(n10749), .A2(n10746), .ZN(n7896) );
  AND2_X1 U8380 ( .A1(n7546), .A2(n7627), .ZN(n7626) );
  NAND2_X1 U8381 ( .A1(n9335), .A2(n9338), .ZN(n7627) );
  NOR2_X1 U8382 ( .A1(n9335), .A2(n9338), .ZN(n7628) );
  NAND2_X1 U8383 ( .A1(n7629), .A2(n8263), .ZN(n9382) );
  OR2_X1 U8384 ( .A1(n8264), .A2(n9357), .ZN(n8263) );
  OAI21_X1 U8385 ( .B1(n9336), .B2(n7628), .A(n7626), .ZN(n7629) );
  INV_X1 U8386 ( .A(n9356), .ZN(n8264) );
  INV_X1 U8387 ( .A(n10768), .ZN(n7897) );
  NOR2_X1 U8388 ( .A1(n10771), .A2(n10768), .ZN(n7898) );
  INV_X1 U8389 ( .A(n9425), .ZN(n7622) );
  NAND2_X1 U8390 ( .A1(n9405), .A2(n9407), .ZN(n8250) );
  NAND2_X1 U8391 ( .A1(n9425), .A2(n7620), .ZN(n7619) );
  INV_X1 U8392 ( .A(n9427), .ZN(n7620) );
  NAND2_X1 U8393 ( .A1(n7618), .A2(n7617), .ZN(n9470) );
  AOI21_X1 U8394 ( .B1(n7456), .B2(n7621), .A(n7452), .ZN(n7617) );
  NAND2_X1 U8395 ( .A1(n9426), .A2(n7456), .ZN(n7618) );
  AND2_X1 U8396 ( .A1(n9427), .A2(n7622), .ZN(n7621) );
  NAND2_X1 U8397 ( .A1(n9494), .A2(n7614), .ZN(n7611) );
  OAI22_X1 U8398 ( .A1(n9529), .A2(n7623), .B1(n9530), .B2(n7624), .ZN(n9554)
         );
  AND2_X1 U8399 ( .A1(n9530), .A2(n7624), .ZN(n7623) );
  INV_X1 U8400 ( .A(n9528), .ZN(n7624) );
  NAND2_X1 U8401 ( .A1(n8364), .A2(n8363), .ZN(n8361) );
  NAND2_X1 U8402 ( .A1(n10802), .A2(n10799), .ZN(n8363) );
  NAND2_X1 U8403 ( .A1(n8255), .A2(n9573), .ZN(n8254) );
  NOR2_X1 U8404 ( .A1(n15159), .A2(n9617), .ZN(n9644) );
  NAND2_X1 U8405 ( .A1(n7869), .A2(n7873), .ZN(n7868) );
  INV_X1 U8406 ( .A(n7870), .ZN(n7869) );
  AOI22_X1 U8407 ( .A1(n7870), .A2(n7871), .B1(n7872), .B2(n7876), .ZN(n7867)
         );
  INV_X1 U8408 ( .A(n7525), .ZN(n7871) );
  NAND2_X1 U8409 ( .A1(n7525), .A2(n10813), .ZN(n7876) );
  NAND2_X1 U8410 ( .A1(n10818), .A2(n10821), .ZN(n7885) );
  OAI21_X1 U8411 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n9705) );
  NAND2_X1 U8412 ( .A1(n9684), .A2(n9686), .ZN(n8242) );
  NOR2_X1 U8413 ( .A1(n9684), .A2(n9686), .ZN(n8243) );
  NAND2_X1 U8414 ( .A1(n9729), .A2(n8252), .ZN(n8251) );
  NAND2_X1 U8415 ( .A1(n9704), .A2(n7633), .ZN(n7632) );
  NAND2_X1 U8416 ( .A1(n8359), .A2(n8358), .ZN(n8356) );
  NAND2_X1 U8417 ( .A1(n14260), .A2(n14261), .ZN(n7659) );
  AOI21_X1 U8418 ( .B1(n7882), .B2(n7459), .A(n7880), .ZN(n7879) );
  NAND2_X1 U8419 ( .A1(n10833), .A2(n7890), .ZN(n7889) );
  INV_X1 U8420 ( .A(n10832), .ZN(n7890) );
  NAND2_X1 U8421 ( .A1(n10580), .A2(n7625), .ZN(n9812) );
  NAND2_X1 U8422 ( .A1(n13032), .A2(n9825), .ZN(n7625) );
  MUX2_X1 U8423 ( .A(n14921), .B(n15686), .S(n7415), .Z(n9774) );
  NAND2_X1 U8424 ( .A1(n9745), .A2(n9744), .ZN(n7637) );
  NAND2_X1 U8425 ( .A1(n9749), .A2(n9748), .ZN(n7636) );
  NOR2_X1 U8426 ( .A1(n7999), .A2(n7995), .ZN(n7994) );
  NOR2_X1 U8427 ( .A1(n10252), .A2(n8830), .ZN(n7999) );
  INV_X1 U8428 ( .A(n9586), .ZN(n7995) );
  AND2_X1 U8429 ( .A1(n9677), .A2(n7998), .ZN(n7997) );
  NAND2_X1 U8430 ( .A1(n10252), .A2(n8830), .ZN(n7998) );
  INV_X1 U8431 ( .A(n7975), .ZN(n7974) );
  OAI21_X1 U8432 ( .B1(n9518), .B2(n7976), .A(n9541), .ZN(n7975) );
  INV_X1 U8433 ( .A(n9521), .ZN(n7976) );
  INV_X1 U8434 ( .A(n9500), .ZN(n7978) );
  OAI21_X1 U8435 ( .B1(n9141), .B2(n7593), .A(n7592), .ZN(n9185) );
  NAND2_X1 U8436 ( .A1(n9141), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U8437 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7677), .ZN(n7676) );
  NAND2_X1 U8438 ( .A1(n15935), .A2(n15934), .ZN(n15936) );
  INV_X1 U8439 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U8440 ( .A1(n8049), .A2(n15949), .ZN(n15960) );
  NOR2_X1 U8441 ( .A1(n7684), .A2(n16031), .ZN(n7683) );
  INV_X1 U8442 ( .A(n7686), .ZN(n7684) );
  INV_X1 U8443 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15543) );
  INV_X1 U8444 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15541) );
  NOR2_X1 U8445 ( .A1(n7967), .A2(n13612), .ZN(n7963) );
  NOR2_X1 U8446 ( .A1(n13507), .A2(n13538), .ZN(n7804) );
  OR2_X1 U8447 ( .A1(n11800), .A2(n7639), .ZN(n11941) );
  AND2_X1 U8448 ( .A1(n11801), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7639) );
  NOR2_X1 U8449 ( .A1(n13782), .A2(n16192), .ZN(n13784) );
  INV_X1 U8450 ( .A(n16266), .ZN(n7829) );
  INV_X1 U8451 ( .A(n8896), .ZN(n7925) );
  NOR2_X1 U8452 ( .A1(n8914), .A2(n7931), .ZN(n7924) );
  NAND2_X1 U8453 ( .A1(n13829), .A2(n13986), .ZN(n7930) );
  OR2_X1 U8454 ( .A1(n13563), .A2(n13897), .ZN(n13471) );
  OR2_X1 U8455 ( .A1(n13570), .A2(n13965), .ZN(n13510) );
  NAND2_X1 U8456 ( .A1(n8573), .A2(n7562), .ZN(n7913) );
  INV_X1 U8457 ( .A(n7913), .ZN(n7910) );
  INV_X1 U8458 ( .A(n8083), .ZN(n8082) );
  OAI21_X1 U8459 ( .B1(n13397), .B2(n8084), .A(n13517), .ZN(n8083) );
  INV_X1 U8460 ( .A(n13399), .ZN(n8084) );
  INV_X1 U8461 ( .A(n12849), .ZN(n13516) );
  NAND2_X1 U8462 ( .A1(n13943), .A2(n8790), .ZN(n7905) );
  NAND2_X1 U8463 ( .A1(n12404), .A2(n13366), .ZN(n13364) );
  NAND2_X1 U8464 ( .A1(n13544), .A2(n13363), .ZN(n13487) );
  INV_X1 U8465 ( .A(n13544), .ZN(n9000) );
  NAND2_X1 U8466 ( .A1(n8411), .A2(n7942), .ZN(n7939) );
  OAI21_X1 U8467 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8863) );
  INV_X1 U8468 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8407) );
  INV_X1 U8469 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8091) );
  NOR2_X1 U8470 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7903) );
  NOR2_X1 U8471 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7902) );
  INV_X1 U8472 ( .A(n8678), .ZN(n7811) );
  INV_X1 U8473 ( .A(n7810), .ZN(n7808) );
  NOR2_X1 U8474 ( .A1(n7811), .A2(n8077), .ZN(n7810) );
  INV_X1 U8475 ( .A(n8623), .ZN(n8060) );
  NAND2_X1 U8476 ( .A1(n7822), .A2(n8061), .ZN(n7821) );
  INV_X1 U8477 ( .A(n7824), .ZN(n7822) );
  INV_X1 U8478 ( .A(n8406), .ZN(n8607) );
  AND2_X1 U8479 ( .A1(n8005), .A2(n8398), .ZN(n8400) );
  AND2_X1 U8480 ( .A1(n10218), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U8481 ( .A1(n14230), .A2(n8139), .ZN(n8138) );
  INV_X1 U8482 ( .A(n13194), .ZN(n8139) );
  OR2_X1 U8483 ( .A1(n14434), .A2(n14438), .ZN(n10905) );
  AND2_X1 U8484 ( .A1(n10905), .A2(n10923), .ZN(n10912) );
  NOR2_X1 U8485 ( .A1(n8337), .A2(n10286), .ZN(n8330) );
  NOR2_X1 U8486 ( .A1(n10220), .A2(n10219), .ZN(n10218) );
  NOR2_X1 U8487 ( .A1(n16575), .A2(n7844), .ZN(n8301) );
  NAND2_X1 U8488 ( .A1(n7846), .A2(n7845), .ZN(n7844) );
  NOR2_X1 U8489 ( .A1(n14720), .A2(n13050), .ZN(n7845) );
  AND2_X1 U8490 ( .A1(n16581), .A2(n10171), .ZN(n8347) );
  NOR2_X1 U8491 ( .A1(n12450), .A2(n12770), .ZN(n12600) );
  INV_X1 U8492 ( .A(n10352), .ZN(n8286) );
  AND2_X1 U8493 ( .A1(n10083), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10095) );
  INV_X1 U8494 ( .A(n10018), .ZN(n8309) );
  NOR2_X1 U8495 ( .A1(n7474), .A2(n7782), .ZN(n7781) );
  OR2_X1 U8496 ( .A1(n8281), .A2(n7485), .ZN(n8279) );
  AND2_X1 U8497 ( .A1(n8277), .A2(n14463), .ZN(n8278) );
  NOR2_X1 U8498 ( .A1(n9511), .A2(n9510), .ZN(n9531) );
  INV_X1 U8499 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U8500 ( .A1(n14877), .A2(n14879), .ZN(n13265) );
  AOI21_X1 U8501 ( .B1(n14807), .B2(n8192), .A(n14867), .ZN(n8191) );
  INV_X1 U8502 ( .A(n14878), .ZN(n8192) );
  INV_X1 U8503 ( .A(n14807), .ZN(n8193) );
  INV_X1 U8504 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9510) );
  NOR2_X2 U8505 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9086) );
  NOR2_X1 U8506 ( .A1(n8238), .A2(n7703), .ZN(n7702) );
  INV_X1 U8507 ( .A(n7705), .ZN(n7703) );
  NAND2_X1 U8508 ( .A1(n15141), .A2(n7487), .ZN(n7704) );
  INV_X1 U8509 ( .A(n10633), .ZN(n8149) );
  NOR2_X1 U8510 ( .A1(n15198), .A2(n15729), .ZN(n15163) );
  OR2_X1 U8511 ( .A1(n9496), .A2(n9495), .ZN(n9511) );
  NOR2_X1 U8512 ( .A1(n9429), .A2(n9428), .ZN(n9454) );
  OR2_X1 U8513 ( .A1(n9410), .A2(n9409), .ZN(n9429) );
  AND2_X1 U8514 ( .A1(n9359), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9390) );
  AND2_X1 U8515 ( .A1(n7946), .A2(n12226), .ZN(n12360) );
  AND2_X1 U8516 ( .A1(n7947), .A2(n12310), .ZN(n7946) );
  INV_X1 U8517 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9339) );
  NOR2_X1 U8518 ( .A1(n12195), .A2(n8246), .ZN(n8245) );
  INV_X1 U8519 ( .A(n10550), .ZN(n8246) );
  OR2_X1 U8520 ( .A1(n9319), .A2(n12568), .ZN(n9340) );
  AND2_X1 U8521 ( .A1(n8392), .A2(n10543), .ZN(n8220) );
  AND2_X1 U8522 ( .A1(n16379), .A2(n9860), .ZN(n12002) );
  NAND2_X1 U8523 ( .A1(n8164), .A2(n8163), .ZN(n15119) );
  AOI21_X1 U8524 ( .B1(n8165), .B2(n15151), .A(n7514), .ZN(n8163) );
  AOI21_X1 U8525 ( .B1(n15257), .B2(n8183), .A(n8180), .ZN(n15201) );
  NAND2_X1 U8526 ( .A1(n8181), .A2(n7493), .ZN(n8180) );
  NOR2_X1 U8527 ( .A1(n8184), .A2(n8186), .ZN(n8183) );
  NAND2_X1 U8528 ( .A1(n7944), .A2(n7943), .ZN(n12186) );
  NOR2_X1 U8529 ( .A1(n11102), .A2(P1_U3086), .ZN(n11419) );
  AOI21_X1 U8530 ( .B1(n10599), .B2(n11238), .A(n11236), .ZN(n11415) );
  INV_X1 U8531 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9077) );
  NOR2_X1 U8532 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9116) );
  INV_X1 U8533 ( .A(n9576), .ZN(n9577) );
  AOI21_X1 U8534 ( .B1(n7981), .B2(n7983), .A(n7567), .ZN(n7980) );
  INV_X1 U8535 ( .A(n7475), .ZN(n7981) );
  INV_X1 U8536 ( .A(n7983), .ZN(n7982) );
  NAND2_X1 U8537 ( .A1(n7766), .A2(n8146), .ZN(n9138) );
  XNOR2_X1 U8538 ( .A(n15943), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n15944) );
  XNOR2_X1 U8539 ( .A(n15946), .B(n8050), .ZN(n15948) );
  INV_X1 U8540 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8050) );
  OAI21_X1 U8541 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(n15971), .A(n15970), .ZN(
        n15972) );
  NAND2_X1 U8542 ( .A1(n7669), .A2(n15980), .ZN(n15991) );
  NAND2_X1 U8543 ( .A1(n15979), .A2(n15978), .ZN(n7669) );
  XNOR2_X1 U8544 ( .A(n15991), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n15993) );
  NOR2_X1 U8545 ( .A1(n16004), .A2(n7587), .ZN(n16010) );
  AND2_X1 U8546 ( .A1(n16005), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n7587) );
  NAND2_X1 U8547 ( .A1(n16018), .A2(n7683), .ZN(n7680) );
  NAND2_X1 U8548 ( .A1(n16060), .A2(n16061), .ZN(n16071) );
  OR2_X1 U8549 ( .A1(n8722), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U8550 ( .A1(n8671), .A2(n15562), .ZN(n8705) );
  INV_X1 U8551 ( .A(n8686), .ZN(n8671) );
  OR2_X2 U8552 ( .A1(n8705), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8755) );
  INV_X1 U8553 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15542) );
  NAND2_X1 U8554 ( .A1(n12821), .A2(n10460), .ZN(n12822) );
  OR2_X1 U8555 ( .A1(n8556), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8575) );
  OR2_X1 U8556 ( .A1(n8593), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8614) );
  OR2_X1 U8557 ( .A1(n8614), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8633) );
  OAI21_X1 U8558 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(n13555) );
  INV_X1 U8559 ( .A(n13358), .ZN(n7798) );
  NAND2_X1 U8560 ( .A1(n7802), .A2(n13508), .ZN(n7801) );
  INV_X1 U8561 ( .A(n7804), .ZN(n7802) );
  NAND2_X1 U8562 ( .A1(n7804), .A2(n16333), .ZN(n7803) );
  NOR4_X1 U8563 ( .A1(n13538), .A2(n13537), .A3(n13536), .A4(n13535), .ZN(
        n13539) );
  NAND2_X1 U8564 ( .A1(n7830), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n11774) );
  INV_X1 U8565 ( .A(n11739), .ZN(n7830) );
  NAND2_X1 U8566 ( .A1(n11774), .A2(n11773), .ZN(n11814) );
  NAND2_X1 U8567 ( .A1(n11814), .A2(n11815), .ZN(n11813) );
  NOR2_X1 U8568 ( .A1(n11769), .A2(n11770), .ZN(n11800) );
  INV_X1 U8569 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15971) );
  XNOR2_X1 U8570 ( .A(n11941), .B(n11927), .ZN(n11802) );
  NAND2_X1 U8571 ( .A1(n7836), .A2(n7835), .ZN(n16109) );
  INV_X1 U8572 ( .A(n16111), .ZN(n7835) );
  INV_X1 U8573 ( .A(n16112), .ZN(n7836) );
  NAND2_X1 U8574 ( .A1(n12284), .A2(n12285), .ZN(n12680) );
  NOR2_X1 U8575 ( .A1(n12689), .A2(n12690), .ZN(n12693) );
  NAND2_X1 U8576 ( .A1(n16127), .A2(n13740), .ZN(n16144) );
  INV_X1 U8577 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15554) );
  NAND2_X1 U8578 ( .A1(n16160), .A2(n13744), .ZN(n16180) );
  NAND2_X1 U8579 ( .A1(n16180), .A2(n16181), .ZN(n16179) );
  NAND2_X1 U8580 ( .A1(n16165), .A2(n13779), .ZN(n16189) );
  XNOR2_X1 U8581 ( .A(n13748), .B(n16197), .ZN(n16199) );
  NAND2_X1 U8582 ( .A1(n8088), .A2(n8090), .ZN(n8737) );
  INV_X1 U8583 ( .A(n8700), .ZN(n8088) );
  NAND2_X1 U8584 ( .A1(n13731), .A2(n7829), .ZN(n7828) );
  NAND2_X1 U8585 ( .A1(n7829), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U8586 ( .A1(n16234), .A2(n13752), .ZN(n16256) );
  OR2_X1 U8587 ( .A1(n8926), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13807) );
  INV_X1 U8588 ( .A(n13480), .ZN(n8098) );
  OAI21_X1 U8589 ( .B1(n13882), .B2(n7521), .A(n7932), .ZN(n13856) );
  OR2_X1 U8590 ( .A1(n7936), .A2(n7933), .ZN(n7932) );
  INV_X1 U8591 ( .A(n8861), .ZN(n7933) );
  NAND2_X1 U8592 ( .A1(n8783), .A2(n15524), .ZN(n8801) );
  AND2_X1 U8593 ( .A1(n13511), .A2(n13510), .ZN(n13950) );
  OR2_X1 U8594 ( .A1(n16517), .A2(n14036), .ZN(n14040) );
  INV_X1 U8595 ( .A(n14053), .ZN(n14051) );
  NAND2_X1 U8596 ( .A1(n16483), .A2(n8630), .ZN(n7906) );
  NOR2_X1 U8597 ( .A1(n8630), .A2(n16483), .ZN(n7907) );
  INV_X1 U8598 ( .A(n13656), .ZN(n14088) );
  AND2_X1 U8599 ( .A1(n13418), .A2(n13424), .ZN(n14091) );
  NAND2_X1 U8600 ( .A1(n7909), .A2(n7911), .ZN(n13074) );
  INV_X1 U8601 ( .A(n7912), .ZN(n7911) );
  NAND2_X1 U8602 ( .A1(n12986), .A2(n7910), .ZN(n7909) );
  OAI22_X1 U8603 ( .A1(n8572), .A2(n7913), .B1(n16462), .B2(n13075), .ZN(n7912) );
  INV_X1 U8604 ( .A(n12986), .ZN(n7914) );
  OR2_X1 U8605 ( .A1(n8518), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8535) );
  AOI21_X1 U8606 ( .B1(n14219), .B2(n13353), .A(n8936), .ZN(n13815) );
  OR2_X1 U8607 ( .A1(n13351), .A2(n15461), .ZN(n8903) );
  AND2_X1 U8608 ( .A1(n13844), .A2(n13843), .ZN(n14110) );
  NAND2_X1 U8609 ( .A1(n13853), .A2(n8993), .ZN(n13844) );
  NAND2_X1 U8610 ( .A1(n8888), .A2(n8887), .ZN(n13686) );
  OR2_X1 U8611 ( .A1(n13351), .A2(n13069), .ZN(n8887) );
  OR2_X1 U8612 ( .A1(n13068), .A2(n8923), .ZN(n8888) );
  NAND2_X1 U8613 ( .A1(n8854), .A2(n8853), .ZN(n13637) );
  OR2_X1 U8614 ( .A1(n13351), .A2(n12905), .ZN(n8853) );
  AND3_X1 U8615 ( .A1(n8822), .A2(n8821), .A3(n8820), .ZN(n13933) );
  NAND2_X1 U8616 ( .A1(n7908), .A2(n10488), .ZN(n13894) );
  NAND2_X1 U8617 ( .A1(n8987), .A2(n8986), .ZN(n13925) );
  AND3_X1 U8618 ( .A1(n8532), .A2(n8531), .A3(n8530), .ZN(n16406) );
  INV_X1 U8619 ( .A(n13987), .ZN(n14087) );
  NAND2_X1 U8620 ( .A1(n8999), .A2(n9048), .ZN(n16428) );
  XNOR2_X1 U8621 ( .A(n8863), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n8862) );
  INV_X1 U8622 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8409) );
  XNOR2_X1 U8623 ( .A(n9036), .B(n9035), .ZN(n11723) );
  OAI21_X1 U8624 ( .B1(n9034), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9036) );
  AND2_X1 U8625 ( .A1(n8824), .A2(n8809), .ZN(n8810) );
  AND2_X1 U8626 ( .A1(n8732), .A2(n8731), .ZN(n8748) );
  AND2_X1 U8627 ( .A1(n8729), .A2(n8696), .ZN(n8697) );
  AND2_X1 U8628 ( .A1(n8656), .A2(n8641), .ZN(n8642) );
  AOI21_X1 U8629 ( .B1(n8073), .B2(n8075), .A(n7523), .ZN(n8071) );
  XNOR2_X1 U8630 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8524) );
  OR2_X1 U8631 ( .A1(n11961), .A2(n11960), .ZN(n8107) );
  NAND2_X1 U8632 ( .A1(n8106), .A2(n8105), .ZN(n8104) );
  INV_X1 U8633 ( .A(n11963), .ZN(n8106) );
  NAND2_X1 U8634 ( .A1(n13195), .A2(n8138), .ZN(n8137) );
  NAND2_X1 U8635 ( .A1(n14257), .A2(n7661), .ZN(n7660) );
  INV_X1 U8636 ( .A(n14258), .ZN(n7661) );
  NAND2_X1 U8637 ( .A1(n8108), .A2(n8111), .ZN(n13186) );
  AOI21_X1 U8638 ( .B1(n13158), .B2(n8113), .A(n8112), .ZN(n8111) );
  INV_X1 U8639 ( .A(n13155), .ZN(n8113) );
  NAND2_X1 U8640 ( .A1(n8099), .A2(n7500), .ZN(n7667) );
  MUX2_X1 U8641 ( .A(n9950), .B(n14793), .S(n11300), .Z(n11492) );
  NOR2_X1 U8642 ( .A1(n8136), .A2(n14278), .ZN(n8135) );
  INV_X1 U8643 ( .A(n14229), .ZN(n8136) );
  INV_X1 U8644 ( .A(n7642), .ZN(n7641) );
  OAI21_X1 U8645 ( .B1(n8117), .B2(n7644), .A(n12870), .ZN(n7642) );
  NAND2_X1 U8646 ( .A1(n11520), .A2(n11497), .ZN(n11528) );
  AND2_X1 U8647 ( .A1(n11498), .A2(n11489), .ZN(n11529) );
  NAND2_X1 U8648 ( .A1(n8145), .A2(n11488), .ZN(n11489) );
  INV_X1 U8649 ( .A(n11486), .ZN(n8145) );
  NAND2_X1 U8650 ( .A1(n11529), .A2(n11528), .ZN(n11527) );
  XNOR2_X1 U8651 ( .A(n14710), .B(n14244), .ZN(n14225) );
  OR2_X1 U8652 ( .A1(n10162), .A2(n9934), .ZN(n10183) );
  CLKBUF_X1 U8653 ( .A(n10091), .Z(n10176) );
  AND2_X1 U8654 ( .A1(n10310), .A2(n10290), .ZN(n14481) );
  OR2_X1 U8655 ( .A1(n14524), .A2(n14676), .ZN(n14514) );
  NAND2_X1 U8656 ( .A1(n8294), .A2(n10368), .ZN(n14496) );
  OR2_X1 U8657 ( .A1(n10255), .A2(n14344), .ZN(n10266) );
  AND3_X1 U8658 ( .A1(n7856), .A2(n14593), .A3(n7857), .ZN(n14550) );
  NAND2_X1 U8659 ( .A1(n14550), .A2(n14752), .ZN(n14524) );
  NAND2_X1 U8660 ( .A1(n14593), .A2(n7857), .ZN(n14562) );
  NAND2_X1 U8661 ( .A1(n14593), .A2(n14587), .ZN(n14583) );
  NOR2_X1 U8662 ( .A1(n14594), .A2(n14617), .ZN(n14593) );
  AOI21_X1 U8663 ( .B1(n7453), .B2(n7780), .A(n7492), .ZN(n7778) );
  NAND2_X1 U8664 ( .A1(n8301), .A2(n8300), .ZN(n14643) );
  INV_X1 U8665 ( .A(n8301), .ZN(n14642) );
  NAND2_X1 U8666 ( .A1(n7843), .A2(n7842), .ZN(n13093) );
  NOR2_X1 U8667 ( .A1(n16600), .A2(n13050), .ZN(n7842) );
  INV_X1 U8668 ( .A(n16575), .ZN(n7843) );
  NAND2_X1 U8669 ( .A1(n12600), .A2(n12882), .ZN(n16575) );
  NOR2_X1 U8670 ( .A1(n16575), .A2(n16600), .ZN(n16578) );
  NAND2_X1 U8671 ( .A1(n12455), .A2(n10352), .ZN(n12594) );
  AND4_X1 U8672 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n12864) );
  NAND2_X1 U8673 ( .A1(n12457), .A2(n12456), .ZN(n12455) );
  NAND2_X1 U8674 ( .A1(n7570), .A2(n7847), .ZN(n12451) );
  AOI21_X1 U8675 ( .B1(n12205), .B2(n8328), .A(n7499), .ZN(n8325) );
  NAND2_X1 U8676 ( .A1(n10077), .A2(n8327), .ZN(n8326) );
  INV_X1 U8677 ( .A(n12375), .ZN(n12371) );
  NAND2_X1 U8678 ( .A1(n7461), .A2(n12087), .ZN(n12206) );
  NAND2_X1 U8679 ( .A1(n12087), .A2(n12153), .ZN(n12138) );
  NAND2_X1 U8680 ( .A1(n8307), .A2(n10851), .ZN(n8305) );
  INV_X1 U8681 ( .A(n16419), .ZN(n7851) );
  NAND2_X1 U8682 ( .A1(n8290), .A2(n8289), .ZN(n12244) );
  OR2_X1 U8683 ( .A1(n11702), .A2(n10345), .ZN(n8290) );
  NOR2_X1 U8684 ( .A1(n11612), .A2(n11684), .ZN(n11698) );
  NAND2_X1 U8685 ( .A1(n11698), .A2(n12071), .ZN(n12257) );
  INV_X1 U8686 ( .A(n10849), .ZN(n11675) );
  NOR2_X1 U8687 ( .A1(n10697), .A2(n11668), .ZN(n11672) );
  NAND2_X1 U8688 ( .A1(n10328), .A2(n13114), .ZN(n14609) );
  INV_X1 U8689 ( .A(n14604), .ZN(n14575) );
  NAND2_X1 U8690 ( .A1(n10668), .A2(n10667), .ZN(n8219) );
  AND2_X1 U8691 ( .A1(n10946), .A2(n10415), .ZN(n16418) );
  OR2_X1 U8692 ( .A1(n14788), .A2(n10396), .ZN(n10413) );
  NAND2_X1 U8693 ( .A1(n10387), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U8694 ( .A1(n10386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10394) );
  OR2_X1 U8695 ( .A1(n10397), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n10386) );
  INV_X1 U8696 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10393) );
  XNOR2_X1 U8697 ( .A(n10399), .B(n10398), .ZN(n11511) );
  INV_X1 U8698 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U8699 ( .A1(n7666), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U8700 ( .A1(n7413), .A2(n10320), .ZN(n7666) );
  NAND2_X1 U8701 ( .A1(n8140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10214) );
  AND2_X1 U8702 ( .A1(n8143), .A2(n8142), .ZN(n8141) );
  AND2_X1 U8703 ( .A1(n10065), .A2(n10079), .ZN(n11423) );
  AND2_X1 U8704 ( .A1(n10021), .A2(n10046), .ZN(n14424) );
  NAND2_X1 U8705 ( .A1(n7491), .A2(n8211), .ZN(n8208) );
  INV_X1 U8706 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n12568) );
  NOR2_X1 U8707 ( .A1(n7730), .A2(n11030), .ZN(n7729) );
  NAND2_X1 U8708 ( .A1(n11016), .A2(n7734), .ZN(n7728) );
  NAND2_X1 U8709 ( .A1(n12883), .A2(n7733), .ZN(n7732) );
  AND2_X1 U8710 ( .A1(n14837), .A2(n13281), .ZN(n14866) );
  NAND2_X1 U8711 ( .A1(n7722), .A2(n8189), .ZN(n14836) );
  AOI21_X1 U8712 ( .B1(n8191), .B2(n8193), .A(n8190), .ZN(n8189) );
  NAND2_X1 U8713 ( .A1(n13265), .A2(n8191), .ZN(n7722) );
  INV_X1 U8714 ( .A(n14866), .ZN(n8190) );
  OAI21_X1 U8715 ( .B1(n11710), .B2(n10984), .A(n10983), .ZN(n11841) );
  INV_X1 U8716 ( .A(n10983), .ZN(n10986) );
  NAND2_X1 U8717 ( .A1(n10969), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10970) );
  OR2_X1 U8718 ( .A1(n9561), .A2(n9560), .ZN(n9618) );
  AND2_X1 U8719 ( .A1(n8194), .A2(n11097), .ZN(n7764) );
  NAND2_X1 U8720 ( .A1(n14857), .A2(n14859), .ZN(n14858) );
  INV_X1 U8721 ( .A(n8209), .ZN(n11115) );
  NOR2_X1 U8722 ( .A1(n11115), .A2(n11114), .ZN(n11113) );
  NOR2_X1 U8723 ( .A1(n9830), .A2(n9829), .ZN(n9883) );
  AOI21_X1 U8724 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9838) );
  AND4_X1 U8725 ( .A1(n9878), .A2(n9837), .A3(n9848), .A4(n9836), .ZN(n9882)
         );
  AND2_X1 U8726 ( .A1(n9599), .A2(n9598), .ZN(n14830) );
  NAND2_X1 U8727 ( .A1(n9248), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9102) );
  INV_X1 U8728 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15947) );
  OR2_X1 U8729 ( .A1(n9352), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U8730 ( .A1(n9111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U8731 ( .A1(n9798), .A2(n9797), .ZN(n15065) );
  OR2_X1 U8732 ( .A1(n13213), .A2(n9796), .ZN(n9798) );
  NOR2_X1 U8733 ( .A1(n15064), .A2(n15065), .ZN(n15066) );
  NAND2_X1 U8734 ( .A1(n10578), .A2(n8160), .ZN(n8159) );
  INV_X1 U8735 ( .A(n10640), .ZN(n8160) );
  AND2_X1 U8736 ( .A1(n8162), .A2(n10578), .ZN(n8156) );
  AND2_X1 U8737 ( .A1(n10639), .A2(n15090), .ZN(n8162) );
  OR2_X1 U8738 ( .A1(n7953), .A2(n15686), .ZN(n7952) );
  NOR2_X1 U8739 ( .A1(n10636), .A2(n8154), .ZN(n8153) );
  INV_X1 U8740 ( .A(n10638), .ZN(n8154) );
  NOR2_X1 U8741 ( .A1(n15131), .A2(n7953), .ZN(n15098) );
  AND2_X1 U8742 ( .A1(n9603), .A2(n9602), .ZN(n15186) );
  NAND2_X1 U8743 ( .A1(n7949), .A2(n7948), .ZN(n15238) );
  INV_X1 U8744 ( .A(n15753), .ZN(n7948) );
  NOR2_X1 U8745 ( .A1(n15238), .A2(n15748), .ZN(n15221) );
  OR2_X1 U8746 ( .A1(n9476), .A2(n14911), .ZN(n9496) );
  NAND2_X1 U8747 ( .A1(n12541), .A2(n10624), .ZN(n12833) );
  NAND2_X1 U8748 ( .A1(n12542), .A2(n12553), .ZN(n12541) );
  NAND2_X1 U8749 ( .A1(n12360), .A2(n16494), .ZN(n12611) );
  INV_X1 U8750 ( .A(n12186), .ZN(n12161) );
  AND2_X1 U8751 ( .A1(n10547), .A2(n10546), .ZN(n8248) );
  NAND2_X1 U8752 ( .A1(n12177), .A2(n10546), .ZN(n12164) );
  AND2_X1 U8753 ( .A1(n16452), .A2(n12808), .ZN(n11100) );
  NOR2_X1 U8754 ( .A1(n16344), .A2(n16365), .ZN(n16379) );
  AND2_X1 U8755 ( .A1(n10644), .A2(n10643), .ZN(n11412) );
  AND2_X1 U8756 ( .A1(n16314), .A2(n16310), .ZN(n16343) );
  INV_X1 U8757 ( .A(n10539), .ZN(n16315) );
  NAND2_X1 U8758 ( .A1(n11595), .A2(n9115), .ZN(n10539) );
  NAND2_X1 U8759 ( .A1(n14786), .A2(n9820), .ZN(n8007) );
  NAND2_X1 U8760 ( .A1(n12954), .A2(n10627), .ZN(n16627) );
  AND2_X1 U8761 ( .A1(n12835), .A2(n10559), .ZN(n12964) );
  INV_X1 U8762 ( .A(n12003), .ZN(n16401) );
  AOI21_X1 U8763 ( .B1(n10599), .B2(n10587), .A(n11242), .ZN(n12157) );
  NAND2_X1 U8764 ( .A1(n9109), .A2(n9112), .ZN(n8256) );
  INV_X1 U8765 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9096) );
  XNOR2_X1 U8766 ( .A(n9741), .B(n9740), .ZN(n14783) );
  NAND2_X1 U8767 ( .A1(n8266), .A2(n7608), .ZN(n8265) );
  AND2_X1 U8768 ( .A1(n15663), .A2(n9082), .ZN(n8266) );
  NAND2_X1 U8769 ( .A1(n9126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U8770 ( .A1(n8009), .A2(n9569), .ZN(n9575) );
  INV_X1 U8771 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U8772 ( .A1(n7973), .A2(n9521), .ZN(n9542) );
  NAND2_X1 U8773 ( .A1(n9519), .A2(n9518), .ZN(n7973) );
  NAND2_X1 U8774 ( .A1(n9351), .A2(n9350), .ZN(n9369) );
  OR2_X1 U8775 ( .A1(n9488), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9352) );
  XNOR2_X1 U8776 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15935) );
  NAND2_X1 U8777 ( .A1(n7586), .A2(n15959), .ZN(n15966) );
  NOR2_X1 U8778 ( .A1(n15985), .A2(n15984), .ZN(n15986) );
  NAND2_X1 U8779 ( .A1(n8037), .A2(n8035), .ZN(n7589) );
  NAND2_X1 U8780 ( .A1(n16023), .A2(n8036), .ZN(n8035) );
  OAI21_X1 U8781 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(n11551), .A(n16038), .ZN(
        n16045) );
  NAND2_X1 U8782 ( .A1(n7680), .A2(n7678), .ZN(n16038) );
  NOR2_X1 U8783 ( .A1(n7681), .A2(n7679), .ZN(n7678) );
  INV_X1 U8784 ( .A(n16037), .ZN(n7679) );
  OAI21_X1 U8785 ( .B1(n8042), .B2(n8041), .A(n16070), .ZN(n16076) );
  INV_X1 U8786 ( .A(n16069), .ZN(n8041) );
  INV_X1 U8787 ( .A(n11540), .ZN(n13075) );
  INV_X1 U8788 ( .A(n12323), .ZN(n10439) );
  AND4_X2 U8789 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n13582)
         );
  NAND2_X1 U8790 ( .A1(n8631), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U8791 ( .A1(n13571), .A2(n13573), .ZN(n13572) );
  AOI21_X1 U8792 ( .B1(n13687), .B2(n13235), .A(n7457), .ZN(n13239) );
  INV_X1 U8793 ( .A(n13681), .ZN(n13692) );
  AND4_X1 U8794 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .ZN(n14028)
         );
  AOI21_X1 U8795 ( .B1(n13640), .B2(n13639), .A(n13638), .ZN(n13642) );
  NAND2_X1 U8796 ( .A1(n12320), .A2(n10443), .ZN(n12386) );
  NAND2_X1 U8797 ( .A1(n7985), .A2(n7988), .ZN(n13649) );
  AOI21_X1 U8798 ( .B1(n13573), .B2(n7989), .A(n7518), .ZN(n7988) );
  AND4_X1 U8799 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n14086)
         );
  NAND2_X1 U8800 ( .A1(n13630), .A2(n10481), .ZN(n13679) );
  OR2_X1 U8801 ( .A1(n10480), .A2(n14012), .ZN(n10481) );
  NAND2_X1 U8802 ( .A1(n13679), .A2(n13678), .ZN(n13677) );
  NAND2_X1 U8803 ( .A1(n13610), .A2(n10504), .ZN(n13688) );
  NAND2_X1 U8804 ( .A1(n10512), .A2(n11722), .ZN(n13675) );
  NAND2_X1 U8805 ( .A1(n10530), .A2(n10529), .ZN(n13681) );
  INV_X1 U8806 ( .A(n13933), .ZN(n13703) );
  INV_X1 U8807 ( .A(n10955), .ZN(n10956) );
  INV_X1 U8808 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n16105) );
  NAND2_X1 U8809 ( .A1(n11756), .A2(n11772), .ZN(n11757) );
  NOR2_X1 U8810 ( .A1(n8458), .A2(n8626), .ZN(n8472) );
  AND2_X1 U8811 ( .A1(n8490), .A2(n8489), .ZN(n11792) );
  NAND2_X1 U8812 ( .A1(n7837), .A2(n8021), .ZN(n11799) );
  NOR2_X1 U8813 ( .A1(n11937), .A2(n8020), .ZN(n11936) );
  INV_X1 U8814 ( .A(n11942), .ZN(n11927) );
  NAND2_X1 U8815 ( .A1(n12102), .A2(n12103), .ZN(n12106) );
  NAND2_X1 U8816 ( .A1(n12106), .A2(n12105), .ZN(n12284) );
  XNOR2_X1 U8817 ( .A(n12680), .B(n12688), .ZN(n12286) );
  INV_X1 U8818 ( .A(n13719), .ZN(n8017) );
  NAND2_X1 U8819 ( .A1(n8019), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U8820 ( .A1(n13719), .A2(n8019), .ZN(n8015) );
  INV_X1 U8821 ( .A(n16142), .ZN(n8019) );
  INV_X1 U8822 ( .A(n7834), .ZN(n16171) );
  INV_X1 U8823 ( .A(n8014), .ZN(n16208) );
  INV_X1 U8824 ( .A(n8013), .ZN(n16225) );
  NOR2_X1 U8825 ( .A1(n16232), .A2(n16233), .ZN(n16231) );
  AND2_X1 U8826 ( .A1(n11742), .A2(n13791), .ZN(n16262) );
  INV_X1 U8827 ( .A(n13795), .ZN(n7606) );
  NAND2_X1 U8828 ( .A1(n9071), .A2(n13496), .ZN(n13327) );
  OAI21_X1 U8829 ( .B1(n8968), .B2(n14084), .A(n8967), .ZN(n13814) );
  INV_X1 U8830 ( .A(n7918), .ZN(n14108) );
  OAI211_X1 U8831 ( .C1(n13836), .C2(n7458), .A(n7920), .B(n7919), .ZN(n7918)
         );
  NAND2_X1 U8832 ( .A1(n7938), .A2(n7936), .ZN(n13868) );
  NAND2_X1 U8833 ( .A1(n8832), .A2(n8831), .ZN(n13903) );
  OR2_X1 U8834 ( .A1(n13351), .A2(n8830), .ZN(n8831) );
  NAND2_X1 U8835 ( .A1(n8800), .A2(n8799), .ZN(n13940) );
  AND2_X1 U8836 ( .A1(n8669), .A2(n8668), .ZN(n16610) );
  NAND2_X1 U8837 ( .A1(n12442), .A2(n12441), .ZN(n14046) );
  AND3_X1 U8838 ( .A1(n8654), .A2(n8653), .A3(n8652), .ZN(n14077) );
  NAND2_X1 U8839 ( .A1(n8973), .A2(n12971), .ZN(n13071) );
  NAND2_X1 U8840 ( .A1(n8081), .A2(n13399), .ZN(n12989) );
  NAND2_X1 U8841 ( .A1(n12738), .A2(n13397), .ZN(n8081) );
  NAND2_X1 U8842 ( .A1(n12848), .A2(n8533), .ZN(n12740) );
  INV_X1 U8843 ( .A(n16406), .ZN(n13391) );
  INV_X1 U8844 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12559) );
  NAND2_X1 U8845 ( .A1(n11722), .A2(n10514), .ZN(n14073) );
  INV_X1 U8846 ( .A(n13892), .ZN(n14098) );
  INV_X1 U8847 ( .A(n14046), .ZN(n14095) );
  AOI21_X1 U8848 ( .B1(n14213), .B2(n13353), .A(n13352), .ZN(n14152) );
  INV_X1 U8849 ( .A(n13686), .ZN(n14160) );
  NAND2_X1 U8850 ( .A1(n8867), .A2(n8866), .ZN(n14164) );
  INV_X1 U8851 ( .A(n13861), .ZN(n14167) );
  INV_X1 U8852 ( .A(n13563), .ZN(n14175) );
  AND2_X1 U8853 ( .A1(n8814), .A2(n8813), .ZN(n14182) );
  INV_X1 U8854 ( .A(n13570), .ZN(n14195) );
  INV_X1 U8855 ( .A(n13449), .ZN(n14203) );
  AND2_X1 U8856 ( .A1(n8704), .A2(n8703), .ZN(n14208) );
  AND2_X1 U8857 ( .A1(n9016), .A2(n9015), .ZN(n14209) );
  INV_X1 U8858 ( .A(n9045), .ZN(n14211) );
  AND2_X1 U8859 ( .A1(n11723), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14210) );
  OR2_X1 U8860 ( .A1(n8414), .A2(n8626), .ZN(n8412) );
  INV_X1 U8861 ( .A(n8417), .ZN(n14222) );
  INV_X1 U8862 ( .A(SI_25_), .ZN(n15466) );
  NOR2_X1 U8863 ( .A1(n11209), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14212) );
  MUX2_X1 U8864 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8949), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8950) );
  NAND2_X1 U8865 ( .A1(n8955), .A2(n8954), .ZN(n12192) );
  OAI21_X1 U8866 ( .B1(n8066), .B2(n7819), .A(n7817), .ZN(n8776) );
  INV_X1 U8867 ( .A(SI_18_), .ZN(n11694) );
  NAND2_X1 U8868 ( .A1(n8735), .A2(n8734), .ZN(n8773) );
  NAND2_X1 U8869 ( .A1(n8066), .A2(n8064), .ZN(n8735) );
  INV_X1 U8870 ( .A(SI_16_), .ZN(n15479) );
  INV_X1 U8871 ( .A(SI_15_), .ZN(n11442) );
  INV_X1 U8872 ( .A(SI_14_), .ZN(n11411) );
  NAND2_X1 U8873 ( .A1(n7813), .A2(n8661), .ZN(n8679) );
  XNOR2_X1 U8874 ( .A(n8682), .B(n8681), .ZN(n16185) );
  INV_X1 U8875 ( .A(SI_13_), .ZN(n15488) );
  OR2_X1 U8876 ( .A1(n7813), .A2(n7812), .ZN(n8714) );
  NAND2_X1 U8877 ( .A1(n8660), .A2(n8661), .ZN(n8712) );
  INV_X1 U8878 ( .A(SI_12_), .ZN(n15487) );
  OAI21_X1 U8879 ( .B1(n8600), .B2(n8603), .A(n8061), .ZN(n8624) );
  NAND2_X1 U8880 ( .A1(n8605), .A2(n8604), .ZN(n8621) );
  NAND2_X1 U8881 ( .A1(n8584), .A2(n8583), .ZN(n8587) );
  NAND2_X1 U8882 ( .A1(n8569), .A2(n8568), .ZN(n8581) );
  NAND2_X1 U8883 ( .A1(n8072), .A2(n8493), .ZN(n8507) );
  NAND2_X1 U8884 ( .A1(n8492), .A2(n8491), .ZN(n8072) );
  INV_X1 U8885 ( .A(n8458), .ZN(n8024) );
  NAND2_X1 U8886 ( .A1(n8457), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n8025) );
  INV_X1 U8887 ( .A(SI_1_), .ZN(n15502) );
  INV_X1 U8888 ( .A(n8439), .ZN(n8436) );
  NAND2_X1 U8889 ( .A1(n8432), .A2(n7839), .ZN(n11738) );
  INV_X1 U8890 ( .A(n7840), .ZN(n7839) );
  OAI22_X1 U8891 ( .A1(n11735), .A2(n7841), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_1__SCAN_IN), .ZN(n7840) );
  AND4_X1 U8892 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n12352) );
  NAND2_X1 U8893 ( .A1(n8104), .A2(n8107), .ZN(n11970) );
  NAND2_X1 U8894 ( .A1(n14349), .A2(n14265), .ZN(n14291) );
  NAND2_X1 U8895 ( .A1(n11527), .A2(n11498), .ZN(n11578) );
  AND2_X1 U8896 ( .A1(n10238), .A2(n10237), .ZN(n14605) );
  NAND2_X1 U8897 ( .A1(n8137), .A2(n14229), .ZN(n14279) );
  INV_X1 U8898 ( .A(n8122), .ZN(n8121) );
  OAI22_X1 U8899 ( .A1(n8123), .A2(n14351), .B1(n14288), .B2(n14289), .ZN(
        n8122) );
  NAND2_X1 U8900 ( .A1(n10243), .A2(n10242), .ZN(n14566) );
  NAND2_X1 U8901 ( .A1(n12780), .A2(n12781), .ZN(n12871) );
  NAND2_X1 U8902 ( .A1(n7645), .A2(n8117), .ZN(n12780) );
  NAND2_X1 U8903 ( .A1(n8115), .A2(n12471), .ZN(n7645) );
  NAND2_X1 U8904 ( .A1(n7662), .A2(n7660), .ZN(n14310) );
  NAND2_X1 U8905 ( .A1(n7652), .A2(n7651), .ZN(n7662) );
  INV_X1 U8906 ( .A(n14319), .ZN(n7651) );
  INV_X1 U8907 ( .A(n14318), .ZN(n7652) );
  NAND2_X1 U8908 ( .A1(n13157), .A2(n13158), .ZN(n13185) );
  NAND2_X1 U8909 ( .A1(n13156), .A2(n13155), .ZN(n13157) );
  NAND2_X1 U8910 ( .A1(n11645), .A2(n11646), .ZN(n11654) );
  AND2_X1 U8911 ( .A1(n8130), .A2(n11576), .ZN(n7646) );
  INV_X1 U8912 ( .A(n11584), .ZN(n8130) );
  OAI21_X1 U8913 ( .B1(n13195), .B2(n8134), .A(n8131), .ZN(n14329) );
  AOI21_X1 U8914 ( .B1(n8135), .B2(n8133), .A(n8132), .ZN(n8131) );
  INV_X1 U8915 ( .A(n8135), .ZN(n8134) );
  INV_X1 U8916 ( .A(n14237), .ZN(n8132) );
  NAND2_X1 U8917 ( .A1(n14329), .A2(n14330), .ZN(n14328) );
  NAND2_X1 U8918 ( .A1(n12629), .A2(n12630), .ZN(n12779) );
  NAND2_X1 U8919 ( .A1(n12628), .A2(n12627), .ZN(n12629) );
  NAND2_X1 U8920 ( .A1(n11654), .A2(n11653), .ZN(n11963) );
  OR2_X1 U8921 ( .A1(n14297), .A2(n14604), .ZN(n14320) );
  NAND2_X1 U8922 ( .A1(n11504), .A2(n11503), .ZN(n14297) );
  INV_X1 U8923 ( .A(n14326), .ZN(n14352) );
  AND2_X1 U8924 ( .A1(n11518), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14332) );
  OR2_X1 U8925 ( .A1(n10840), .A2(n10841), .ZN(n10842) );
  OAI21_X1 U8926 ( .B1(n10932), .B2(n8231), .A(n8230), .ZN(n8229) );
  NAND2_X1 U8927 ( .A1(n10930), .A2(n10925), .ZN(n8231) );
  AOI21_X1 U8928 ( .B1(n10930), .B2(n7504), .A(n13001), .ZN(n8230) );
  AND4_X1 U8929 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n12247) );
  NAND2_X1 U8930 ( .A1(n9966), .A2(n9965), .ZN(n14387) );
  AND2_X1 U8931 ( .A1(n9995), .A2(n10006), .ZN(n14391) );
  OAI21_X1 U8932 ( .B1(n13213), .B2(n10845), .A(n10844), .ZN(n14447) );
  NAND2_X1 U8933 ( .A1(n7784), .A2(n7786), .ZN(n10665) );
  NAND2_X1 U8934 ( .A1(n7787), .A2(n7792), .ZN(n7786) );
  AND2_X1 U8935 ( .A1(n10332), .A2(n10688), .ZN(n14455) );
  NAND2_X1 U8936 ( .A1(n14489), .A2(n10369), .ZN(n14474) );
  AND2_X1 U8937 ( .A1(n8336), .A2(n8334), .ZN(n14487) );
  NAND2_X1 U8938 ( .A1(n8336), .A2(n8340), .ZN(n14488) );
  NOR2_X1 U8939 ( .A1(n8275), .A2(n8274), .ZN(n14507) );
  NAND2_X1 U8940 ( .A1(n8276), .A2(n10367), .ZN(n14508) );
  OR2_X1 U8941 ( .A1(n14545), .A2(n14544), .ZN(n14686) );
  NAND2_X1 U8942 ( .A1(n14623), .A2(n8343), .ZN(n14591) );
  OAI21_X1 U8943 ( .B1(n13090), .B2(n7780), .A(n7453), .ZN(n14635) );
  NAND2_X1 U8944 ( .A1(n13088), .A2(n10187), .ZN(n14637) );
  AND2_X1 U8945 ( .A1(n8292), .A2(n7495), .ZN(n13086) );
  NAND2_X1 U8946 ( .A1(n10356), .A2(n10355), .ZN(n12908) );
  AND2_X1 U8947 ( .A1(n16574), .A2(n10156), .ZN(n12913) );
  NAND2_X1 U8948 ( .A1(n8311), .A2(n10135), .ZN(n12706) );
  NAND2_X1 U8949 ( .A1(n7771), .A2(n10115), .ZN(n12593) );
  NAND2_X1 U8950 ( .A1(n10094), .A2(n10093), .ZN(n12463) );
  NAND2_X1 U8951 ( .A1(n12125), .A2(n10078), .ZN(n12204) );
  INV_X1 U8952 ( .A(n14621), .ZN(n16599) );
  NAND2_X1 U8953 ( .A1(n11695), .A2(n11703), .ZN(n11697) );
  NAND2_X1 U8954 ( .A1(n11610), .A2(n10018), .ZN(n11695) );
  NAND2_X1 U8955 ( .A1(n11670), .A2(n9991), .ZN(n11682) );
  AND2_X1 U8956 ( .A1(n16591), .A2(n14654), .ZN(n7854) );
  AOI22_X1 U8957 ( .A1(n10215), .A2(n15846), .B1(n7522), .B2(n11300), .ZN(
        n9983) );
  INV_X1 U8958 ( .A(n14434), .ZN(n14728) );
  AND2_X1 U8959 ( .A1(n16595), .A2(n14654), .ZN(n7855) );
  INV_X1 U8960 ( .A(n14447), .ZN(n14732) );
  INV_X1 U8961 ( .A(n14527), .ZN(n14752) );
  INV_X1 U8962 ( .A(n11701), .ZN(n12071) );
  NAND2_X1 U8963 ( .A1(n16595), .A2(n16418), .ZN(n14764) );
  INV_X1 U8964 ( .A(n15823), .ZN(n15820) );
  INV_X1 U8965 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14770) );
  INV_X1 U8966 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9938) );
  INV_X1 U8967 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U8968 ( .A1(n9928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8270) );
  XNOR2_X1 U8969 ( .A(n10389), .B(n10388), .ZN(n14788) );
  NAND2_X1 U8970 ( .A1(n10390), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10389) );
  OAI21_X1 U8971 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(n14790) );
  INV_X1 U8972 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13003) );
  INV_X1 U8973 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12807) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11902) );
  INV_X1 U8975 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11719) );
  INV_X1 U8976 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11547) );
  INV_X1 U8977 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11440) );
  INV_X1 U8978 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n11213) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n11252) );
  INV_X1 U8980 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n11211) );
  INV_X1 U8981 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n11249) );
  INV_X1 U8982 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8454) );
  INV_X1 U8983 ( .A(n14938), .ZN(n12166) );
  NAND2_X1 U8984 ( .A1(n14795), .A2(n7755), .ZN(n14797) );
  NAND2_X1 U8985 ( .A1(n14894), .A2(n7756), .ZN(n7755) );
  NOR2_X1 U8986 ( .A1(n14796), .A2(n13301), .ZN(n7756) );
  INV_X1 U8987 ( .A(n11016), .ZN(n7740) );
  NAND2_X1 U8988 ( .A1(n12883), .A2(n12884), .ZN(n7741) );
  NOR2_X1 U8989 ( .A1(n11711), .A2(n11712), .ZN(n11710) );
  AOI21_X1 U8990 ( .B1(n8199), .B2(n13301), .A(n13312), .ZN(n8197) );
  NAND2_X1 U8991 ( .A1(n13253), .A2(n13252), .ZN(n14828) );
  CLKBUF_X1 U8992 ( .A(n11882), .Z(n11887) );
  INV_X1 U8993 ( .A(n14936), .ZN(n12888) );
  NAND2_X1 U8994 ( .A1(n7713), .A2(n9450), .ZN(n13176) );
  NAND2_X1 U8995 ( .A1(n7714), .A2(n9820), .ZN(n7713) );
  NAND2_X1 U8996 ( .A1(n11016), .A2(n7742), .ZN(n7739) );
  NAND2_X1 U8997 ( .A1(n11592), .A2(n7477), .ZN(n11599) );
  NOR2_X1 U8998 ( .A1(n11108), .A2(n11107), .ZN(n14899) );
  NAND2_X1 U8999 ( .A1(n11095), .A2(n11094), .ZN(n16549) );
  INV_X1 U9000 ( .A(n14937), .ZN(n12570) );
  NAND2_X1 U9001 ( .A1(n14895), .A2(n14896), .ZN(n14894) );
  NOR2_X1 U9002 ( .A1(n7484), .A2(n7750), .ZN(n7745) );
  INV_X1 U9003 ( .A(n14830), .ZN(n14925) );
  NAND4_X1 U9004 ( .A1(n9397), .A2(n9396), .A3(n9395), .A4(n9394), .ZN(n14933)
         );
  OR2_X1 U9005 ( .A1(n7439), .A2(n11153), .ZN(n9195) );
  OR2_X1 U9006 ( .A1(n7433), .A2(n14962), .ZN(n9176) );
  NAND2_X1 U9007 ( .A1(n9822), .A2(n9821), .ZN(n15262) );
  INV_X1 U9008 ( .A(n15065), .ZN(n15674) );
  AOI21_X1 U9009 ( .B1(n10660), .B2(n16498), .A(n10659), .ZN(n10661) );
  AOI21_X1 U9010 ( .B1(n15081), .B2(n16631), .A(n15080), .ZN(n15688) );
  NAND2_X1 U9011 ( .A1(n8241), .A2(n10573), .ZN(n15095) );
  NAND2_X1 U9012 ( .A1(n14789), .A2(n9820), .ZN(n9703) );
  NAND2_X1 U9013 ( .A1(n8166), .A2(n8165), .ZN(n15128) );
  AND2_X1 U9014 ( .A1(n8166), .A2(n7472), .ZN(n15129) );
  INV_X1 U9015 ( .A(n10572), .ZN(n7706) );
  NAND2_X1 U9016 ( .A1(n15141), .A2(n15151), .ZN(n7707) );
  INV_X1 U9017 ( .A(n10645), .ZN(n15726) );
  NAND2_X1 U9018 ( .A1(n15177), .A2(n10569), .ZN(n15158) );
  NAND2_X1 U9019 ( .A1(n15183), .A2(n10633), .ZN(n15155) );
  AND2_X1 U9020 ( .A1(n15210), .A2(n10568), .ZN(n15193) );
  NAND2_X1 U9021 ( .A1(n15229), .A2(n10567), .ZN(n15212) );
  NAND2_X1 U9022 ( .A1(n8179), .A2(n10631), .ZN(n15209) );
  NAND2_X1 U9023 ( .A1(n15257), .A2(n8185), .ZN(n8179) );
  NAND2_X1 U9024 ( .A1(n15257), .A2(n10629), .ZN(n15228) );
  INV_X1 U9025 ( .A(n7951), .ZN(n15253) );
  NAND2_X1 U9026 ( .A1(n7694), .A2(n7698), .ZN(n15249) );
  NAND2_X1 U9027 ( .A1(n16620), .A2(n7700), .ZN(n7694) );
  OAI21_X1 U9028 ( .B1(n12954), .B2(n8174), .A(n8170), .ZN(n13120) );
  NAND2_X1 U9029 ( .A1(n8169), .A2(n8177), .ZN(n13121) );
  NAND2_X1 U9030 ( .A1(n16619), .A2(n10562), .ZN(n13119) );
  NAND2_X1 U9031 ( .A1(n9467), .A2(n9466), .ZN(n16561) );
  INV_X1 U9032 ( .A(n16498), .ZN(n16644) );
  INV_X1 U9033 ( .A(n16493), .ZN(n16389) );
  NAND2_X1 U9034 ( .A1(n11412), .A2(n13032), .ZN(n16324) );
  NAND2_X1 U9035 ( .A1(n15683), .A2(n7507), .ZN(n15773) );
  AND2_X1 U9036 ( .A1(n10957), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10600) );
  NOR2_X1 U9037 ( .A1(n9111), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n9108) );
  XNOR2_X1 U9038 ( .A(n9784), .B(n9783), .ZN(n15796) );
  AOI21_X1 U9039 ( .B1(n7759), .B2(n7761), .A(n7530), .ZN(n7757) );
  NAND2_X1 U9040 ( .A1(n9899), .A2(n9898), .ZN(n15807) );
  NAND2_X1 U9041 ( .A1(n9904), .A2(n9903), .ZN(n13205) );
  NAND2_X1 U9042 ( .A1(n9657), .A2(n8267), .ZN(n9681) );
  NAND2_X1 U9043 ( .A1(n9588), .A2(n10252), .ZN(n8267) );
  XNOR2_X1 U9044 ( .A(n9589), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15811) );
  INV_X1 U9045 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12810) );
  INV_X1 U9046 ( .A(n10646), .ZN(n12808) );
  AOI21_X1 U9047 ( .B1(n9125), .B2(n15663), .A(n7761), .ZN(n8201) );
  INV_X1 U9048 ( .A(n9126), .ZN(n9125) );
  NAND2_X1 U9049 ( .A1(n8008), .A2(n9569), .ZN(n9570) );
  NAND2_X1 U9050 ( .A1(n8222), .A2(n9569), .ZN(n9545) );
  INV_X1 U9051 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11900) );
  INV_X1 U9052 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11717) );
  INV_X1 U9053 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11545) );
  AOI21_X1 U9054 ( .B1(n7718), .B2(n7720), .A(n7717), .ZN(n7716) );
  INV_X1 U9055 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n11346) );
  INV_X1 U9056 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n11291) );
  OAI21_X1 U9057 ( .B1(n9372), .B2(n9373), .A(n9399), .ZN(n11287) );
  INV_X1 U9058 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n11246) );
  INV_X1 U9059 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n11288) );
  AND2_X1 U9060 ( .A1(n9225), .A2(n9235), .ZN(n9210) );
  NOR2_X1 U9061 ( .A1(n15938), .A2(n15937), .ZN(n15940) );
  XNOR2_X1 U9062 ( .A(n15956), .B(n14402), .ZN(n15958) );
  INV_X1 U9063 ( .A(n8038), .ZN(n16026) );
  OR2_X1 U9064 ( .A1(n16020), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8034) );
  AND2_X1 U9065 ( .A1(n16020), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9066 ( .A1(n7685), .A2(n7686), .ZN(n16030) );
  OR2_X1 U9067 ( .A1(n16018), .A2(n16019), .ZN(n7685) );
  OAI21_X1 U9068 ( .B1(n16035), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7478), .ZN(
        n8029) );
  XNOR2_X1 U9069 ( .A(n16076), .B(n8040), .ZN(n16075) );
  INV_X1 U9070 ( .A(n16077), .ZN(n8040) );
  OR2_X1 U9071 ( .A1(n13546), .A2(n13545), .ZN(n7794) );
  INV_X1 U9072 ( .A(n8018), .ZN(n16124) );
  AND2_X1 U9073 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  NAND2_X1 U9074 ( .A1(n10423), .A2(n16615), .ZN(n9076) );
  AOI21_X1 U9075 ( .B1(n10423), .B2(n16618), .A(n10422), .ZN(n10424) );
  OAI21_X1 U9076 ( .B1(n13823), .B2(n14207), .A(n10421), .ZN(n10422) );
  AOI211_X1 U9077 ( .C1(n14676), .C2(n14324), .A(n14323), .B(n14322), .ZN(
        n14325) );
  INV_X1 U9078 ( .A(n10693), .ZN(n10694) );
  OR2_X1 U9079 ( .A1(n16591), .A2(n10379), .ZN(n7772) );
  NAND2_X1 U9080 ( .A1(n7774), .A2(n16591), .ZN(n7773) );
  NAND2_X1 U9081 ( .A1(n8319), .A2(n7590), .ZN(n7774) );
  NOR2_X1 U9082 ( .A1(n10418), .A2(n10417), .ZN(n10419) );
  NOR2_X1 U9083 ( .A1(n7596), .A2(n7595), .ZN(n7594) );
  NOR2_X1 U9084 ( .A1(n16591), .A2(n14663), .ZN(n7595) );
  OAI211_X1 U9085 ( .C1(n8319), .C2(n16592), .A(n8317), .B(n8320), .ZN(
        P2_U3496) );
  INV_X1 U9086 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8321) );
  OR4_X1 U9087 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(
        P1_U3233) );
  OAI211_X1 U9088 ( .C1(n15694), .C2(n15247), .A(n8011), .B(n8010), .ZN(
        P1_U3266) );
  AOI21_X1 U9089 ( .B1(n15690), .B2(n16498), .A(n13230), .ZN(n8011) );
  OR2_X1 U9090 ( .A1(n15693), .A2(n16398), .ZN(n8010) );
  NAND2_X1 U9091 ( .A1(n15268), .A2(n15267), .ZN(n15672) );
  NAND2_X1 U9092 ( .A1(n7693), .A2(n7692), .ZN(P1_U3525) );
  NAND2_X1 U9093 ( .A1(n16636), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9094 ( .A1(n15773), .A2(n16638), .ZN(n7693) );
  NOR2_X1 U9095 ( .A1(n16092), .A2(n16091), .ZN(n16090) );
  INV_X1 U9096 ( .A(n8026), .ZN(n16000) );
  AND2_X1 U9097 ( .A1(n8033), .A2(n8039), .ZN(n16021) );
  OAI21_X1 U9098 ( .B1(n8039), .B2(n16020), .A(n8030), .ZN(n16022) );
  INV_X1 U9099 ( .A(n8042), .ZN(n16068) );
  MUX2_X2 U9100 ( .A(n10646), .B(n7436), .S(n9812), .Z(n9260) );
  OAI21_X1 U9101 ( .B1(n9260), .B2(n7943), .A(n7616), .ZN(n9287) );
  INV_X1 U9102 ( .A(n9287), .ZN(n8259) );
  AND2_X1 U9103 ( .A1(n13471), .A2(n13472), .ZN(n13881) );
  INV_X1 U9104 ( .A(n13881), .ZN(n7935) );
  AND2_X1 U9105 ( .A1(n10809), .A2(n7875), .ZN(n7451) );
  AND2_X1 U9106 ( .A1(n9451), .A2(n9453), .ZN(n7452) );
  NAND2_X2 U9107 ( .A1(n14609), .A2(n11485), .ZN(n11490) );
  AND2_X1 U9108 ( .A1(n14636), .A2(n7779), .ZN(n7453) );
  INV_X1 U9109 ( .A(n15256), .ZN(n7696) );
  INV_X1 U9110 ( .A(n10563), .ZN(n8228) );
  OAI211_X1 U9111 ( .C1(P3_IR_REG_2__SCAN_IN), .C2(P3_IR_REG_31__SCAN_IN), .A(
        n8025), .B(n8024), .ZN(n11771) );
  AND2_X1 U9112 ( .A1(n14736), .A2(n10920), .ZN(n7454) );
  AND2_X1 U9113 ( .A1(n11083), .A2(n8195), .ZN(n7455) );
  AND2_X1 U9114 ( .A1(n7527), .A2(n7619), .ZN(n7456) );
  NOR2_X1 U9115 ( .A1(n13231), .A2(n13234), .ZN(n7457) );
  INV_X1 U9116 ( .A(n14498), .ZN(n10368) );
  INV_X1 U9117 ( .A(n15213), .ZN(n8184) );
  OR2_X1 U9118 ( .A1(n7926), .A2(n14084), .ZN(n7458) );
  AND2_X1 U9119 ( .A1(n10820), .A2(n7886), .ZN(n7459) );
  OR2_X1 U9120 ( .A1(n15711), .A2(n14843), .ZN(n7460) );
  XNOR2_X1 U9121 ( .A(n13176), .B(n14931), .ZN(n12836) );
  INV_X1 U9122 ( .A(n12836), .ZN(n8236) );
  AND2_X1 U9123 ( .A1(n12153), .A2(n8299), .ZN(n7461) );
  OR2_X1 U9124 ( .A1(n15966), .A2(n15965), .ZN(n7462) );
  NAND2_X1 U9125 ( .A1(n7765), .A2(n8194), .ZN(n11096) );
  NAND2_X1 U9126 ( .A1(n13265), .A2(n14878), .ZN(n14805) );
  INV_X1 U9127 ( .A(n14467), .ZN(n14740) );
  NAND2_X1 U9128 ( .A1(n14467), .A2(n14367), .ZN(n7792) );
  INV_X1 U9129 ( .A(n7792), .ZN(n7782) );
  NAND2_X1 U9130 ( .A1(n12189), .A2(n14938), .ZN(n7463) );
  NAND2_X1 U9131 ( .A1(n10306), .A2(n10305), .ZN(n14453) );
  INV_X1 U9132 ( .A(n14453), .ZN(n14736) );
  INV_X1 U9133 ( .A(n9493), .ZN(n7614) );
  AND2_X1 U9134 ( .A1(n9728), .A2(n9730), .ZN(n7465) );
  INV_X1 U9135 ( .A(n10811), .ZN(n7875) );
  INV_X1 U9136 ( .A(n10560), .ZN(n12963) );
  AND2_X1 U9137 ( .A1(n13924), .A2(n8791), .ZN(n7466) );
  OR2_X2 U9138 ( .A1(n11491), .A2(n10848), .ZN(n11533) );
  OAI211_X1 U9139 ( .C1(n8558), .C2(n8838), .A(n8837), .B(n8836), .ZN(n13914)
         );
  NAND2_X1 U9140 ( .A1(n13140), .A2(n13142), .ZN(n13141) );
  NAND2_X1 U9141 ( .A1(n13040), .A2(n13042), .ZN(n13041) );
  NAND2_X1 U9142 ( .A1(n7951), .A2(n7950), .ZN(n15252) );
  INV_X1 U9143 ( .A(n15252), .ZN(n7949) );
  INV_X1 U9144 ( .A(n12463), .ZN(n7847) );
  INV_X1 U9145 ( .A(n12928), .ZN(n7947) );
  OR2_X1 U9146 ( .A1(n16595), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7467) );
  OR2_X1 U9147 ( .A1(n16591), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7468) );
  AND2_X1 U9148 ( .A1(n10551), .A2(n10550), .ZN(n7469) );
  INV_X1 U9149 ( .A(n12189), .ZN(n7943) );
  INV_X1 U9150 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7761) );
  INV_X1 U9151 ( .A(n10643), .ZN(n13305) );
  NAND2_X2 U9152 ( .A1(n10958), .A2(n10642), .ZN(n10643) );
  INV_X1 U9153 ( .A(n7849), .ZN(n12421) );
  OAI21_X2 U9154 ( .B1(n11251), .B2(n10845), .A(n10081), .ZN(n7849) );
  INV_X2 U9155 ( .A(n8558), .ZN(n8833) );
  AND4_X1 U9156 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n8463), .ZN(n10438)
         );
  NAND2_X1 U9157 ( .A1(n11977), .A2(n11978), .ZN(n7470) );
  AND4_X1 U9159 ( .A1(n9116), .A2(n9085), .A3(n9084), .A4(n9890), .ZN(n7471)
         );
  NAND2_X1 U9160 ( .A1(n14858), .A2(n11072), .ZN(n14816) );
  INV_X2 U9161 ( .A(n7439), .ZN(n9248) );
  NAND2_X1 U9162 ( .A1(n15718), .A2(n14924), .ZN(n7472) );
  AND2_X1 U9163 ( .A1(n8241), .A2(n8239), .ZN(n7473) );
  INV_X1 U9164 ( .A(n9854), .ZN(n15175) );
  NOR2_X1 U9165 ( .A1(n14736), .A2(n10920), .ZN(n7474) );
  AND2_X1 U9166 ( .A1(n9443), .A2(n9438), .ZN(n7475) );
  AND2_X1 U9167 ( .A1(n8237), .A2(n10574), .ZN(n7476) );
  OR2_X1 U9168 ( .A1(n10967), .A2(n10966), .ZN(n7477) );
  INV_X1 U9169 ( .A(n13050), .ZN(n13067) );
  NAND2_X1 U9170 ( .A1(n10160), .A2(n10159), .ZN(n13050) );
  OR2_X1 U9171 ( .A1(n15150), .A2(n15151), .ZN(n8166) );
  OR2_X1 U9172 ( .A1(n16034), .A2(n16033), .ZN(n7478) );
  XNOR2_X1 U9173 ( .A(n15123), .B(n14923), .ZN(n15118) );
  INV_X1 U9174 ( .A(n15118), .ZN(n10636) );
  AND2_X1 U9175 ( .A1(n12849), .A2(n8517), .ZN(n7479) );
  AND2_X1 U9176 ( .A1(n16550), .A2(n11054), .ZN(n7480) );
  AND3_X1 U9177 ( .A1(n9102), .A2(n9101), .A3(n9100), .ZN(n7481) );
  NAND2_X1 U9178 ( .A1(n13903), .A2(n13914), .ZN(n7482) );
  AND2_X1 U9179 ( .A1(n9968), .A2(n9967), .ZN(n7483) );
  NAND2_X1 U9180 ( .A1(n9984), .A2(n9983), .ZN(n11679) );
  AND2_X1 U9181 ( .A1(n11054), .A2(n7751), .ZN(n7484) );
  OAI21_X1 U9182 ( .B1(n8178), .B2(n9796), .A(n9215), .ZN(n16390) );
  INV_X1 U9183 ( .A(n16390), .ZN(n9860) );
  AND2_X1 U9184 ( .A1(n14467), .A2(n14266), .ZN(n7485) );
  NAND2_X1 U9185 ( .A1(n14676), .A2(n14535), .ZN(n7486) );
  AND2_X1 U9186 ( .A1(n7460), .A2(n15151), .ZN(n7487) );
  NAND2_X1 U9187 ( .A1(n14826), .A2(n13258), .ZN(n14877) );
  OR2_X1 U9188 ( .A1(n16197), .A2(n13726), .ZN(n7488) );
  AND2_X1 U9189 ( .A1(n9895), .A2(n7762), .ZN(n7489) );
  AND2_X1 U9190 ( .A1(n8251), .A2(n7632), .ZN(n7490) );
  INV_X1 U9191 ( .A(n14922), .ZN(n15112) );
  NAND2_X1 U9192 ( .A1(n11006), .A2(n11005), .ZN(n7491) );
  INV_X1 U9193 ( .A(n13496), .ZN(n8054) );
  AND2_X1 U9194 ( .A1(n14716), .A2(n14373), .ZN(n7492) );
  INV_X1 U9195 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7942) );
  INV_X1 U9196 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9082) );
  AND2_X1 U9197 ( .A1(n13481), .A2(n13482), .ZN(n13360) );
  NAND2_X1 U9198 ( .A1(n10288), .A2(n10287), .ZN(n14480) );
  INV_X1 U9199 ( .A(n14480), .ZN(n14744) );
  NAND2_X1 U9200 ( .A1(n10875), .A2(n10874), .ZN(n14434) );
  NAND2_X1 U9201 ( .A1(n10228), .A2(n10227), .ZN(n14698) );
  OR2_X1 U9202 ( .A1(n15748), .A2(n15235), .ZN(n7493) );
  OR2_X1 U9203 ( .A1(n15131), .A2(n15123), .ZN(n7494) );
  NAND2_X1 U9204 ( .A1(n13050), .A2(n10357), .ZN(n7495) );
  INV_X1 U9205 ( .A(n11962), .ZN(n8105) );
  INV_X1 U9206 ( .A(n9706), .ZN(n7633) );
  NAND2_X1 U9207 ( .A1(n12891), .A2(n12925), .ZN(n7496) );
  INV_X1 U9208 ( .A(n9509), .ZN(n8262) );
  INV_X1 U9209 ( .A(n10759), .ZN(n7602) );
  AND2_X1 U9210 ( .A1(n15711), .A2(n14843), .ZN(n7497) );
  INV_X1 U9211 ( .A(n9775), .ZN(n8224) );
  AND2_X1 U9212 ( .A1(n13639), .A2(n7963), .ZN(n7498) );
  AND2_X1 U9213 ( .A1(n7849), .A2(n14379), .ZN(n7499) );
  AND2_X1 U9214 ( .A1(n8100), .A2(n7470), .ZN(n7500) );
  OR2_X1 U9215 ( .A1(n13050), .A2(n10357), .ZN(n7501) );
  AND2_X1 U9216 ( .A1(n16419), .A2(n12079), .ZN(n7502) );
  INV_X1 U9217 ( .A(n12920), .ZN(n7742) );
  INV_X1 U9218 ( .A(n8177), .ZN(n8174) );
  AND2_X1 U9219 ( .A1(n13521), .A2(n12971), .ZN(n7503) );
  AND2_X1 U9220 ( .A1(n10926), .A2(n10937), .ZN(n7504) );
  NAND2_X1 U9221 ( .A1(n8294), .A2(n7859), .ZN(n7861) );
  INV_X1 U9222 ( .A(n7701), .ZN(n7700) );
  NAND2_X1 U9223 ( .A1(n10565), .A2(n16625), .ZN(n7701) );
  INV_X1 U9224 ( .A(n7658), .ZN(n7655) );
  NAND2_X1 U9225 ( .A1(n7659), .A2(n7660), .ZN(n7658) );
  AND2_X1 U9226 ( .A1(n12289), .A2(n12288), .ZN(n7505) );
  NAND2_X1 U9227 ( .A1(n10697), .A2(n14387), .ZN(n7506) );
  INV_X1 U9228 ( .A(n7873), .ZN(n7872) );
  OAI21_X1 U9229 ( .B1(n7874), .B2(n8376), .A(n10812), .ZN(n7873) );
  INV_X1 U9230 ( .A(n9574), .ZN(n8255) );
  AND2_X1 U9231 ( .A1(n15682), .A2(n8395), .ZN(n7507) );
  AND2_X1 U9232 ( .A1(n14594), .A2(n14579), .ZN(n7508) );
  NAND2_X1 U9233 ( .A1(n7765), .A2(n7764), .ZN(n13253) );
  NOR2_X1 U9234 ( .A1(n16231), .A2(n13731), .ZN(n7509) );
  AND2_X1 U9235 ( .A1(n13639), .A2(n10500), .ZN(n7510) );
  INV_X1 U9236 ( .A(n7791), .ZN(n7790) );
  NOR2_X1 U9237 ( .A1(n14744), .A2(n14312), .ZN(n7791) );
  AND2_X1 U9238 ( .A1(n8396), .A2(n9195), .ZN(n7511) );
  INV_X1 U9239 ( .A(n7938), .ZN(n13883) );
  NAND2_X1 U9240 ( .A1(n7934), .A2(n7935), .ZN(n7938) );
  INV_X1 U9241 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7608) );
  AND2_X1 U9242 ( .A1(n8146), .A2(n15502), .ZN(n7512) );
  OR2_X1 U9243 ( .A1(n12111), .A2(n12110), .ZN(n7513) );
  INV_X1 U9244 ( .A(SI_2_), .ZN(n15308) );
  NOR2_X1 U9245 ( .A1(n15711), .A2(n15114), .ZN(n7514) );
  NOR2_X1 U9246 ( .A1(n11090), .A2(n11089), .ZN(n7515) );
  NAND2_X1 U9247 ( .A1(n10211), .A2(n10210), .ZN(n14623) );
  NAND2_X1 U9248 ( .A1(n7481), .A2(n9106), .ZN(n14943) );
  AND2_X1 U9249 ( .A1(n12770), .A2(n12702), .ZN(n7516) );
  INV_X1 U9250 ( .A(n10504), .ZN(n7967) );
  AND2_X1 U9251 ( .A1(n7881), .A2(n7879), .ZN(n7517) );
  NOR2_X1 U9252 ( .A1(n10484), .A2(n13965), .ZN(n7518) );
  INV_X1 U9253 ( .A(n8389), .ZN(n7931) );
  INV_X1 U9254 ( .A(n7738), .ZN(n7737) );
  NAND2_X1 U9255 ( .A1(n7742), .A2(n12884), .ZN(n7738) );
  INV_X1 U9256 ( .A(n10286), .ZN(n8333) );
  OR2_X1 U9257 ( .A1(n8902), .A2(n8901), .ZN(n7519) );
  INV_X1 U9258 ( .A(n7860), .ZN(n7859) );
  NAND2_X1 U9259 ( .A1(n10368), .A2(n14744), .ZN(n7860) );
  AND2_X1 U9260 ( .A1(n8323), .A2(n8322), .ZN(n7520) );
  NAND2_X1 U9261 ( .A1(n10254), .A2(n10253), .ZN(n14551) );
  INV_X1 U9262 ( .A(n14551), .ZN(n7856) );
  INV_X1 U9263 ( .A(n8186), .ZN(n8185) );
  OR2_X1 U9264 ( .A1(n10630), .A2(n8187), .ZN(n8186) );
  NAND2_X1 U9265 ( .A1(n8861), .A2(n7935), .ZN(n7521) );
  AND2_X1 U9266 ( .A1(n9930), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7522) );
  AND2_X1 U9267 ( .A1(n11249), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7523) );
  AND2_X1 U9268 ( .A1(n13458), .A2(n13906), .ZN(n13931) );
  INV_X1 U9269 ( .A(n13931), .ZN(n13924) );
  NAND2_X1 U9270 ( .A1(n14805), .A2(n14807), .ZN(n14806) );
  AND2_X1 U9271 ( .A1(n7787), .A2(n7781), .ZN(n7524) );
  OR2_X1 U9272 ( .A1(n7875), .A2(n10809), .ZN(n7525) );
  INV_X1 U9273 ( .A(n10809), .ZN(n8376) );
  AND2_X1 U9274 ( .A1(n13360), .A2(n8896), .ZN(n7526) );
  OR2_X1 U9275 ( .A1(n9453), .A2(n9451), .ZN(n7527) );
  OR2_X1 U9276 ( .A1(n9508), .A2(n8262), .ZN(n7528) );
  OR2_X1 U9277 ( .A1(n10572), .A2(n7497), .ZN(n7529) );
  AND2_X1 U9278 ( .A1(n7763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U9279 ( .A1(n15210), .A2(n7712), .ZN(n15173) );
  AND2_X1 U9280 ( .A1(n10619), .A2(n7496), .ZN(n7531) );
  INV_X1 U9281 ( .A(n8171), .ZN(n8170) );
  NAND2_X1 U9282 ( .A1(n8228), .A2(n8172), .ZN(n8171) );
  INV_X1 U9283 ( .A(n9494), .ZN(n7612) );
  INV_X1 U9284 ( .A(n10833), .ZN(n7892) );
  AND2_X1 U9285 ( .A1(n8582), .A2(n8568), .ZN(n7532) );
  INV_X1 U9286 ( .A(n10723), .ZN(n8380) );
  OR2_X1 U9287 ( .A1(n14480), .A2(n14312), .ZN(n7533) );
  OR2_X1 U9288 ( .A1(n16159), .A2(n13722), .ZN(n7534) );
  AND2_X1 U9289 ( .A1(n12770), .A2(n12772), .ZN(n7535) );
  AND2_X1 U9290 ( .A1(n7707), .A2(n7706), .ZN(n7536) );
  NAND2_X1 U9291 ( .A1(n9773), .A2(n9772), .ZN(n15686) );
  AND2_X1 U9292 ( .A1(n7526), .A2(n13979), .ZN(n7537) );
  NOR2_X1 U9293 ( .A1(n13873), .A2(n13477), .ZN(n7538) );
  INV_X1 U9294 ( .A(n16310), .ZN(n9115) );
  NAND2_X1 U9295 ( .A1(n9462), .A2(n9461), .ZN(n9484) );
  AND2_X1 U9296 ( .A1(n7858), .A2(n14736), .ZN(n7539) );
  NOR2_X1 U9297 ( .A1(n11969), .A2(n8103), .ZN(n8102) );
  AND2_X1 U9298 ( .A1(n8296), .A2(n8295), .ZN(n7540) );
  NOR2_X1 U9299 ( .A1(n15213), .A2(n8225), .ZN(n7541) );
  OR2_X1 U9300 ( .A1(n11724), .A2(n11772), .ZN(n7542) );
  AND2_X1 U9301 ( .A1(n10570), .A2(n10569), .ZN(n7543) );
  AND2_X1 U9302 ( .A1(n12071), .A2(n7851), .ZN(n7544) );
  INV_X1 U9303 ( .A(n12781), .ZN(n7644) );
  INV_X1 U9304 ( .A(n9418), .ZN(n7720) );
  AND2_X1 U9305 ( .A1(n7482), .A2(n10488), .ZN(n7545) );
  OR2_X1 U9306 ( .A1(n9358), .A2(n9356), .ZN(n7546) );
  AND2_X1 U9307 ( .A1(n12349), .A2(n12348), .ZN(n7547) );
  AND2_X1 U9308 ( .A1(n14623), .A2(n10212), .ZN(n7548) );
  INV_X1 U9309 ( .A(n7719), .ZN(n7718) );
  OAI21_X1 U9310 ( .B1(n7721), .B2(n7720), .A(n9435), .ZN(n7719) );
  AND2_X1 U9311 ( .A1(n13255), .A2(n13252), .ZN(n7549) );
  NOR2_X1 U9312 ( .A1(n12189), .A2(n14938), .ZN(n7550) );
  OR2_X1 U9313 ( .A1(n8255), .A2(n9573), .ZN(n7551) );
  OR2_X1 U9314 ( .A1(n10745), .A2(n10743), .ZN(n7552) );
  OR2_X1 U9315 ( .A1(n9407), .A2(n9405), .ZN(n7553) );
  OR2_X1 U9316 ( .A1(n7602), .A2(n10758), .ZN(n7554) );
  OR2_X1 U9317 ( .A1(n15175), .A2(n8149), .ZN(n7555) );
  AND2_X1 U9318 ( .A1(n7528), .A2(n7613), .ZN(n7556) );
  OR2_X1 U9319 ( .A1(n8224), .A2(n9774), .ZN(n7557) );
  INV_X1 U9320 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9922) );
  INV_X1 U9321 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8401) );
  INV_X1 U9322 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U9323 ( .A1(n15696), .A2(n14922), .ZN(n7558) );
  INV_X1 U9324 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n15437) );
  NAND2_X1 U9325 ( .A1(n12835), .A2(n8232), .ZN(n12965) );
  INV_X1 U9326 ( .A(n8498), .ZN(n8558) );
  OR2_X1 U9327 ( .A1(n8700), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7559) );
  NAND3_X1 U9328 ( .A1(n10320), .A2(n8144), .A3(n10178), .ZN(n7560) );
  OAI21_X1 U9329 ( .B1(n14082), .B2(n7907), .A(n7906), .ZN(n14067) );
  NAND2_X1 U9330 ( .A1(n13195), .A2(n13194), .ZN(n14231) );
  NAND2_X1 U9331 ( .A1(n13141), .A2(n11037), .ZN(n13167) );
  AND2_X1 U9332 ( .A1(n7741), .A2(n7740), .ZN(n12919) );
  INV_X1 U9333 ( .A(n9824), .ZN(n9825) );
  AND2_X1 U9334 ( .A1(n12551), .A2(n10558), .ZN(n12834) );
  AND2_X1 U9335 ( .A1(n8400), .A2(n8458), .ZN(n8563) );
  NOR2_X1 U9336 ( .A1(n8373), .A2(n10091), .ZN(n10384) );
  NAND2_X1 U9337 ( .A1(n7914), .A2(n8572), .ZN(n12984) );
  NAND2_X1 U9338 ( .A1(n14906), .A2(n11061), .ZN(n14848) );
  NAND2_X1 U9339 ( .A1(n12610), .A2(n10621), .ZN(n12609) );
  NAND2_X1 U9340 ( .A1(n16574), .A2(n8348), .ZN(n12911) );
  INV_X1 U9341 ( .A(n13985), .ZN(n13946) );
  NAND2_X1 U9342 ( .A1(n7905), .A2(n8791), .ZN(n13930) );
  NAND2_X1 U9343 ( .A1(n7736), .A2(n7739), .ZN(n13040) );
  NAND2_X1 U9344 ( .A1(n13677), .A2(n10483), .ZN(n13571) );
  NAND2_X1 U9345 ( .A1(n13958), .A2(n13957), .ZN(n7561) );
  OR2_X1 U9346 ( .A1(n11540), .A2(n12828), .ZN(n7562) );
  AND4_X1 U9347 ( .A1(n8806), .A2(n8805), .A3(n8804), .A4(n8803), .ZN(n13945)
         );
  INV_X1 U9348 ( .A(n13945), .ZN(n13915) );
  AND2_X1 U9349 ( .A1(n8137), .A2(n8135), .ZN(n7563) );
  AND2_X1 U9350 ( .A1(n16619), .A2(n8226), .ZN(n7564) );
  OR2_X1 U9351 ( .A1(n10176), .A2(n10175), .ZN(n7565) );
  AND2_X1 U9352 ( .A1(n9543), .A2(n15480), .ZN(n7566) );
  AND2_X1 U9353 ( .A1(n9482), .A2(n11411), .ZN(n7567) );
  INV_X1 U9354 ( .A(n10495), .ZN(n7958) );
  AND2_X1 U9355 ( .A1(n7958), .A2(n13596), .ZN(n7568) );
  INV_X1 U9356 ( .A(n10687), .ZN(n8322) );
  OAI21_X1 U9357 ( .B1(n10920), .B2(n14602), .A(n10686), .ZN(n10687) );
  AND2_X1 U9358 ( .A1(n8316), .A2(n8318), .ZN(n7569) );
  NAND2_X2 U9359 ( .A1(n12440), .A2(n14073), .ZN(n16340) );
  INV_X1 U9360 ( .A(n12142), .ZN(n8299) );
  NAND2_X1 U9361 ( .A1(n10151), .A2(n10150), .ZN(n16600) );
  INV_X1 U9362 ( .A(n16600), .ZN(n7846) );
  NAND2_X1 U9363 ( .A1(n9424), .A2(n9423), .ZN(n12813) );
  INV_X1 U9364 ( .A(n12813), .ZN(n7945) );
  NAND2_X1 U9365 ( .A1(n9527), .A2(n9526), .ZN(n15757) );
  INV_X1 U9366 ( .A(n15757), .ZN(n7950) );
  INV_X1 U9367 ( .A(n7850), .ZN(n12087) );
  INV_X1 U9368 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n8077) );
  INV_X2 U9369 ( .A(n16592), .ZN(n16595) );
  AND2_X1 U9370 ( .A1(n7461), .A2(n7848), .ZN(n7570) );
  NAND2_X1 U9371 ( .A1(n11993), .A2(n11994), .ZN(n11992) );
  NAND2_X1 U9372 ( .A1(n8099), .A2(n8100), .ZN(n12347) );
  NAND2_X1 U9373 ( .A1(n10544), .A2(n10543), .ZN(n16380) );
  INV_X1 U9374 ( .A(n10554), .ZN(n12615) );
  NAND2_X1 U9375 ( .A1(n10193), .A2(n10192), .ZN(n14716) );
  INV_X1 U9376 ( .A(n14716), .ZN(n8300) );
  AND2_X1 U9377 ( .A1(n11022), .A2(n11021), .ZN(n7571) );
  NAND2_X1 U9378 ( .A1(n10545), .A2(n12176), .ZN(n12177) );
  AND2_X1 U9379 ( .A1(n8104), .A2(n8102), .ZN(n7572) );
  OR2_X1 U9380 ( .A1(n11710), .A2(n10987), .ZN(n7573) );
  AND2_X1 U9381 ( .A1(n8018), .A2(n8017), .ZN(n7574) );
  NAND2_X1 U9382 ( .A1(n8247), .A2(n7496), .ZN(n7575) );
  OR2_X1 U9383 ( .A1(n13747), .A2(n16538), .ZN(n7576) );
  AND2_X1 U9384 ( .A1(n12226), .A2(n12310), .ZN(n7577) );
  AND2_X1 U9385 ( .A1(n12492), .A2(n8517), .ZN(n7578) );
  AND2_X1 U9386 ( .A1(n8290), .A2(n10346), .ZN(n7579) );
  AND2_X1 U9387 ( .A1(n7667), .A2(n12348), .ZN(n7580) );
  OR2_X1 U9388 ( .A1(n12158), .A2(n12157), .ZN(n16636) );
  INV_X2 U9389 ( .A(n16636), .ZN(n16638) );
  INV_X1 U9390 ( .A(n14084), .ZN(n13979) );
  AND2_X1 U9391 ( .A1(n9031), .A2(n13358), .ZN(n14084) );
  AOI21_X1 U9392 ( .B1(n13315), .B2(n14943), .A(n7726), .ZN(n11461) );
  NOR2_X1 U9393 ( .A1(n8384), .A2(n11927), .ZN(n11937) );
  INV_X1 U9394 ( .A(n11937), .ZN(n7837) );
  XNOR2_X1 U9395 ( .A(n10967), .B(n8188), .ZN(n11591) );
  NAND2_X1 U9396 ( .A1(n12002), .A2(n16401), .ZN(n12185) );
  INV_X1 U9397 ( .A(n12185), .ZN(n7944) );
  AND2_X1 U9398 ( .A1(n14609), .A2(n12148), .ZN(n14723) );
  INV_X1 U9399 ( .A(n14723), .ZN(n16588) );
  AND2_X1 U9400 ( .A1(n16032), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n7581) );
  INV_X1 U9401 ( .A(n7682), .ZN(n7681) );
  AOI21_X1 U9402 ( .B1(n7683), .B2(n16019), .A(n7581), .ZN(n7682) );
  XNOR2_X1 U9403 ( .A(n8778), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13736) );
  INV_X1 U9404 ( .A(n13736), .ZN(n13799) );
  INV_X1 U9405 ( .A(n8178), .ZN(n11191) );
  NAND2_X1 U9406 ( .A1(n9212), .A2(n9213), .ZN(n8178) );
  INV_X1 U9407 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U9408 ( .A1(n12413), .A2(n9030), .ZN(n13541) );
  INV_X1 U9409 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7593) );
  INV_X1 U9410 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7668) );
  INV_X1 U9411 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7687) );
  INV_X1 U9412 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7688) );
  INV_X1 U9413 ( .A(n16631), .ZN(n16351) );
  INV_X1 U9414 ( .A(n16560), .ZN(n16624) );
  NAND2_X1 U9415 ( .A1(n15262), .A2(n16560), .ZN(n15263) );
  OAI21_X2 U9416 ( .B1(n11092), .B2(n13032), .A(n16640), .ZN(n16560) );
  NAND3_X1 U9417 ( .A1(n7598), .A2(n10912), .A3(n7582), .ZN(n10882) );
  NAND2_X1 U9418 ( .A1(n10869), .A2(n7600), .ZN(n7599) );
  NAND2_X1 U9419 ( .A1(n8273), .A2(n8272), .ZN(n14491) );
  NAND2_X1 U9420 ( .A1(n7689), .A2(n9269), .ZN(n9273) );
  NAND2_X1 U9421 ( .A1(n9326), .A2(n9325), .ZN(n9330) );
  AOI21_X1 U9422 ( .B1(n8284), .B2(n8286), .A(n7535), .ZN(n8282) );
  OAI21_X1 U9423 ( .B1(n12456), .B2(n8286), .A(n10353), .ZN(n8285) );
  INV_X1 U9424 ( .A(n9142), .ZN(n9156) );
  NAND2_X1 U9425 ( .A1(n8283), .A2(n8282), .ZN(n12701) );
  NAND2_X1 U9426 ( .A1(n9232), .A2(n9233), .ZN(n9227) );
  NAND2_X1 U9427 ( .A1(n14341), .A2(n14340), .ZN(n14339) );
  XNOR2_X1 U9428 ( .A(n14252), .B(n14250), .ZN(n14341) );
  NOR2_X1 U9429 ( .A1(n15953), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n15954) );
  XNOR2_X1 U9430 ( .A(n15952), .B(n15951), .ZN(n15953) );
  NOR2_X1 U9431 ( .A1(n15988), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n15989) );
  XNOR2_X1 U9432 ( .A(n15986), .B(n15987), .ZN(n15988) );
  INV_X1 U9433 ( .A(n16014), .ZN(n7588) );
  INV_X1 U9434 ( .A(n8138), .ZN(n8133) );
  NOR2_X1 U9435 ( .A1(n16041), .A2(n16040), .ZN(n16042) );
  NOR2_X1 U9436 ( .A1(n16053), .A2(n16052), .ZN(n16054) );
  NOR2_X1 U9437 ( .A1(n16026), .A2(n16025), .ZN(n16029) );
  NAND2_X1 U9438 ( .A1(n15998), .A2(n15999), .ZN(n8028) );
  NAND2_X1 U9439 ( .A1(n7647), .A2(n7653), .ZN(n14350) );
  XNOR2_X1 U9440 ( .A(n8124), .B(n14294), .ZN(n14301) );
  NAND2_X1 U9441 ( .A1(n15948), .A2(n15947), .ZN(n8049) );
  INV_X1 U9442 ( .A(n16064), .ZN(n8044) );
  OAI21_X1 U9443 ( .B1(n10494), .B2(n10495), .A(n7956), .ZN(n10496) );
  INV_X1 U9444 ( .A(n13668), .ZN(n7957) );
  NAND2_X1 U9445 ( .A1(n8271), .A2(n16584), .ZN(n8323) );
  NAND2_X1 U9446 ( .A1(n10373), .A2(n10372), .ZN(n10677) );
  INV_X1 U9447 ( .A(n8285), .ZN(n8284) );
  NAND2_X1 U9448 ( .A1(n7773), .A2(n7772), .ZN(P2_U3528) );
  INV_X1 U9449 ( .A(n12081), .ZN(n10348) );
  NAND2_X1 U9450 ( .A1(n7597), .A2(n7594), .ZN(P2_U3526) );
  OR2_X1 U9451 ( .A1(n14737), .A2(n16589), .ZN(n7597) );
  NAND2_X1 U9452 ( .A1(n9227), .A2(n9236), .ZN(n9231) );
  INV_X1 U9453 ( .A(n8000), .ZN(n7996) );
  NAND2_X1 U9454 ( .A1(n7884), .A2(n7885), .ZN(n10823) );
  NAND3_X1 U9455 ( .A1(n10757), .A2(n10756), .A3(n7554), .ZN(n7603) );
  NAND2_X1 U9456 ( .A1(n10741), .A2(n10739), .ZN(n7894) );
  OAI22_X2 U9457 ( .A1(n10769), .A2(n7898), .B1(n10770), .B2(n7897), .ZN(
        n10774) );
  NAND2_X1 U9458 ( .A1(n7863), .A2(n7862), .ZN(n10793) );
  NAND2_X1 U9459 ( .A1(n8380), .A2(n10724), .ZN(n8378) );
  OAI22_X1 U9460 ( .A1(n10815), .A2(n8354), .B1(n10816), .B2(n8353), .ZN(
        n10819) );
  OAI22_X1 U9461 ( .A1(n8371), .A2(n8370), .B1(n10744), .B2(n8372), .ZN(n10747) );
  AND4_X2 U9462 ( .A1(n8006), .A2(n8401), .A3(n8005), .A4(n8458), .ZN(n8406)
         );
  XNOR2_X1 U9463 ( .A(n7607), .B(n7606), .ZN(n13796) );
  OAI21_X1 U9464 ( .B1(n13794), .B2(n13793), .A(n16257), .ZN(n7607) );
  INV_X2 U9465 ( .A(n13542), .ZN(n13791) );
  NOR2_X2 U9466 ( .A1(n9485), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U9467 ( .A1(n7610), .A2(n7556), .ZN(n8260) );
  NAND3_X1 U9468 ( .A1(n9475), .A2(n7611), .A3(n9474), .ZN(n7610) );
  NAND3_X1 U9469 ( .A1(n9268), .A2(n9267), .A3(n7615), .ZN(n8257) );
  NAND2_X1 U9470 ( .A1(n9554), .A2(n9555), .ZN(n9553) );
  NAND2_X1 U9471 ( .A1(n9705), .A2(n7490), .ZN(n7630) );
  NAND2_X1 U9472 ( .A1(n7630), .A2(n7631), .ZN(n9746) );
  NAND3_X1 U9473 ( .A1(n7637), .A2(n7636), .A3(n7557), .ZN(n7635) );
  NAND2_X1 U9474 ( .A1(n7643), .A2(n7641), .ZN(n12872) );
  NAND3_X1 U9475 ( .A1(n8127), .A2(n8125), .A3(n7646), .ZN(n11644) );
  NAND2_X1 U9476 ( .A1(n14271), .A2(n14272), .ZN(n7664) );
  NAND2_X1 U9477 ( .A1(n14256), .A2(n14255), .ZN(n7663) );
  NAND2_X1 U9478 ( .A1(n7667), .A2(n7547), .ZN(n12470) );
  XNOR2_X1 U9479 ( .A(n12045), .B(n14244), .ZN(n11572) );
  NAND2_X1 U9480 ( .A1(n9242), .A2(n7689), .ZN(n11210) );
  NAND2_X1 U9481 ( .A1(n9231), .A2(n9230), .ZN(n7689) );
  NAND3_X1 U9482 ( .A1(n7691), .A2(n7690), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7960) );
  NAND2_X1 U9483 ( .A1(n7704), .A2(n7705), .ZN(n15110) );
  NAND2_X1 U9484 ( .A1(n7704), .A2(n7702), .ZN(n7708) );
  NAND2_X1 U9485 ( .A1(n15074), .A2(n15073), .ZN(n10576) );
  NAND2_X1 U9486 ( .A1(n9420), .A2(n9418), .ZN(n7715) );
  OAI21_X1 U9487 ( .B1(n9420), .B2(n7719), .A(n7716), .ZN(n9445) );
  OAI21_X1 U9488 ( .B1(n9420), .B2(n9419), .A(n9418), .ZN(n9436) );
  NAND2_X1 U9489 ( .A1(n14836), .A2(n14837), .ZN(n13291) );
  NAND2_X1 U9490 ( .A1(n11591), .A2(n11593), .ZN(n11592) );
  NAND2_X1 U9491 ( .A1(n7723), .A2(n7725), .ZN(n11593) );
  OAI21_X1 U9492 ( .B1(n11059), .B2(n16310), .A(n10970), .ZN(n7726) );
  OAI21_X1 U9493 ( .B1(n11059), .B2(n11602), .A(n10965), .ZN(n7727) );
  NAND3_X1 U9494 ( .A1(n7732), .A2(n7729), .A3(n7728), .ZN(n13140) );
  OAI21_X1 U9495 ( .B1(n16550), .B2(n7751), .A(n7743), .ZN(n14908) );
  AOI21_X1 U9496 ( .B1(n16550), .B2(n7484), .A(n7750), .ZN(n7743) );
  NAND2_X1 U9497 ( .A1(n16550), .A2(n7745), .ZN(n7744) );
  INV_X1 U9498 ( .A(n7747), .ZN(n7746) );
  INV_X1 U9499 ( .A(n11060), .ZN(n7751) );
  NAND2_X1 U9500 ( .A1(n9900), .A2(n9895), .ZN(n9904) );
  NAND2_X1 U9501 ( .A1(n7758), .A2(n7757), .ZN(n9896) );
  NAND2_X1 U9502 ( .A1(n9900), .A2(n7759), .ZN(n7758) );
  NAND2_X1 U9503 ( .A1(n9900), .A2(n7489), .ZN(n9899) );
  NAND2_X1 U9504 ( .A1(n7512), .A2(n7766), .ZN(n9155) );
  INV_X1 U9505 ( .A(n9160), .ZN(n7767) );
  NAND3_X1 U9506 ( .A1(n7768), .A2(n9162), .A3(n9159), .ZN(n9166) );
  NAND2_X1 U9507 ( .A1(n7767), .A2(SI_2_), .ZN(n7768) );
  AND2_X1 U9508 ( .A1(n7768), .A2(n9159), .ZN(n9161) );
  INV_X1 U9509 ( .A(n9166), .ZN(n9163) );
  NAND2_X1 U9510 ( .A1(n7776), .A2(n9349), .ZN(n7775) );
  INV_X1 U9511 ( .A(n9351), .ZN(n7776) );
  NAND2_X1 U9512 ( .A1(n13090), .A2(n7453), .ZN(n7777) );
  NAND2_X1 U9513 ( .A1(n7777), .A2(n7778), .ZN(n14625) );
  XNOR2_X1 U9514 ( .A(n12421), .B(n14379), .ZN(n12205) );
  NAND2_X1 U9515 ( .A1(n14478), .A2(n7788), .ZN(n7784) );
  OAI21_X1 U9516 ( .B1(n14478), .B2(n14477), .A(n7790), .ZN(n14464) );
  NAND2_X1 U9517 ( .A1(n7795), .A2(n7794), .ZN(P3_U3296) );
  NAND2_X1 U9518 ( .A1(n7796), .A2(n11721), .ZN(n7795) );
  NAND3_X1 U9519 ( .A1(n7805), .A2(n7800), .A3(n7797), .ZN(n7796) );
  NAND2_X1 U9520 ( .A1(n7799), .A2(n7798), .ZN(n7797) );
  XNOR2_X1 U9521 ( .A(n13357), .B(n13799), .ZN(n7799) );
  NAND2_X1 U9522 ( .A1(n13540), .A2(n10425), .ZN(n7805) );
  OR2_X1 U9523 ( .A1(n8658), .A2(n7808), .ZN(n7807) );
  AOI22_X1 U9524 ( .A1(n8659), .A2(n7809), .B1(n11444), .B2(n7810), .ZN(n7806)
         );
  NAND2_X1 U9525 ( .A1(n8659), .A2(n11444), .ZN(n8661) );
  NOR2_X1 U9526 ( .A1(n7811), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U9527 ( .A1(n8066), .A2(n7817), .ZN(n7814) );
  NAND2_X1 U9528 ( .A1(n7814), .A2(n7815), .ZN(n8793) );
  NAND2_X1 U9529 ( .A1(n8880), .A2(n8879), .ZN(n8882) );
  NAND2_X1 U9530 ( .A1(n7519), .A2(n8918), .ZN(n13130) );
  OAI211_X1 U9531 ( .C1(n13486), .C2(n13485), .A(n13484), .B(n13492), .ZN(
        n13488) );
  NAND3_X1 U9532 ( .A1(n13359), .A2(n13360), .A3(n7538), .ZN(n13492) );
  NAND2_X1 U9533 ( .A1(n7828), .A2(n7826), .ZN(n16267) );
  NAND2_X1 U9534 ( .A1(n7544), .A2(n11698), .ZN(n7850) );
  NAND2_X1 U9535 ( .A1(n7852), .A2(n7468), .ZN(n14653) );
  NAND2_X1 U9536 ( .A1(n14651), .A2(n7854), .ZN(n7852) );
  NAND2_X1 U9537 ( .A1(n7853), .A2(n7467), .ZN(n14727) );
  NAND2_X1 U9538 ( .A1(n14651), .A2(n7855), .ZN(n7853) );
  NAND2_X1 U9539 ( .A1(n8294), .A2(n7539), .ZN(n10688) );
  INV_X1 U9540 ( .A(n7861), .ZN(n14479) );
  NAND3_X1 U9541 ( .A1(n10790), .A2(n10788), .A3(n10789), .ZN(n7862) );
  NAND2_X1 U9542 ( .A1(n7864), .A2(n10786), .ZN(n7863) );
  NAND2_X1 U9543 ( .A1(n7865), .A2(n10787), .ZN(n7864) );
  NAND2_X1 U9544 ( .A1(n10790), .A2(n10788), .ZN(n7865) );
  INV_X2 U9545 ( .A(n10873), .ZN(n10005) );
  NAND2_X1 U9546 ( .A1(n10810), .A2(n7868), .ZN(n7866) );
  NAND2_X1 U9547 ( .A1(n7866), .A2(n7867), .ZN(n10815) );
  NAND2_X1 U9548 ( .A1(n10819), .A2(n7882), .ZN(n7881) );
  NAND2_X1 U9549 ( .A1(n7888), .A2(n7891), .ZN(n10835) );
  NAND3_X1 U9550 ( .A1(n10830), .A2(n7889), .A3(n10831), .ZN(n7888) );
  OAI22_X1 U9551 ( .A1(n10747), .A2(n7896), .B1(n10748), .B2(n7895), .ZN(
        n10752) );
  NAND2_X1 U9552 ( .A1(n10752), .A2(n10753), .ZN(n10751) );
  NAND2_X1 U9553 ( .A1(n10774), .A2(n10775), .ZN(n10773) );
  NAND2_X1 U9554 ( .A1(n13367), .A2(n13366), .ZN(n12405) );
  OAI211_X1 U9555 ( .C1(n13367), .C2(n7901), .A(n7899), .B(n8449), .ZN(n12331)
         );
  NAND2_X1 U9556 ( .A1(n7900), .A2(n12393), .ZN(n7899) );
  INV_X1 U9557 ( .A(n13366), .ZN(n7900) );
  INV_X1 U9558 ( .A(n12393), .ZN(n7901) );
  NAND4_X1 U9559 ( .A1(n8090), .A2(n7904), .A3(n7903), .A4(n7902), .ZN(n8089)
         );
  NAND2_X1 U9560 ( .A1(n7905), .A2(n7466), .ZN(n13929) );
  NAND2_X1 U9561 ( .A1(n7908), .A2(n7545), .ZN(n8840) );
  NAND2_X1 U9562 ( .A1(n13836), .A2(n7537), .ZN(n7920) );
  NAND2_X1 U9563 ( .A1(n13836), .A2(n8896), .ZN(n7922) );
  AOI21_X1 U9564 ( .B1(n7927), .B2(n7925), .A(n7924), .ZN(n7923) );
  INV_X1 U9565 ( .A(n7927), .ZN(n7926) );
  INV_X1 U9566 ( .A(n13882), .ZN(n7934) );
  NOR2_X1 U9567 ( .A1(n13883), .A2(n8385), .ZN(n13869) );
  NOR2_X1 U9568 ( .A1(n8430), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n8426) );
  OR2_X2 U9569 ( .A1(n8430), .A2(n7939), .ZN(n8423) );
  NOR2_X1 U9570 ( .A1(n8430), .A2(n7940), .ZN(n8414) );
  NAND3_X1 U9571 ( .A1(n8411), .A2(n7942), .A3(n7941), .ZN(n7940) );
  NAND3_X1 U9572 ( .A1(n7945), .A2(n12360), .A3(n16494), .ZN(n12548) );
  NOR2_X2 U9573 ( .A1(n16621), .A2(n15762), .ZN(n7951) );
  NAND2_X1 U9574 ( .A1(n7957), .A2(n13596), .ZN(n7959) );
  NOR2_X2 U9575 ( .A1(n10496), .A2(n7954), .ZN(n13564) );
  NAND2_X1 U9576 ( .A1(n7957), .A2(n7568), .ZN(n7956) );
  INV_X1 U9577 ( .A(n7959), .ZN(n13667) );
  NAND2_X2 U9578 ( .A1(n8434), .A2(n8435), .ZN(n9141) );
  NAND2_X1 U9579 ( .A1(n13640), .A2(n7498), .ZN(n7964) );
  NAND2_X1 U9580 ( .A1(n7510), .A2(n13640), .ZN(n7970) );
  NAND2_X1 U9581 ( .A1(n9519), .A2(n7974), .ZN(n7971) );
  NAND2_X1 U9582 ( .A1(n7971), .A2(n7972), .ZN(n9544) );
  OAI21_X1 U9583 ( .B1(n9439), .B2(n7982), .A(n7980), .ZN(n9501) );
  NAND2_X1 U9584 ( .A1(n7979), .A2(n7977), .ZN(n9504) );
  NAND2_X1 U9585 ( .A1(n9439), .A2(n7980), .ZN(n7979) );
  NAND2_X1 U9586 ( .A1(n13679), .A2(n7986), .ZN(n7985) );
  NAND2_X1 U9587 ( .A1(n12320), .A2(n7991), .ZN(n12384) );
  NAND2_X1 U9588 ( .A1(n10440), .A2(n10439), .ZN(n12320) );
  NAND2_X1 U9589 ( .A1(n12384), .A2(n10446), .ZN(n12529) );
  NAND2_X1 U9590 ( .A1(n9587), .A2(n9586), .ZN(n8000) );
  NAND2_X1 U9591 ( .A1(n9587), .A2(n7994), .ZN(n7993) );
  OR2_X2 U9592 ( .A1(n13227), .A2(n13226), .ZN(n13225) );
  NAND3_X1 U9593 ( .A1(n8002), .A2(n8001), .A3(n7558), .ZN(n13227) );
  NAND2_X1 U9594 ( .A1(n8151), .A2(n8154), .ZN(n8001) );
  NAND2_X1 U9595 ( .A1(n8151), .A2(n10637), .ZN(n8002) );
  NAND2_X1 U9596 ( .A1(n12822), .A2(n8003), .ZN(n12897) );
  NAND2_X2 U9597 ( .A1(n8007), .A2(n9727), .ZN(n15696) );
  NOR2_X2 U9598 ( .A1(n13228), .A2(n13229), .ZN(n15694) );
  NOR2_X1 U9599 ( .A1(n8153), .A2(n8152), .ZN(n8151) );
  AND2_X4 U9600 ( .A1(n10428), .A2(n10427), .ZN(n10507) );
  XNOR2_X1 U9601 ( .A(n13718), .B(n13768), .ZN(n16125) );
  NAND2_X1 U9602 ( .A1(n8384), .A2(n11927), .ZN(n8021) );
  NOR2_X2 U9603 ( .A1(n15989), .A2(n15990), .ZN(n15998) );
  OR2_X1 U9604 ( .A1(n16020), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U9605 ( .A1(n16091), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8045) );
  OAI211_X1 U9606 ( .C1(n16091), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n8047), .B(
        n7462), .ZN(n8046) );
  AOI21_X1 U9607 ( .B1(n13356), .B2(n8051), .A(n13355), .ZN(n13357) );
  OAI21_X2 U9608 ( .B1(n8055), .B2(n8057), .A(n13390), .ZN(n12847) );
  NOR2_X2 U9609 ( .A1(n12480), .A2(n8058), .ZN(n8055) );
  NAND2_X1 U9610 ( .A1(n8056), .A2(n13381), .ZN(n12494) );
  NAND2_X1 U9611 ( .A1(n12480), .A2(n13518), .ZN(n8056) );
  OAI21_X1 U9612 ( .B1(n13518), .B2(n8058), .A(n13512), .ZN(n8057) );
  INV_X1 U9613 ( .A(n13381), .ZN(n8058) );
  NAND2_X1 U9614 ( .A1(n8698), .A2(n8697), .ZN(n8730) );
  OAI21_X1 U9615 ( .B1(n8698), .B2(n8069), .A(n8067), .ZN(n8751) );
  NAND2_X1 U9616 ( .A1(n8698), .A2(n8067), .ZN(n8066) );
  NAND2_X1 U9617 ( .A1(n8730), .A2(n8729), .ZN(n8749) );
  NAND2_X1 U9618 ( .A1(n8492), .A2(n8073), .ZN(n8070) );
  NAND2_X1 U9619 ( .A1(n8070), .A2(n8071), .ZN(n8525) );
  NAND2_X1 U9620 ( .A1(n12738), .A2(n8082), .ZN(n8078) );
  NAND2_X1 U9621 ( .A1(n8078), .A2(n8079), .ZN(n12972) );
  NAND2_X1 U9622 ( .A1(n8987), .A2(n8085), .ZN(n13927) );
  NAND2_X1 U9623 ( .A1(n8406), .A2(n8405), .ZN(n8700) );
  NAND2_X1 U9624 ( .A1(n8569), .A2(n7532), .ZN(n8584) );
  NAND2_X1 U9625 ( .A1(n8794), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8093) );
  NAND3_X1 U9626 ( .A1(n8094), .A2(n8092), .A3(n8093), .ZN(n8808) );
  NAND2_X1 U9627 ( .A1(n8094), .A2(n8093), .ZN(n8797) );
  NAND2_X1 U9628 ( .A1(n8808), .A2(n8093), .ZN(n8811) );
  INV_X1 U9629 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U9630 ( .A1(n8796), .A2(n8795), .ZN(n8094) );
  NAND3_X1 U9631 ( .A1(n8400), .A2(n8458), .A3(n8401), .ZN(n8566) );
  NAND2_X1 U9632 ( .A1(n8096), .A2(n8095), .ZN(n13830) );
  AOI21_X1 U9633 ( .B1(n8993), .B2(n13855), .A(n8098), .ZN(n8095) );
  NAND2_X1 U9634 ( .A1(n13874), .A2(n8097), .ZN(n8096) );
  NAND2_X1 U9635 ( .A1(n13874), .A2(n13485), .ZN(n13851) );
  NAND2_X1 U9636 ( .A1(n11963), .A2(n8102), .ZN(n8099) );
  NAND2_X1 U9637 ( .A1(n13058), .A2(n8109), .ZN(n8108) );
  OAI21_X1 U9638 ( .B1(n14350), .B2(n8123), .A(n8121), .ZN(n8124) );
  INV_X1 U9639 ( .A(n11577), .ZN(n8128) );
  INV_X1 U9640 ( .A(n11529), .ZN(n8129) );
  NAND3_X1 U9641 ( .A1(n8127), .A2(n8125), .A3(n11576), .ZN(n11585) );
  NAND3_X1 U9642 ( .A1(n8128), .A2(n11498), .A3(n8126), .ZN(n8125) );
  NAND3_X1 U9643 ( .A1(n8129), .A2(n8128), .A3(n11498), .ZN(n8127) );
  NAND3_X1 U9644 ( .A1(n10320), .A2(n8141), .A3(n8144), .ZN(n8140) );
  NAND3_X1 U9645 ( .A1(n10320), .A2(n8144), .A3(n8143), .ZN(n10213) );
  AND2_X2 U9646 ( .A1(n12609), .A2(n10622), .ZN(n12542) );
  NAND3_X1 U9647 ( .A1(n8435), .A2(n8434), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n8146) );
  NAND2_X1 U9648 ( .A1(n15181), .A2(n10633), .ZN(n8147) );
  NAND2_X1 U9649 ( .A1(n8147), .A2(n8148), .ZN(n10635) );
  INV_X1 U9650 ( .A(n15181), .ZN(n8150) );
  NAND2_X1 U9651 ( .A1(n13225), .A2(n8156), .ZN(n8155) );
  NAND2_X1 U9652 ( .A1(n13225), .A2(n8162), .ZN(n15092) );
  OAI211_X1 U9653 ( .C1(n13225), .C2(n8161), .A(n8157), .B(n8155), .ZN(n15675)
         );
  AND2_X1 U9654 ( .A1(n13225), .A2(n10639), .ZN(n15091) );
  NAND2_X1 U9655 ( .A1(n15150), .A2(n8165), .ZN(n8164) );
  OR2_X1 U9656 ( .A1(n11055), .A2(n14929), .ZN(n8177) );
  INV_X1 U9657 ( .A(n10966), .ZN(n8188) );
  OAI21_X1 U9658 ( .B1(n14895), .B2(n13301), .A(n8199), .ZN(n14795) );
  NAND2_X1 U9659 ( .A1(n8198), .A2(n8197), .ZN(n13320) );
  NAND2_X1 U9660 ( .A1(n14895), .A2(n8199), .ZN(n8198) );
  NAND2_X1 U9661 ( .A1(n13253), .A2(n7549), .ZN(n14826) );
  NAND2_X1 U9662 ( .A1(n13141), .A2(n8202), .ZN(n16547) );
  AOI21_X1 U9663 ( .B1(n11115), .B2(n8211), .A(n8207), .ZN(n8205) );
  NAND2_X1 U9664 ( .A1(n8207), .A2(n7491), .ZN(n8206) );
  AND2_X1 U9665 ( .A1(n10999), .A2(n11000), .ZN(n8212) );
  NAND2_X1 U9666 ( .A1(n9079), .A2(n9135), .ZN(n8216) );
  NAND2_X1 U9667 ( .A1(n8216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9214) );
  INV_X1 U9668 ( .A(n8219), .ZN(n10891) );
  NAND2_X1 U9669 ( .A1(n14365), .A2(n10702), .ZN(n8217) );
  NAND2_X1 U9670 ( .A1(n8219), .A2(n10714), .ZN(n8218) );
  AOI21_X1 U9671 ( .B1(n8219), .B2(n16418), .A(n10687), .ZN(n8295) );
  NOR2_X1 U9672 ( .A1(n10688), .A2(n8219), .ZN(n14443) );
  AOI21_X1 U9673 ( .B1(n10688), .B2(n8219), .A(n11533), .ZN(n8298) );
  AOI21_X1 U9674 ( .B1(n10544), .B2(n8220), .A(n8391), .ZN(n11993) );
  NAND2_X1 U9675 ( .A1(n15229), .A2(n7541), .ZN(n15210) );
  NAND2_X1 U9676 ( .A1(n15110), .A2(n15118), .ZN(n8241) );
  NAND2_X1 U9677 ( .A1(n8239), .A2(n10636), .ZN(n8237) );
  INV_X1 U9678 ( .A(n8239), .ZN(n8238) );
  NAND2_X1 U9679 ( .A1(n9668), .A2(n9667), .ZN(n8244) );
  NAND2_X1 U9680 ( .A1(n15177), .A2(n7543), .ZN(n15156) );
  NAND2_X1 U9681 ( .A1(n8247), .A2(n7531), .ZN(n12358) );
  NAND2_X1 U9682 ( .A1(n10551), .A2(n8245), .ZN(n8247) );
  NAND2_X1 U9683 ( .A1(n12177), .A2(n8248), .ZN(n12165) );
  NAND3_X1 U9684 ( .A1(n9387), .A2(n9386), .A3(n7553), .ZN(n8249) );
  NAND2_X1 U9685 ( .A1(n8249), .A2(n8250), .ZN(n9426) );
  INV_X1 U9686 ( .A(n9728), .ZN(n8252) );
  NAND3_X1 U9687 ( .A1(n9637), .A2(n8254), .A3(n8253), .ZN(n9646) );
  NAND3_X1 U9688 ( .A1(n9559), .A2(n9558), .A3(n7551), .ZN(n8253) );
  NOR2_X2 U9689 ( .A1(n9111), .A2(n8256), .ZN(n9095) );
  NAND2_X1 U9690 ( .A1(n8257), .A2(n8258), .ZN(n9312) );
  NAND2_X1 U9691 ( .A1(n8260), .A2(n8261), .ZN(n9529) );
  MUX2_X1 U9692 ( .A(n14942), .B(n16358), .S(n9260), .Z(n9197) );
  INV_X1 U9693 ( .A(n9117), .ZN(n9118) );
  XNOR2_X1 U9694 ( .A(n10679), .B(n10678), .ZN(n8271) );
  NAND3_X1 U9695 ( .A1(n14533), .A2(n7486), .A3(n8383), .ZN(n8273) );
  NAND2_X1 U9696 ( .A1(n12457), .A2(n8284), .ZN(n8283) );
  AOI21_X1 U9697 ( .B1(n8288), .B2(n12245), .A(n7502), .ZN(n8287) );
  NAND2_X1 U9698 ( .A1(n8292), .A2(n8291), .ZN(n13084) );
  NAND3_X1 U9699 ( .A1(n10320), .A2(n7413), .A3(n9921), .ZN(n8302) );
  OAI21_X1 U9700 ( .B1(n11610), .B2(n10851), .A(n8307), .ZN(n12251) );
  NAND3_X1 U9701 ( .A1(n8306), .A2(n8305), .A3(n12250), .ZN(n12253) );
  NAND2_X1 U9702 ( .A1(n8307), .A2(n11610), .ZN(n8306) );
  NAND3_X1 U9703 ( .A1(n8314), .A2(n8312), .A3(n8316), .ZN(n14659) );
  NAND3_X1 U9704 ( .A1(n8314), .A2(n8312), .A3(n7569), .ZN(n8317) );
  OR2_X1 U9705 ( .A1(n16595), .A2(n8321), .ZN(n8320) );
  NAND2_X1 U9706 ( .A1(n8326), .A2(n8325), .ZN(n12370) );
  NAND2_X1 U9707 ( .A1(n8331), .A2(n8333), .ZN(n8329) );
  INV_X1 U9708 ( .A(n8331), .ZN(n8334) );
  NAND2_X1 U9709 ( .A1(n10275), .A2(n10274), .ZN(n14506) );
  OR2_X1 U9710 ( .A1(n14676), .A2(n14492), .ZN(n8340) );
  NAND2_X1 U9711 ( .A1(n16572), .A2(n8347), .ZN(n8346) );
  NAND2_X1 U9712 ( .A1(n8352), .A2(n10734), .ZN(n8351) );
  NAND2_X1 U9713 ( .A1(n10732), .A2(n10731), .ZN(n8352) );
  NAND3_X1 U9714 ( .A1(n10732), .A2(n10731), .A3(n10735), .ZN(n10739) );
  NAND2_X1 U9715 ( .A1(n10762), .A2(n10763), .ZN(n10761) );
  NAND2_X1 U9716 ( .A1(n10823), .A2(n8358), .ZN(n8357) );
  NAND2_X1 U9717 ( .A1(n8357), .A2(n8355), .ZN(n10827) );
  AND2_X1 U9718 ( .A1(n8356), .A2(n10828), .ZN(n8355) );
  NAND2_X1 U9719 ( .A1(n10800), .A2(n8363), .ZN(n8362) );
  NAND2_X1 U9720 ( .A1(n8362), .A2(n8360), .ZN(n10804) );
  AND2_X1 U9721 ( .A1(n10805), .A2(n8361), .ZN(n8360) );
  NAND2_X1 U9722 ( .A1(n10835), .A2(n8368), .ZN(n8365) );
  OAI21_X1 U9723 ( .B1(n10835), .B2(n8369), .A(n8368), .ZN(n10840) );
  NAND2_X1 U9724 ( .A1(n8365), .A2(n8366), .ZN(n10839) );
  NAND2_X1 U9725 ( .A1(n10742), .A2(n7552), .ZN(n8370) );
  NAND2_X1 U9726 ( .A1(n8375), .A2(n8374), .ZN(n8373) );
  NOR2_X1 U9727 ( .A1(n10384), .A2(n9939), .ZN(n10323) );
  NAND2_X1 U9728 ( .A1(n8377), .A2(n8379), .ZN(n10727) );
  NAND3_X1 U9729 ( .A1(n10722), .A2(n10721), .A3(n8378), .ZN(n8377) );
  OR2_X1 U9730 ( .A1(n10873), .A2(n8454), .ZN(n9975) );
  NAND2_X1 U9731 ( .A1(n10696), .A2(n10329), .ZN(n11852) );
  INV_X1 U9732 ( .A(n10696), .ZN(n13114) );
  NAND2_X1 U9733 ( .A1(n13114), .A2(n10329), .ZN(n10946) );
  NAND2_X1 U9734 ( .A1(n11780), .A2(n11781), .ZN(n11797) );
  AOI21_X1 U9735 ( .B1(n15675), .B2(n16394), .A(n10662), .ZN(n10663) );
  NAND2_X1 U9736 ( .A1(n8527), .A2(n8526), .ZN(n8543) );
  AND2_X1 U9737 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  OAI21_X1 U9738 ( .B1(n14302), .B2(n14303), .A(n14249), .ZN(n14252) );
  INV_X1 U9739 ( .A(n7414), .ZN(n13542) );
  XNOR2_X1 U9740 ( .A(n13327), .B(n8994), .ZN(n13813) );
  OR2_X1 U9741 ( .A1(n10650), .A2(n9824), .ZN(n16640) );
  NAND2_X1 U9742 ( .A1(n9155), .A2(n9157), .ZN(n9144) );
  OR2_X1 U9743 ( .A1(n8863), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U9744 ( .A1(n8430), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8431) );
  INV_X1 U9745 ( .A(n13328), .ZN(n8962) );
  OAI211_X1 U9746 ( .C1(n9141), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n9140), .B(
        SI_0_), .ZN(n9142) );
  NAND2_X1 U9747 ( .A1(n9141), .A2(n9948), .ZN(n9140) );
  NAND2_X1 U9748 ( .A1(n10607), .A2(n10606), .ZN(n12037) );
  NAND2_X1 U9749 ( .A1(n14546), .A2(n10263), .ZN(n14523) );
  AOI211_X1 U9750 ( .C1(n16358), .C2(n16346), .A(n16345), .B(n16566), .ZN(
        n16359) );
  NAND2_X1 U9751 ( .A1(n9196), .A2(n16358), .ZN(n10541) );
  NAND2_X1 U9752 ( .A1(n12358), .A2(n10552), .ZN(n10554) );
  NAND2_X1 U9753 ( .A1(n9174), .A2(n9173), .ZN(n16358) );
  NAND2_X1 U9754 ( .A1(n9118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U9755 ( .A1(n10325), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U9756 ( .A1(n10322), .A2(n10321), .ZN(n10325) );
  NAND2_X2 U9757 ( .A1(n15201), .A2(n15200), .ZN(n15741) );
  INV_X1 U9758 ( .A(n10708), .ZN(n10711) );
  AND2_X1 U9759 ( .A1(n9522), .A2(n7471), .ZN(n9900) );
  OAI222_X1 U9760 ( .A1(n14792), .A2(n13039), .B1(P2_U3088), .B2(n10695), .C1(
        n14775), .C2(n13038), .ZN(P2_U3305) );
  NAND2_X1 U9761 ( .A1(n10695), .A2(n10331), .ZN(n11491) );
  NAND2_X4 U9762 ( .A1(n9941), .A2(n9963), .ZN(n9999) );
  XNOR2_X1 U9763 ( .A(n11015), .B(n11012), .ZN(n12883) );
  OR2_X1 U9764 ( .A1(n13656), .A2(n14077), .ZN(n8381) );
  INV_X1 U9765 ( .A(n13245), .ZN(n13823) );
  AND2_X2 U9766 ( .A1(n9040), .A2(n11722), .ZN(n16618) );
  OR2_X1 U9767 ( .A1(n16615), .A2(n9057), .ZN(n8382) );
  INV_X2 U9768 ( .A(n16340), .ZN(n14100) );
  AND3_X2 U9769 ( .A1(n12402), .A2(n9055), .A3(n9054), .ZN(n16615) );
  INV_X1 U9770 ( .A(n16615), .ZN(n9060) );
  INV_X1 U9771 ( .A(n14149), .ZN(n9056) );
  AND2_X2 U9772 ( .A1(n10954), .A2(n11146), .ZN(P1_U4016) );
  AND2_X1 U9773 ( .A1(n11797), .A2(n11796), .ZN(n8384) );
  AND2_X1 U9774 ( .A1(n11501), .A2(n10374), .ZN(n14578) );
  AND2_X1 U9775 ( .A1(n13563), .A2(n13871), .ZN(n8385) );
  INV_X1 U9776 ( .A(n9999), .ZN(n10375) );
  OR2_X1 U9777 ( .A1(n10479), .A2(n14028), .ZN(n8386) );
  AND2_X1 U9778 ( .A1(n10476), .A2(n14039), .ZN(n8387) );
  INV_X1 U9779 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9137) );
  INV_X1 U9780 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8402) );
  AND2_X1 U9781 ( .A1(n10317), .A2(n10316), .ZN(n10920) );
  INV_X1 U9782 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9207) );
  INV_X1 U9783 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15950) );
  INV_X1 U9784 ( .A(n13873), .ZN(n8991) );
  INV_X1 U9785 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8411) );
  INV_X4 U9786 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U9787 ( .A(n10858), .ZN(n12705) );
  AND2_X1 U9788 ( .A1(n13686), .A2(n13857), .ZN(n8389) );
  OR3_X1 U9789 ( .A1(n15218), .A2(n15060), .A3(n15059), .ZN(n8390) );
  AND2_X1 U9790 ( .A1(n9860), .A2(n14940), .ZN(n8391) );
  OR2_X1 U9791 ( .A1(n9860), .A2(n14940), .ZN(n8392) );
  NOR2_X1 U9792 ( .A1(n10945), .A2(n10944), .ZN(n8393) );
  XNOR2_X1 U9793 ( .A(n9819), .B(n9818), .ZN(n10872) );
  OR2_X1 U9794 ( .A1(n14659), .A2(n14648), .ZN(n8394) );
  AND2_X1 U9795 ( .A1(n15681), .A2(n15680), .ZN(n8395) );
  NAND2_X2 U9796 ( .A1(n10673), .A2(n14640), .ZN(n14610) );
  NAND2_X2 U9797 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11302), .ZN(n14385) );
  AND2_X1 U9798 ( .A1(n9193), .A2(n9192), .ZN(n8396) );
  OR2_X1 U9799 ( .A1(n12158), .A2(n11420), .ZN(n16633) );
  AND2_X2 U9800 ( .A1(n10655), .A2(n16653), .ZN(n16398) );
  NAND2_X1 U9801 ( .A1(n7435), .A2(n10714), .ZN(n10704) );
  NAND2_X1 U9802 ( .A1(n10704), .A2(n10703), .ZN(n10709) );
  INV_X1 U9803 ( .A(n10709), .ZN(n10710) );
  INV_X1 U9804 ( .A(n10718), .ZN(n10719) );
  MUX2_X1 U9805 ( .A(n14924), .B(n15718), .S(n7415), .Z(n9664) );
  MUX2_X1 U9806 ( .A(n14922), .B(n15696), .S(n7415), .Z(n9728) );
  NOR2_X1 U9807 ( .A1(n13491), .A2(n13466), .ZN(n13493) );
  INV_X1 U9808 ( .A(n12163), .ZN(n10547) );
  INV_X1 U9809 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8408) );
  INV_X1 U9810 ( .A(n13512), .ZN(n8515) );
  INV_X1 U9811 ( .A(n10901), .ZN(n11485) );
  INV_X1 U9812 ( .A(n10984), .ZN(n10985) );
  OR4_X1 U9813 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U9814 ( .A1(n13245), .A2(n13829), .ZN(n8933) );
  INV_X1 U9815 ( .A(n13001), .ZN(n10942) );
  INV_X1 U9816 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10202) );
  NAND2_X1 U9817 ( .A1(n10368), .A2(n14368), .ZN(n10369) );
  NOR2_X1 U9818 ( .A1(n10266), .A2(n14273), .ZN(n9935) );
  AND2_X1 U9819 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n9933) );
  INV_X1 U9820 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10069) );
  AND2_X1 U9821 ( .A1(n11015), .A2(n11014), .ZN(n11016) );
  NAND2_X1 U9822 ( .A1(n11008), .A2(n11009), .ZN(n11010) );
  OR2_X1 U9823 ( .A1(n11036), .A2(n11035), .ZN(n11037) );
  NAND2_X1 U9824 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  AND2_X1 U9825 ( .A1(n9591), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9647) );
  AND2_X1 U9826 ( .A1(n9600), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9591) );
  INV_X1 U9827 ( .A(n15159), .ZN(n10570) );
  INV_X1 U9828 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9560) );
  INV_X1 U9829 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n15449) );
  INV_X1 U9830 ( .A(n12616), .ZN(n10621) );
  AND4_X1 U9831 ( .A1(n9091), .A2(n9090), .A3(n15449), .A4(n8215), .ZN(n9092)
         );
  INV_X1 U9832 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n15651) );
  INV_X1 U9833 ( .A(n8755), .ZN(n8741) );
  OR2_X1 U9834 ( .A1(n10474), .A2(n13655), .ZN(n10475) );
  OR2_X1 U9835 ( .A1(n8889), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8906) );
  INV_X1 U9836 ( .A(n13729), .ZN(n13730) );
  INV_X1 U9837 ( .A(n13360), .ZN(n8914) );
  INV_X1 U9838 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15532) );
  INV_X1 U9839 ( .A(n8423), .ZN(n8425) );
  INV_X1 U9840 ( .A(n8605), .ZN(n8602) );
  NAND2_X1 U9841 ( .A1(n10943), .A2(n10942), .ZN(n10944) );
  OR2_X1 U9842 ( .A1(n10289), .A2(n14354), .ZN(n10310) );
  OR2_X1 U9843 ( .A1(n10203), .A2(n10202), .ZN(n10220) );
  OR2_X1 U9844 ( .A1(n12727), .A2(n12726), .ZN(n15870) );
  AND2_X1 U9845 ( .A1(n14498), .A2(n14368), .ZN(n10286) );
  INV_X1 U9846 ( .A(n10331), .ZN(n10902) );
  OR2_X1 U9847 ( .A1(n10070), .A2(n10069), .ZN(n10085) );
  AND2_X1 U9848 ( .A1(n15823), .A2(n10671), .ZN(n11499) );
  INV_X1 U9849 ( .A(n10867), .ZN(n10678) );
  INV_X2 U9850 ( .A(n10845), .ZN(n10871) );
  NAND2_X1 U9851 ( .A1(n10384), .A2(n10385), .ZN(n10397) );
  INV_X1 U9852 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U9853 ( .A1(n9708), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9750) );
  AND2_X1 U9854 ( .A1(n9647), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9669) );
  INV_X1 U9855 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9495) );
  INV_X1 U9856 ( .A(n15163), .ZN(n15185) );
  OAI21_X1 U9857 ( .B1(n10602), .B2(n10539), .A(n10538), .ZN(n16350) );
  INV_X1 U9858 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15512) );
  OR2_X1 U9859 ( .A1(n8845), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U9860 ( .A1(n10486), .A2(n13915), .ZN(n10487) );
  NAND2_X1 U9861 ( .A1(n10530), .A2(n10517), .ZN(n13671) );
  INV_X1 U9862 ( .A(n12101), .ZN(n12111) );
  INV_X1 U9863 ( .A(n12681), .ZN(n12688) );
  INV_X1 U9864 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15335) );
  INV_X1 U9865 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15562) );
  AND2_X1 U9866 ( .A1(n11732), .A2(n11730), .ZN(n11742) );
  NAND2_X1 U9867 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  OR2_X1 U9868 ( .A1(n8834), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8845) );
  OR2_X1 U9869 ( .A1(n13351), .A2(n12193), .ZN(n8799) );
  INV_X1 U9870 ( .A(n13704), .ZN(n13965) );
  NOR2_X1 U9871 ( .A1(n16609), .A2(n12397), .ZN(n10514) );
  INV_X1 U9872 ( .A(n14209), .ZN(n12399) );
  OR2_X1 U9873 ( .A1(n13351), .A2(n12608), .ZN(n8843) );
  INV_X1 U9874 ( .A(n13625), .ZN(n14039) );
  AND2_X1 U9875 ( .A1(n13426), .A2(n13423), .ZN(n14068) );
  AND2_X1 U9876 ( .A1(n12192), .A2(n13736), .ZN(n16333) );
  INV_X1 U9877 ( .A(n12482), .ZN(n13518) );
  NAND2_X1 U9878 ( .A1(n9000), .A2(n12413), .ZN(n16609) );
  NAND2_X1 U9879 ( .A1(n10517), .A2(n13466), .ZN(n14089) );
  INV_X1 U9880 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9035) );
  AND2_X1 U9881 ( .A1(n8841), .A2(n8826), .ZN(n8827) );
  AND2_X1 U9882 ( .A1(n8772), .A2(n8733), .ZN(n8734) );
  OR2_X1 U9883 ( .A1(n8715), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U9884 ( .A1(n8456), .A2(n8455), .ZN(n8469) );
  INV_X1 U9885 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n12876) );
  INV_X1 U9886 ( .A(n14333), .ZN(n14281) );
  OR2_X1 U9887 ( .A1(n15822), .A2(n11500), .ZN(n11506) );
  OR2_X1 U9888 ( .A1(n14451), .A2(n9999), .ZN(n10317) );
  NOR3_X1 U9889 ( .A1(n14788), .A2(n13204), .A3(n14790), .ZN(n10953) );
  INV_X1 U9890 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15867) );
  XNOR2_X1 U9891 ( .A(n14480), .B(n14493), .ZN(n14477) );
  AND2_X1 U9892 ( .A1(n10948), .A2(n10902), .ZN(n11501) );
  INV_X1 U9893 ( .A(n14578), .ZN(n14602) );
  OR2_X1 U9894 ( .A1(n16598), .A2(n11505), .ZN(n14621) );
  INV_X1 U9895 ( .A(n16584), .ZN(n14510) );
  OR2_X1 U9896 ( .A1(n10137), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n10157) );
  INV_X1 U9897 ( .A(n14931), .ZN(n16544) );
  AND2_X1 U9898 ( .A1(n13292), .A2(n13290), .ZN(n14838) );
  OR2_X1 U9899 ( .A1(n15167), .A2(n9689), .ZN(n9599) );
  INV_X1 U9900 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15992) );
  INV_X1 U9901 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n16017) );
  INV_X1 U9902 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n16032) );
  INV_X1 U9903 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U9904 ( .A1(n14922), .A2(n15233), .ZN(n13217) );
  INV_X1 U9905 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14911) );
  INV_X1 U9906 ( .A(n12360), .ZN(n12613) );
  INV_X1 U9907 ( .A(n16377), .ZN(n16381) );
  NAND2_X1 U9908 ( .A1(n9168), .A2(n9820), .ZN(n9174) );
  INV_X1 U9909 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n15663) );
  NAND2_X1 U9910 ( .A1(n9889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9891) );
  INV_X1 U9911 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9109) );
  INV_X1 U9912 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9895) );
  INV_X1 U9913 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15973) );
  OR2_X1 U9914 ( .A1(n11722), .A2(n11721), .ZN(n11732) );
  OAI21_X1 U9915 ( .B1(n13833), .B2(n13700), .A(n10534), .ZN(n10535) );
  AND3_X1 U9916 ( .A1(n8611), .A2(n8610), .A3(n8609), .ZN(n12901) );
  AND3_X1 U9917 ( .A1(n8592), .A2(n8591), .A3(n8590), .ZN(n12828) );
  INV_X1 U9918 ( .A(n13694), .ZN(n13683) );
  NAND2_X1 U9919 ( .A1(n10515), .A2(n14073), .ZN(n13673) );
  AND2_X1 U9920 ( .A1(n8913), .A2(n8912), .ZN(n13839) );
  AND4_X1 U9921 ( .A1(n8761), .A2(n8760), .A3(n8759), .A4(n8758), .ZN(n14012)
         );
  INV_X1 U9922 ( .A(n16244), .ZN(n16254) );
  INV_X1 U9923 ( .A(n14089), .ZN(n13986) );
  INV_X1 U9924 ( .A(n14073), .ZN(n16337) );
  AND3_X1 U9925 ( .A1(n11722), .A2(n9047), .A3(n9046), .ZN(n12402) );
  NOR2_X1 U9926 ( .A1(n16618), .A2(n9041), .ZN(n9042) );
  INV_X1 U9927 ( .A(n16609), .ZN(n14105) );
  AND2_X1 U9928 ( .A1(n9000), .A2(n16333), .ZN(n16521) );
  OR2_X1 U9929 ( .A1(n16428), .A2(n16521), .ZN(n16614) );
  NOR2_X1 U9930 ( .A1(n11377), .A2(n11376), .ZN(n11382) );
  XNOR2_X1 U9931 ( .A(n8947), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13544) );
  AND2_X1 U9932 ( .A1(n8694), .A2(n8664), .ZN(n8665) );
  NOR2_X1 U9933 ( .A1(n8651), .A2(n8650), .ZN(n13741) );
  INV_X1 U9934 ( .A(n14320), .ZN(n14331) );
  INV_X1 U9935 ( .A(n11506), .ZN(n11504) );
  INV_X1 U9936 ( .A(n10695), .ZN(n10948) );
  OR2_X1 U9937 ( .A1(n14517), .A2(n9999), .ZN(n9947) );
  AND4_X1 U9938 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n12634) );
  INV_X1 U9939 ( .A(n15922), .ZN(n14418) );
  AND2_X1 U9940 ( .A1(n11310), .A2(n11309), .ZN(n15922) );
  INV_X1 U9941 ( .A(n14648), .ZN(n16604) );
  INV_X1 U9942 ( .A(n16601), .ZN(n14645) );
  INV_X1 U9943 ( .A(n12148), .ZN(n16514) );
  NOR2_X1 U9944 ( .A1(n15815), .A2(n10411), .ZN(n11690) );
  OR2_X1 U9945 ( .A1(n10670), .A2(n15820), .ZN(n15815) );
  NAND2_X1 U9946 ( .A1(n10392), .A2(n10391), .ZN(n10390) );
  AND2_X1 U9947 ( .A1(n10138), .A2(n10157), .ZN(n12583) );
  INV_X1 U9948 ( .A(n14775), .ZN(n14779) );
  INV_X1 U9949 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n11105) );
  INV_X1 U9950 ( .A(n16549), .ZN(n14905) );
  OR2_X1 U9951 ( .A1(n15134), .A2(n9689), .ZN(n9676) );
  AND4_X2 U9952 ( .A1(n9219), .A2(n9218), .A3(n9217), .A4(n9216), .ZN(n11996)
         );
  INV_X1 U9953 ( .A(n13028), .ZN(n16277) );
  INV_X1 U9954 ( .A(n13026), .ZN(n16285) );
  INV_X1 U9955 ( .A(n16566), .ZN(n16622) );
  NAND2_X1 U9956 ( .A1(n15079), .A2(n15078), .ZN(n15080) );
  INV_X1 U9957 ( .A(n15216), .ZN(n15233) );
  INV_X1 U9958 ( .A(n16646), .ZN(n16394) );
  AND2_X1 U9959 ( .A1(n7416), .A2(n13032), .ZN(n16498) );
  INV_X1 U9960 ( .A(n15218), .ZN(n15234) );
  NAND2_X1 U9961 ( .A1(n15263), .A2(n8390), .ZN(n15264) );
  INV_X1 U9962 ( .A(n16568), .ZN(n16628) );
  OR2_X1 U9963 ( .A1(n10582), .A2(n10581), .ZN(n16631) );
  AND2_X1 U9964 ( .A1(n9825), .A2(n16295), .ZN(n16452) );
  AND3_X2 U9965 ( .A1(n9124), .A2(n9123), .A3(n9122), .ZN(n9824) );
  AND2_X1 U9966 ( .A1(n11732), .A2(n11731), .ZN(n16252) );
  INV_X1 U9967 ( .A(n10535), .ZN(n10536) );
  AND2_X1 U9968 ( .A1(n10528), .A2(n10527), .ZN(n13694) );
  INV_X1 U9969 ( .A(n13839), .ZN(n13702) );
  NAND2_X1 U9970 ( .A1(n14210), .A2(n10956), .ZN(n13711) );
  INV_X1 U9971 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n16123) );
  INV_X1 U9972 ( .A(n16265), .ZN(n16250) );
  INV_X1 U9973 ( .A(n13928), .ZN(n14189) );
  NAND2_X1 U9974 ( .A1(n16340), .A2(n16335), .ZN(n14080) );
  AND2_X1 U9975 ( .A1(n9058), .A2(n8382), .ZN(n9059) );
  NAND2_X1 U9976 ( .A1(n16615), .A2(n14105), .ZN(n14149) );
  INV_X1 U9977 ( .A(n13637), .ZN(n14171) );
  NAND2_X1 U9978 ( .A1(n16618), .A2(n14105), .ZN(n14207) );
  INV_X1 U9979 ( .A(SI_26_), .ZN(n13069) );
  INV_X1 U9980 ( .A(SI_17_), .ZN(n15480) );
  INV_X1 U9981 ( .A(SI_11_), .ZN(n15493) );
  INV_X1 U9982 ( .A(n12644), .ZN(n12646) );
  NAND2_X1 U9983 ( .A1(n11504), .A2(n11502), .ZN(n14326) );
  INV_X1 U9984 ( .A(n10920), .ZN(n14366) );
  INV_X1 U9985 ( .A(n14512), .ZN(n14369) );
  INV_X1 U9986 ( .A(n10357), .ZN(n14375) );
  OR2_X1 U9987 ( .A1(n11310), .A2(P2_U3088), .ZN(n15928) );
  OR2_X1 U9988 ( .A1(n16598), .A2(n10696), .ZN(n16601) );
  AND2_X1 U9989 ( .A1(n12256), .A2(n12255), .ZN(n16425) );
  NAND2_X1 U9990 ( .A1(n16591), .A2(n16418), .ZN(n14708) );
  INV_X1 U9991 ( .A(n16591), .ZN(n16589) );
  AND2_X2 U9992 ( .A1(n11690), .A2(n10414), .ZN(n16591) );
  NAND2_X1 U9993 ( .A1(n11690), .A2(n15822), .ZN(n16592) );
  OR2_X1 U9994 ( .A1(n15820), .A2(n15818), .ZN(n15819) );
  AND2_X1 U9995 ( .A1(n11511), .A2(n10400), .ZN(n15823) );
  XNOR2_X1 U9996 ( .A(n10394), .B(n10393), .ZN(n13204) );
  INV_X1 U9997 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U9998 ( .A1(n11464), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16558) );
  INV_X1 U9999 ( .A(n11055), .ZN(n16641) );
  NAND2_X1 U10000 ( .A1(n9676), .A2(n9675), .ZN(n15114) );
  OR2_X1 U10001 ( .A1(n9434), .A2(n9433), .ZN(n14931) );
  INV_X1 U10002 ( .A(n11996), .ZN(n14940) );
  NAND2_X1 U10003 ( .A1(n11177), .A2(n11176), .ZN(n15046) );
  INV_X1 U10004 ( .A(n10601), .ZN(n10664) );
  AND2_X1 U10005 ( .A1(n15251), .A2(n15250), .ZN(n15759) );
  NAND2_X1 U10006 ( .A1(n11100), .A2(n11237), .ZN(n16653) );
  NAND2_X1 U10007 ( .A1(n7416), .A2(n11412), .ZN(n16646) );
  INV_X2 U10008 ( .A(n16633), .ZN(n16635) );
  AND2_X1 U10009 ( .A1(n10600), .A2(n11146), .ZN(n11237) );
  INV_X1 U10010 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15798) );
  INV_X1 U10011 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n12064) );
  INV_X1 U10012 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n11438) );
  INV_X2 U10013 ( .A(n13711), .ZN(P3_U3897) );
  NAND2_X1 U10014 ( .A1(n9076), .A2(n9075), .ZN(P3_U3487) );
  INV_X1 U10015 ( .A(n10424), .ZN(P3_U3455) );
  INV_X1 U10016 ( .A(n14385), .ZN(P2_U3947) );
  NAND2_X1 U10017 ( .A1(n8394), .A2(n10694), .ZN(P2_U3236) );
  NAND2_X1 U10018 ( .A1(n10664), .A2(n10663), .ZN(P1_U3356) );
  NOR2_X1 U10019 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n8404) );
  NOR2_X2 U10020 ( .A1(n9005), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n9008) );
  INV_X1 U10021 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10022 ( .A1(n9008), .A2(n8410), .ZN(n8430) );
  XNOR2_X2 U10023 ( .A(n8412), .B(n14215), .ZN(n8418) );
  INV_X1 U10024 ( .A(n8418), .ZN(n8416) );
  NAND2_X1 U10025 ( .A1(n8423), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8413) );
  MUX2_X1 U10026 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8413), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8415) );
  INV_X1 U10027 ( .A(n8414), .ZN(n14214) );
  AND2_X2 U10028 ( .A1(n8415), .A2(n14214), .ZN(n8417) );
  AND2_X2 U10029 ( .A1(n8416), .A2(n14222), .ZN(n8498) );
  NAND2_X1 U10030 ( .A1(n8498), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8422) );
  AND2_X2 U10031 ( .A1(n8416), .A2(n8417), .ZN(n8631) );
  NAND2_X1 U10032 ( .A1(n8631), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8421) );
  AND2_X2 U10033 ( .A1(n8418), .A2(n14222), .ZN(n8481) );
  NAND2_X1 U10034 ( .A1(n7437), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8420) );
  AND2_X4 U10035 ( .A1(n8418), .A2(n8417), .ZN(n13328) );
  NAND2_X1 U10036 ( .A1(n13328), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8419) );
  AND4_X4 U10037 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n12330)
         );
  INV_X1 U10038 ( .A(n12330), .ZN(n13715) );
  OR2_X1 U10039 ( .A1(n8426), .A2(n8626), .ZN(n8427) );
  NAND2_X2 U10040 ( .A1(n8429), .A2(n8428), .ZN(n8956) );
  NAND2_X4 U10041 ( .A1(n8956), .A2(n7414), .ZN(n11724) );
  INV_X1 U10042 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11735) );
  INV_X1 U10043 ( .A(n11736), .ZN(n8432) );
  INV_X2 U10044 ( .A(n9141), .ZN(n11208) );
  INV_X8 U10045 ( .A(n11208), .ZN(n11209) );
  NAND2_X1 U10046 ( .A1(n9948), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10047 ( .A1(n8436), .A2(n8437), .ZN(n8440) );
  INV_X1 U10048 ( .A(n8437), .ZN(n8438) );
  NAND2_X1 U10049 ( .A1(n8439), .A2(n8438), .ZN(n8456) );
  AND2_X1 U10050 ( .A1(n8440), .A2(n8456), .ZN(n11195) );
  OR2_X1 U10051 ( .A1(n8467), .A2(n11195), .ZN(n8442) );
  OR2_X1 U10052 ( .A1(n8494), .A2(n15502), .ZN(n8441) );
  OAI211_X1 U10053 ( .C1(n11724), .C2(n11738), .A(n8442), .B(n8441), .ZN(
        n10429) );
  INV_X1 U10054 ( .A(n10429), .ZN(n8448) );
  NAND2_X1 U10055 ( .A1(n13328), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10056 ( .A1(n8481), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10057 ( .A1(n8631), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10058 ( .A1(n8498), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8443) );
  XNOR2_X1 U10059 ( .A(n9948), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n8447) );
  MUX2_X1 U10060 ( .A(n8447), .B(SI_0_), .S(n11209), .Z(n14224) );
  MUX2_X1 U10061 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14224), .S(n11724), .Z(n12443) );
  NAND2_X1 U10062 ( .A1(n13585), .A2(n12443), .ZN(n12393) );
  NAND2_X1 U10063 ( .A1(n12330), .A2(n8448), .ZN(n8449) );
  NAND2_X1 U10064 ( .A1(n7437), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10065 ( .A1(n8498), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10066 ( .A1(n13328), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8450) );
  OR2_X1 U10067 ( .A1(n8494), .A2(SI_2_), .ZN(n8460) );
  NAND2_X1 U10068 ( .A1(n8454), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8455) );
  XNOR2_X1 U10069 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8468) );
  XNOR2_X1 U10070 ( .A(n8469), .B(n8468), .ZN(n11224) );
  OR2_X1 U10071 ( .A1(n8467), .A2(n11224), .ZN(n8459) );
  NOR2_X1 U10072 ( .A1(n11736), .A2(n8626), .ZN(n8457) );
  NAND2_X1 U10073 ( .A1(n13582), .A2(n11919), .ZN(n13374) );
  INV_X1 U10074 ( .A(n13582), .ZN(n13714) );
  INV_X1 U10075 ( .A(n11919), .ZN(n12335) );
  NAND2_X1 U10076 ( .A1(n13714), .A2(n12335), .ZN(n13370) );
  NAND2_X1 U10077 ( .A1(n13374), .A2(n13370), .ZN(n12328) );
  NAND2_X1 U10078 ( .A1(n12331), .A2(n12328), .ZN(n8462) );
  NAND2_X1 U10079 ( .A1(n13582), .A2(n12335), .ZN(n8461) );
  NAND2_X1 U10080 ( .A1(n8462), .A2(n8461), .ZN(n12428) );
  INV_X1 U10081 ( .A(n12428), .ZN(n8479) );
  NAND2_X1 U10082 ( .A1(n7437), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10083 ( .A1(n8498), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U10084 ( .A1(n8631), .A2(n12559), .ZN(n8464) );
  NAND2_X1 U10085 ( .A1(n13328), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8463) );
  OR2_X1 U10086 ( .A1(n13351), .A2(SI_3_), .ZN(n8478) );
  NAND2_X1 U10087 ( .A1(n8469), .A2(n8468), .ZN(n8471) );
  INV_X1 U10088 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U10089 ( .A1(n11217), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10090 ( .A1(n8471), .A2(n8470), .ZN(n8492) );
  XNOR2_X1 U10091 ( .A(n8492), .B(n8491), .ZN(n11226) );
  OR2_X1 U10092 ( .A1(n8923), .A2(n11226), .ZN(n8477) );
  MUX2_X1 U10093 ( .A(n8626), .B(n8472), .S(P3_IR_REG_3__SCAN_IN), .Z(n8475)
         );
  INV_X1 U10094 ( .A(n8487), .ZN(n8474) );
  OR2_X1 U10095 ( .A1(n11724), .A2(n11838), .ZN(n8476) );
  AND3_X2 U10096 ( .A1(n8478), .A2(n8477), .A3(n8476), .ZN(n12560) );
  INV_X1 U10097 ( .A(n12560), .ZN(n12436) );
  NAND2_X1 U10098 ( .A1(n13713), .A2(n12436), .ZN(n13378) );
  NAND2_X1 U10099 ( .A1(n10438), .A2(n12560), .ZN(n13376) );
  NAND2_X1 U10100 ( .A1(n8479), .A2(n13515), .ZN(n12426) );
  NAND2_X1 U10101 ( .A1(n13713), .A2(n12560), .ZN(n8480) );
  NAND2_X1 U10102 ( .A1(n12426), .A2(n8480), .ZN(n12483) );
  NAND2_X1 U10103 ( .A1(n7437), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10104 ( .A1(n13328), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10105 ( .A1(n12559), .A2(n15542), .ZN(n8500) );
  NAND2_X1 U10106 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8482) );
  NAND2_X1 U10107 ( .A1(n8500), .A2(n8482), .ZN(n12653) );
  NAND2_X1 U10108 ( .A1(n8631), .A2(n12653), .ZN(n8484) );
  NAND2_X1 U10109 ( .A1(n8498), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8483) );
  NAND4_X1 U10110 ( .A1(n8486), .A2(n8485), .A3(n8484), .A4(n8483), .ZN(n13712) );
  NOR2_X1 U10111 ( .A1(n8487), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8510) );
  INV_X1 U10112 ( .A(n8510), .ZN(n8490) );
  NAND2_X1 U10113 ( .A1(n8487), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8488) );
  MUX2_X1 U10114 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8488), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8489) );
  INV_X1 U10115 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U10116 ( .A1(n11215), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10117 ( .A(n8507), .B(n8506), .ZN(n11221) );
  OR2_X1 U10118 ( .A1(n8923), .A2(n11221), .ZN(n8496) );
  OR2_X1 U10119 ( .A1(n13351), .A2(SI_4_), .ZN(n8495) );
  OAI211_X1 U10120 ( .C1(n11792), .C2(n11724), .A(n8496), .B(n8495), .ZN(
        n13379) );
  XNOR2_X1 U10121 ( .A(n13712), .B(n13379), .ZN(n12482) );
  NAND2_X1 U10122 ( .A1(n12483), .A2(n12482), .ZN(n12481) );
  INV_X1 U10123 ( .A(n13379), .ZN(n12654) );
  NAND2_X1 U10124 ( .A1(n13712), .A2(n12654), .ZN(n8497) );
  NAND2_X1 U10125 ( .A1(n12481), .A2(n8497), .ZN(n12490) );
  INV_X1 U10126 ( .A(n12490), .ZN(n8516) );
  NAND2_X1 U10127 ( .A1(n7437), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10128 ( .A1(n8833), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8504) );
  INV_X1 U10129 ( .A(n8500), .ZN(n8499) );
  INV_X1 U10130 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n11803) );
  NAND2_X1 U10131 ( .A1(n8499), .A2(n11803), .ZN(n8518) );
  NAND2_X1 U10132 ( .A1(n8500), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10133 ( .A1(n8518), .A2(n8501), .ZN(n12669) );
  NAND2_X1 U10134 ( .A1(n8631), .A2(n12669), .ZN(n8503) );
  NAND2_X1 U10135 ( .A1(n13328), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8502) );
  OR2_X1 U10136 ( .A1(n13351), .A2(SI_5_), .ZN(n8514) );
  XNOR2_X1 U10137 ( .A(n8525), .B(n8524), .ZN(n11218) );
  OR2_X1 U10138 ( .A1(n8923), .A2(n11218), .ZN(n8513) );
  OR2_X1 U10139 ( .A1(n8510), .A2(n8626), .ZN(n8508) );
  MUX2_X1 U10140 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8508), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8511) );
  NAND2_X1 U10141 ( .A1(n8510), .A2(n8509), .ZN(n8549) );
  NAND2_X1 U10142 ( .A1(n8511), .A2(n8549), .ZN(n11942) );
  OR2_X1 U10143 ( .A1(n11724), .A2(n11927), .ZN(n8512) );
  NAND2_X1 U10144 ( .A1(n12850), .A2(n12670), .ZN(n13390) );
  INV_X1 U10145 ( .A(n12850), .ZN(n13710) );
  INV_X1 U10146 ( .A(n12670), .ZN(n12499) );
  NAND2_X1 U10147 ( .A1(n13710), .A2(n12499), .ZN(n13387) );
  NAND2_X1 U10148 ( .A1(n8516), .A2(n8515), .ZN(n12492) );
  NAND2_X1 U10149 ( .A1(n12850), .A2(n12499), .ZN(n8517) );
  NAND2_X1 U10150 ( .A1(n13328), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10151 ( .A1(n7437), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10152 ( .A1(n8518), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10153 ( .A1(n8535), .A2(n8519), .ZN(n12857) );
  NAND2_X1 U10154 ( .A1(n8631), .A2(n12857), .ZN(n8521) );
  NAND2_X1 U10155 ( .A1(n8833), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8520) );
  NAND4_X1 U10156 ( .A1(n8523), .A2(n8522), .A3(n8521), .A4(n8520), .ZN(n13709) );
  INV_X1 U10157 ( .A(SI_6_), .ZN(n11196) );
  OR2_X1 U10158 ( .A1(n13351), .A2(n11196), .ZN(n8532) );
  NAND2_X1 U10159 ( .A1(n8525), .A2(n8524), .ZN(n8527) );
  NAND2_X1 U10160 ( .A1(n11211), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8526) );
  XNOR2_X1 U10161 ( .A(n11252), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8541) );
  XNOR2_X1 U10162 ( .A(n8543), .B(n8541), .ZN(n11197) );
  OR2_X1 U10163 ( .A1(n8923), .A2(n11197), .ZN(n8531) );
  NAND2_X1 U10164 ( .A1(n8549), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8529) );
  XNOR2_X1 U10165 ( .A(n8529), .B(n8528), .ZN(n16108) );
  OR2_X1 U10166 ( .A1(n11724), .A2(n16108), .ZN(n8530) );
  XNOR2_X1 U10167 ( .A(n13709), .B(n16406), .ZN(n12849) );
  NAND2_X1 U10168 ( .A1(n13709), .A2(n13391), .ZN(n8533) );
  NAND2_X1 U10169 ( .A1(n7437), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10170 ( .A1(n13328), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8539) );
  INV_X1 U10171 ( .A(n8535), .ZN(n8534) );
  NAND2_X1 U10172 ( .A1(n8534), .A2(n15512), .ZN(n8556) );
  NAND2_X1 U10173 ( .A1(n8535), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10174 ( .A1(n8556), .A2(n8536), .ZN(n12658) );
  NAND2_X1 U10175 ( .A1(n8631), .A2(n12658), .ZN(n8538) );
  NAND2_X1 U10176 ( .A1(n8833), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8537) );
  OR2_X1 U10177 ( .A1(n13351), .A2(SI_7_), .ZN(n8554) );
  INV_X1 U10178 ( .A(n8541), .ZN(n8542) );
  NAND2_X1 U10179 ( .A1(n11252), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10180 ( .A1(n11288), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10181 ( .A1(n11213), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10182 ( .A1(n8568), .A2(n8545), .ZN(n8546) );
  NAND2_X1 U10183 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  AND2_X1 U10184 ( .A1(n8569), .A2(n8548), .ZN(n11201) );
  OR2_X1 U10185 ( .A1(n8923), .A2(n11201), .ZN(n8553) );
  OAI21_X1 U10186 ( .B1(n8549), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8551) );
  INV_X1 U10187 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8550) );
  XNOR2_X1 U10188 ( .A(n8551), .B(n8550), .ZN(n12101) );
  OR2_X1 U10189 ( .A1(n11724), .A2(n12111), .ZN(n8552) );
  NAND2_X1 U10190 ( .A1(n12988), .A2(n12663), .ZN(n13399) );
  INV_X1 U10191 ( .A(n12988), .ZN(n13708) );
  INV_X1 U10192 ( .A(n12663), .ZN(n16430) );
  NAND2_X1 U10193 ( .A1(n13708), .A2(n16430), .ZN(n13400) );
  NAND2_X1 U10194 ( .A1(n13399), .A2(n13400), .ZN(n13514) );
  NAND2_X1 U10195 ( .A1(n13708), .A2(n12663), .ZN(n8555) );
  NAND2_X1 U10196 ( .A1(n12739), .A2(n8555), .ZN(n12986) );
  NAND2_X1 U10197 ( .A1(n13328), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10198 ( .A1(n8958), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10199 ( .A1(n8556), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10200 ( .A1(n8575), .A2(n8557), .ZN(n12990) );
  NAND2_X1 U10201 ( .A1(n8631), .A2(n12990), .ZN(n8560) );
  NAND2_X1 U10202 ( .A1(n8833), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8559) );
  NAND4_X1 U10203 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n13707) );
  NOR2_X1 U10204 ( .A1(n8563), .A2(n8626), .ZN(n8564) );
  MUX2_X1 U10205 ( .A(n8626), .B(n8564), .S(P3_IR_REG_8__SCAN_IN), .Z(n8565)
         );
  INV_X1 U10206 ( .A(n8565), .ZN(n8567) );
  NAND2_X1 U10207 ( .A1(n8567), .A2(n8566), .ZN(n12283) );
  INV_X1 U10208 ( .A(SI_8_), .ZN(n11206) );
  OR2_X1 U10209 ( .A1(n13351), .A2(n11206), .ZN(n8571) );
  XNOR2_X1 U10210 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8582) );
  XNOR2_X1 U10211 ( .A(n8581), .B(n8582), .ZN(n11207) );
  OR2_X1 U10212 ( .A1(n8923), .A2(n11207), .ZN(n8570) );
  OAI211_X1 U10213 ( .C1(n11724), .C2(n12283), .A(n8571), .B(n8570), .ZN(
        n12991) );
  XNOR2_X1 U10214 ( .A(n13707), .B(n12991), .ZN(n13517) );
  INV_X1 U10215 ( .A(n13517), .ZN(n8572) );
  INV_X1 U10216 ( .A(n13707), .ZN(n12974) );
  INV_X1 U10217 ( .A(n12991), .ZN(n16439) );
  NAND2_X1 U10218 ( .A1(n12974), .A2(n16439), .ZN(n8573) );
  NAND2_X1 U10219 ( .A1(n13328), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U10220 ( .A1(n7437), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8579) );
  INV_X1 U10221 ( .A(n8575), .ZN(n8574) );
  NAND2_X1 U10222 ( .A1(n8574), .A2(n15543), .ZN(n8593) );
  NAND2_X1 U10223 ( .A1(n8575), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U10224 ( .A1(n8593), .A2(n8576), .ZN(n12978) );
  NAND2_X1 U10225 ( .A1(n8631), .A2(n12978), .ZN(n8578) );
  NAND2_X1 U10226 ( .A1(n8833), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8577) );
  NAND4_X1 U10227 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n11540) );
  OR2_X1 U10228 ( .A1(n13351), .A2(SI_9_), .ZN(n8592) );
  INV_X1 U10229 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n11247) );
  NAND2_X1 U10230 ( .A1(n11247), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U10231 ( .A1(n11246), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8599) );
  INV_X1 U10232 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n11250) );
  NAND2_X1 U10233 ( .A1(n11250), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U10234 ( .A1(n8599), .A2(n8585), .ZN(n8586) );
  NAND2_X1 U10235 ( .A1(n8587), .A2(n8586), .ZN(n8588) );
  AND2_X1 U10236 ( .A1(n8600), .A2(n8588), .ZN(n11203) );
  OR2_X1 U10237 ( .A1(n8923), .A2(n11203), .ZN(n8591) );
  NAND2_X1 U10238 ( .A1(n8566), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10239 ( .A(n8589), .B(n8402), .ZN(n12681) );
  OR2_X1 U10240 ( .A1(n11724), .A2(n12688), .ZN(n8590) );
  NAND2_X1 U10241 ( .A1(n13328), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10242 ( .A1(n7437), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10243 ( .A1(n8593), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10244 ( .A1(n8614), .A2(n8594), .ZN(n12894) );
  NAND2_X1 U10245 ( .A1(n8932), .A2(n12894), .ZN(n8596) );
  NAND2_X1 U10246 ( .A1(n8833), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10247 ( .A1(n11291), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8620) );
  INV_X1 U10248 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n11285) );
  NAND2_X1 U10249 ( .A1(n11285), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10250 ( .A1(n8620), .A2(n8601), .ZN(n8603) );
  NAND2_X1 U10251 ( .A1(n8602), .A2(n8603), .ZN(n8606) );
  INV_X1 U10252 ( .A(n8603), .ZN(n8604) );
  AND2_X1 U10253 ( .A1(n8606), .A2(n8621), .ZN(n11228) );
  OR2_X1 U10254 ( .A1(n8923), .A2(n11228), .ZN(n8611) );
  OR2_X1 U10255 ( .A1(n13351), .A2(SI_10_), .ZN(n8610) );
  NAND2_X1 U10256 ( .A1(n8607), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8608) );
  XNOR2_X1 U10257 ( .A(n8608), .B(P3_IR_REG_10__SCAN_IN), .ZN(n13762) );
  OR2_X1 U10258 ( .A1(n11724), .A2(n13762), .ZN(n8609) );
  NAND2_X1 U10259 ( .A1(n14086), .A2(n12901), .ZN(n13412) );
  INV_X1 U10260 ( .A(n14086), .ZN(n11619) );
  INV_X1 U10261 ( .A(n12901), .ZN(n16469) );
  NAND2_X1 U10262 ( .A1(n11619), .A2(n16469), .ZN(n13413) );
  NAND2_X1 U10263 ( .A1(n13412), .A2(n13413), .ZN(n13403) );
  NAND2_X1 U10264 ( .A1(n13074), .A2(n13403), .ZN(n8613) );
  NAND2_X1 U10265 ( .A1(n11619), .A2(n12901), .ZN(n8612) );
  NAND2_X1 U10266 ( .A1(n8613), .A2(n8612), .ZN(n14082) );
  NAND2_X1 U10267 ( .A1(n13328), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U10268 ( .A1(n7437), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U10269 ( .A1(n8614), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10270 ( .A1(n8633), .A2(n8615), .ZN(n14093) );
  NAND2_X1 U10271 ( .A1(n8631), .A2(n14093), .ZN(n8617) );
  NAND2_X1 U10272 ( .A1(n8833), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8616) );
  NAND4_X1 U10273 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n13706) );
  NAND2_X1 U10274 ( .A1(n11346), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8639) );
  INV_X1 U10275 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n11348) );
  NAND2_X1 U10276 ( .A1(n11348), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8622) );
  OR2_X1 U10277 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  AND2_X1 U10278 ( .A1(n8625), .A2(n8640), .ZN(n11243) );
  OR2_X1 U10279 ( .A1(n13351), .A2(SI_11_), .ZN(n8629) );
  NOR2_X1 U10280 ( .A1(n8607), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8646) );
  OR2_X1 U10281 ( .A1(n8646), .A2(n8626), .ZN(n8627) );
  XNOR2_X1 U10282 ( .A(n8627), .B(n8645), .ZN(n16134) );
  OR2_X1 U10283 ( .A1(n11724), .A2(n13768), .ZN(n8628) );
  OAI211_X1 U10284 ( .C1(n8923), .C2(n11243), .A(n8629), .B(n8628), .ZN(n16483) );
  INV_X1 U10285 ( .A(n13706), .ZN(n8630) );
  NAND2_X1 U10286 ( .A1(n13328), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10287 ( .A1(n8958), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8637) );
  INV_X1 U10288 ( .A(n8633), .ZN(n8632) );
  NAND2_X1 U10289 ( .A1(n8632), .A2(n15335), .ZN(n8720) );
  NAND2_X1 U10290 ( .A1(n8633), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U10291 ( .A1(n8720), .A2(n8634), .ZN(n13600) );
  NAND2_X1 U10292 ( .A1(n8932), .A2(n13600), .ZN(n8636) );
  NAND2_X1 U10293 ( .A1(n8833), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8635) );
  NAND4_X1 U10294 ( .A1(n8638), .A2(n8637), .A3(n8636), .A4(n8635), .ZN(n13656) );
  NAND2_X1 U10295 ( .A1(n8640), .A2(n8639), .ZN(n8643) );
  NAND2_X1 U10296 ( .A1(n11438), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U10297 ( .A1(n11440), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U10298 ( .A1(n8643), .A2(n8642), .ZN(n8657) );
  OR2_X1 U10299 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  NAND2_X1 U10300 ( .A1(n8657), .A2(n8644), .ZN(n11254) );
  NAND2_X1 U10301 ( .A1(n13353), .A2(n11254), .ZN(n8654) );
  OR2_X1 U10302 ( .A1(n13351), .A2(SI_12_), .ZN(n8653) );
  AND2_X1 U10303 ( .A1(n8646), .A2(n8645), .ZN(n8649) );
  NOR2_X1 U10304 ( .A1(n8649), .A2(n8626), .ZN(n8647) );
  MUX2_X1 U10305 ( .A(n8626), .B(n8647), .S(P3_IR_REG_12__SCAN_IN), .Z(n8651)
         );
  NAND2_X1 U10306 ( .A1(n8649), .A2(n8648), .ZN(n8715) );
  INV_X1 U10307 ( .A(n8715), .ZN(n8650) );
  OR2_X1 U10308 ( .A1(n11724), .A2(n13741), .ZN(n8652) );
  NAND2_X1 U10309 ( .A1(n8655), .A2(n8381), .ZN(n14002) );
  NAND2_X1 U10310 ( .A1(n13656), .A2(n14077), .ZN(n14001) );
  NAND2_X1 U10311 ( .A1(n8657), .A2(n8656), .ZN(n8659) );
  INV_X1 U10312 ( .A(n8659), .ZN(n8658) );
  INV_X1 U10313 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U10314 ( .A1(n11545), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U10315 ( .A1(n11547), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U10316 ( .A1(n8677), .A2(n8663), .ZN(n8666) );
  NAND2_X1 U10317 ( .A1(n11717), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U10318 ( .A1(n11719), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U10319 ( .A1(n8666), .A2(n8665), .ZN(n8695) );
  OAI21_X1 U10320 ( .B1(n8666), .B2(n8665), .A(n8695), .ZN(n11441) );
  OR2_X1 U10321 ( .A1(n11441), .A2(n8923), .ZN(n8669) );
  INV_X1 U10322 ( .A(n11724), .ZN(n8779) );
  OAI21_X1 U10323 ( .B1(n8680), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8667) );
  XNOR2_X1 U10324 ( .A(n8667), .B(P3_IR_REG_15__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U10325 ( .A1(n8780), .A2(SI_15_), .B1(n8779), .B2(n16197), .ZN(
        n8668) );
  NAND2_X1 U10326 ( .A1(n13328), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U10327 ( .A1(n8958), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8675) );
  INV_X1 U10328 ( .A(n8720), .ZN(n8670) );
  NAND2_X1 U10329 ( .A1(n8670), .A2(n15554), .ZN(n8722) );
  NAND2_X1 U10330 ( .A1(n8686), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U10331 ( .A1(n8705), .A2(n8672), .ZN(n14031) );
  NAND2_X1 U10332 ( .A1(n8631), .A2(n14031), .ZN(n8674) );
  NAND2_X1 U10333 ( .A1(n8833), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8673) );
  NAND4_X1 U10334 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n13625) );
  NAND2_X1 U10335 ( .A1(n16610), .A2(n13625), .ZN(n13430) );
  NAND2_X1 U10336 ( .A1(n13137), .A2(n14039), .ZN(n13947) );
  NAND2_X1 U10337 ( .A1(n13430), .A2(n13947), .ZN(n14025) );
  INV_X1 U10338 ( .A(n14025), .ZN(n8691) );
  OAI21_X1 U10339 ( .B1(n8679), .B2(n8678), .A(n8677), .ZN(n11410) );
  NAND2_X1 U10340 ( .A1(n11410), .A2(n13353), .ZN(n8684) );
  NAND2_X1 U10341 ( .A1(n8680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8682) );
  INV_X1 U10342 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8681) );
  AOI22_X1 U10343 ( .A1(n8780), .A2(n11411), .B1(n8779), .B2(n16185), .ZN(
        n8683) );
  NAND2_X1 U10344 ( .A1(n13328), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U10345 ( .A1(n8958), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U10346 ( .A1(n8722), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U10347 ( .A1(n8686), .A2(n8685), .ZN(n14044) );
  NAND2_X1 U10348 ( .A1(n8631), .A2(n14044), .ZN(n8688) );
  NAND2_X1 U10349 ( .A1(n8833), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8687) );
  NAND4_X1 U10350 ( .A1(n8690), .A2(n8689), .A3(n8688), .A4(n8687), .ZN(n13655) );
  INV_X1 U10351 ( .A(n13655), .ZN(n14055) );
  OR2_X1 U10352 ( .A1(n16534), .A2(n14055), .ZN(n14023) );
  OR2_X1 U10353 ( .A1(n8691), .A2(n14023), .ZN(n8693) );
  NAND2_X1 U10354 ( .A1(n13137), .A2(n13625), .ZN(n8692) );
  AND2_X1 U10355 ( .A1(n8693), .A2(n8692), .ZN(n14006) );
  NAND2_X1 U10356 ( .A1(n8695), .A2(n8694), .ZN(n8698) );
  NAND2_X1 U10357 ( .A1(n11900), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U10358 ( .A1(n11902), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8696) );
  OR2_X1 U10359 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  AND2_X1 U10360 ( .A1(n8730), .A2(n8699), .ZN(n11548) );
  NAND2_X1 U10361 ( .A1(n11548), .A2(n13353), .ZN(n8704) );
  NAND2_X1 U10362 ( .A1(n8700), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8701) );
  MUX2_X1 U10363 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8701), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8702) );
  AND2_X1 U10364 ( .A1(n8702), .A2(n7559), .ZN(n16213) );
  AOI22_X1 U10365 ( .A1(n8780), .A2(SI_16_), .B1(n8779), .B2(n16213), .ZN(
        n8703) );
  NAND2_X1 U10366 ( .A1(n7437), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U10367 ( .A1(n13328), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U10368 ( .A1(n8705), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U10369 ( .A1(n8755), .A2(n8706), .ZN(n14016) );
  NAND2_X1 U10370 ( .A1(n8932), .A2(n14016), .ZN(n8708) );
  NAND2_X1 U10371 ( .A1(n8833), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U10372 ( .A1(n14208), .A2(n14028), .ZN(n13984) );
  INV_X1 U10373 ( .A(n14208), .ZN(n8976) );
  INV_X1 U10374 ( .A(n14028), .ZN(n13988) );
  NAND2_X1 U10375 ( .A1(n8976), .A2(n13988), .ZN(n13438) );
  NAND2_X1 U10376 ( .A1(n13984), .A2(n13438), .ZN(n14014) );
  INV_X1 U10377 ( .A(n14014), .ZN(n8711) );
  AND2_X1 U10378 ( .A1(n14006), .A2(n8711), .ZN(n8728) );
  XNOR2_X1 U10379 ( .A(n16534), .B(n13655), .ZN(n14041) );
  AND2_X1 U10380 ( .A1(n14041), .A2(n14025), .ZN(n8766) );
  INV_X1 U10381 ( .A(n8766), .ZN(n8727) );
  NAND2_X1 U10382 ( .A1(n8712), .A2(n8077), .ZN(n8713) );
  NAND2_X1 U10383 ( .A1(n8714), .A2(n8713), .ZN(n11343) );
  NAND2_X1 U10384 ( .A1(n11343), .A2(n13353), .ZN(n8719) );
  NAND2_X1 U10385 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8717) );
  INV_X1 U10386 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8716) );
  XNOR2_X1 U10387 ( .A(n8717), .B(n8716), .ZN(n13776) );
  AOI22_X1 U10388 ( .A1(n8780), .A2(n15488), .B1(n8779), .B2(n13776), .ZN(
        n8718) );
  NAND2_X1 U10389 ( .A1(n8719), .A2(n8718), .ZN(n16517) );
  INV_X1 U10390 ( .A(n16517), .ZN(n14061) );
  NAND2_X1 U10391 ( .A1(n13328), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U10392 ( .A1(n7437), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U10393 ( .A1(n8720), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U10394 ( .A1(n8722), .A2(n8721), .ZN(n13654) );
  NAND2_X1 U10395 ( .A1(n8631), .A2(n13654), .ZN(n8724) );
  NAND2_X1 U10396 ( .A1(n8833), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8723) );
  NAND4_X1 U10397 ( .A1(n8726), .A2(n8725), .A3(n8724), .A4(n8723), .ZN(n14036) );
  NAND2_X1 U10398 ( .A1(n14061), .A2(n14036), .ZN(n14021) );
  OR2_X1 U10399 ( .A1(n8727), .A2(n14021), .ZN(n14004) );
  AND2_X1 U10400 ( .A1(n8728), .A2(n14004), .ZN(n8764) );
  AND2_X1 U10401 ( .A1(n14001), .A2(n8764), .ZN(n13959) );
  NAND2_X1 U10402 ( .A1(n12064), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U10403 ( .A1(n12066), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U10404 ( .A1(n12340), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10405 ( .A1(n12338), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8733) );
  OR2_X1 U10406 ( .A1(n8735), .A2(n8734), .ZN(n8736) );
  NAND2_X1 U10407 ( .A1(n8773), .A2(n8736), .ZN(n11693) );
  OR2_X1 U10408 ( .A1(n11693), .A2(n8923), .ZN(n8740) );
  NAND2_X1 U10409 ( .A1(n8737), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8738) );
  XNOR2_X1 U10410 ( .A(n8738), .B(P3_IR_REG_18__SCAN_IN), .ZN(n16253) );
  AOI22_X1 U10411 ( .A1(n8780), .A2(SI_18_), .B1(n8779), .B2(n16253), .ZN(
        n8739) );
  NAND2_X1 U10412 ( .A1(n13328), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U10413 ( .A1(n8958), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U10414 ( .A1(n8757), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U10415 ( .A1(n8784), .A2(n8742), .ZN(n13974) );
  NAND2_X1 U10416 ( .A1(n8932), .A2(n13974), .ZN(n8744) );
  NAND2_X1 U10417 ( .A1(n8833), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8743) );
  NAND4_X1 U10418 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(n13985) );
  NAND2_X1 U10419 ( .A1(n14199), .A2(n13985), .ZN(n13452) );
  INV_X1 U10420 ( .A(n14199), .ZN(n8747) );
  NAND2_X1 U10421 ( .A1(n8747), .A2(n13946), .ZN(n13450) );
  NAND2_X1 U10422 ( .A1(n13452), .A2(n13450), .ZN(n13961) );
  OR2_X1 U10423 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  NAND2_X1 U10424 ( .A1(n8751), .A2(n8750), .ZN(n11637) );
  OR2_X1 U10425 ( .A1(n11637), .A2(n8923), .ZN(n8754) );
  NAND2_X1 U10426 ( .A1(n7559), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8752) );
  XNOR2_X1 U10427 ( .A(n8752), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U10428 ( .A1(n8780), .A2(SI_17_), .B1(n8779), .B2(n13756), .ZN(
        n8753) );
  NAND2_X1 U10429 ( .A1(n13328), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U10430 ( .A1(n8958), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U10431 ( .A1(n8755), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U10432 ( .A1(n8757), .A2(n8756), .ZN(n13996) );
  NAND2_X1 U10433 ( .A1(n8932), .A2(n13996), .ZN(n8759) );
  NAND2_X1 U10434 ( .A1(n8833), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8758) );
  INV_X1 U10435 ( .A(n14012), .ZN(n13705) );
  NAND2_X1 U10436 ( .A1(n13449), .A2(n13705), .ZN(n13962) );
  AND2_X1 U10437 ( .A1(n13961), .A2(n13962), .ZN(n8763) );
  AND2_X1 U10438 ( .A1(n13959), .A2(n8763), .ZN(n8762) );
  NAND2_X1 U10439 ( .A1(n14002), .A2(n8762), .ZN(n13958) );
  NAND2_X1 U10440 ( .A1(n14199), .A2(n13946), .ZN(n8770) );
  INV_X1 U10441 ( .A(n8763), .ZN(n8769) );
  AND2_X1 U10442 ( .A1(n13983), .A2(n13984), .ZN(n8768) );
  INV_X1 U10443 ( .A(n8764), .ZN(n8767) );
  NAND2_X1 U10444 ( .A1(n16517), .A2(n14036), .ZN(n8765) );
  NAND2_X1 U10445 ( .A1(n14040), .A2(n8765), .ZN(n14053) );
  AND2_X1 U10446 ( .A1(n14053), .A2(n8766), .ZN(n14003) );
  OR2_X1 U10447 ( .A1(n8767), .A2(n14003), .ZN(n13981) );
  AND2_X1 U10448 ( .A1(n8768), .A2(n13981), .ZN(n13960) );
  OR2_X1 U10449 ( .A1(n8769), .A2(n13960), .ZN(n13957) );
  AND2_X1 U10450 ( .A1(n8770), .A2(n13957), .ZN(n8771) );
  NAND2_X1 U10451 ( .A1(n13958), .A2(n8771), .ZN(n13943) );
  INV_X1 U10452 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U10453 ( .A1(n12538), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8792) );
  INV_X1 U10454 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12540) );
  NAND2_X1 U10455 ( .A1(n12540), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8774) );
  OR2_X1 U10456 ( .A1(n8776), .A2(n8775), .ZN(n8777) );
  NAND2_X1 U10457 ( .A1(n8793), .A2(n8777), .ZN(n11881) );
  OR2_X1 U10458 ( .A1(n11881), .A2(n8923), .ZN(n8782) );
  NAND2_X1 U10459 ( .A1(n8944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8778) );
  AOI22_X1 U10460 ( .A1(n8780), .A2(SI_19_), .B1(n13736), .B2(n8779), .ZN(
        n8781) );
  NAND2_X1 U10461 ( .A1(n8958), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8789) );
  INV_X1 U10462 ( .A(n8784), .ZN(n8783) );
  NAND2_X1 U10463 ( .A1(n8784), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U10464 ( .A1(n8801), .A2(n8785), .ZN(n13952) );
  NAND2_X1 U10465 ( .A1(n8932), .A2(n13952), .ZN(n8788) );
  NAND2_X1 U10466 ( .A1(n13328), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U10467 ( .A1(n8833), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8786) );
  NAND4_X1 U10468 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n13704) );
  NAND2_X1 U10469 ( .A1(n13570), .A2(n13704), .ZN(n8790) );
  OR2_X1 U10470 ( .A1(n13570), .A2(n13704), .ZN(n8791) );
  NAND2_X1 U10471 ( .A1(n8793), .A2(n8792), .ZN(n8794) );
  INV_X1 U10472 ( .A(n8794), .ZN(n8796) );
  INV_X1 U10473 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U10474 ( .A1(n8797), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U10475 ( .A1(n8808), .A2(n8798), .ZN(n12194) );
  OR2_X1 U10476 ( .A1(n12194), .A2(n8923), .ZN(n8800) );
  INV_X1 U10477 ( .A(SI_20_), .ZN(n12193) );
  NAND2_X1 U10478 ( .A1(n8958), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U10479 ( .A1(n8498), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U10480 ( .A1(n8801), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U10481 ( .A1(n8818), .A2(n8802), .ZN(n13939) );
  NAND2_X1 U10482 ( .A1(n8932), .A2(n13939), .ZN(n8804) );
  NAND2_X1 U10483 ( .A1(n13328), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8803) );
  OR2_X1 U10484 ( .A1(n13940), .A2(n13945), .ZN(n13458) );
  NAND2_X1 U10485 ( .A1(n13940), .A2(n13945), .ZN(n13906) );
  NAND2_X1 U10486 ( .A1(n13940), .A2(n13915), .ZN(n8807) );
  NAND2_X1 U10487 ( .A1(n12810), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U10488 ( .A1(n12807), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U10489 ( .A1(n8811), .A2(n8810), .ZN(n8825) );
  OR2_X1 U10490 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  NAND2_X1 U10491 ( .A1(n8825), .A2(n8812), .ZN(n12415) );
  OR2_X1 U10492 ( .A1(n12415), .A2(n8923), .ZN(n8814) );
  INV_X1 U10493 ( .A(SI_21_), .ZN(n12414) );
  OR2_X1 U10494 ( .A1(n13351), .A2(n12414), .ZN(n8813) );
  NAND2_X1 U10495 ( .A1(n13328), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U10496 ( .A1(n8958), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8815) );
  AND2_X1 U10497 ( .A1(n8816), .A2(n8815), .ZN(n8822) );
  NAND2_X1 U10498 ( .A1(n8818), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U10499 ( .A1(n8834), .A2(n8819), .ZN(n13920) );
  NAND2_X1 U10500 ( .A1(n13920), .A2(n8932), .ZN(n8821) );
  NAND2_X1 U10501 ( .A1(n8498), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U10502 ( .A1(n14182), .A2(n13933), .ZN(n8823) );
  NAND2_X1 U10503 ( .A1(n13921), .A2(n13703), .ZN(n10488) );
  NAND2_X1 U10504 ( .A1(n8825), .A2(n8824), .ZN(n8828) );
  INV_X1 U10505 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U10506 ( .A1(n9655), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8841) );
  INV_X1 U10507 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U10508 ( .A1(n13039), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U10509 ( .A1(n8828), .A2(n8827), .ZN(n8842) );
  OR2_X1 U10510 ( .A1(n8828), .A2(n8827), .ZN(n8829) );
  NAND2_X1 U10511 ( .A1(n8842), .A2(n8829), .ZN(n12447) );
  OR2_X1 U10512 ( .A1(n12447), .A2(n8923), .ZN(n8832) );
  INV_X1 U10513 ( .A(SI_22_), .ZN(n8830) );
  INV_X1 U10514 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U10515 ( .A1(n8834), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U10516 ( .A1(n8845), .A2(n8835), .ZN(n13902) );
  NAND2_X1 U10517 ( .A1(n13902), .A2(n8932), .ZN(n8837) );
  AOI22_X1 U10518 ( .A1(n13328), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n8958), 
        .B2(P3_REG0_REG_22__SCAN_IN), .ZN(n8836) );
  INV_X1 U10519 ( .A(n13903), .ZN(n14177) );
  INV_X1 U10520 ( .A(n13914), .ZN(n13596) );
  NAND2_X1 U10521 ( .A1(n14177), .A2(n13596), .ZN(n8839) );
  NAND2_X1 U10522 ( .A1(n8840), .A2(n8839), .ZN(n13882) );
  NAND2_X1 U10523 ( .A1(n8842), .A2(n8841), .ZN(n8852) );
  XNOR2_X1 U10524 ( .A(n13003), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8851) );
  XNOR2_X1 U10525 ( .A(n8852), .B(n8851), .ZN(n12606) );
  NAND2_X1 U10526 ( .A1(n12606), .A2(n13353), .ZN(n8844) );
  INV_X1 U10527 ( .A(SI_23_), .ZN(n12608) );
  NAND2_X1 U10528 ( .A1(n8845), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U10529 ( .A1(n8856), .A2(n8846), .ZN(n13887) );
  NAND2_X1 U10530 ( .A1(n13887), .A2(n8932), .ZN(n8849) );
  AOI22_X1 U10531 ( .A1(n13328), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n7437), 
        .B2(P3_REG0_REG_23__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U10532 ( .A1(n8498), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U10533 ( .A1(n13563), .A2(n13897), .ZN(n13472) );
  INV_X1 U10534 ( .A(n13897), .ZN(n13871) );
  NAND2_X1 U10535 ( .A1(n13003), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8850) );
  XNOR2_X1 U10536 ( .A(n8862), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U10537 ( .A1(n12904), .A2(n13353), .ZN(n8854) );
  INV_X1 U10538 ( .A(SI_24_), .ZN(n12905) );
  INV_X1 U10539 ( .A(n8856), .ZN(n8855) );
  INV_X1 U10540 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15544) );
  NAND2_X1 U10541 ( .A1(n8855), .A2(n15544), .ZN(n8869) );
  NAND2_X1 U10542 ( .A1(n8856), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U10543 ( .A1(n8869), .A2(n8857), .ZN(n13876) );
  INV_X1 U10544 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U10545 ( .A1(n8498), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U10546 ( .A1(n7437), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8858) );
  OAI211_X1 U10547 ( .C1(n8962), .C2(n14120), .A(n8859), .B(n8858), .ZN(n8860)
         );
  AOI21_X1 U10548 ( .B1(n13876), .B2(n8932), .A(n8860), .ZN(n13859) );
  OR2_X1 U10549 ( .A1(n13637), .A2(n13859), .ZN(n13490) );
  NAND2_X1 U10550 ( .A1(n13637), .A2(n13859), .ZN(n13485) );
  NAND2_X1 U10551 ( .A1(n13490), .A2(n13485), .ZN(n13873) );
  INV_X1 U10552 ( .A(n13859), .ZN(n13884) );
  OR2_X1 U10553 ( .A1(n13637), .A2(n13884), .ZN(n8861) );
  INV_X1 U10554 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15809) );
  NAND2_X1 U10555 ( .A1(n15809), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8881) );
  INV_X1 U10556 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U10557 ( .A1(n14791), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U10558 ( .A1(n8881), .A2(n8865), .ZN(n8878) );
  XNOR2_X1 U10559 ( .A(n8880), .B(n8878), .ZN(n13011) );
  NAND2_X1 U10560 ( .A1(n13011), .A2(n13353), .ZN(n8867) );
  OR2_X1 U10561 ( .A1(n13351), .A2(n15466), .ZN(n8866) );
  INV_X1 U10562 ( .A(n8869), .ZN(n8868) );
  INV_X1 U10563 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15533) );
  NAND2_X1 U10564 ( .A1(n8868), .A2(n15533), .ZN(n8889) );
  NAND2_X1 U10565 ( .A1(n8869), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U10566 ( .A1(n8889), .A2(n8870), .ZN(n13865) );
  NAND2_X1 U10567 ( .A1(n13865), .A2(n8932), .ZN(n8875) );
  INV_X1 U10568 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U10569 ( .A1(n8498), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U10570 ( .A1(n8958), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8871) );
  OAI211_X1 U10571 ( .C1(n8962), .C2(n14114), .A(n8872), .B(n8871), .ZN(n8873)
         );
  INV_X1 U10572 ( .A(n8873), .ZN(n8874) );
  NAND2_X1 U10573 ( .A1(n14164), .A2(n13838), .ZN(n13840) );
  OR2_X1 U10574 ( .A1(n14164), .A2(n13838), .ZN(n8876) );
  NAND2_X1 U10575 ( .A1(n13840), .A2(n8876), .ZN(n13855) );
  NAND2_X1 U10576 ( .A1(n13856), .A2(n13855), .ZN(n13854) );
  NAND2_X1 U10577 ( .A1(n14164), .A2(n13870), .ZN(n8877) );
  NAND2_X1 U10578 ( .A1(n13854), .A2(n8877), .ZN(n13836) );
  INV_X1 U10579 ( .A(n8878), .ZN(n8879) );
  NAND2_X1 U10580 ( .A1(n8882), .A2(n8881), .ZN(n8885) );
  INV_X1 U10581 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U10582 ( .A1(n9726), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8897) );
  INV_X1 U10583 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14787) );
  NAND2_X1 U10584 ( .A1(n14787), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8883) );
  AND2_X1 U10585 ( .A1(n8897), .A2(n8883), .ZN(n8884) );
  NAND2_X1 U10586 ( .A1(n8885), .A2(n8884), .ZN(n8898) );
  OR2_X1 U10587 ( .A1(n8885), .A2(n8884), .ZN(n8886) );
  NAND2_X1 U10588 ( .A1(n8898), .A2(n8886), .ZN(n13068) );
  NAND2_X1 U10589 ( .A1(n8889), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U10590 ( .A1(n8906), .A2(n8890), .ZN(n13845) );
  NAND2_X1 U10591 ( .A1(n13845), .A2(n8932), .ZN(n8895) );
  INV_X1 U10592 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U10593 ( .A1(n8498), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U10594 ( .A1(n8958), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8891) );
  OAI211_X1 U10595 ( .C1(n8962), .C2(n14111), .A(n8892), .B(n8891), .ZN(n8893)
         );
  INV_X1 U10596 ( .A(n8893), .ZN(n8894) );
  NAND2_X2 U10597 ( .A1(n8895), .A2(n8894), .ZN(n13857) );
  OR2_X1 U10598 ( .A1(n13686), .A2(n13857), .ZN(n8896) );
  NAND2_X1 U10599 ( .A1(n8898), .A2(n8897), .ZN(n8902) );
  INV_X1 U10600 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U10601 ( .A1(n8899), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8917) );
  INV_X1 U10602 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14785) );
  NAND2_X1 U10603 ( .A1(n14785), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8900) );
  AND2_X1 U10604 ( .A1(n8917), .A2(n8900), .ZN(n8901) );
  NAND2_X1 U10605 ( .A1(n8902), .A2(n8901), .ZN(n8918) );
  INV_X1 U10606 ( .A(SI_27_), .ZN(n15461) );
  INV_X1 U10607 ( .A(n8906), .ZN(n8905) );
  INV_X1 U10608 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U10609 ( .A1(n8905), .A2(n8904), .ZN(n8926) );
  NAND2_X1 U10610 ( .A1(n8906), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U10611 ( .A1(n8926), .A2(n8907), .ZN(n13831) );
  NAND2_X1 U10612 ( .A1(n13831), .A2(n8932), .ZN(n8913) );
  INV_X1 U10613 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U10614 ( .A1(n8498), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U10615 ( .A1(n7437), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8908) );
  OAI211_X1 U10616 ( .C1(n8962), .C2(n8910), .A(n8909), .B(n8908), .ZN(n8911)
         );
  INV_X1 U10617 ( .A(n8911), .ZN(n8912) );
  NAND2_X1 U10618 ( .A1(n8915), .A2(n13839), .ZN(n13482) );
  OR2_X1 U10619 ( .A1(n8915), .A2(n13702), .ZN(n8916) );
  NAND2_X1 U10620 ( .A1(n8918), .A2(n8917), .ZN(n8921) );
  NAND2_X1 U10621 ( .A1(n15798), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8934) );
  INV_X1 U10622 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U10623 ( .A1(n14782), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8919) );
  AND2_X1 U10624 ( .A1(n8934), .A2(n8919), .ZN(n8920) );
  NAND2_X1 U10625 ( .A1(n8921), .A2(n8920), .ZN(n8935) );
  OR2_X1 U10626 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  NAND2_X1 U10627 ( .A1(n8935), .A2(n8922), .ZN(n13248) );
  OR2_X1 U10628 ( .A1(n13248), .A2(n8923), .ZN(n8925) );
  INV_X1 U10629 ( .A(SI_28_), .ZN(n15459) );
  OR2_X1 U10630 ( .A1(n13351), .A2(n15459), .ZN(n8924) );
  NAND2_X1 U10631 ( .A1(n8926), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8927) );
  NAND2_X1 U10632 ( .A1(n13807), .A2(n8927), .ZN(n13821) );
  INV_X1 U10633 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U10634 ( .A1(n8498), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U10635 ( .A1(n8958), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8928) );
  OAI211_X1 U10636 ( .C1(n8962), .C2(n8930), .A(n8929), .B(n8928), .ZN(n8931)
         );
  AOI21_X1 U10637 ( .B1(n13821), .B2(n8932), .A(n8931), .ZN(n8957) );
  OR2_X1 U10638 ( .A1(n13245), .A2(n8957), .ZN(n13497) );
  NAND2_X1 U10639 ( .A1(n13245), .A2(n8957), .ZN(n13496) );
  NAND2_X1 U10640 ( .A1(n13497), .A2(n13496), .ZN(n13237) );
  NAND2_X1 U10641 ( .A1(n9062), .A2(n13237), .ZN(n9066) );
  NAND2_X1 U10642 ( .A1(n9066), .A2(n8933), .ZN(n8943) );
  NAND2_X1 U10643 ( .A1(n8935), .A2(n8934), .ZN(n13336) );
  INV_X1 U10644 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13337) );
  XNOR2_X1 U10645 ( .A(n13337), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n13334) );
  XNOR2_X1 U10646 ( .A(n13336), .B(n13334), .ZN(n14219) );
  INV_X1 U10647 ( .A(SI_29_), .ZN(n15460) );
  NOR2_X1 U10648 ( .A1(n13351), .A2(n15460), .ZN(n8936) );
  INV_X1 U10649 ( .A(n13807), .ZN(n8937) );
  NAND2_X1 U10650 ( .A1(n8937), .A2(n8932), .ZN(n13333) );
  INV_X1 U10651 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10652 ( .A1(n8958), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U10653 ( .A1(n8498), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8938) );
  OAI211_X1 U10654 ( .C1(n8962), .C2(n9057), .A(n8939), .B(n8938), .ZN(n8940)
         );
  INV_X1 U10655 ( .A(n8940), .ZN(n8941) );
  NAND2_X1 U10656 ( .A1(n13333), .A2(n8941), .ZN(n12512) );
  NAND2_X1 U10657 ( .A1(n13815), .A2(n12512), .ZN(n13498) );
  INV_X1 U10658 ( .A(n13815), .ZN(n8942) );
  INV_X1 U10659 ( .A(n12512), .ZN(n13242) );
  NAND2_X1 U10660 ( .A1(n8942), .A2(n13242), .ZN(n13343) );
  NAND2_X1 U10661 ( .A1(n13498), .A2(n13343), .ZN(n13509) );
  XNOR2_X1 U10662 ( .A(n8943), .B(n13509), .ZN(n8968) );
  NAND2_X1 U10663 ( .A1(n9034), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U10664 ( .A1(n13544), .A2(n13736), .ZN(n9031) );
  INV_X1 U10665 ( .A(n8948), .ZN(n8954) );
  NAND2_X1 U10666 ( .A1(n8954), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8949) );
  INV_X1 U10667 ( .A(n8951), .ZN(n8952) );
  NAND2_X1 U10668 ( .A1(n8952), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8953) );
  MUX2_X1 U10669 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8953), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8955) );
  INV_X1 U10670 ( .A(n12192), .ZN(n9030) );
  NAND2_X1 U10671 ( .A1(n13363), .A2(n9030), .ZN(n13358) );
  OR2_X1 U10672 ( .A1(n8956), .A2(n7414), .ZN(n11740) );
  NAND2_X1 U10673 ( .A1(n11740), .A2(n11724), .ZN(n10517) );
  INV_X1 U10674 ( .A(n10517), .ZN(n10529) );
  INV_X1 U10675 ( .A(n8957), .ZN(n13829) );
  INV_X1 U10676 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U10677 ( .A1(n8498), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U10678 ( .A1(n8958), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8959) );
  OAI211_X1 U10679 ( .C1(n8962), .C2(n8961), .A(n8960), .B(n8959), .ZN(n8963)
         );
  INV_X1 U10680 ( .A(n8963), .ZN(n8964) );
  NAND2_X1 U10681 ( .A1(n13333), .A2(n8964), .ZN(n13701) );
  INV_X1 U10682 ( .A(P3_B_REG_SCAN_IN), .ZN(n8965) );
  NOR2_X1 U10683 ( .A1(n8956), .A2(n8965), .ZN(n8966) );
  NOR2_X1 U10684 ( .A1(n14089), .A2(n8966), .ZN(n13805) );
  AOI22_X1 U10685 ( .A1(n13987), .A2(n13829), .B1(n13701), .B2(n13805), .ZN(
        n8967) );
  INV_X1 U10686 ( .A(n13585), .ZN(n8969) );
  NAND2_X1 U10687 ( .A1(n8969), .A2(n12443), .ZN(n12404) );
  NAND2_X1 U10688 ( .A1(n8388), .A2(n8970), .ZN(n12329) );
  NAND2_X1 U10689 ( .A1(n12329), .A2(n13374), .ZN(n12425) );
  INV_X1 U10690 ( .A(n13515), .ZN(n12429) );
  NAND2_X1 U10691 ( .A1(n12425), .A2(n12429), .ZN(n8971) );
  NAND2_X2 U10692 ( .A1(n8971), .A2(n13376), .ZN(n12480) );
  INV_X1 U10693 ( .A(n13712), .ZN(n12531) );
  NAND2_X1 U10694 ( .A1(n12531), .A2(n12654), .ZN(n13381) );
  NAND2_X1 U10695 ( .A1(n12847), .A2(n13516), .ZN(n8972) );
  INV_X1 U10696 ( .A(n13709), .ZN(n13392) );
  NAND2_X1 U10697 ( .A1(n13392), .A2(n13391), .ZN(n13388) );
  INV_X1 U10698 ( .A(n13514), .ZN(n13397) );
  NAND2_X1 U10699 ( .A1(n12974), .A2(n12991), .ZN(n13405) );
  NOR2_X1 U10700 ( .A1(n11540), .A2(n16462), .ZN(n13409) );
  NAND2_X1 U10701 ( .A1(n11540), .A2(n16462), .ZN(n12971) );
  INV_X1 U10702 ( .A(n16483), .ZN(n14094) );
  NAND2_X1 U10703 ( .A1(n8630), .A2(n14094), .ZN(n13418) );
  NAND2_X1 U10704 ( .A1(n13706), .A2(n16483), .ZN(n13424) );
  NAND2_X1 U10705 ( .A1(n14092), .A2(n14091), .ZN(n14090) );
  NAND2_X1 U10706 ( .A1(n14090), .A2(n13418), .ZN(n14066) );
  NAND2_X1 U10707 ( .A1(n14088), .A2(n14077), .ZN(n13426) );
  INV_X1 U10708 ( .A(n14077), .ZN(n16502) );
  NAND2_X1 U10709 ( .A1(n13656), .A2(n16502), .ZN(n13423) );
  NAND2_X1 U10710 ( .A1(n14066), .A2(n14068), .ZN(n14065) );
  NAND2_X1 U10711 ( .A1(n14065), .A2(n13426), .ZN(n14052) );
  NAND2_X1 U10712 ( .A1(n14052), .A2(n14051), .ZN(n14050) );
  NAND2_X1 U10713 ( .A1(n14050), .A2(n14040), .ZN(n8974) );
  INV_X1 U10714 ( .A(n14041), .ZN(n13527) );
  NAND2_X1 U10715 ( .A1(n8974), .A2(n13527), .ZN(n14043) );
  OR2_X1 U10716 ( .A1(n16534), .A2(n13655), .ZN(n13431) );
  NAND2_X1 U10717 ( .A1(n14043), .A2(n13431), .ZN(n14030) );
  INV_X1 U10718 ( .A(n13510), .ZN(n8980) );
  AND2_X1 U10719 ( .A1(n13570), .A2(n13965), .ZN(n13447) );
  INV_X1 U10720 ( .A(n13447), .ZN(n13511) );
  NAND2_X1 U10721 ( .A1(n13449), .A2(n14012), .ZN(n13445) );
  INV_X1 U10722 ( .A(n13445), .ZN(n8975) );
  OR2_X1 U10723 ( .A1(n8975), .A2(n13994), .ZN(n8983) );
  INV_X1 U10724 ( .A(n8983), .ZN(n8978) );
  NAND2_X1 U10725 ( .A1(n8976), .A2(n14028), .ZN(n13992) );
  AND2_X1 U10726 ( .A1(n13992), .A2(n13445), .ZN(n8977) );
  OR2_X1 U10727 ( .A1(n13961), .A2(n13967), .ZN(n13969) );
  AND2_X1 U10728 ( .A1(n13450), .A2(n13969), .ZN(n13949) );
  AND2_X1 U10729 ( .A1(n13511), .A2(n13949), .ZN(n8979) );
  OR2_X2 U10730 ( .A1(n8980), .A2(n8979), .ZN(n8982) );
  AND2_X1 U10731 ( .A1(n8982), .A2(n13947), .ZN(n8981) );
  NAND2_X1 U10732 ( .A1(n14029), .A2(n8981), .ZN(n8987) );
  INV_X1 U10733 ( .A(n8982), .ZN(n8985) );
  AND2_X1 U10734 ( .A1(n8983), .A2(n14014), .ZN(n13966) );
  INV_X1 U10735 ( .A(n13961), .ZN(n13972) );
  AND2_X1 U10736 ( .A1(n13966), .A2(n13972), .ZN(n13948) );
  AND2_X1 U10737 ( .A1(n13948), .A2(n13510), .ZN(n8984) );
  NAND2_X1 U10738 ( .A1(n14182), .A2(n13703), .ZN(n13463) );
  NAND2_X1 U10739 ( .A1(n13921), .A2(n13933), .ZN(n13462) );
  NAND2_X1 U10740 ( .A1(n13463), .A2(n13462), .ZN(n13907) );
  INV_X1 U10741 ( .A(n13906), .ZN(n8988) );
  NOR2_X1 U10742 ( .A1(n13907), .A2(n8988), .ZN(n8989) );
  NOR2_X1 U10743 ( .A1(n13903), .A2(n13596), .ZN(n13467) );
  NAND2_X1 U10744 ( .A1(n13903), .A2(n13596), .ZN(n13461) );
  OR2_X1 U10745 ( .A1(n13880), .A2(n7935), .ZN(n8990) );
  AND2_X2 U10746 ( .A1(n8990), .A2(n13471), .ZN(n13875) );
  NAND2_X1 U10747 ( .A1(n13875), .A2(n8991), .ZN(n13874) );
  INV_X1 U10748 ( .A(n13855), .ZN(n13850) );
  INV_X1 U10749 ( .A(n13857), .ZN(n13616) );
  OR2_X2 U10750 ( .A1(n13686), .A2(n13616), .ZN(n13480) );
  NAND2_X1 U10751 ( .A1(n13686), .A2(n13616), .ZN(n13478) );
  NAND2_X1 U10752 ( .A1(n13480), .A2(n13478), .ZN(n13841) );
  INV_X1 U10753 ( .A(n13840), .ZN(n8992) );
  NOR2_X1 U10754 ( .A1(n13841), .A2(n8992), .ZN(n8993) );
  OAI21_X2 U10755 ( .B1(n13830), .B2(n8914), .A(n13482), .ZN(n9069) );
  AND2_X1 U10756 ( .A1(n12413), .A2(n12192), .ZN(n9053) );
  INV_X1 U10757 ( .A(n9053), .ZN(n8995) );
  XNOR2_X1 U10758 ( .A(n13544), .B(n8995), .ZN(n8997) );
  NAND2_X1 U10759 ( .A1(n12413), .A2(n13799), .ZN(n8996) );
  NAND2_X1 U10760 ( .A1(n8997), .A2(n8996), .ZN(n10510) );
  NAND2_X1 U10761 ( .A1(n12192), .A2(n13799), .ZN(n9049) );
  INV_X1 U10762 ( .A(n9049), .ZN(n13508) );
  AND2_X1 U10763 ( .A1(n16609), .A2(n13508), .ZN(n8998) );
  NAND2_X1 U10764 ( .A1(n10510), .A2(n8998), .ZN(n8999) );
  NAND2_X1 U10765 ( .A1(n9031), .A2(n9049), .ZN(n9051) );
  AND2_X1 U10766 ( .A1(n13813), .A2(n16614), .ZN(n9001) );
  NOR2_X2 U10767 ( .A1(n13814), .A2(n9001), .ZN(n9061) );
  INV_X1 U10768 ( .A(n9002), .ZN(n9003) );
  NAND2_X1 U10769 ( .A1(n9003), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9004) );
  MUX2_X1 U10770 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9004), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9006) );
  NAND2_X1 U10771 ( .A1(n9006), .A2(n9005), .ZN(n12907) );
  XNOR2_X1 U10772 ( .A(n12907), .B(P3_B_REG_SCAN_IN), .ZN(n9010) );
  NAND2_X1 U10773 ( .A1(n9005), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9007) );
  MUX2_X1 U10774 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9007), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9009) );
  INV_X1 U10775 ( .A(n9008), .ZN(n9011) );
  INV_X1 U10776 ( .A(n9038), .ZN(n13013) );
  NAND2_X1 U10777 ( .A1(n9010), .A2(n13013), .ZN(n9013) );
  NAND2_X1 U10778 ( .A1(n9011), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9012) );
  INV_X1 U10779 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U10780 ( .A1(n11376), .A2(n9014), .ZN(n9016) );
  INV_X1 U10781 ( .A(n9039), .ZN(n13070) );
  NAND2_X1 U10782 ( .A1(n13070), .A2(n13013), .ZN(n9015) );
  INV_X1 U10783 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U10784 ( .A1(n11376), .A2(n9017), .ZN(n9019) );
  NAND2_X1 U10785 ( .A1(n13070), .A2(n12907), .ZN(n9018) );
  NOR2_X1 U10786 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9023) );
  NOR4_X1 U10787 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9022) );
  NOR4_X1 U10788 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9021) );
  NOR4_X1 U10789 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9020) );
  NAND4_X1 U10790 ( .A1(n9023), .A2(n9022), .A3(n9021), .A4(n9020), .ZN(n9029)
         );
  NOR4_X1 U10791 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9027) );
  NOR4_X1 U10792 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9026) );
  NOR4_X1 U10793 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9025) );
  NOR4_X1 U10794 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9024) );
  NAND4_X1 U10795 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(n9028)
         );
  OAI21_X1 U10796 ( .B1(n9029), .B2(n9028), .A(n11376), .ZN(n9046) );
  NAND3_X1 U10797 ( .A1(n12399), .A2(n9045), .A3(n9046), .ZN(n10521) );
  INV_X1 U10798 ( .A(n10510), .ZN(n10524) );
  AND3_X1 U10799 ( .A1(n14211), .A2(n14209), .A3(n9046), .ZN(n10525) );
  OR2_X1 U10800 ( .A1(n13487), .A2(n9049), .ZN(n11893) );
  OR2_X1 U10801 ( .A1(n13541), .A2(n9031), .ZN(n10519) );
  NAND2_X1 U10802 ( .A1(n11893), .A2(n10519), .ZN(n9032) );
  NAND2_X1 U10803 ( .A1(n10525), .A2(n9032), .ZN(n9033) );
  OAI21_X1 U10804 ( .B1(n10521), .B2(n10524), .A(n9033), .ZN(n9040) );
  INV_X1 U10805 ( .A(n12907), .ZN(n9037) );
  INV_X1 U10806 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9041) );
  AOI21_X1 U10807 ( .B1(n8942), .B2(n14163), .A(n9042), .ZN(n9043) );
  OAI21_X1 U10808 ( .B1(n9061), .B2(n9044), .A(n9043), .ZN(P3_U3456) );
  XNOR2_X1 U10809 ( .A(n14209), .B(n9045), .ZN(n9047) );
  NAND2_X1 U10810 ( .A1(n9048), .A2(n13487), .ZN(n12403) );
  NAND2_X1 U10811 ( .A1(n13466), .A2(n9049), .ZN(n12398) );
  NAND2_X1 U10812 ( .A1(n12403), .A2(n12398), .ZN(n9050) );
  NAND2_X1 U10813 ( .A1(n9050), .A2(n14209), .ZN(n9055) );
  NAND2_X1 U10814 ( .A1(n9051), .A2(n12413), .ZN(n9052) );
  OAI211_X1 U10815 ( .C1(n13544), .C2(n9053), .A(n9052), .B(n12399), .ZN(n9054) );
  NAND2_X1 U10816 ( .A1(n8942), .A2(n9056), .ZN(n9058) );
  OAI21_X1 U10817 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(P3_U3488) );
  INV_X1 U10818 ( .A(n9062), .ZN(n9064) );
  INV_X1 U10819 ( .A(n13237), .ZN(n9063) );
  NAND3_X1 U10820 ( .A1(n9066), .A2(n13979), .A3(n9065), .ZN(n9068) );
  AOI22_X1 U10821 ( .A1(n13702), .A2(n13987), .B1(n12512), .B2(n13986), .ZN(
        n9067) );
  OR2_X1 U10822 ( .A1(n9069), .A2(n9063), .ZN(n9070) );
  NAND2_X1 U10823 ( .A1(n9071), .A2(n9070), .ZN(n13825) );
  NAND2_X1 U10824 ( .A1(n13825), .A2(n16614), .ZN(n9072) );
  NAND2_X1 U10825 ( .A1(n13827), .A2(n9072), .ZN(n10423) );
  NAND2_X1 U10826 ( .A1(n13245), .A2(n9056), .ZN(n9074) );
  NAND2_X1 U10827 ( .A1(n9060), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9073) );
  NOR2_X2 U10828 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9087) );
  NOR2_X2 U10829 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9089) );
  NOR2_X2 U10830 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9088) );
  NAND4_X1 U10831 ( .A1(n9087), .A2(n9089), .A3(n9088), .A4(n9086), .ZN(n9078)
         );
  INV_X2 U10832 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n15637) );
  NAND3_X1 U10833 ( .A1(n9077), .A2(n15636), .A3(n15637), .ZN(n9083) );
  NOR2_X1 U10834 ( .A1(n9078), .A2(n9083), .ZN(n9080) );
  NOR2_X4 U10835 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9135) );
  NOR2_X1 U10836 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9079) );
  NAND2_X1 U10837 ( .A1(n9080), .A2(n9243), .ZN(n9485) );
  NAND2_X1 U10838 ( .A1(n9135), .A2(n15631), .ZN(n9171) );
  NOR2_X2 U10839 ( .A1(n9171), .A2(n9083), .ZN(n9093) );
  NOR2_X1 U10840 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9085) );
  NOR2_X1 U10841 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9091) );
  NOR2_X1 U10842 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n9090) );
  NAND4_X2 U10843 ( .A1(n9093), .A2(n7471), .A3(n9486), .A4(n9092), .ZN(n9111)
         );
  NAND2_X1 U10844 ( .A1(n9095), .A2(n9096), .ZN(n15792) );
  XNOR2_X2 U10845 ( .A(n9094), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9103) );
  INV_X1 U10846 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9098) );
  OR2_X1 U10847 ( .A1(n7449), .A2(n9098), .ZN(n9101) );
  INV_X1 U10848 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9099) );
  OR2_X1 U10849 ( .A1(n9249), .A2(n9099), .ZN(n9100) );
  INV_X1 U10850 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9105) );
  OR2_X1 U10851 ( .A1(n7434), .A2(n9105), .ZN(n9106) );
  INV_X1 U10852 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9114) );
  INV_X1 U10853 ( .A(SI_0_), .ZN(n9139) );
  NOR2_X1 U10854 ( .A1(n11209), .A2(n9139), .ZN(n9107) );
  XNOR2_X1 U10855 ( .A(n9107), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15812) );
  XNOR2_X2 U10856 ( .A(n9110), .B(n9109), .ZN(n9908) );
  NAND2_X2 U10857 ( .A1(n9908), .A2(n14954), .ZN(n9147) );
  MUX2_X1 U10858 ( .A(n9114), .B(n15812), .S(n9590), .Z(n16310) );
  AND2_X1 U10859 ( .A1(n14943), .A2(n16310), .ZN(n9857) );
  AOI21_X1 U10860 ( .B1(n10958), .B2(n10539), .A(n9857), .ZN(n9128) );
  NAND2_X1 U10861 ( .A1(n9117), .A2(n9888), .ZN(n9124) );
  NAND3_X1 U10862 ( .A1(n9118), .A2(P1_IR_REG_22__SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9123) );
  INV_X1 U10863 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U10864 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9119) );
  NAND2_X1 U10865 ( .A1(n9119), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9120) );
  OAI21_X1 U10866 ( .B1(n9121), .B2(P1_IR_REG_31__SCAN_IN), .A(n9120), .ZN(
        n9122) );
  NAND2_X1 U10867 ( .A1(n9824), .A2(n9874), .ZN(n10580) );
  NAND2_X1 U10868 ( .A1(n9128), .A2(n9260), .ZN(n9153) );
  INV_X1 U10869 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9129) );
  OR2_X1 U10870 ( .A1(n9754), .A2(n9129), .ZN(n9133) );
  INV_X1 U10871 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9130) );
  OR2_X1 U10872 ( .A1(n9191), .A2(n9130), .ZN(n9132) );
  INV_X1 U10873 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U10874 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9134) );
  MUX2_X1 U10875 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9134), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9136) );
  INV_X1 U10876 ( .A(n9135), .ZN(n9169) );
  NAND2_X1 U10877 ( .A1(n9136), .A2(n9169), .ZN(n11190) );
  INV_X1 U10878 ( .A(n11190), .ZN(n14949) );
  NAND2_X1 U10879 ( .A1(n7441), .A2(n14949), .ZN(n9150) );
  NAND2_X1 U10880 ( .A1(n9138), .A2(SI_1_), .ZN(n9157) );
  INV_X1 U10881 ( .A(n9144), .ZN(n9143) );
  NAND2_X1 U10882 ( .A1(n9143), .A2(n9156), .ZN(n9146) );
  NAND2_X1 U10883 ( .A1(n9144), .A2(n9142), .ZN(n9145) );
  AND2_X1 U10884 ( .A1(n9146), .A2(n9145), .ZN(n11189) );
  NAND2_X1 U10885 ( .A1(n7440), .A2(n11189), .ZN(n9149) );
  NAND2_X1 U10886 ( .A1(n7445), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U10887 ( .A1(n10603), .A2(n16314), .ZN(n9856) );
  NAND2_X1 U10888 ( .A1(n16315), .A2(n9856), .ZN(n9151) );
  NAND2_X1 U10889 ( .A1(n7415), .A2(n9151), .ZN(n9152) );
  NAND2_X1 U10890 ( .A1(n9153), .A2(n9152), .ZN(n9183) );
  INV_X2 U10891 ( .A(n10603), .ZN(n11602) );
  NAND2_X2 U10892 ( .A1(n11602), .A2(n9154), .ZN(n10538) );
  INV_X1 U10893 ( .A(n10538), .ZN(n9182) );
  MUX2_X1 U10894 ( .A(n9856), .B(n10538), .S(n7415), .Z(n9181) );
  NAND2_X1 U10895 ( .A1(n9156), .A2(n9155), .ZN(n9160) );
  NAND3_X1 U10896 ( .A1(n9160), .A2(n15308), .A3(n9157), .ZN(n9162) );
  INV_X1 U10897 ( .A(n9157), .ZN(n9158) );
  NAND2_X1 U10898 ( .A1(n9158), .A2(SI_2_), .ZN(n9159) );
  MUX2_X1 U10899 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9141), .Z(n9164) );
  INV_X1 U10900 ( .A(n9164), .ZN(n9165) );
  NAND2_X1 U10901 ( .A1(n9166), .A2(n9165), .ZN(n9167) );
  NAND2_X1 U10902 ( .A1(n9184), .A2(n9167), .ZN(n11216) );
  INV_X1 U10903 ( .A(n11216), .ZN(n9168) );
  NAND2_X1 U10904 ( .A1(n9169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9170) );
  MUX2_X1 U10905 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9170), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9172) );
  NAND2_X1 U10906 ( .A1(n9172), .A2(n9171), .ZN(n11185) );
  INV_X1 U10907 ( .A(n11185), .ZN(n14965) );
  AOI22_X1 U10908 ( .A1(n7445), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n7443), .B2(
        n14965), .ZN(n9173) );
  INV_X2 U10909 ( .A(n16358), .ZN(n16348) );
  INV_X1 U10910 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9175) );
  OR2_X1 U10911 ( .A1(n9191), .A2(n9175), .ZN(n9179) );
  INV_X1 U10912 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11152) );
  OR2_X1 U10913 ( .A1(n7439), .A2(n11152), .ZN(n9178) );
  NAND2_X1 U10914 ( .A1(n7447), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9177) );
  INV_X1 U10915 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14962) );
  NAND4_X1 U10916 ( .A1(n9179), .A2(n9178), .A3(n9177), .A4(n9176), .ZN(n14942) );
  NAND2_X1 U10917 ( .A1(n16348), .A2(n14942), .ZN(n9855) );
  INV_X2 U10918 ( .A(n14942), .ZN(n9196) );
  MUX2_X1 U10919 ( .A(n9855), .B(n10541), .S(n7415), .Z(n9180) );
  OAI211_X1 U10920 ( .C1(n9183), .C2(n9182), .A(n9181), .B(n9180), .ZN(n9199)
         );
  NAND2_X1 U10921 ( .A1(n9185), .A2(SI_3_), .ZN(n9226) );
  OAI21_X1 U10922 ( .B1(n9185), .B2(SI_3_), .A(n9226), .ZN(n9205) );
  XNOR2_X1 U10923 ( .A(n9232), .B(n9205), .ZN(n11187) );
  NAND2_X1 U10924 ( .A1(n11187), .A2(n9820), .ZN(n9189) );
  NAND2_X1 U10925 ( .A1(n9171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9187) );
  XNOR2_X1 U10926 ( .A(n9187), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14979) );
  AOI22_X1 U10927 ( .A1(n9186), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n7443), .B2(
        n14979), .ZN(n9188) );
  NAND2_X1 U10928 ( .A1(n9189), .A2(n9188), .ZN(n16365) );
  INV_X1 U10929 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U10930 ( .A1(n9318), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9194) );
  OR2_X1 U10931 ( .A1(n7434), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9193) );
  INV_X1 U10932 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11129) );
  OR2_X1 U10933 ( .A1(n9249), .A2(n11129), .ZN(n9192) );
  NAND2_X1 U10934 ( .A1(n16365), .A2(n11846), .ZN(n10543) );
  OAI21_X1 U10935 ( .B1(n9196), .B2(n16348), .A(n9197), .ZN(n9198) );
  OR2_X1 U10936 ( .A1(n16365), .A2(n11846), .ZN(n9200) );
  NAND4_X1 U10937 ( .A1(n9199), .A2(n10543), .A3(n9198), .A4(n9200), .ZN(n9204) );
  INV_X1 U10938 ( .A(n9200), .ZN(n9202) );
  NAND2_X1 U10939 ( .A1(n7415), .A2(n10543), .ZN(n9201) );
  OAI21_X1 U10940 ( .B1(n7415), .B2(n9202), .A(n9201), .ZN(n9203) );
  NAND2_X1 U10941 ( .A1(n9204), .A2(n9203), .ZN(n9222) );
  INV_X1 U10942 ( .A(n9205), .ZN(n9233) );
  NAND2_X1 U10943 ( .A1(n9227), .A2(n9226), .ZN(n9211) );
  NAND2_X1 U10944 ( .A1(n9208), .A2(SI_4_), .ZN(n9225) );
  NAND2_X1 U10945 ( .A1(n9211), .A2(n9210), .ZN(n9213) );
  OR2_X1 U10946 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  XNOR2_X1 U10947 ( .A(n9214), .B(P1_IR_REG_4__SCAN_IN), .ZN(n16284) );
  AOI22_X1 U10948 ( .A1(n9186), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7442), .B2(
        n16284), .ZN(n9215) );
  NAND2_X1 U10949 ( .A1(n9318), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9219) );
  INV_X1 U10950 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11156) );
  OR2_X1 U10951 ( .A1(n7438), .A2(n11156), .ZN(n9218) );
  AND2_X1 U10952 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9251) );
  INV_X1 U10953 ( .A(n9251), .ZN(n9253) );
  OAI21_X1 U10954 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9253), .ZN(n11844) );
  OR2_X1 U10955 ( .A1(n9689), .A2(n11844), .ZN(n9217) );
  INV_X1 U10956 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11132) );
  OR2_X1 U10957 ( .A1(n9805), .A2(n11132), .ZN(n9216) );
  MUX2_X1 U10958 ( .A(n9860), .B(n11996), .S(n7415), .Z(n9221) );
  MUX2_X1 U10959 ( .A(n16390), .B(n14940), .S(n9260), .Z(n9220) );
  OAI21_X1 U10960 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(n9224) );
  NAND2_X1 U10961 ( .A1(n9222), .A2(n9221), .ZN(n9223) );
  NAND2_X1 U10962 ( .A1(n9224), .A2(n9223), .ZN(n9263) );
  AND2_X1 U10963 ( .A1(n9226), .A2(n9225), .ZN(n9236) );
  MUX2_X1 U10964 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9141), .Z(n9228) );
  NAND2_X1 U10965 ( .A1(n9228), .A2(SI_5_), .ZN(n9269) );
  OAI21_X1 U10966 ( .B1(n9228), .B2(SI_5_), .A(n9269), .ZN(n9229) );
  INV_X1 U10967 ( .A(n9229), .ZN(n9240) );
  AND2_X1 U10968 ( .A1(n9240), .A2(n9235), .ZN(n9230) );
  AND2_X1 U10969 ( .A1(n9233), .A2(n9235), .ZN(n9234) );
  NAND2_X1 U10970 ( .A1(n9232), .A2(n9234), .ZN(n9239) );
  INV_X1 U10971 ( .A(n9235), .ZN(n9237) );
  OR2_X1 U10972 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  NAND2_X1 U10973 ( .A1(n9239), .A2(n9238), .ZN(n9241) );
  OR2_X1 U10974 ( .A1(n9241), .A2(n9240), .ZN(n9242) );
  OR2_X1 U10975 ( .A1(n11210), .A2(n9796), .ZN(n9247) );
  INV_X1 U10976 ( .A(n9243), .ZN(n9244) );
  NAND2_X1 U10977 ( .A1(n9244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9245) );
  XNOR2_X1 U10978 ( .A(n9245), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U10979 ( .A1(n9186), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7443), .B2(
        n14994), .ZN(n9246) );
  NAND2_X1 U10980 ( .A1(n9247), .A2(n9246), .ZN(n12003) );
  NAND2_X1 U10981 ( .A1(n9248), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9259) );
  INV_X1 U10982 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9250) );
  OR2_X1 U10983 ( .A1(n9805), .A2(n9250), .ZN(n9258) );
  NAND2_X1 U10984 ( .A1(n9251), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9280) );
  INV_X1 U10985 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U10986 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  NAND2_X1 U10987 ( .A1(n9280), .A2(n9254), .ZN(n12007) );
  OR2_X1 U10988 ( .A1(n7433), .A2(n12007), .ZN(n9257) );
  INV_X1 U10989 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9255) );
  OR2_X1 U10990 ( .A1(n7449), .A2(n9255), .ZN(n9256) );
  NAND4_X1 U10991 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n14939) );
  MUX2_X1 U10992 ( .A(n12003), .B(n14939), .S(n9260), .Z(n9264) );
  NAND2_X1 U10993 ( .A1(n9263), .A2(n9264), .ZN(n9262) );
  MUX2_X1 U10994 ( .A(n14939), .B(n12003), .S(n9260), .Z(n9261) );
  NAND2_X1 U10995 ( .A1(n9262), .A2(n9261), .ZN(n9268) );
  INV_X1 U10996 ( .A(n9263), .ZN(n9266) );
  INV_X1 U10997 ( .A(n9264), .ZN(n9265) );
  NAND2_X1 U10998 ( .A1(n9266), .A2(n9265), .ZN(n9267) );
  MUX2_X1 U10999 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11209), .Z(n9270) );
  NAND2_X1 U11000 ( .A1(n9270), .A2(SI_6_), .ZN(n9298) );
  OAI21_X1 U11001 ( .B1(SI_6_), .B2(n9270), .A(n9298), .ZN(n9271) );
  INV_X1 U11002 ( .A(n9271), .ZN(n9272) );
  NAND2_X1 U11003 ( .A1(n9273), .A2(n9272), .ZN(n9299) );
  OR2_X1 U11004 ( .A1(n9273), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U11005 ( .A1(n9299), .A2(n9274), .ZN(n11253) );
  OR2_X1 U11006 ( .A1(n11253), .A2(n9796), .ZN(n9278) );
  AND2_X1 U11007 ( .A1(n9243), .A2(n15637), .ZN(n9306) );
  INV_X1 U11008 ( .A(n9306), .ZN(n9275) );
  NAND2_X1 U11009 ( .A1(n9275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9276) );
  XNOR2_X1 U11010 ( .A(n9276), .B(P1_IR_REG_6__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U11011 ( .A1(n9186), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7442), .B2(
        n15006), .ZN(n9277) );
  NAND2_X1 U11012 ( .A1(n9278), .A2(n9277), .ZN(n12189) );
  NAND2_X1 U11013 ( .A1(n7447), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9286) );
  INV_X1 U11014 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11161) );
  OR2_X1 U11015 ( .A1(n7439), .A2(n11161), .ZN(n9285) );
  INV_X1 U11016 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9279) );
  NOR2_X1 U11017 ( .A1(n9280), .A2(n9279), .ZN(n9289) );
  INV_X1 U11018 ( .A(n9289), .ZN(n9291) );
  NAND2_X1 U11019 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  NAND2_X1 U11020 ( .A1(n9291), .A2(n9281), .ZN(n12184) );
  OR2_X1 U11021 ( .A1(n9689), .A2(n12184), .ZN(n9284) );
  INV_X1 U11022 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9282) );
  OR2_X1 U11023 ( .A1(n7450), .A2(n9282), .ZN(n9283) );
  NAND4_X1 U11024 ( .A1(n9286), .A2(n9285), .A3(n9284), .A4(n9283), .ZN(n14938) );
  MUX2_X1 U11025 ( .A(n12189), .B(n14938), .S(n7415), .Z(n9288) );
  NAND2_X1 U11026 ( .A1(n7447), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9297) );
  INV_X1 U11027 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11164) );
  OR2_X1 U11028 ( .A1(n7439), .A2(n11164), .ZN(n9296) );
  NAND2_X1 U11029 ( .A1(n9289), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9319) );
  INV_X1 U11030 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11031 ( .A1(n9291), .A2(n9290), .ZN(n9292) );
  NAND2_X1 U11032 ( .A1(n9319), .A2(n9292), .ZN(n12234) );
  OR2_X1 U11033 ( .A1(n7434), .A2(n12234), .ZN(n9295) );
  INV_X1 U11034 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9293) );
  OR2_X1 U11035 ( .A1(n7450), .A2(n9293), .ZN(n9294) );
  NAND4_X1 U11036 ( .A1(n9297), .A2(n9296), .A3(n9295), .A4(n9294), .ZN(n14937) );
  NAND2_X1 U11037 ( .A1(n9299), .A2(n9298), .ZN(n9304) );
  MUX2_X1 U11038 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11209), .Z(n9300) );
  NAND2_X1 U11039 ( .A1(n9300), .A2(SI_7_), .ZN(n9325) );
  INV_X1 U11040 ( .A(n9300), .ZN(n9301) );
  INV_X1 U11041 ( .A(SI_7_), .ZN(n15306) );
  NAND2_X1 U11042 ( .A1(n9301), .A2(n15306), .ZN(n9302) );
  AND2_X1 U11043 ( .A1(n9325), .A2(n9302), .ZN(n9303) );
  NAND2_X1 U11044 ( .A1(n9304), .A2(n9303), .ZN(n9326) );
  OR2_X1 U11045 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  NAND2_X1 U11046 ( .A1(n9326), .A2(n9305), .ZN(n11212) );
  OR2_X1 U11047 ( .A1(n11212), .A2(n9796), .ZN(n9309) );
  NAND2_X1 U11048 ( .A1(n9306), .A2(n15636), .ZN(n9488) );
  NAND2_X1 U11049 ( .A1(n9488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9307) );
  XNOR2_X1 U11050 ( .A(n9307), .B(P1_IR_REG_7__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U11051 ( .A1(n9186), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7443), .B2(
        n15021), .ZN(n9308) );
  NAND2_X1 U11052 ( .A1(n9309), .A2(n9308), .ZN(n12236) );
  MUX2_X1 U11053 ( .A(n14937), .B(n12236), .S(n7415), .Z(n9313) );
  NAND2_X1 U11054 ( .A1(n9312), .A2(n9313), .ZN(n9311) );
  MUX2_X1 U11055 ( .A(n12236), .B(n14937), .S(n7415), .Z(n9310) );
  NAND2_X1 U11056 ( .A1(n9311), .A2(n9310), .ZN(n9317) );
  INV_X1 U11057 ( .A(n9312), .ZN(n9315) );
  INV_X1 U11058 ( .A(n9313), .ZN(n9314) );
  NAND2_X1 U11059 ( .A1(n9315), .A2(n9314), .ZN(n9316) );
  NAND2_X1 U11060 ( .A1(n9317), .A2(n9316), .ZN(n9336) );
  NAND2_X1 U11061 ( .A1(n9318), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9324) );
  INV_X1 U11062 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11141) );
  OR2_X1 U11063 ( .A1(n9805), .A2(n11141), .ZN(n9323) );
  INV_X1 U11064 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11167) );
  OR2_X1 U11065 ( .A1(n7438), .A2(n11167), .ZN(n9322) );
  NAND2_X1 U11066 ( .A1(n9319), .A2(n12568), .ZN(n9320) );
  NAND2_X1 U11067 ( .A1(n9340), .A2(n9320), .ZN(n12569) );
  OR2_X1 U11068 ( .A1(n9689), .A2(n12569), .ZN(n9321) );
  NAND4_X1 U11069 ( .A1(n9324), .A2(n9323), .A3(n9322), .A4(n9321), .ZN(n14936) );
  MUX2_X1 U11070 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11209), .Z(n9327) );
  NAND2_X1 U11071 ( .A1(n9327), .A2(SI_8_), .ZN(n9346) );
  OAI21_X1 U11072 ( .B1(SI_8_), .B2(n9327), .A(n9346), .ZN(n9328) );
  INV_X1 U11073 ( .A(n9328), .ZN(n9329) );
  NAND2_X1 U11074 ( .A1(n9330), .A2(n9329), .ZN(n9347) );
  OR2_X1 U11075 ( .A1(n9330), .A2(n9329), .ZN(n9331) );
  NAND2_X1 U11076 ( .A1(n9347), .A2(n9331), .ZN(n11248) );
  OR2_X1 U11077 ( .A1(n11248), .A2(n9796), .ZN(n9334) );
  NAND2_X1 U11078 ( .A1(n9352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9332) );
  XNOR2_X1 U11079 ( .A(n9332), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U11080 ( .A1(n7442), .A2(n11260), .B1(n9186), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11081 ( .A1(n9334), .A2(n9333), .ZN(n12573) );
  MUX2_X1 U11082 ( .A(n14936), .B(n12573), .S(n9260), .Z(n9337) );
  MUX2_X1 U11083 ( .A(n14936), .B(n12573), .S(n7415), .Z(n9335) );
  INV_X1 U11084 ( .A(n9337), .ZN(n9338) );
  NAND2_X1 U11085 ( .A1(n9318), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9345) );
  OR2_X1 U11086 ( .A1(n9805), .A2(n12316), .ZN(n9344) );
  INV_X1 U11087 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12199) );
  OR2_X1 U11088 ( .A1(n7438), .A2(n12199), .ZN(n9343) );
  NOR2_X1 U11089 ( .A1(n9340), .A2(n9339), .ZN(n9359) );
  INV_X1 U11090 ( .A(n9359), .ZN(n9361) );
  NAND2_X1 U11091 ( .A1(n9340), .A2(n9339), .ZN(n9341) );
  NAND2_X1 U11092 ( .A1(n9361), .A2(n9341), .ZN(n12886) );
  OR2_X1 U11093 ( .A1(n7433), .A2(n12886), .ZN(n9342) );
  NAND4_X1 U11094 ( .A1(n9345), .A2(n9344), .A3(n9343), .A4(n9342), .ZN(n14935) );
  NAND2_X1 U11095 ( .A1(n9347), .A2(n9346), .ZN(n9351) );
  MUX2_X1 U11096 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11209), .Z(n9348) );
  NAND2_X1 U11097 ( .A1(n9348), .A2(SI_9_), .ZN(n9368) );
  OAI21_X1 U11098 ( .B1(n9348), .B2(SI_9_), .A(n9368), .ZN(n9349) );
  INV_X1 U11099 ( .A(n9349), .ZN(n9350) );
  OR2_X1 U11100 ( .A1(n11251), .A2(n9796), .ZN(n9355) );
  NAND2_X1 U11101 ( .A1(n9374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  XNOR2_X1 U11102 ( .A(n9353), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U11103 ( .A1(n11275), .A2(n7443), .B1(n9186), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9354) );
  NAND2_X2 U11104 ( .A1(n9355), .A2(n9354), .ZN(n12891) );
  MUX2_X1 U11105 ( .A(n14935), .B(n12891), .S(n7415), .Z(n9357) );
  MUX2_X1 U11106 ( .A(n14935), .B(n12891), .S(n9260), .Z(n9356) );
  INV_X1 U11107 ( .A(n9357), .ZN(n9358) );
  NAND2_X1 U11108 ( .A1(n7447), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9367) );
  INV_X1 U11109 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12362) );
  OR2_X1 U11110 ( .A1(n7439), .A2(n12362), .ZN(n9366) );
  INV_X1 U11111 ( .A(n9390), .ZN(n9392) );
  INV_X1 U11112 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11113 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  NAND2_X1 U11114 ( .A1(n9392), .A2(n9362), .ZN(n12923) );
  OR2_X1 U11115 ( .A1(n9689), .A2(n12923), .ZN(n9365) );
  INV_X1 U11116 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9363) );
  OR2_X1 U11117 ( .A1(n7450), .A2(n9363), .ZN(n9364) );
  NAND4_X1 U11118 ( .A1(n9367), .A2(n9366), .A3(n9365), .A4(n9364), .ZN(n14934) );
  MUX2_X1 U11119 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11209), .Z(n9370) );
  NAND2_X1 U11120 ( .A1(n9370), .A2(SI_10_), .ZN(n9398) );
  OAI21_X1 U11121 ( .B1(n9370), .B2(SI_10_), .A(n9398), .ZN(n9371) );
  INV_X1 U11122 ( .A(n9371), .ZN(n9372) );
  OR2_X1 U11123 ( .A1(n11287), .A2(n9796), .ZN(n9379) );
  INV_X1 U11124 ( .A(n9374), .ZN(n9376) );
  INV_X1 U11125 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U11126 ( .A1(n9376), .A2(n9375), .ZN(n9400) );
  NAND2_X1 U11127 ( .A1(n9400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9377) );
  XNOR2_X1 U11128 ( .A(n9377), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U11129 ( .A1(n11353), .A2(n7442), .B1(n9186), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9378) );
  MUX2_X1 U11130 ( .A(n14934), .B(n12928), .S(n9260), .Z(n9383) );
  NAND2_X1 U11131 ( .A1(n9382), .A2(n9383), .ZN(n9381) );
  MUX2_X1 U11132 ( .A(n14934), .B(n12928), .S(n7415), .Z(n9380) );
  NAND2_X1 U11133 ( .A1(n9381), .A2(n9380), .ZN(n9387) );
  INV_X1 U11134 ( .A(n9382), .ZN(n9385) );
  INV_X1 U11135 ( .A(n9383), .ZN(n9384) );
  NAND2_X1 U11136 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U11137 ( .A1(n9318), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9397) );
  INV_X1 U11138 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9388) );
  OR2_X1 U11139 ( .A1(n9805), .A2(n9388), .ZN(n9396) );
  INV_X1 U11140 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9389) );
  OR2_X1 U11141 ( .A1(n7438), .A2(n9389), .ZN(n9395) );
  NAND2_X1 U11142 ( .A1(n9390), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9410) );
  INV_X1 U11143 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U11144 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  NAND2_X1 U11145 ( .A1(n9410), .A2(n9393), .ZN(n13044) );
  OR2_X1 U11146 ( .A1(n7434), .A2(n13044), .ZN(n9394) );
  MUX2_X1 U11147 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11209), .Z(n9416) );
  XNOR2_X1 U11148 ( .A(n9416), .B(SI_11_), .ZN(n9419) );
  NAND2_X1 U11149 ( .A1(n11344), .A2(n9820), .ZN(n9404) );
  INV_X1 U11150 ( .A(n9400), .ZN(n9401) );
  INV_X1 U11151 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15438) );
  NAND2_X1 U11152 ( .A1(n9401), .A2(n15438), .ZN(n9402) );
  NAND2_X1 U11153 ( .A1(n9402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9421) );
  XNOR2_X1 U11154 ( .A(n9421), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U11155 ( .A1(n11450), .A2(n7443), .B1(n9186), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9403) );
  MUX2_X1 U11156 ( .A(n14933), .B(n12614), .S(n7415), .Z(n9406) );
  MUX2_X1 U11157 ( .A(n14933), .B(n12614), .S(n9260), .Z(n9405) );
  INV_X1 U11158 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U11159 ( .A1(n9318), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9415) );
  INV_X1 U11160 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9408) );
  OR2_X1 U11161 ( .A1(n9805), .A2(n9408), .ZN(n9414) );
  INV_X1 U11162 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12546) );
  OR2_X1 U11163 ( .A1(n7439), .A2(n12546), .ZN(n9413) );
  NAND2_X1 U11164 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U11165 ( .A1(n9429), .A2(n9411), .ZN(n12543) );
  OR2_X1 U11166 ( .A1(n9689), .A2(n12543), .ZN(n9412) );
  NAND4_X1 U11167 ( .A1(n9415), .A2(n9414), .A3(n9413), .A4(n9412), .ZN(n14932) );
  INV_X1 U11168 ( .A(n9416), .ZN(n9417) );
  NAND2_X1 U11169 ( .A1(n9417), .A2(n15493), .ZN(n9418) );
  MUX2_X1 U11170 ( .A(n11438), .B(n11440), .S(n11209), .Z(n9437) );
  XNOR2_X1 U11171 ( .A(n9437), .B(SI_12_), .ZN(n9435) );
  XNOR2_X1 U11172 ( .A(n9436), .B(n9435), .ZN(n11436) );
  NAND2_X1 U11173 ( .A1(n11436), .A2(n9820), .ZN(n9424) );
  NAND2_X1 U11174 ( .A1(n9421), .A2(n15437), .ZN(n9422) );
  NAND2_X1 U11175 ( .A1(n9422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9447) );
  XNOR2_X1 U11176 ( .A(n9447), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U11177 ( .A1(n11558), .A2(n7443), .B1(n9186), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9423) );
  MUX2_X1 U11178 ( .A(n14932), .B(n12813), .S(n9260), .Z(n9427) );
  MUX2_X1 U11179 ( .A(n14932), .B(n12813), .S(n7415), .Z(n9425) );
  INV_X1 U11180 ( .A(n9454), .ZN(n9456) );
  NAND2_X1 U11181 ( .A1(n9429), .A2(n9428), .ZN(n9430) );
  NAND2_X1 U11182 ( .A1(n9456), .A2(n9430), .ZN(n13171) );
  NAND2_X1 U11183 ( .A1(n9318), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9431) );
  OAI21_X1 U11184 ( .B1(n13171), .B2(n9689), .A(n9431), .ZN(n9434) );
  INV_X1 U11185 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U11186 ( .A1(n9248), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9432) );
  OAI21_X1 U11187 ( .B1(n11561), .B2(n9805), .A(n9432), .ZN(n9433) );
  NAND2_X1 U11188 ( .A1(n9437), .A2(n15487), .ZN(n9438) );
  MUX2_X1 U11189 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n11209), .Z(n9440) );
  NAND2_X1 U11190 ( .A1(n9440), .A2(SI_13_), .ZN(n9461) );
  INV_X1 U11191 ( .A(n9440), .ZN(n9441) );
  NAND2_X1 U11192 ( .A1(n9441), .A2(n15488), .ZN(n9442) );
  NAND2_X1 U11193 ( .A1(n9461), .A2(n9442), .ZN(n9444) );
  NAND2_X1 U11194 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  NAND2_X1 U11195 ( .A1(n9462), .A2(n9446), .ZN(n11445) );
  NAND2_X1 U11196 ( .A1(n9447), .A2(n15651), .ZN(n9448) );
  NAND2_X1 U11197 ( .A1(n9448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U11198 ( .A(n9463), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11627) );
  NOR2_X1 U11199 ( .A1(n7446), .A2(n11444), .ZN(n9449) );
  AOI21_X1 U11200 ( .B1(n11627), .B2(n7443), .A(n9449), .ZN(n9450) );
  MUX2_X1 U11201 ( .A(n14931), .B(n13176), .S(n7415), .Z(n9452) );
  MUX2_X1 U11202 ( .A(n14931), .B(n13176), .S(n9260), .Z(n9451) );
  INV_X1 U11203 ( .A(n9452), .ZN(n9453) );
  INV_X1 U11204 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U11205 ( .A1(n9454), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9476) );
  INV_X1 U11206 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U11207 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  NAND2_X1 U11208 ( .A1(n9476), .A2(n9457), .ZN(n16557) );
  OR2_X1 U11209 ( .A1(n16557), .A2(n7434), .ZN(n9459) );
  AOI22_X1 U11210 ( .A1(n7447), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9248), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n9458) );
  OAI211_X1 U11211 ( .C1(n7450), .C2(n9460), .A(n9459), .B(n9458), .ZN(n14930)
         );
  MUX2_X1 U11212 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n11209), .Z(n9481) );
  XNOR2_X1 U11213 ( .A(n9481), .B(SI_14_), .ZN(n9483) );
  XNOR2_X1 U11214 ( .A(n9484), .B(n9483), .ZN(n11544) );
  NAND2_X1 U11215 ( .A1(n11544), .A2(n9820), .ZN(n9467) );
  INV_X1 U11216 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n15652) );
  NAND2_X1 U11217 ( .A1(n9463), .A2(n15652), .ZN(n9464) );
  NAND2_X1 U11218 ( .A1(n9464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9465) );
  XNOR2_X1 U11219 ( .A(n9465), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U11220 ( .A1(n11904), .A2(n7442), .B1(n7444), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U11221 ( .A(n14930), .B(n16561), .S(n9260), .Z(n9471) );
  NAND2_X1 U11222 ( .A1(n9470), .A2(n9471), .ZN(n9469) );
  MUX2_X1 U11223 ( .A(n14930), .B(n16561), .S(n7415), .Z(n9468) );
  NAND2_X1 U11224 ( .A1(n9469), .A2(n9468), .ZN(n9475) );
  INV_X1 U11225 ( .A(n9470), .ZN(n9473) );
  INV_X1 U11226 ( .A(n9471), .ZN(n9472) );
  NAND2_X1 U11227 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  INV_X1 U11228 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U11229 ( .A1(n9476), .A2(n14911), .ZN(n9477) );
  NAND2_X1 U11230 ( .A1(n9496), .A2(n9477), .ZN(n16652) );
  OR2_X1 U11231 ( .A1(n16652), .A2(n9689), .ZN(n9479) );
  AOI22_X1 U11232 ( .A1(n7447), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9248), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n9478) );
  OAI211_X1 U11233 ( .C1(n7450), .C2(n9480), .A(n9479), .B(n9478), .ZN(n14929)
         );
  INV_X1 U11234 ( .A(n9481), .ZN(n9482) );
  MUX2_X1 U11235 ( .A(n11717), .B(n11719), .S(n11209), .Z(n9502) );
  XNOR2_X1 U11236 ( .A(n9502), .B(SI_15_), .ZN(n9500) );
  XNOR2_X1 U11237 ( .A(n9501), .B(n9500), .ZN(n11716) );
  NAND2_X1 U11238 ( .A1(n11716), .A2(n9820), .ZN(n9492) );
  INV_X1 U11239 ( .A(n9486), .ZN(n9487) );
  OAI21_X1 U11240 ( .B1(n9488), .B2(n9487), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9489) );
  MUX2_X1 U11241 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9489), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9490) );
  AND2_X1 U11242 ( .A1(n9485), .A2(n9490), .ZN(n12758) );
  AOI22_X1 U11243 ( .A1(n12758), .A2(n7442), .B1(n7444), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n9491) );
  MUX2_X1 U11244 ( .A(n14929), .B(n11055), .S(n7415), .Z(n9494) );
  MUX2_X1 U11245 ( .A(n14929), .B(n11055), .S(n9260), .Z(n9493) );
  NAND2_X1 U11246 ( .A1(n9496), .A2(n9495), .ZN(n9497) );
  NAND2_X1 U11247 ( .A1(n9511), .A2(n9497), .ZN(n14852) );
  AOI22_X1 U11248 ( .A1(n7447), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9248), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U11249 ( .A1(n9318), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9498) );
  OAI211_X1 U11250 ( .C1(n14852), .C2(n7433), .A(n9499), .B(n9498), .ZN(n14928) );
  NAND2_X1 U11251 ( .A1(n9502), .A2(n11442), .ZN(n9503) );
  NAND2_X1 U11252 ( .A1(n9504), .A2(n9503), .ZN(n9519) );
  MUX2_X1 U11253 ( .A(n11900), .B(n11902), .S(n11209), .Z(n9520) );
  XNOR2_X1 U11254 ( .A(n9520), .B(SI_16_), .ZN(n9518) );
  XNOR2_X1 U11255 ( .A(n9519), .B(n9518), .ZN(n11899) );
  NAND2_X1 U11256 ( .A1(n11899), .A2(n9820), .ZN(n9507) );
  NAND2_X1 U11257 ( .A1(n9485), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9505) );
  XNOR2_X1 U11258 ( .A(n9505), .B(P1_IR_REG_16__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U11259 ( .A1(n7444), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7443), 
        .B2(n15037), .ZN(n9506) );
  MUX2_X1 U11260 ( .A(n14928), .B(n15762), .S(n9260), .Z(n9509) );
  MUX2_X1 U11261 ( .A(n14928), .B(n15762), .S(n7415), .Z(n9508) );
  INV_X1 U11262 ( .A(n9531), .ZN(n9533) );
  NAND2_X1 U11263 ( .A1(n9511), .A2(n9510), .ZN(n9512) );
  NAND2_X1 U11264 ( .A1(n9533), .A2(n9512), .ZN(n14861) );
  OR2_X1 U11265 ( .A1(n14861), .A2(n9689), .ZN(n9517) );
  INV_X1 U11266 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U11267 ( .A1(n9318), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9514) );
  INV_X1 U11268 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12755) );
  OR2_X1 U11269 ( .A1(n7438), .A2(n12755), .ZN(n9513) );
  OAI211_X1 U11270 ( .C1(n9805), .C2(n12753), .A(n9514), .B(n9513), .ZN(n9515)
         );
  INV_X1 U11271 ( .A(n9515), .ZN(n9516) );
  NAND2_X1 U11272 ( .A1(n9517), .A2(n9516), .ZN(n15232) );
  NAND2_X1 U11273 ( .A1(n9520), .A2(n15479), .ZN(n9521) );
  MUX2_X1 U11274 ( .A(n12064), .B(n12066), .S(n11209), .Z(n9543) );
  XNOR2_X1 U11275 ( .A(n9543), .B(SI_17_), .ZN(n9541) );
  XNOR2_X1 U11276 ( .A(n9542), .B(n9541), .ZN(n12063) );
  NAND2_X1 U11277 ( .A1(n12063), .A2(n9820), .ZN(n9527) );
  INV_X1 U11278 ( .A(n9522), .ZN(n9523) );
  NAND2_X1 U11279 ( .A1(n9523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9524) );
  XNOR2_X1 U11280 ( .A(n9524), .B(n9081), .ZN(n15044) );
  OAI22_X1 U11281 ( .A1(n7446), .A2(n12064), .B1(n15044), .B2(n9590), .ZN(
        n9525) );
  INV_X1 U11282 ( .A(n9525), .ZN(n9526) );
  MUX2_X1 U11283 ( .A(n15232), .B(n15757), .S(n7415), .Z(n9530) );
  MUX2_X1 U11284 ( .A(n15232), .B(n15757), .S(n9260), .Z(n9528) );
  NAND2_X1 U11285 ( .A1(n9531), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9561) );
  INV_X1 U11286 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U11287 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NAND2_X1 U11288 ( .A1(n9561), .A2(n9534), .ZN(n15240) );
  OR2_X1 U11289 ( .A1(n15240), .A2(n7434), .ZN(n9540) );
  INV_X1 U11290 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U11291 ( .A1(n9318), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9536) );
  INV_X1 U11292 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15241) );
  OR2_X1 U11293 ( .A1(n7439), .A2(n15241), .ZN(n9535) );
  OAI211_X1 U11294 ( .C1(n9805), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9538)
         );
  INV_X1 U11295 ( .A(n9538), .ZN(n9539) );
  NAND2_X1 U11296 ( .A1(n9540), .A2(n9539), .ZN(n14927) );
  MUX2_X1 U11297 ( .A(n12340), .B(n12338), .S(n11209), .Z(n9546) );
  NAND2_X1 U11298 ( .A1(n9545), .A2(n9546), .ZN(n9547) );
  NAND2_X1 U11299 ( .A1(n9570), .A2(n9547), .ZN(n12341) );
  OR2_X1 U11300 ( .A1(n12341), .A2(n9796), .ZN(n9551) );
  NAND2_X1 U11301 ( .A1(n9548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9549) );
  XNOR2_X1 U11302 ( .A(n9549), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U11303 ( .A1(n7442), .A2(n13019), .B1(n7444), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n9550) );
  MUX2_X1 U11304 ( .A(n14927), .B(n15753), .S(n9260), .Z(n9555) );
  MUX2_X1 U11305 ( .A(n14927), .B(n15753), .S(n7415), .Z(n9552) );
  NAND2_X1 U11306 ( .A1(n9553), .A2(n9552), .ZN(n9559) );
  INV_X1 U11307 ( .A(n9554), .ZN(n9557) );
  INV_X1 U11308 ( .A(n9555), .ZN(n9556) );
  NAND2_X1 U11309 ( .A1(n9557), .A2(n9556), .ZN(n9558) );
  NAND2_X1 U11310 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  NAND2_X1 U11311 ( .A1(n9618), .A2(n9562), .ZN(n15219) );
  OR2_X1 U11312 ( .A1(n15219), .A2(n9689), .ZN(n9568) );
  INV_X1 U11313 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U11314 ( .A1(n9318), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U11315 ( .A1(n9248), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9563) );
  OAI211_X1 U11316 ( .C1(n9805), .C2(n9565), .A(n9564), .B(n9563), .ZN(n9566)
         );
  INV_X1 U11317 ( .A(n9566), .ZN(n9567) );
  NAND2_X1 U11318 ( .A1(n9568), .A2(n9567), .ZN(n15235) );
  MUX2_X1 U11319 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n11209), .Z(n9578) );
  XNOR2_X1 U11320 ( .A(n9578), .B(SI_19_), .ZN(n9576) );
  XNOR2_X1 U11321 ( .A(n9575), .B(n9576), .ZN(n12537) );
  NAND2_X1 U11322 ( .A1(n12537), .A2(n9820), .ZN(n9572) );
  AOI22_X1 U11323 ( .A1(n9874), .A2(n7443), .B1(n7444), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n9571) );
  MUX2_X1 U11324 ( .A(n15235), .B(n15748), .S(n7415), .Z(n9574) );
  MUX2_X1 U11325 ( .A(n15235), .B(n15748), .S(n9260), .Z(n9573) );
  MUX2_X1 U11326 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n11209), .Z(n9629) );
  OR2_X1 U11327 ( .A1(n9629), .A2(SI_20_), .ZN(n9580) );
  INV_X1 U11328 ( .A(n9578), .ZN(n9579) );
  INV_X1 U11329 ( .A(SI_19_), .ZN(n15474) );
  NAND2_X1 U11330 ( .A1(n9579), .A2(n15474), .ZN(n9627) );
  NAND2_X1 U11331 ( .A1(n9628), .A2(n9581), .ZN(n9583) );
  NAND2_X1 U11332 ( .A1(n9629), .A2(SI_20_), .ZN(n9582) );
  NAND2_X1 U11333 ( .A1(n9583), .A2(n9582), .ZN(n9610) );
  MUX2_X1 U11334 ( .A(n12810), .B(n12807), .S(n11209), .Z(n9584) );
  XNOR2_X1 U11335 ( .A(n9584), .B(SI_21_), .ZN(n9611) );
  NAND2_X1 U11336 ( .A1(n9610), .A2(n9611), .ZN(n9587) );
  INV_X1 U11337 ( .A(n9584), .ZN(n9585) );
  NAND2_X1 U11338 ( .A1(n9585), .A2(SI_21_), .ZN(n9586) );
  NAND2_X1 U11339 ( .A1(n9656), .A2(n9930), .ZN(n9589) );
  INV_X1 U11340 ( .A(n9647), .ZN(n9593) );
  INV_X1 U11341 ( .A(n9591), .ZN(n9603) );
  INV_X1 U11342 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14881) );
  NAND2_X1 U11343 ( .A1(n9603), .A2(n14881), .ZN(n9592) );
  NAND2_X1 U11344 ( .A1(n9593), .A2(n9592), .ZN(n15167) );
  INV_X1 U11345 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11346 ( .A1(n9318), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U11347 ( .A1(n9248), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9594) );
  OAI211_X1 U11348 ( .C1(n9805), .C2(n9596), .A(n9595), .B(n9594), .ZN(n9597)
         );
  INV_X1 U11349 ( .A(n9597), .ZN(n9598) );
  NAND2_X1 U11350 ( .A1(n15726), .A2(n14830), .ZN(n10571) );
  INV_X1 U11351 ( .A(n9600), .ZN(n9620) );
  INV_X1 U11352 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U11353 ( .A1(n9620), .A2(n9601), .ZN(n9602) );
  INV_X1 U11354 ( .A(n9689), .ZN(n9604) );
  NAND2_X1 U11355 ( .A1(n15186), .A2(n9604), .ZN(n9609) );
  INV_X1 U11356 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15736) );
  NAND2_X1 U11357 ( .A1(n9318), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U11358 ( .A1(n9248), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9605) );
  OAI211_X1 U11359 ( .C1(n9805), .C2(n15736), .A(n9606), .B(n9605), .ZN(n9607)
         );
  INV_X1 U11360 ( .A(n9607), .ZN(n9608) );
  AND2_X1 U11361 ( .A1(n15194), .A2(n7415), .ZN(n9616) );
  NOR2_X1 U11362 ( .A1(n15194), .A2(n7415), .ZN(n9615) );
  INV_X1 U11363 ( .A(n9611), .ZN(n9612) );
  XNOR2_X1 U11364 ( .A(n9610), .B(n9612), .ZN(n12806) );
  NAND2_X1 U11365 ( .A1(n12806), .A2(n9820), .ZN(n9614) );
  NAND2_X1 U11366 ( .A1(n7444), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9613) );
  MUX2_X1 U11367 ( .A(n9616), .B(n9615), .S(n15729), .Z(n9617) );
  NAND2_X1 U11368 ( .A1(n9618), .A2(n11105), .ZN(n9619) );
  NAND2_X1 U11369 ( .A1(n9620), .A2(n9619), .ZN(n15202) );
  OR2_X1 U11370 ( .A1(n15202), .A2(n7433), .ZN(n9626) );
  INV_X1 U11371 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U11372 ( .A1(n9318), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U11373 ( .A1(n9248), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9621) );
  OAI211_X1 U11374 ( .C1(n9805), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9624)
         );
  INV_X1 U11375 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U11376 ( .A1(n9626), .A2(n9625), .ZN(n14926) );
  NAND2_X1 U11377 ( .A1(n9628), .A2(n9627), .ZN(n9632) );
  INV_X1 U11378 ( .A(n9629), .ZN(n9630) );
  XNOR2_X1 U11379 ( .A(n9630), .B(SI_20_), .ZN(n9631) );
  XNOR2_X1 U11380 ( .A(n9632), .B(n9631), .ZN(n12666) );
  NAND2_X1 U11381 ( .A1(n12666), .A2(n9820), .ZN(n9634) );
  NAND2_X1 U11382 ( .A1(n7444), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9633) );
  MUX2_X1 U11383 ( .A(n14926), .B(n15739), .S(n9260), .Z(n9638) );
  AND2_X1 U11384 ( .A1(n14926), .A2(n9260), .ZN(n9635) );
  AOI21_X1 U11385 ( .B1(n15739), .B2(n7415), .A(n9635), .ZN(n9639) );
  NAND2_X1 U11386 ( .A1(n9638), .A2(n9639), .ZN(n9636) );
  XNOR2_X1 U11387 ( .A(n15729), .B(n15194), .ZN(n9854) );
  OAI21_X1 U11388 ( .B1(n9639), .B2(n9638), .A(n9854), .ZN(n9643) );
  OR2_X1 U11389 ( .A1(n9640), .A2(n7415), .ZN(n9641) );
  OAI21_X1 U11390 ( .B1(n10571), .B2(n9260), .A(n9641), .ZN(n9642) );
  AOI21_X1 U11391 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9645) );
  NAND2_X1 U11392 ( .A1(n9646), .A2(n9645), .ZN(n9663) );
  NOR2_X1 U11393 ( .A1(n9647), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9648) );
  OR2_X1 U11394 ( .A1(n9669), .A2(n9648), .ZN(n15145) );
  OR2_X1 U11395 ( .A1(n15145), .A2(n7434), .ZN(n9654) );
  INV_X1 U11396 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U11397 ( .A1(n9248), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U11398 ( .A1(n9318), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9649) );
  OAI211_X1 U11399 ( .C1(n9805), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9652)
         );
  INV_X1 U11400 ( .A(n9652), .ZN(n9653) );
  MUX2_X1 U11401 ( .A(n9655), .B(n13039), .S(n11209), .Z(n10252) );
  INV_X1 U11402 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9658) );
  MUX2_X1 U11403 ( .A(n9658), .B(n13003), .S(n11209), .Z(n9678) );
  XNOR2_X1 U11404 ( .A(n9678), .B(SI_23_), .ZN(n9677) );
  XNOR2_X1 U11405 ( .A(n9681), .B(n9677), .ZN(n13000) );
  NAND2_X1 U11406 ( .A1(n13000), .A2(n9820), .ZN(n9660) );
  NAND2_X1 U11407 ( .A1(n7444), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U11408 ( .A1(n9663), .A2(n9664), .ZN(n9662) );
  MUX2_X1 U11409 ( .A(n15718), .B(n14924), .S(n7415), .Z(n9661) );
  NAND2_X1 U11410 ( .A1(n9662), .A2(n9661), .ZN(n9668) );
  INV_X1 U11411 ( .A(n9663), .ZN(n9666) );
  INV_X1 U11412 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U11413 ( .A1(n9666), .A2(n9665), .ZN(n9667) );
  OR2_X1 U11414 ( .A1(n9669), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U11415 ( .A1(n9669), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U11416 ( .A1(n9670), .A2(n9687), .ZN(n15134) );
  INV_X1 U11417 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U11418 ( .A1(n9318), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U11419 ( .A1(n9248), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9671) );
  OAI211_X1 U11420 ( .C1(n9805), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9674)
         );
  INV_X1 U11421 ( .A(n9674), .ZN(n9675) );
  INV_X1 U11422 ( .A(n9678), .ZN(n9679) );
  NAND2_X1 U11423 ( .A1(n9679), .A2(SI_23_), .ZN(n9680) );
  XNOR2_X1 U11424 ( .A(n9725), .B(SI_24_), .ZN(n9694) );
  MUX2_X1 U11425 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n11209), .Z(n9718) );
  XNOR2_X1 U11426 ( .A(n9694), .B(n9718), .ZN(n13203) );
  NAND2_X1 U11427 ( .A1(n13203), .A2(n9820), .ZN(n9683) );
  NAND2_X1 U11428 ( .A1(n7444), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9682) );
  NAND2_X2 U11429 ( .A1(n9683), .A2(n9682), .ZN(n15711) );
  MUX2_X1 U11430 ( .A(n15114), .B(n15711), .S(n9260), .Z(n9685) );
  MUX2_X1 U11431 ( .A(n15114), .B(n15711), .S(n7415), .Z(n9684) );
  INV_X1 U11432 ( .A(n9685), .ZN(n9686) );
  NAND2_X1 U11433 ( .A1(n9248), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9693) );
  INV_X1 U11434 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15778) );
  OR2_X1 U11435 ( .A1(n7450), .A2(n15778), .ZN(n9692) );
  INV_X1 U11436 ( .A(n9687), .ZN(n9688) );
  NAND2_X1 U11437 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9688), .ZN(n9710) );
  OAI21_X1 U11438 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9688), .A(n9710), .ZN(
        n15120) );
  OR2_X1 U11439 ( .A1(n9689), .A2(n15120), .ZN(n9691) );
  INV_X1 U11440 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15707) );
  OR2_X1 U11441 ( .A1(n9805), .A2(n15707), .ZN(n9690) );
  NAND4_X1 U11442 ( .A1(n9693), .A2(n9692), .A3(n9691), .A4(n9690), .ZN(n14923) );
  INV_X1 U11443 ( .A(n9694), .ZN(n9695) );
  NAND2_X1 U11444 ( .A1(n9695), .A2(n9718), .ZN(n9697) );
  NAND2_X1 U11445 ( .A1(n9725), .A2(SI_24_), .ZN(n9696) );
  NAND2_X1 U11446 ( .A1(n9697), .A2(n9696), .ZN(n9701) );
  MUX2_X1 U11447 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n11209), .Z(n9698) );
  NAND2_X1 U11448 ( .A1(n9698), .A2(SI_25_), .ZN(n9721) );
  INV_X1 U11449 ( .A(n9698), .ZN(n9699) );
  NAND2_X1 U11450 ( .A1(n9699), .A2(n15466), .ZN(n9719) );
  NAND2_X1 U11451 ( .A1(n9721), .A2(n9719), .ZN(n9700) );
  NAND2_X1 U11452 ( .A1(n7444), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9702) );
  NAND2_X2 U11453 ( .A1(n9703), .A2(n9702), .ZN(n15123) );
  MUX2_X1 U11454 ( .A(n14923), .B(n15123), .S(n7415), .Z(n9706) );
  MUX2_X1 U11455 ( .A(n14923), .B(n15123), .S(n9260), .Z(n9704) );
  NAND2_X1 U11456 ( .A1(n7447), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9716) );
  INV_X1 U11457 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9707) );
  OR2_X1 U11458 ( .A1(n7439), .A2(n9707), .ZN(n9715) );
  INV_X1 U11459 ( .A(n9710), .ZN(n9708) );
  INV_X1 U11460 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U11461 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  NAND2_X1 U11462 ( .A1(n9750), .A2(n9711), .ZN(n15099) );
  OR2_X1 U11463 ( .A1(n7433), .A2(n15099), .ZN(n9714) );
  INV_X1 U11464 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9712) );
  OR2_X1 U11465 ( .A1(n7450), .A2(n9712), .ZN(n9713) );
  NAND4_X1 U11466 ( .A1(n9716), .A2(n9715), .A3(n9714), .A4(n9713), .ZN(n14922) );
  INV_X1 U11467 ( .A(n9718), .ZN(n9717) );
  OAI21_X1 U11468 ( .B1(n12905), .B2(n9717), .A(n9721), .ZN(n9724) );
  NOR2_X1 U11469 ( .A1(n9718), .A2(SI_24_), .ZN(n9722) );
  INV_X1 U11470 ( .A(n9719), .ZN(n9720) );
  AOI21_X1 U11471 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9723) );
  XNOR2_X1 U11472 ( .A(n9768), .B(SI_26_), .ZN(n9737) );
  MUX2_X1 U11473 ( .A(n9726), .B(n14787), .S(n11209), .Z(n9762) );
  XNOR2_X1 U11474 ( .A(n9737), .B(n9762), .ZN(n14786) );
  NAND2_X1 U11475 ( .A1(n7444), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9727) );
  MUX2_X1 U11476 ( .A(n14922), .B(n15696), .S(n9260), .Z(n9729) );
  INV_X1 U11477 ( .A(n9729), .ZN(n9730) );
  NAND2_X1 U11478 ( .A1(n7447), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9736) );
  INV_X1 U11479 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9731) );
  OR2_X1 U11480 ( .A1(n7438), .A2(n9731), .ZN(n9735) );
  INV_X1 U11481 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14798) );
  XNOR2_X1 U11482 ( .A(n9750), .B(n14798), .ZN(n14799) );
  OR2_X1 U11483 ( .A1(n7433), .A2(n14799), .ZN(n9734) );
  INV_X1 U11484 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9732) );
  OR2_X1 U11485 ( .A1(n7450), .A2(n9732), .ZN(n9733) );
  NAND4_X1 U11486 ( .A1(n9736), .A2(n9735), .A3(n9734), .A4(n9733), .ZN(n15076) );
  INV_X1 U11487 ( .A(n9762), .ZN(n9761) );
  NAND2_X1 U11488 ( .A1(n9737), .A2(n9761), .ZN(n9739) );
  OR2_X1 U11489 ( .A1(n9768), .A2(n13069), .ZN(n9738) );
  NAND2_X1 U11490 ( .A1(n9739), .A2(n9738), .ZN(n9741) );
  MUX2_X1 U11491 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n11209), .Z(n9763) );
  XNOR2_X1 U11492 ( .A(n9763), .B(SI_27_), .ZN(n9740) );
  NAND2_X1 U11493 ( .A1(n14783), .A2(n9820), .ZN(n9743) );
  NAND2_X1 U11494 ( .A1(n7444), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9742) );
  NAND2_X2 U11495 ( .A1(n9743), .A2(n9742), .ZN(n15691) );
  MUX2_X1 U11496 ( .A(n15076), .B(n15691), .S(n7415), .Z(n9747) );
  NAND2_X1 U11497 ( .A1(n9746), .A2(n9747), .ZN(n9745) );
  MUX2_X1 U11498 ( .A(n15076), .B(n15691), .S(n9260), .Z(n9744) );
  INV_X1 U11499 ( .A(n9746), .ZN(n9749) );
  INV_X1 U11500 ( .A(n9747), .ZN(n9748) );
  NAND2_X1 U11501 ( .A1(n7447), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9759) );
  INV_X1 U11502 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n15087) );
  OR2_X1 U11503 ( .A1(n7439), .A2(n15087), .ZN(n9758) );
  INV_X1 U11504 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13321) );
  OAI21_X1 U11505 ( .B1(n9750), .B2(n14798), .A(n13321), .ZN(n9753) );
  INV_X1 U11506 ( .A(n9750), .ZN(n9752) );
  AND2_X1 U11507 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9751) );
  NAND2_X1 U11508 ( .A1(n9752), .A2(n9751), .ZN(n10654) );
  NAND2_X1 U11509 ( .A1(n9753), .A2(n10654), .ZN(n15086) );
  OR2_X1 U11510 ( .A1(n7434), .A2(n15086), .ZN(n9757) );
  INV_X1 U11511 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9755) );
  OR2_X1 U11512 ( .A1(n7450), .A2(n9755), .ZN(n9756) );
  NAND4_X1 U11513 ( .A1(n9759), .A2(n9758), .A3(n9757), .A4(n9756), .ZN(n14921) );
  INV_X1 U11514 ( .A(n9763), .ZN(n9760) );
  NAND2_X1 U11515 ( .A1(n9760), .A2(n15461), .ZN(n9764) );
  OAI21_X1 U11516 ( .B1(SI_26_), .B2(n9761), .A(n9764), .ZN(n9767) );
  NOR2_X1 U11517 ( .A1(n9762), .A2(n13069), .ZN(n9765) );
  AOI22_X1 U11518 ( .A1(n9765), .A2(n9764), .B1(n9763), .B2(SI_27_), .ZN(n9766) );
  MUX2_X1 U11519 ( .A(n15798), .B(n14782), .S(n11209), .Z(n9769) );
  NAND2_X1 U11520 ( .A1(n9769), .A2(n15459), .ZN(n9782) );
  INV_X1 U11521 ( .A(n9769), .ZN(n9770) );
  NAND2_X1 U11522 ( .A1(n9770), .A2(SI_28_), .ZN(n9771) );
  NAND2_X1 U11523 ( .A1(n9782), .A2(n9771), .ZN(n9783) );
  NAND2_X1 U11524 ( .A1(n15796), .A2(n9820), .ZN(n9773) );
  NAND2_X1 U11525 ( .A1(n7444), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9772) );
  MUX2_X1 U11526 ( .A(n14921), .B(n15686), .S(n9260), .Z(n9775) );
  NAND2_X1 U11527 ( .A1(n7447), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9781) );
  INV_X1 U11528 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9776) );
  OR2_X1 U11529 ( .A1(n7438), .A2(n9776), .ZN(n9780) );
  OR2_X1 U11530 ( .A1(n9689), .A2(n10654), .ZN(n9779) );
  INV_X1 U11531 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9777) );
  OR2_X1 U11532 ( .A1(n7450), .A2(n9777), .ZN(n9778) );
  NAND4_X1 U11533 ( .A1(n9781), .A2(n9780), .A3(n9779), .A4(n9778), .ZN(n15077) );
  INV_X1 U11534 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14778) );
  MUX2_X1 U11535 ( .A(n13337), .B(n14778), .S(n11209), .Z(n9789) );
  XNOR2_X1 U11536 ( .A(n9789), .B(SI_29_), .ZN(n9787) );
  NAND2_X1 U11537 ( .A1(n13208), .A2(n9820), .ZN(n9786) );
  NAND2_X1 U11538 ( .A1(n7444), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9785) );
  MUX2_X1 U11539 ( .A(n15077), .B(n15679), .S(n7415), .Z(n9829) );
  NAND2_X1 U11540 ( .A1(n9788), .A2(n9787), .ZN(n9791) );
  NAND2_X1 U11541 ( .A1(n9789), .A2(n15460), .ZN(n9790) );
  NAND2_X1 U11542 ( .A1(n9791), .A2(n9790), .ZN(n9794) );
  MUX2_X1 U11543 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11209), .Z(n9792) );
  NAND2_X1 U11544 ( .A1(n9792), .A2(SI_30_), .ZN(n9815) );
  OAI21_X1 U11545 ( .B1(n9792), .B2(SI_30_), .A(n9815), .ZN(n9793) );
  NAND2_X1 U11546 ( .A1(n9794), .A2(n9793), .ZN(n9795) );
  NAND2_X1 U11547 ( .A1(n7444), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9797) );
  INV_X1 U11548 ( .A(n7436), .ZN(n9823) );
  AND2_X1 U11549 ( .A1(n10646), .A2(n9823), .ZN(n10582) );
  INV_X1 U11550 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15266) );
  NOR2_X1 U11551 ( .A1(n9805), .A2(n15266), .ZN(n9803) );
  INV_X1 U11552 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9799) );
  NOR2_X1 U11553 ( .A1(n7438), .A2(n9799), .ZN(n9802) );
  INV_X1 U11554 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U11555 ( .A1(n7450), .A2(n9800), .ZN(n9801) );
  OR3_X1 U11556 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(n14919) );
  INV_X1 U11557 ( .A(n14919), .ZN(n15059) );
  INV_X1 U11558 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9804) );
  OR2_X1 U11559 ( .A1(n9805), .A2(n9804), .ZN(n9810) );
  INV_X1 U11560 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9806) );
  OR2_X1 U11561 ( .A1(n7439), .A2(n9806), .ZN(n9809) );
  INV_X1 U11562 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9807) );
  OR2_X1 U11563 ( .A1(n7450), .A2(n9807), .ZN(n9808) );
  AND3_X1 U11564 ( .A1(n9810), .A2(n9809), .A3(n9808), .ZN(n10652) );
  AOI21_X1 U11565 ( .B1(n10582), .B2(n15059), .A(n10652), .ZN(n9811) );
  MUX2_X1 U11566 ( .A(n15065), .B(n9811), .S(n9260), .Z(n9834) );
  INV_X1 U11567 ( .A(n9834), .ZN(n9814) );
  AOI21_X1 U11568 ( .B1(n9812), .B2(n15059), .A(n10652), .ZN(n9813) );
  MUX2_X1 U11569 ( .A(n15065), .B(n9813), .S(n7415), .Z(n9833) );
  NAND2_X1 U11570 ( .A1(n9814), .A2(n9833), .ZN(n9841) );
  NAND2_X1 U11571 ( .A1(n9816), .A2(n9815), .ZN(n9819) );
  MUX2_X1 U11572 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11209), .Z(n9817) );
  XNOR2_X1 U11573 ( .A(n9817), .B(SI_31_), .ZN(n9818) );
  NAND2_X1 U11574 ( .A1(n10872), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U11575 ( .A1(n7444), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9821) );
  XNOR2_X1 U11576 ( .A(n15262), .B(n14919), .ZN(n9871) );
  NAND2_X1 U11577 ( .A1(n12808), .A2(n9823), .ZN(n10650) );
  NAND2_X1 U11578 ( .A1(n9824), .A2(n10646), .ZN(n11093) );
  NAND2_X1 U11579 ( .A1(n9825), .A2(n7436), .ZN(n9826) );
  NAND2_X1 U11580 ( .A1(n11093), .A2(n9826), .ZN(n9827) );
  NAND2_X1 U11581 ( .A1(n10646), .A2(n16295), .ZN(n16323) );
  NAND2_X1 U11582 ( .A1(n9827), .A2(n16323), .ZN(n9842) );
  NAND4_X1 U11583 ( .A1(n9841), .A2(n9871), .A3(n10650), .A4(n9842), .ZN(n9877) );
  NOR2_X1 U11584 ( .A1(n9883), .A2(n9877), .ZN(n9832) );
  INV_X1 U11585 ( .A(n15077), .ZN(n13322) );
  INV_X1 U11586 ( .A(n15679), .ZN(n10658) );
  MUX2_X1 U11587 ( .A(n13322), .B(n10658), .S(n9260), .Z(n9828) );
  INV_X1 U11588 ( .A(n9838), .ZN(n9831) );
  NAND2_X1 U11589 ( .A1(n9832), .A2(n9831), .ZN(n9886) );
  INV_X1 U11590 ( .A(n9833), .ZN(n9835) );
  NAND2_X1 U11591 ( .A1(n9835), .A2(n9834), .ZN(n9878) );
  OR2_X1 U11592 ( .A1(n15262), .A2(n9260), .ZN(n9847) );
  OR2_X1 U11593 ( .A1(n9847), .A2(n15059), .ZN(n9837) );
  INV_X1 U11594 ( .A(n9842), .ZN(n9848) );
  NAND2_X1 U11595 ( .A1(n15262), .A2(n9260), .ZN(n9849) );
  OR2_X1 U11596 ( .A1(n9849), .A2(n14919), .ZN(n9836) );
  NAND2_X1 U11597 ( .A1(n9838), .A2(n9882), .ZN(n9885) );
  NAND2_X1 U11598 ( .A1(n9848), .A2(n14919), .ZN(n9840) );
  INV_X1 U11599 ( .A(n9847), .ZN(n9839) );
  AOI211_X1 U11600 ( .C1(n15262), .C2(n9841), .A(n9840), .B(n9839), .ZN(n9852)
         );
  NAND2_X1 U11601 ( .A1(n9842), .A2(n14919), .ZN(n9846) );
  INV_X1 U11602 ( .A(n9841), .ZN(n9844) );
  NOR2_X1 U11603 ( .A1(n9842), .A2(n14919), .ZN(n9843) );
  OAI211_X1 U11604 ( .C1(n9844), .C2(n15262), .A(n9843), .B(n9849), .ZN(n9845)
         );
  OAI211_X1 U11605 ( .C1(n9847), .C2(n9846), .A(n9845), .B(n10650), .ZN(n9851)
         );
  NOR3_X1 U11606 ( .A1(n9849), .A2(n9848), .A3(n14919), .ZN(n9850) );
  NOR3_X1 U11607 ( .A1(n9852), .A2(n9851), .A3(n9850), .ZN(n9880) );
  INV_X1 U11608 ( .A(n10652), .ZN(n14920) );
  XOR2_X1 U11609 ( .A(n14920), .B(n15065), .Z(n9869) );
  NAND2_X1 U11610 ( .A1(n15686), .A2(n14921), .ZN(n10640) );
  OR2_X1 U11611 ( .A1(n15686), .A2(n14921), .ZN(n9853) );
  XNOR2_X1 U11612 ( .A(n15711), .B(n14843), .ZN(n15130) );
  XNOR2_X1 U11613 ( .A(n15718), .B(n14924), .ZN(n15151) );
  INV_X1 U11614 ( .A(n14927), .ZN(n15215) );
  XNOR2_X1 U11615 ( .A(n15753), .B(n15215), .ZN(n15227) );
  XNOR2_X1 U11616 ( .A(n15748), .B(n14888), .ZN(n15213) );
  XNOR2_X1 U11617 ( .A(n15757), .B(n15232), .ZN(n15256) );
  INV_X1 U11618 ( .A(n14930), .ZN(n13172) );
  XNOR2_X1 U11619 ( .A(n16561), .B(n13172), .ZN(n10560) );
  INV_X1 U11620 ( .A(n14932), .ZN(n13173) );
  XNOR2_X1 U11621 ( .A(n12813), .B(n13173), .ZN(n12553) );
  XNOR2_X1 U11622 ( .A(n12614), .B(n14933), .ZN(n12616) );
  XNOR2_X1 U11623 ( .A(n12573), .B(n12888), .ZN(n12221) );
  XNOR2_X1 U11624 ( .A(n12236), .B(n12570), .ZN(n12163) );
  XNOR2_X1 U11625 ( .A(n12189), .B(n12166), .ZN(n12179) );
  XNOR2_X2 U11626 ( .A(n16365), .B(n14941), .ZN(n12036) );
  NAND2_X2 U11627 ( .A1(n10538), .A2(n9856), .ZN(n10602) );
  INV_X1 U11628 ( .A(n9857), .ZN(n9858) );
  NAND2_X1 U11629 ( .A1(n10539), .A2(n9858), .ZN(n16296) );
  NOR3_X1 U11630 ( .A1(n16349), .A2(n10602), .A3(n16296), .ZN(n9861) );
  NAND2_X1 U11631 ( .A1(n16401), .A2(n14939), .ZN(n9859) );
  INV_X1 U11632 ( .A(n14939), .ZN(n11845) );
  NAND2_X1 U11633 ( .A1(n12003), .A2(n11845), .ZN(n12178) );
  XNOR2_X2 U11634 ( .A(n14940), .B(n9860), .ZN(n16377) );
  NAND4_X1 U11635 ( .A1(n12036), .A2(n9861), .A3(n11994), .A4(n16381), .ZN(
        n9862) );
  NOR4_X1 U11636 ( .A1(n12221), .A2(n12163), .A3(n12179), .A4(n9862), .ZN(
        n9863) );
  XNOR2_X1 U11637 ( .A(n12928), .B(n14934), .ZN(n10619) );
  XNOR2_X1 U11638 ( .A(n12891), .B(n14935), .ZN(n12197) );
  NAND4_X1 U11639 ( .A1(n12616), .A2(n9863), .A3(n10619), .A4(n12197), .ZN(
        n9864) );
  NOR4_X1 U11640 ( .A1(n10560), .A2(n8236), .A3(n12553), .A4(n9864), .ZN(n9865) );
  XNOR2_X1 U11641 ( .A(n15762), .B(n14928), .ZN(n10563) );
  XNOR2_X1 U11642 ( .A(n11055), .B(n14929), .ZN(n16625) );
  NAND4_X1 U11643 ( .A1(n15256), .A2(n9865), .A3(n10563), .A4(n16625), .ZN(
        n9866) );
  NOR4_X1 U11644 ( .A1(n15175), .A2(n15227), .A3(n15213), .A4(n9866), .ZN(
        n9867) );
  XNOR2_X1 U11645 ( .A(n15739), .B(n14926), .ZN(n15192) );
  NAND4_X1 U11646 ( .A1(n15151), .A2(n10570), .A3(n9867), .A4(n15192), .ZN(
        n9868) );
  NOR4_X1 U11647 ( .A1(n9869), .A2(n15090), .A3(n15130), .A4(n9868), .ZN(n9873) );
  XNOR2_X1 U11648 ( .A(n15679), .B(n13322), .ZN(n10641) );
  NAND2_X1 U11649 ( .A1(n15691), .A2(n14897), .ZN(n15073) );
  OR2_X1 U11650 ( .A1(n15691), .A2(n14897), .ZN(n9870) );
  NAND2_X1 U11651 ( .A1(n15073), .A2(n9870), .ZN(n13214) );
  NOR3_X1 U11652 ( .A1(n10641), .A2(n13214), .A3(n15103), .ZN(n9872) );
  NAND4_X1 U11653 ( .A1(n9873), .A2(n9872), .A3(n15118), .A4(n9871), .ZN(n9875) );
  XNOR2_X1 U11654 ( .A(n9875), .B(n9874), .ZN(n9876) );
  NOR2_X1 U11655 ( .A1(n9876), .A2(n10650), .ZN(n9879) );
  OAI22_X1 U11656 ( .A1(n9880), .A2(n9879), .B1(n9878), .B2(n9877), .ZN(n9881)
         );
  AOI21_X1 U11657 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9884) );
  NAND3_X1 U11658 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(n9894) );
  NAND2_X1 U11659 ( .A1(n9887), .A2(n9888), .ZN(n9889) );
  INV_X1 U11660 ( .A(n11146), .ZN(n9892) );
  NAND2_X1 U11661 ( .A1(n9892), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12998) );
  INV_X1 U11662 ( .A(n12998), .ZN(n9893) );
  NAND2_X1 U11663 ( .A1(n9894), .A2(n9893), .ZN(n9912) );
  NAND2_X1 U11664 ( .A1(n9904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9897) );
  MUX2_X1 U11665 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9897), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9898) );
  INV_X1 U11666 ( .A(n9900), .ZN(n9901) );
  NAND2_X1 U11667 ( .A1(n9901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9902) );
  MUX2_X1 U11668 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9902), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9903) );
  NOR2_X1 U11669 ( .A1(n15807), .A2(n13205), .ZN(n9905) );
  AND2_X1 U11670 ( .A1(n11146), .A2(n10957), .ZN(n9907) );
  AND2_X1 U11671 ( .A1(n7436), .A2(n13032), .ZN(n9906) );
  OR2_X1 U11672 ( .A1(n11093), .A2(n9906), .ZN(n11106) );
  NAND2_X1 U11673 ( .A1(n9907), .A2(n11106), .ZN(n11102) );
  INV_X1 U11674 ( .A(n14954), .ZN(n13024) );
  NAND2_X1 U11675 ( .A1(n13024), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15799) );
  NOR3_X1 U11676 ( .A1(n11102), .A2(n15216), .A3(n15799), .ZN(n9910) );
  OAI21_X1 U11677 ( .B1(n12998), .B2(n9824), .A(P1_B_REG_SCAN_IN), .ZN(n9909)
         );
  OR2_X1 U11678 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  NAND2_X1 U11679 ( .A1(n9912), .A2(n9911), .ZN(P1_U3242) );
  NOR2_X1 U11680 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9924) );
  NOR2_X1 U11681 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9914) );
  NAND2_X1 U11682 ( .A1(n9924), .A2(n9914), .ZN(n9915) );
  NAND4_X1 U11683 ( .A1(n10326), .A2(n10398), .A3(n10391), .A4(n10388), .ZN(
        n9923) );
  NOR2_X1 U11684 ( .A1(n9915), .A2(n9923), .ZN(n9921) );
  NOR2_X2 U11685 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n10173) );
  NOR2_X1 U11686 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n9917) );
  NOR2_X1 U11687 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n9916) );
  NAND3_X1 U11688 ( .A1(n10173), .A2(n9917), .A3(n9916), .ZN(n9920) );
  INV_X1 U11689 ( .A(n9923), .ZN(n9927) );
  INV_X1 U11690 ( .A(n9924), .ZN(n9925) );
  NOR2_X1 U11691 ( .A1(n9925), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9926) );
  NAND4_X1 U11692 ( .A1(n7413), .A2(n10320), .A3(n9927), .A4(n9926), .ZN(n9928) );
  NAND2_X1 U11693 ( .A1(n13203), .A2(n10871), .ZN(n9932) );
  OR2_X1 U11694 ( .A1(n10873), .A2(n8076), .ZN(n9931) );
  AND2_X1 U11695 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10013) );
  NAND2_X1 U11696 ( .A1(n10013), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10039) );
  INV_X1 U11697 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U11698 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U11699 ( .A1(n10037), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10070) );
  INV_X1 U11700 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U11701 ( .A1(n10085), .A2(n10084), .ZN(n10083) );
  NAND2_X1 U11702 ( .A1(n10095), .A2(n9933), .ZN(n10142) );
  NAND2_X1 U11703 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n9934) );
  NAND2_X1 U11704 ( .A1(n10182), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10203) );
  INV_X1 U11705 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U11706 ( .A1(n10229), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n10255) );
  INV_X1 U11707 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14344) );
  INV_X1 U11708 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14273) );
  NAND2_X1 U11709 ( .A1(n9935), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n10279) );
  INV_X1 U11710 ( .A(n9935), .ZN(n10268) );
  INV_X1 U11711 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U11712 ( .A1(n10268), .A2(n9936), .ZN(n9937) );
  NAND2_X1 U11713 ( .A1(n10279), .A2(n9937), .ZN(n14517) );
  INV_X2 U11714 ( .A(n9942), .ZN(n9941) );
  INV_X1 U11715 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9939) );
  XNOR2_X2 U11716 ( .A(n9940), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9963) );
  INV_X1 U11717 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14516) );
  NAND2_X4 U11718 ( .A1(n9941), .A2(n14776), .ZN(n10877) );
  BUF_X2 U11719 ( .A(n9942), .Z(n13212) );
  NAND2_X1 U11720 ( .A1(n10682), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U11721 ( .A1(n13212), .A2(n14776), .ZN(n10035) );
  NAND2_X1 U11722 ( .A1(n10683), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9943) );
  OAI211_X1 U11723 ( .C1(n14516), .C2(n10877), .A(n9944), .B(n9943), .ZN(n9945) );
  INV_X1 U11724 ( .A(n9945), .ZN(n9946) );
  NAND2_X1 U11725 ( .A1(n9947), .A2(n9946), .ZN(n14492) );
  INV_X1 U11726 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U11727 ( .A1(n11209), .A2(SI_0_), .ZN(n9949) );
  XNOR2_X1 U11728 ( .A(n9949), .B(n9948), .ZN(n14793) );
  INV_X1 U11729 ( .A(n11492), .ZN(n10697) );
  AOI22_X1 U11730 ( .A1(n14770), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n9956) );
  INV_X1 U11731 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U11732 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_30__SCAN_IN), 
        .ZN(n9952) );
  OAI21_X1 U11733 ( .B1(n9953), .B2(P2_IR_REG_30__SCAN_IN), .A(n9952), .ZN(
        n9954) );
  NAND2_X1 U11734 ( .A1(n9951), .A2(n9954), .ZN(n9955) );
  OAI21_X1 U11735 ( .B1(n9951), .B2(n9956), .A(n9955), .ZN(n9957) );
  NAND2_X1 U11736 ( .A1(n9957), .A2(n14776), .ZN(n9966) );
  AOI22_X1 U11737 ( .A1(n14770), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n9962) );
  INV_X1 U11738 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U11739 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n9958) );
  OAI21_X1 U11740 ( .B1(n9959), .B2(P2_IR_REG_30__SCAN_IN), .A(n9958), .ZN(
        n9960) );
  NAND2_X1 U11741 ( .A1(n9951), .A2(n9960), .ZN(n9961) );
  OAI21_X1 U11742 ( .B1(n9951), .B2(n9962), .A(n9961), .ZN(n9964) );
  NAND2_X1 U11743 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  INV_X1 U11744 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U11745 ( .A1(n9998), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9967) );
  INV_X1 U11746 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9969) );
  OR2_X1 U11747 ( .A1(n10876), .A2(n9969), .ZN(n9971) );
  INV_X1 U11748 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n12058) );
  OR2_X1 U11749 ( .A1(n10877), .A2(n12058), .ZN(n9970) );
  NAND2_X1 U11750 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9972) );
  MUX2_X1 U11751 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9972), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9973) );
  INV_X1 U11752 ( .A(n9981), .ZN(n9978) );
  NAND2_X1 U11753 ( .A1(n9973), .A2(n9978), .ZN(n11313) );
  INV_X1 U11754 ( .A(n11189), .ZN(n9974) );
  OR2_X1 U11755 ( .A1(n9974), .A2(n10845), .ZN(n9976) );
  OAI211_X2 U11756 ( .C1(n11300), .C2(n11313), .A(n9976), .B(n9975), .ZN(
        n11668) );
  INV_X1 U11757 ( .A(n10333), .ZN(n11662) );
  NAND2_X1 U11758 ( .A1(n7506), .A2(n11662), .ZN(n11661) );
  OR2_X1 U11759 ( .A1(n7435), .A2(n11668), .ZN(n9977) );
  OR2_X1 U11760 ( .A1(n11216), .A2(n10845), .ZN(n9984) );
  INV_X2 U11761 ( .A(n11300), .ZN(n10215) );
  NAND2_X1 U11762 ( .A1(n9978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9979) );
  MUX2_X1 U11763 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9979), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n9982) );
  AND2_X1 U11764 ( .A1(n9981), .A2(n9980), .ZN(n10061) );
  INV_X1 U11765 ( .A(n10061), .ZN(n9992) );
  NAND2_X1 U11766 ( .A1(n9982), .A2(n9992), .ZN(n11316) );
  INV_X1 U11767 ( .A(n11316), .ZN(n15846) );
  NAND2_X1 U11768 ( .A1(n9998), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9990) );
  INV_X1 U11769 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9985) );
  OR2_X1 U11770 ( .A1(n9999), .A2(n9985), .ZN(n9989) );
  INV_X1 U11771 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11315) );
  OR2_X1 U11772 ( .A1(n10877), .A2(n11315), .ZN(n9988) );
  INV_X1 U11773 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9986) );
  OR2_X1 U11774 ( .A1(n10876), .A2(n9986), .ZN(n9987) );
  XNOR2_X1 U11775 ( .A(n11679), .B(n14386), .ZN(n10849) );
  INV_X1 U11776 ( .A(n11679), .ZN(n12271) );
  INV_X1 U11777 ( .A(n14386), .ZN(n10337) );
  NAND2_X1 U11778 ( .A1(n12271), .A2(n10337), .ZN(n9991) );
  NAND2_X1 U11779 ( .A1(n11187), .A2(n10871), .ZN(n9997) );
  NAND2_X1 U11780 ( .A1(n9992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9993) );
  INV_X1 U11781 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9994) );
  MUX2_X1 U11782 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9993), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9995) );
  AND2_X1 U11783 ( .A1(n10061), .A2(n9994), .ZN(n10009) );
  INV_X1 U11784 ( .A(n10009), .ZN(n10006) );
  AOI22_X1 U11785 ( .A1(n10005), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10215), 
        .B2(n14391), .ZN(n9996) );
  NAND2_X1 U11786 ( .A1(n10683), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n10003) );
  OR2_X1 U11787 ( .A1(n9999), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10002) );
  INV_X1 U11788 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n12044) );
  OR2_X1 U11789 ( .A1(n10877), .A2(n12044), .ZN(n10001) );
  INV_X1 U11790 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11293) );
  OR2_X1 U11791 ( .A1(n10876), .A2(n11293), .ZN(n10000) );
  XNOR2_X1 U11792 ( .A(n12045), .B(n14384), .ZN(n10852) );
  INV_X1 U11793 ( .A(n10852), .ZN(n11686) );
  OR2_X1 U11794 ( .A1(n12045), .A2(n14384), .ZN(n10004) );
  NAND2_X1 U11795 ( .A1(n11681), .A2(n10004), .ZN(n11611) );
  NAND2_X1 U11796 ( .A1(n11191), .A2(n10871), .ZN(n10012) );
  NAND2_X1 U11797 ( .A1(n10006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10007) );
  MUX2_X1 U11798 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10007), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n10010) );
  INV_X1 U11799 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U11800 ( .A1(n10009), .A2(n10008), .ZN(n10020) );
  NAND2_X1 U11801 ( .A1(n10010), .A2(n10020), .ZN(n11319) );
  INV_X1 U11802 ( .A(n11319), .ZN(n14404) );
  AOI22_X1 U11803 ( .A1(n10005), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10215), 
        .B2(n14404), .ZN(n10011) );
  NAND2_X1 U11804 ( .A1(n10012), .A2(n10011), .ZN(n11612) );
  NAND2_X1 U11805 ( .A1(n10683), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n10017) );
  INV_X1 U11806 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11294) );
  OR2_X1 U11807 ( .A1(n10876), .A2(n11294), .ZN(n10016) );
  INV_X1 U11808 ( .A(n10013), .ZN(n10025) );
  OAI21_X1 U11809 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n10025), .ZN(n11568) );
  OR2_X1 U11810 ( .A1(n9999), .A2(n11568), .ZN(n10015) );
  INV_X1 U11811 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11318) );
  OR2_X1 U11812 ( .A1(n10877), .A2(n11318), .ZN(n10014) );
  NAND2_X1 U11813 ( .A1(n11611), .A2(n11614), .ZN(n11610) );
  INV_X1 U11814 ( .A(n11612), .ZN(n12303) );
  NAND2_X1 U11815 ( .A1(n12303), .A2(n11647), .ZN(n10018) );
  OR2_X1 U11816 ( .A1(n11210), .A2(n10845), .ZN(n10023) );
  NAND2_X1 U11817 ( .A1(n10020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10019) );
  MUX2_X1 U11818 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10019), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n10021) );
  AOI22_X1 U11819 ( .A1(n10005), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10215), 
        .B2(n14424), .ZN(n10022) );
  NAND2_X1 U11820 ( .A1(n10023), .A2(n10022), .ZN(n11701) );
  NAND2_X1 U11821 ( .A1(n10683), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n10030) );
  INV_X1 U11822 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U11823 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  NAND2_X1 U11824 ( .A1(n10039), .A2(n10026), .ZN(n12070) );
  OR2_X1 U11825 ( .A1(n9999), .A2(n12070), .ZN(n10029) );
  INV_X1 U11826 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11320) );
  OR2_X1 U11827 ( .A1(n10877), .A2(n11320), .ZN(n10028) );
  INV_X1 U11828 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11295) );
  OR2_X1 U11829 ( .A1(n10876), .A2(n11295), .ZN(n10027) );
  NAND4_X1 U11830 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        n14382) );
  XNOR2_X1 U11831 ( .A(n11701), .B(n14382), .ZN(n10851) );
  INV_X1 U11832 ( .A(n10851), .ZN(n11703) );
  INV_X1 U11833 ( .A(n14382), .ZN(n11656) );
  NAND2_X1 U11834 ( .A1(n12071), .A2(n11656), .ZN(n10031) );
  OR2_X1 U11835 ( .A1(n11253), .A2(n10845), .ZN(n10034) );
  NAND2_X1 U11836 ( .A1(n10046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10032) );
  XNOR2_X1 U11837 ( .A(n10032), .B(P2_IR_REG_6__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U11838 ( .A1(n10005), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10215), 
        .B2(n11297), .ZN(n10033) );
  NAND2_X1 U11839 ( .A1(n10034), .A2(n10033), .ZN(n16419) );
  NAND2_X1 U11840 ( .A1(n10682), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10044) );
  INV_X1 U11841 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10036) );
  OR2_X1 U11842 ( .A1(n10878), .A2(n10036), .ZN(n10043) );
  INV_X1 U11843 ( .A(n10037), .ZN(n10052) );
  NAND2_X1 U11844 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  NAND2_X1 U11845 ( .A1(n10052), .A2(n10040), .ZN(n12259) );
  OR2_X1 U11846 ( .A1(n9999), .A2(n12259), .ZN(n10042) );
  INV_X1 U11847 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n12260) );
  OR2_X1 U11848 ( .A1(n10877), .A2(n12260), .ZN(n10041) );
  NAND4_X1 U11849 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n14381) );
  XNOR2_X1 U11850 ( .A(n16419), .B(n14381), .ZN(n12245) );
  INV_X1 U11851 ( .A(n12245), .ZN(n12250) );
  OR2_X1 U11852 ( .A1(n16419), .A2(n14381), .ZN(n10045) );
  NAND2_X1 U11853 ( .A1(n12253), .A2(n10045), .ZN(n12078) );
  OR2_X1 U11854 ( .A1(n11212), .A2(n10845), .ZN(n10049) );
  OAI21_X1 U11855 ( .B1(n10046), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10047) );
  XNOR2_X1 U11856 ( .A(n10047), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U11857 ( .A1(n10005), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11366), 
        .B2(n10215), .ZN(n10048) );
  NAND2_X1 U11858 ( .A1(n10049), .A2(n10048), .ZN(n12088) );
  NAND2_X1 U11859 ( .A1(n10682), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10057) );
  INV_X1 U11860 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10050) );
  OR2_X1 U11861 ( .A1(n10878), .A2(n10050), .ZN(n10056) );
  INV_X1 U11862 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U11863 ( .A1(n10052), .A2(n10051), .ZN(n10053) );
  NAND2_X1 U11864 ( .A1(n10070), .A2(n10053), .ZN(n12090) );
  OR2_X1 U11865 ( .A1(n9999), .A2(n12090), .ZN(n10055) );
  INV_X1 U11866 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n12086) );
  OR2_X1 U11867 ( .A1(n10877), .A2(n12086), .ZN(n10054) );
  XNOR2_X1 U11868 ( .A(n12088), .B(n12247), .ZN(n12082) );
  NAND2_X1 U11869 ( .A1(n12078), .A2(n12082), .ZN(n12077) );
  INV_X1 U11870 ( .A(n12247), .ZN(n12126) );
  OR2_X1 U11871 ( .A1(n12088), .A2(n12126), .ZN(n10058) );
  NAND2_X1 U11872 ( .A1(n12077), .A2(n10058), .ZN(n12123) );
  INV_X1 U11873 ( .A(n12123), .ZN(n10077) );
  OR2_X1 U11874 ( .A1(n11248), .A2(n10845), .ZN(n10067) );
  INV_X1 U11875 ( .A(n10059), .ZN(n10060) );
  NOR2_X1 U11876 ( .A1(n10060), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U11877 ( .A1(n10062), .A2(n10061), .ZN(n10064) );
  NAND2_X1 U11878 ( .A1(n10064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10063) );
  MUX2_X1 U11879 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10063), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n10065) );
  AOI22_X1 U11880 ( .A1(n10005), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10215), 
        .B2(n11423), .ZN(n10066) );
  NAND2_X1 U11881 ( .A1(n10067), .A2(n10066), .ZN(n12142) );
  NAND2_X1 U11882 ( .A1(n10683), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10075) );
  INV_X1 U11883 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10068) );
  OR2_X1 U11884 ( .A1(n10876), .A2(n10068), .ZN(n10074) );
  NAND2_X1 U11885 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  NAND2_X1 U11886 ( .A1(n10085), .A2(n10071), .ZN(n12136) );
  OR2_X1 U11887 ( .A1(n9999), .A2(n12136), .ZN(n10073) );
  INV_X1 U11888 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12137) );
  OR2_X1 U11889 ( .A1(n10877), .A2(n12137), .ZN(n10072) );
  NAND2_X1 U11890 ( .A1(n12142), .A2(n12352), .ZN(n10350) );
  OR2_X1 U11891 ( .A1(n12142), .A2(n12352), .ZN(n10076) );
  NAND2_X1 U11892 ( .A1(n10350), .A2(n10076), .ZN(n10855) );
  INV_X1 U11893 ( .A(n10855), .ZN(n12128) );
  INV_X1 U11894 ( .A(n12352), .ZN(n14380) );
  NAND2_X1 U11895 ( .A1(n12142), .A2(n14380), .ZN(n10078) );
  NAND2_X1 U11896 ( .A1(n10079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10080) );
  XNOR2_X1 U11897 ( .A(n10080), .B(P2_IR_REG_9__SCAN_IN), .ZN(n15923) );
  AOI22_X1 U11898 ( .A1(n10005), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10215), 
        .B2(n15923), .ZN(n10081) );
  NAND2_X1 U11899 ( .A1(n10682), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10090) );
  INV_X1 U11900 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10082) );
  OR2_X1 U11901 ( .A1(n10878), .A2(n10082), .ZN(n10089) );
  INV_X1 U11902 ( .A(n10083), .ZN(n10097) );
  NAND2_X1 U11903 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  NAND2_X1 U11904 ( .A1(n10097), .A2(n10086), .ZN(n12351) );
  OR2_X1 U11905 ( .A1(n9999), .A2(n12351), .ZN(n10088) );
  INV_X1 U11906 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n12207) );
  OR2_X1 U11907 ( .A1(n10877), .A2(n12207), .ZN(n10087) );
  NAND4_X1 U11908 ( .A1(n10090), .A2(n10089), .A3(n10088), .A4(n10087), .ZN(
        n14379) );
  OR2_X1 U11909 ( .A1(n11287), .A2(n10845), .ZN(n10094) );
  NAND2_X1 U11910 ( .A1(n10176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10092) );
  XNOR2_X1 U11911 ( .A(n10092), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U11912 ( .A1(n10005), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10215), 
        .B2(n11474), .ZN(n10093) );
  NAND2_X1 U11913 ( .A1(n10682), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10102) );
  OR2_X1 U11914 ( .A1(n10878), .A2(n16481), .ZN(n10101) );
  INV_X1 U11915 ( .A(n10095), .ZN(n10129) );
  INV_X1 U11916 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U11917 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NAND2_X1 U11918 ( .A1(n10129), .A2(n10098), .ZN(n12474) );
  OR2_X1 U11919 ( .A1(n9999), .A2(n12474), .ZN(n10100) );
  INV_X1 U11920 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n12379) );
  OR2_X1 U11921 ( .A1(n10877), .A2(n12379), .ZN(n10099) );
  OR2_X1 U11922 ( .A1(n12463), .A2(n12634), .ZN(n10351) );
  NAND2_X1 U11923 ( .A1(n12463), .A2(n12634), .ZN(n10103) );
  NAND2_X1 U11924 ( .A1(n12370), .A2(n12371), .ZN(n10105) );
  INV_X1 U11925 ( .A(n12634), .ZN(n12355) );
  NAND2_X1 U11926 ( .A1(n12463), .A2(n12355), .ZN(n10104) );
  NAND2_X1 U11927 ( .A1(n10105), .A2(n10104), .ZN(n12448) );
  NAND2_X1 U11928 ( .A1(n11344), .A2(n10871), .ZN(n10109) );
  NOR2_X1 U11929 ( .A1(n10176), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n10116) );
  INV_X1 U11930 ( .A(n10116), .ZN(n10106) );
  NAND2_X1 U11931 ( .A1(n10106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10107) );
  XNOR2_X1 U11932 ( .A(n10107), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U11933 ( .A1(n10005), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10215), 
        .B2(n11874), .ZN(n10108) );
  NAND2_X1 U11934 ( .A1(n10682), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10114) );
  INV_X1 U11935 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10110) );
  OR2_X1 U11936 ( .A1(n10878), .A2(n10110), .ZN(n10113) );
  INV_X1 U11937 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10128) );
  XNOR2_X1 U11938 ( .A(n10129), .B(n10128), .ZN(n12633) );
  OR2_X1 U11939 ( .A1(n9999), .A2(n12633), .ZN(n10112) );
  INV_X1 U11940 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12452) );
  OR2_X1 U11941 ( .A1(n10877), .A2(n12452), .ZN(n10111) );
  NAND4_X1 U11942 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n14378) );
  XNOR2_X1 U11943 ( .A(n12644), .B(n14378), .ZN(n12456) );
  INV_X1 U11944 ( .A(n12456), .ZN(n12449) );
  NAND2_X1 U11945 ( .A1(n12644), .A2(n14378), .ZN(n10115) );
  NAND2_X1 U11946 ( .A1(n11436), .A2(n10871), .ZN(n10125) );
  AND2_X1 U11947 ( .A1(n10117), .A2(n10116), .ZN(n10121) );
  INV_X1 U11948 ( .A(n10121), .ZN(n10118) );
  NAND2_X1 U11949 ( .A1(n10118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U11950 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10119), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n10122) );
  NAND2_X1 U11951 ( .A1(n10121), .A2(n10120), .ZN(n10137) );
  NAND2_X1 U11952 ( .A1(n10122), .A2(n10137), .ZN(n15896) );
  OAI22_X1 U11953 ( .A1(n10873), .A2(n11440), .B1(n11300), .B2(n15896), .ZN(
        n10123) );
  INV_X1 U11954 ( .A(n10123), .ZN(n10124) );
  NAND2_X1 U11955 ( .A1(n10682), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10134) );
  INV_X1 U11956 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10126) );
  OR2_X1 U11957 ( .A1(n10878), .A2(n10126), .ZN(n10133) );
  INV_X1 U11958 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10127) );
  OAI21_X1 U11959 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(n10130) );
  NAND2_X1 U11960 ( .A1(n10130), .A2(n10142), .ZN(n12783) );
  OR2_X1 U11961 ( .A1(n9999), .A2(n12783), .ZN(n10132) );
  INV_X1 U11962 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12599) );
  OR2_X1 U11963 ( .A1(n10877), .A2(n12599), .ZN(n10131) );
  INV_X1 U11964 ( .A(n12772), .ZN(n12702) );
  OR2_X1 U11965 ( .A1(n12770), .A2(n12702), .ZN(n10135) );
  OR2_X1 U11966 ( .A1(n11445), .A2(n10845), .ZN(n10140) );
  NAND2_X1 U11967 ( .A1(n10137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10136) );
  MUX2_X1 U11968 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10136), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n10138) );
  AOI22_X1 U11969 ( .A1(n12583), .A2(n10215), .B1(n10005), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U11970 ( .A1(n10682), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10147) );
  INV_X1 U11971 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10141) );
  OR2_X1 U11972 ( .A1(n10878), .A2(n10141), .ZN(n10146) );
  NAND2_X1 U11973 ( .A1(n10142), .A2(n12876), .ZN(n10143) );
  NAND2_X1 U11974 ( .A1(n10162), .A2(n10143), .ZN(n12875) );
  OR2_X1 U11975 ( .A1(n9999), .A2(n12875), .ZN(n10145) );
  INV_X1 U11976 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11872) );
  OR2_X1 U11977 ( .A1(n10877), .A2(n11872), .ZN(n10144) );
  XNOR2_X1 U11978 ( .A(n12863), .B(n12864), .ZN(n10858) );
  INV_X1 U11979 ( .A(n12864), .ZN(n14377) );
  NAND2_X1 U11980 ( .A1(n12863), .A2(n14377), .ZN(n10148) );
  NAND2_X1 U11981 ( .A1(n12708), .A2(n10148), .ZN(n16572) );
  NAND2_X1 U11982 ( .A1(n11544), .A2(n10871), .ZN(n10151) );
  NAND2_X1 U11983 ( .A1(n10157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10149) );
  XNOR2_X1 U11984 ( .A(n10149), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15859) );
  AOI22_X1 U11985 ( .A1(n15859), .A2(n10215), .B1(n10005), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n10150) );
  XNOR2_X1 U11986 ( .A(n10162), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n16597) );
  NAND2_X1 U11987 ( .A1(n16597), .A2(n10375), .ZN(n10155) );
  NAND2_X1 U11988 ( .A1(n10683), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10154) );
  NAND2_X1 U11989 ( .A1(n10682), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10153) );
  INV_X1 U11990 ( .A(n10877), .ZN(n10376) );
  NAND2_X1 U11991 ( .A1(n10376), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10152) );
  AND4_X1 U11992 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n12931) );
  XNOR2_X1 U11993 ( .A(n16600), .B(n12931), .ZN(n16581) );
  INV_X1 U11994 ( .A(n12931), .ZN(n14376) );
  NAND2_X1 U11995 ( .A1(n16600), .A2(n14376), .ZN(n10156) );
  NAND2_X1 U11996 ( .A1(n11716), .A2(n10871), .ZN(n10160) );
  OAI21_X1 U11997 ( .B1(n10157), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10158) );
  XNOR2_X1 U11998 ( .A(n10158), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U11999 ( .A1(n12718), .A2(n10215), .B1(n10005), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n10159) );
  INV_X1 U12000 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12942) );
  INV_X1 U12001 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10161) );
  OAI21_X1 U12002 ( .B1(n10162), .B2(n12942), .A(n10161), .ZN(n10163) );
  AND2_X1 U12003 ( .A1(n10163), .A2(n10183), .ZN(n13064) );
  NAND2_X1 U12004 ( .A1(n13064), .A2(n10375), .ZN(n10170) );
  INV_X1 U12005 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10164) );
  OR2_X1 U12006 ( .A1(n10876), .A2(n10164), .ZN(n10167) );
  INV_X1 U12007 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10165) );
  OR2_X1 U12008 ( .A1(n10878), .A2(n10165), .ZN(n10166) );
  AND2_X1 U12009 ( .A1(n10167), .A2(n10166), .ZN(n10169) );
  NAND2_X1 U12010 ( .A1(n10376), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n10168) );
  AND3_X1 U12011 ( .A1(n10170), .A2(n10169), .A3(n10168), .ZN(n10357) );
  XNOR2_X1 U12012 ( .A(n13050), .B(n10357), .ZN(n12912) );
  INV_X1 U12013 ( .A(n12912), .ZN(n12909) );
  OR2_X1 U12014 ( .A1(n13050), .A2(n14375), .ZN(n10171) );
  NAND2_X1 U12015 ( .A1(n11899), .A2(n10871), .ZN(n10181) );
  INV_X1 U12016 ( .A(n10172), .ZN(n10174) );
  NAND2_X1 U12017 ( .A1(n10174), .A2(n10173), .ZN(n10175) );
  NAND2_X1 U12018 ( .A1(n7565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10177) );
  MUX2_X1 U12019 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10177), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n10179) );
  AND2_X1 U12020 ( .A1(n10179), .A2(n7560), .ZN(n15874) );
  AOI22_X1 U12021 ( .A1(n10005), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10215), 
        .B2(n15874), .ZN(n10180) );
  INV_X1 U12022 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12729) );
  INV_X1 U12023 ( .A(n10182), .ZN(n10195) );
  NAND2_X1 U12024 ( .A1(n10183), .A2(n15867), .ZN(n10184) );
  NAND2_X1 U12025 ( .A1(n10195), .A2(n10184), .ZN(n13160) );
  OR2_X1 U12026 ( .A1(n13160), .A2(n9999), .ZN(n10186) );
  AOI22_X1 U12027 ( .A1(n10682), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n10683), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n10185) );
  OAI211_X1 U12028 ( .C1(n10877), .C2(n12729), .A(n10186), .B(n10185), .ZN(
        n14374) );
  XNOR2_X1 U12029 ( .A(n14720), .B(n14374), .ZN(n13085) );
  INV_X1 U12030 ( .A(n13085), .ZN(n13089) );
  NAND2_X1 U12031 ( .A1(n14720), .A2(n14374), .ZN(n10187) );
  NAND2_X1 U12032 ( .A1(n12063), .A2(n10871), .ZN(n10193) );
  NAND2_X1 U12033 ( .A1(n7560), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10188) );
  MUX2_X1 U12034 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10188), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n10190) );
  NAND2_X1 U12035 ( .A1(n10190), .A2(n10213), .ZN(n13105) );
  OAI22_X1 U12036 ( .A1(n10873), .A2(n12066), .B1(n11300), .B2(n13105), .ZN(
        n10191) );
  INV_X1 U12037 ( .A(n10191), .ZN(n10192) );
  INV_X1 U12038 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13100) );
  INV_X1 U12039 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U12040 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  NAND2_X1 U12041 ( .A1(n10203), .A2(n10196), .ZN(n14639) );
  OR2_X1 U12042 ( .A1(n14639), .A2(n9999), .ZN(n10198) );
  AOI22_X1 U12043 ( .A1(n10682), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n10683), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n10197) );
  OAI211_X1 U12044 ( .C1(n10877), .C2(n13100), .A(n10198), .B(n10197), .ZN(
        n14373) );
  XNOR2_X1 U12045 ( .A(n14716), .B(n14373), .ZN(n14632) );
  INV_X1 U12046 ( .A(n14632), .ZN(n14636) );
  INV_X1 U12047 ( .A(n14625), .ZN(n10211) );
  NAND2_X1 U12048 ( .A1(n10213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10199) );
  XNOR2_X1 U12049 ( .A(n10199), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15885) );
  AOI22_X1 U12050 ( .A1(n10005), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n15885), 
        .B2(n10215), .ZN(n10200) );
  NAND2_X1 U12051 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  AND2_X1 U12052 ( .A1(n10220), .A2(n10204), .ZN(n14619) );
  NAND2_X1 U12053 ( .A1(n14619), .A2(n10375), .ZN(n10209) );
  INV_X1 U12054 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15882) );
  NAND2_X1 U12055 ( .A1(n10682), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U12056 ( .A1(n10683), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n10205) );
  OAI211_X1 U12057 ( .C1(n15882), .C2(n10877), .A(n10206), .B(n10205), .ZN(
        n10207) );
  INV_X1 U12058 ( .A(n10207), .ZN(n10208) );
  NAND2_X1 U12059 ( .A1(n10209), .A2(n10208), .ZN(n14372) );
  XNOR2_X1 U12060 ( .A(n14710), .B(n14372), .ZN(n14626) );
  INV_X1 U12061 ( .A(n14626), .ZN(n10210) );
  OR2_X1 U12062 ( .A1(n14710), .A2(n14372), .ZN(n10212) );
  NAND2_X1 U12063 ( .A1(n12537), .A2(n10871), .ZN(n10217) );
  XNOR2_X2 U12064 ( .A(n10214), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U12065 ( .A1(n10696), .A2(n10215), .B1(n10005), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n10216) );
  INV_X1 U12066 ( .A(n10218), .ZN(n10231) );
  NAND2_X1 U12067 ( .A1(n10220), .A2(n10219), .ZN(n10221) );
  NAND2_X1 U12068 ( .A1(n10231), .A2(n10221), .ZN(n14595) );
  OR2_X1 U12069 ( .A1(n14595), .A2(n9999), .ZN(n10226) );
  INV_X1 U12070 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U12071 ( .A1(n10682), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U12072 ( .A1(n10683), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n10222) );
  OAI211_X1 U12073 ( .C1(n14596), .C2(n10877), .A(n10223), .B(n10222), .ZN(
        n10224) );
  INV_X1 U12074 ( .A(n10224), .ZN(n10225) );
  NAND2_X1 U12075 ( .A1(n10226), .A2(n10225), .ZN(n14579) );
  XNOR2_X1 U12076 ( .A(n14594), .B(n14579), .ZN(n14600) );
  INV_X1 U12077 ( .A(n14600), .ZN(n14592) );
  NAND2_X1 U12078 ( .A1(n12666), .A2(n10871), .ZN(n10228) );
  OR2_X1 U12079 ( .A1(n10873), .A2(n8795), .ZN(n10227) );
  INV_X1 U12080 ( .A(n10229), .ZN(n10245) );
  INV_X1 U12081 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U12082 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  AND2_X1 U12083 ( .A1(n10245), .A2(n10232), .ZN(n14584) );
  NAND2_X1 U12084 ( .A1(n14584), .A2(n10375), .ZN(n10238) );
  INV_X1 U12085 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U12086 ( .A1(n10683), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U12087 ( .A1(n10682), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n10233) );
  OAI211_X1 U12088 ( .C1(n10235), .C2(n10877), .A(n10234), .B(n10233), .ZN(
        n10236) );
  INV_X1 U12089 ( .A(n10236), .ZN(n10237) );
  INV_X1 U12090 ( .A(n14605), .ZN(n14371) );
  OR2_X1 U12091 ( .A1(n14698), .A2(n14371), .ZN(n10239) );
  NAND2_X1 U12092 ( .A1(n14581), .A2(n10239), .ZN(n10241) );
  NAND2_X1 U12093 ( .A1(n14698), .A2(n14371), .ZN(n10240) );
  NAND2_X1 U12094 ( .A1(n10241), .A2(n10240), .ZN(n14569) );
  NAND2_X1 U12095 ( .A1(n12806), .A2(n10871), .ZN(n10243) );
  OR2_X1 U12096 ( .A1(n10873), .A2(n12807), .ZN(n10242) );
  INV_X1 U12097 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U12098 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  NAND2_X1 U12099 ( .A1(n10255), .A2(n10246), .ZN(n14564) );
  OR2_X1 U12100 ( .A1(n14564), .A2(n9999), .ZN(n10251) );
  INV_X1 U12101 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U12102 ( .A1(n10682), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U12103 ( .A1(n10683), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n10247) );
  OAI211_X1 U12104 ( .C1(n14565), .C2(n10877), .A(n10248), .B(n10247), .ZN(
        n10249) );
  INV_X1 U12105 ( .A(n10249), .ZN(n10250) );
  NAND2_X1 U12106 ( .A1(n10251), .A2(n10250), .ZN(n14576) );
  XNOR2_X1 U12107 ( .A(n14566), .B(n14576), .ZN(n14570) );
  OAI22_X1 U12108 ( .A1(n14569), .A2(n14570), .B1(n14566), .B2(n14576), .ZN(
        n14548) );
  XNOR2_X1 U12109 ( .A(n9656), .B(n10252), .ZN(n13037) );
  NAND2_X1 U12110 ( .A1(n13037), .A2(n10871), .ZN(n10254) );
  OR2_X1 U12111 ( .A1(n10873), .A2(n13039), .ZN(n10253) );
  NAND2_X1 U12112 ( .A1(n10255), .A2(n14344), .ZN(n10256) );
  AND2_X1 U12113 ( .A1(n10266), .A2(n10256), .ZN(n14552) );
  NAND2_X1 U12114 ( .A1(n14552), .A2(n10375), .ZN(n10262) );
  INV_X1 U12115 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12116 ( .A1(n10682), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U12117 ( .A1(n10683), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n10257) );
  OAI211_X1 U12118 ( .C1(n10259), .C2(n10877), .A(n10258), .B(n10257), .ZN(
        n10260) );
  INV_X1 U12119 ( .A(n10260), .ZN(n10261) );
  NAND2_X1 U12120 ( .A1(n10262), .A2(n10261), .ZN(n14370) );
  NAND2_X1 U12121 ( .A1(n14551), .A2(n14370), .ZN(n10263) );
  NAND2_X1 U12122 ( .A1(n13000), .A2(n10871), .ZN(n10265) );
  OR2_X1 U12123 ( .A1(n10873), .A2(n13003), .ZN(n10264) );
  NAND2_X1 U12124 ( .A1(n10266), .A2(n14273), .ZN(n10267) );
  NAND2_X1 U12125 ( .A1(n10268), .A2(n10267), .ZN(n14529) );
  OR2_X1 U12126 ( .A1(n14529), .A2(n9999), .ZN(n10273) );
  INV_X1 U12127 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14528) );
  NAND2_X1 U12128 ( .A1(n10683), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U12129 ( .A1(n10682), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n10269) );
  OAI211_X1 U12130 ( .C1(n14528), .C2(n10877), .A(n10270), .B(n10269), .ZN(
        n10271) );
  INV_X1 U12131 ( .A(n10271), .ZN(n10272) );
  XNOR2_X1 U12132 ( .A(n14527), .B(n14512), .ZN(n14532) );
  NAND2_X1 U12133 ( .A1(n14523), .A2(n14532), .ZN(n10275) );
  NAND2_X1 U12134 ( .A1(n14527), .A2(n14369), .ZN(n10274) );
  NAND2_X1 U12135 ( .A1(n14789), .A2(n10871), .ZN(n10277) );
  OR2_X1 U12136 ( .A1(n10873), .A2(n14791), .ZN(n10276) );
  INV_X1 U12137 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U12138 ( .A1(n10279), .A2(n10278), .ZN(n10280) );
  NAND2_X1 U12139 ( .A1(n10289), .A2(n10280), .ZN(n14500) );
  OR2_X1 U12140 ( .A1(n14500), .A2(n9999), .ZN(n10285) );
  INV_X1 U12141 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n14499) );
  NAND2_X1 U12142 ( .A1(n10682), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12143 ( .A1(n10683), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10281) );
  OAI211_X1 U12144 ( .C1(n14499), .C2(n10877), .A(n10282), .B(n10281), .ZN(
        n10283) );
  INV_X1 U12145 ( .A(n10283), .ZN(n10284) );
  NAND2_X1 U12146 ( .A1(n10285), .A2(n10284), .ZN(n14368) );
  XNOR2_X1 U12147 ( .A(n14498), .B(n14368), .ZN(n14490) );
  NAND2_X1 U12148 ( .A1(n14786), .A2(n10871), .ZN(n10288) );
  OR2_X1 U12149 ( .A1(n10873), .A2(n14787), .ZN(n10287) );
  INV_X1 U12150 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n14354) );
  NAND2_X1 U12151 ( .A1(n10289), .A2(n14354), .ZN(n10290) );
  NAND2_X1 U12152 ( .A1(n14481), .A2(n10375), .ZN(n10296) );
  INV_X1 U12153 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12154 ( .A1(n10683), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U12155 ( .A1(n10682), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n10291) );
  OAI211_X1 U12156 ( .C1(n10293), .C2(n10877), .A(n10292), .B(n10291), .ZN(
        n10294) );
  INV_X1 U12157 ( .A(n10294), .ZN(n10295) );
  INV_X1 U12158 ( .A(n14493), .ZN(n14312) );
  NAND2_X1 U12159 ( .A1(n14783), .A2(n10871), .ZN(n10298) );
  OR2_X1 U12160 ( .A1(n10873), .A2(n14785), .ZN(n10297) );
  XNOR2_X1 U12161 ( .A(n10310), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U12162 ( .A1(n14468), .A2(n10375), .ZN(n10304) );
  INV_X1 U12163 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U12164 ( .A1(n10683), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U12165 ( .A1(n10682), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n10299) );
  OAI211_X1 U12166 ( .C1(n10301), .C2(n10877), .A(n10300), .B(n10299), .ZN(
        n10302) );
  INV_X1 U12167 ( .A(n10302), .ZN(n10303) );
  XNOR2_X1 U12168 ( .A(n14467), .B(n14367), .ZN(n14463) );
  INV_X1 U12169 ( .A(n14463), .ZN(n14460) );
  NAND2_X1 U12170 ( .A1(n15796), .A2(n10871), .ZN(n10306) );
  OR2_X1 U12171 ( .A1(n10873), .A2(n14782), .ZN(n10305) );
  NAND2_X1 U12172 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n10307) );
  NOR2_X1 U12173 ( .A1(n10310), .A2(n10307), .ZN(n10689) );
  INV_X1 U12174 ( .A(n10689), .ZN(n10312) );
  INV_X1 U12175 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10309) );
  INV_X1 U12176 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10308) );
  OAI21_X1 U12177 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(n10311) );
  NAND2_X1 U12178 ( .A1(n10312), .A2(n10311), .ZN(n14451) );
  INV_X1 U12179 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14450) );
  NAND2_X1 U12180 ( .A1(n10682), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U12181 ( .A1(n10683), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10313) );
  OAI211_X1 U12182 ( .C1(n14450), .C2(n10877), .A(n10314), .B(n10313), .ZN(
        n10315) );
  INV_X1 U12183 ( .A(n10315), .ZN(n10316) );
  OR2_X1 U12184 ( .A1(n14453), .A2(n10920), .ZN(n10676) );
  NAND2_X1 U12185 ( .A1(n14453), .A2(n10920), .ZN(n10318) );
  NAND2_X1 U12186 ( .A1(n10676), .A2(n10318), .ZN(n10865) );
  XNOR2_X1 U12187 ( .A(n10665), .B(n10865), .ZN(n14454) );
  INV_X1 U12188 ( .A(n10323), .ZN(n10322) );
  NAND2_X1 U12189 ( .A1(n10323), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U12190 ( .A1(n10325), .A2(n10324), .ZN(n10331) );
  XNOR2_X2 U12191 ( .A(n10327), .B(n10326), .ZN(n10695) );
  XNOR2_X1 U12192 ( .A(n10901), .B(n10695), .ZN(n10328) );
  OR2_X1 U12193 ( .A1(n11852), .A2(n10948), .ZN(n12148) );
  INV_X1 U12194 ( .A(n14698), .ZN(n14587) );
  NAND2_X1 U12195 ( .A1(n12271), .A2(n11672), .ZN(n11683) );
  OR2_X1 U12196 ( .A1(n11683), .A2(n12045), .ZN(n11684) );
  INV_X1 U12197 ( .A(n12088), .ZN(n12153) );
  INV_X1 U12198 ( .A(n12451), .ZN(n10330) );
  NAND2_X1 U12199 ( .A1(n12646), .A2(n10330), .ZN(n12450) );
  INV_X1 U12200 ( .A(n12863), .ZN(n12882) );
  OR2_X1 U12201 ( .A1(n14710), .A2(n14643), .ZN(n14617) );
  AOI21_X1 U12202 ( .B1(n14465), .B2(n14453), .A(n11533), .ZN(n10332) );
  INV_X1 U12203 ( .A(n11614), .ZN(n10343) );
  OR2_X1 U12204 ( .A1(n11492), .A2(n14387), .ZN(n11665) );
  INV_X1 U12205 ( .A(n11665), .ZN(n10334) );
  INV_X1 U12206 ( .A(n11668), .ZN(n12054) );
  OR2_X1 U12207 ( .A1(n7435), .A2(n12054), .ZN(n10335) );
  NAND2_X1 U12208 ( .A1(n10336), .A2(n10335), .ZN(n11676) );
  NAND2_X1 U12209 ( .A1(n11676), .A2(n10849), .ZN(n10339) );
  NAND2_X1 U12210 ( .A1(n10337), .A2(n11679), .ZN(n10338) );
  INV_X1 U12211 ( .A(n14384), .ZN(n10340) );
  NAND2_X1 U12212 ( .A1(n12045), .A2(n10340), .ZN(n10341) );
  NAND2_X1 U12213 ( .A1(n10342), .A2(n10341), .ZN(n11613) );
  NAND2_X1 U12214 ( .A1(n11612), .A2(n11647), .ZN(n10344) );
  AND2_X1 U12215 ( .A1(n11701), .A2(n11656), .ZN(n10345) );
  NAND2_X1 U12216 ( .A1(n12071), .A2(n14382), .ZN(n10346) );
  INV_X1 U12217 ( .A(n14381), .ZN(n12079) );
  INV_X1 U12218 ( .A(n12082), .ZN(n10347) );
  NOR2_X1 U12219 ( .A1(n12088), .A2(n12247), .ZN(n12127) );
  NOR2_X1 U12220 ( .A1(n10855), .A2(n12127), .ZN(n10349) );
  INV_X1 U12221 ( .A(n14379), .ZN(n12475) );
  NAND2_X1 U12222 ( .A1(n7849), .A2(n12475), .ZN(n12372) );
  INV_X1 U12223 ( .A(n14378), .ZN(n12784) );
  NAND2_X1 U12224 ( .A1(n12644), .A2(n12784), .ZN(n10352) );
  OR2_X1 U12225 ( .A1(n12770), .A2(n12772), .ZN(n10353) );
  NAND2_X1 U12226 ( .A1(n12863), .A2(n12864), .ZN(n10354) );
  OR2_X1 U12227 ( .A1(n16600), .A2(n12931), .ZN(n10355) );
  INV_X1 U12228 ( .A(n14374), .ZN(n10358) );
  OR2_X1 U12229 ( .A1(n14720), .A2(n10358), .ZN(n10359) );
  NAND2_X1 U12230 ( .A1(n13084), .A2(n10359), .ZN(n14630) );
  NAND2_X1 U12231 ( .A1(n14630), .A2(n14632), .ZN(n14631) );
  INV_X1 U12232 ( .A(n14373), .ZN(n13196) );
  OR2_X1 U12233 ( .A1(n14716), .A2(n13196), .ZN(n10360) );
  INV_X1 U12234 ( .A(n14372), .ZN(n14603) );
  INV_X1 U12235 ( .A(n14579), .ZN(n13197) );
  NAND2_X1 U12236 ( .A1(n14594), .A2(n13197), .ZN(n10363) );
  NAND2_X1 U12237 ( .A1(n14698), .A2(n14605), .ZN(n10846) );
  INV_X1 U12238 ( .A(n10846), .ZN(n10364) );
  OR2_X1 U12239 ( .A1(n14698), .A2(n14605), .ZN(n10847) );
  INV_X1 U12240 ( .A(n14576), .ZN(n14343) );
  INV_X1 U12241 ( .A(n14370), .ZN(n14534) );
  INV_X1 U12242 ( .A(n14492), .ZN(n14535) );
  INV_X1 U12243 ( .A(n14368), .ZN(n14513) );
  INV_X1 U12244 ( .A(n14367), .ZN(n14266) );
  INV_X1 U12245 ( .A(n10865), .ZN(n10372) );
  NAND2_X1 U12246 ( .A1(n10948), .A2(n10696), .ZN(n10371) );
  NOR2_X1 U12247 ( .A1(n10331), .A2(n10329), .ZN(n10884) );
  INV_X1 U12248 ( .A(n10884), .ZN(n10370) );
  OAI211_X1 U12249 ( .C1(n10373), .C2(n10372), .A(n10677), .B(n16584), .ZN(
        n10383) );
  INV_X1 U12250 ( .A(n11308), .ZN(n10374) );
  NAND2_X1 U12251 ( .A1(n10689), .A2(n10375), .ZN(n10382) );
  INV_X1 U12252 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U12253 ( .A1(n10376), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U12254 ( .A1(n10683), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10377) );
  OAI211_X1 U12255 ( .C1(n10379), .C2(n10876), .A(n10378), .B(n10377), .ZN(
        n10380) );
  INV_X1 U12256 ( .A(n10380), .ZN(n10381) );
  NAND2_X1 U12257 ( .A1(n10382), .A2(n10381), .ZN(n14365) );
  AOI22_X1 U12258 ( .A1(n14367), .A2(n14578), .B1(n14365), .B2(n14575), .ZN(
        n14298) );
  NAND2_X1 U12259 ( .A1(n10394), .A2(n10393), .ZN(n10387) );
  XNOR2_X1 U12260 ( .A(P2_B_REG_SCAN_IN), .B(n13204), .ZN(n10395) );
  AND2_X1 U12261 ( .A1(n14790), .A2(n10395), .ZN(n10396) );
  INV_X1 U12262 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15817) );
  AOI22_X1 U12263 ( .A1(n15818), .A2(n15817), .B1(n14788), .B2(n14790), .ZN(
        n10670) );
  NAND2_X1 U12264 ( .A1(n10397), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10399) );
  INV_X1 U12265 ( .A(n10953), .ZN(n11510) );
  AND2_X1 U12266 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11510), .ZN(n10400) );
  NOR4_X1 U12267 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10404) );
  NOR4_X1 U12268 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10403) );
  NOR4_X1 U12269 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10402) );
  NOR4_X1 U12270 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10401) );
  NAND4_X1 U12271 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10410) );
  NOR2_X1 U12272 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n10408) );
  NOR4_X1 U12273 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10407) );
  NOR4_X1 U12274 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10406) );
  NOR4_X1 U12275 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U12276 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10409) );
  OAI21_X1 U12277 ( .B1(n10410), .B2(n10409), .A(n15818), .ZN(n10669) );
  NAND2_X1 U12278 ( .A1(n10946), .A2(n11501), .ZN(n11512) );
  OR2_X1 U12279 ( .A1(n11852), .A2(n11491), .ZN(n11508) );
  NAND3_X1 U12280 ( .A1(n10669), .A2(n11512), .A3(n11508), .ZN(n10411) );
  NAND2_X1 U12281 ( .A1(n14788), .A2(n13204), .ZN(n10412) );
  INV_X1 U12282 ( .A(n15822), .ZN(n10414) );
  OR2_X1 U12283 ( .A1(n14733), .A2(n16589), .ZN(n10420) );
  INV_X1 U12284 ( .A(n11491), .ZN(n10415) );
  INV_X1 U12285 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10416) );
  NOR2_X1 U12286 ( .A1(n16591), .A2(n10416), .ZN(n10417) );
  NAND2_X1 U12287 ( .A1(n10420), .A2(n10419), .ZN(P2_U3527) );
  NAND2_X1 U12288 ( .A1(n9044), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10421) );
  INV_X1 U12289 ( .A(n13541), .ZN(n10425) );
  NAND2_X1 U12290 ( .A1(n14211), .A2(n10425), .ZN(n10428) );
  NAND2_X1 U12291 ( .A1(n12413), .A2(n13736), .ZN(n10426) );
  NAND2_X1 U12292 ( .A1(n10426), .A2(n12192), .ZN(n10427) );
  XNOR2_X1 U12293 ( .A(n10431), .B(n12330), .ZN(n13579) );
  OR2_X1 U12294 ( .A1(n12443), .A2(n10507), .ZN(n10430) );
  AND2_X1 U12295 ( .A1(n12393), .A2(n10430), .ZN(n13580) );
  NAND2_X1 U12296 ( .A1(n13579), .A2(n13580), .ZN(n13578) );
  INV_X1 U12297 ( .A(n10431), .ZN(n10432) );
  NAND2_X1 U12298 ( .A1(n12330), .A2(n10432), .ZN(n10433) );
  NAND2_X1 U12299 ( .A1(n13578), .A2(n10433), .ZN(n11917) );
  XNOR2_X1 U12300 ( .A(n11919), .B(n10507), .ZN(n10434) );
  XNOR2_X1 U12301 ( .A(n10434), .B(n13582), .ZN(n11918) );
  NAND2_X1 U12302 ( .A1(n11917), .A2(n11918), .ZN(n10437) );
  INV_X1 U12303 ( .A(n10434), .ZN(n10435) );
  NAND2_X1 U12304 ( .A1(n10435), .A2(n13582), .ZN(n10436) );
  NAND2_X1 U12305 ( .A1(n10437), .A2(n10436), .ZN(n12322) );
  INV_X1 U12306 ( .A(n12322), .ZN(n10440) );
  INV_X4 U12307 ( .A(n10507), .ZN(n13236) );
  XNOR2_X1 U12308 ( .A(n12560), .B(n13236), .ZN(n10441) );
  XNOR2_X1 U12309 ( .A(n10441), .B(n10438), .ZN(n12323) );
  INV_X1 U12310 ( .A(n10441), .ZN(n10442) );
  NAND2_X1 U12311 ( .A1(n13713), .A2(n10442), .ZN(n10443) );
  XNOR2_X1 U12312 ( .A(n13379), .B(n13236), .ZN(n10444) );
  XNOR2_X1 U12313 ( .A(n10444), .B(n13712), .ZN(n12387) );
  INV_X1 U12314 ( .A(n10444), .ZN(n10445) );
  NAND2_X1 U12315 ( .A1(n12531), .A2(n10445), .ZN(n10446) );
  XNOR2_X1 U12316 ( .A(n12670), .B(n10507), .ZN(n10447) );
  XNOR2_X1 U12317 ( .A(n10447), .B(n12850), .ZN(n12530) );
  INV_X1 U12318 ( .A(n10447), .ZN(n10448) );
  AND2_X1 U12319 ( .A1(n10448), .A2(n12850), .ZN(n10449) );
  XNOR2_X1 U12320 ( .A(n16406), .B(n13236), .ZN(n10450) );
  XNOR2_X1 U12321 ( .A(n10450), .B(n13392), .ZN(n12519) );
  NAND2_X1 U12322 ( .A1(n12520), .A2(n12519), .ZN(n12518) );
  NAND2_X1 U12323 ( .A1(n10450), .A2(n13709), .ZN(n10451) );
  NAND2_X1 U12324 ( .A1(n12518), .A2(n10451), .ZN(n12660) );
  XNOR2_X1 U12325 ( .A(n12663), .B(n10507), .ZN(n10455) );
  XNOR2_X1 U12326 ( .A(n10455), .B(n12988), .ZN(n12659) );
  XNOR2_X1 U12327 ( .A(n12991), .B(n13236), .ZN(n10453) );
  XNOR2_X1 U12328 ( .A(n10453), .B(n13707), .ZN(n12793) );
  AND2_X1 U12329 ( .A1(n12659), .A2(n12793), .ZN(n10452) );
  NAND2_X1 U12330 ( .A1(n12660), .A2(n10452), .ZN(n12821) );
  XNOR2_X1 U12331 ( .A(n12828), .B(n13236), .ZN(n10461) );
  XNOR2_X1 U12332 ( .A(n10461), .B(n13075), .ZN(n12825) );
  INV_X1 U12333 ( .A(n12825), .ZN(n10459) );
  INV_X1 U12334 ( .A(n10453), .ZN(n10454) );
  NAND2_X1 U12335 ( .A1(n10454), .A2(n13707), .ZN(n10458) );
  INV_X1 U12336 ( .A(n12793), .ZN(n10457) );
  INV_X1 U12337 ( .A(n10455), .ZN(n10456) );
  OR2_X1 U12338 ( .A1(n12988), .A2(n10456), .ZN(n12789) );
  OR2_X1 U12339 ( .A1(n10457), .A2(n12789), .ZN(n12791) );
  AND2_X1 U12340 ( .A1(n10458), .A2(n12791), .ZN(n12820) );
  AND2_X1 U12341 ( .A1(n10459), .A2(n12820), .ZN(n10460) );
  NAND2_X1 U12342 ( .A1(n10461), .A2(n13075), .ZN(n10462) );
  XNOR2_X1 U12343 ( .A(n12901), .B(n13236), .ZN(n10463) );
  XNOR2_X1 U12344 ( .A(n10463), .B(n14086), .ZN(n12895) );
  OR2_X1 U12345 ( .A1(n14086), .A2(n10463), .ZN(n10464) );
  NAND2_X1 U12346 ( .A1(n12897), .A2(n10464), .ZN(n12946) );
  INV_X1 U12347 ( .A(n12946), .ZN(n10473) );
  XNOR2_X1 U12348 ( .A(n14053), .B(n10507), .ZN(n13551) );
  XNOR2_X1 U12349 ( .A(n14077), .B(n13236), .ZN(n10467) );
  NAND2_X1 U12350 ( .A1(n10467), .A2(n14088), .ZN(n10466) );
  XNOR2_X1 U12351 ( .A(n14091), .B(n13236), .ZN(n12947) );
  NAND3_X1 U12352 ( .A1(n13551), .A2(n10466), .A3(n12947), .ZN(n10472) );
  INV_X1 U12353 ( .A(n12947), .ZN(n10465) );
  NAND2_X1 U12354 ( .A1(n10465), .A2(n13706), .ZN(n13552) );
  INV_X1 U12355 ( .A(n10466), .ZN(n13659) );
  INV_X1 U12356 ( .A(n10467), .ZN(n10468) );
  NAND2_X1 U12357 ( .A1(n10468), .A2(n13656), .ZN(n13554) );
  OAI211_X1 U12358 ( .C1(n13552), .C2(n13659), .A(n13551), .B(n13554), .ZN(
        n10469) );
  OAI21_X1 U12359 ( .B1(n13551), .B2(n14036), .A(n10469), .ZN(n10470) );
  XNOR2_X1 U12360 ( .A(n16534), .B(n13236), .ZN(n10474) );
  XNOR2_X1 U12361 ( .A(n10474), .B(n14055), .ZN(n13556) );
  AND2_X1 U12362 ( .A1(n10470), .A2(n13556), .ZN(n10471) );
  NAND2_X1 U12363 ( .A1(n13555), .A2(n10475), .ZN(n13131) );
  XNOR2_X1 U12364 ( .A(n16610), .B(n13236), .ZN(n13132) );
  NAND2_X1 U12365 ( .A1(n13132), .A2(n13625), .ZN(n10477) );
  INV_X1 U12366 ( .A(n13132), .ZN(n10476) );
  XNOR2_X1 U12367 ( .A(n14208), .B(n13236), .ZN(n10478) );
  XNOR2_X1 U12368 ( .A(n10478), .B(n14028), .ZN(n13622) );
  NAND2_X1 U12369 ( .A1(n13623), .A2(n13622), .ZN(n13621) );
  INV_X1 U12370 ( .A(n10478), .ZN(n10479) );
  NAND2_X1 U12371 ( .A1(n13621), .A2(n8386), .ZN(n13632) );
  XNOR2_X1 U12372 ( .A(n13449), .B(n13236), .ZN(n10480) );
  XNOR2_X1 U12373 ( .A(n10480), .B(n13705), .ZN(n13631) );
  NAND2_X1 U12374 ( .A1(n13632), .A2(n13631), .ZN(n13630) );
  XNOR2_X1 U12375 ( .A(n14199), .B(n13236), .ZN(n10482) );
  XNOR2_X1 U12376 ( .A(n10482), .B(n13946), .ZN(n13678) );
  NAND2_X1 U12377 ( .A1(n10482), .A2(n13985), .ZN(n10483) );
  XNOR2_X1 U12378 ( .A(n13570), .B(n13236), .ZN(n10484) );
  XNOR2_X1 U12379 ( .A(n10484), .B(n13704), .ZN(n13573) );
  XNOR2_X1 U12380 ( .A(n13940), .B(n13236), .ZN(n10485) );
  XNOR2_X1 U12381 ( .A(n10485), .B(n13915), .ZN(n13648) );
  NAND2_X1 U12382 ( .A1(n13649), .A2(n13648), .ZN(n13647) );
  INV_X1 U12383 ( .A(n10485), .ZN(n10486) );
  NAND2_X1 U12384 ( .A1(n13647), .A2(n10487), .ZN(n13592) );
  MUX2_X1 U12385 ( .A(n10488), .B(n13463), .S(n13236), .Z(n13591) );
  INV_X1 U12386 ( .A(n13591), .ZN(n10490) );
  XNOR2_X1 U12387 ( .A(n13921), .B(n13236), .ZN(n10489) );
  NAND2_X1 U12388 ( .A1(n10489), .A2(n13933), .ZN(n13590) );
  OAI21_X1 U12389 ( .B1(n13592), .B2(n10490), .A(n13590), .ZN(n10492) );
  XNOR2_X1 U12390 ( .A(n13903), .B(n13236), .ZN(n10491) );
  NAND2_X1 U12391 ( .A1(n10492), .A2(n10491), .ZN(n10493) );
  OAI21_X1 U12392 ( .B1(n10492), .B2(n10491), .A(n10493), .ZN(n13668) );
  XOR2_X1 U12393 ( .A(n13236), .B(n13563), .Z(n10495) );
  NAND2_X1 U12394 ( .A1(n13564), .A2(n13897), .ZN(n13640) );
  INV_X1 U12395 ( .A(n10496), .ZN(n13639) );
  XNOR2_X1 U12396 ( .A(n13637), .B(n13236), .ZN(n10497) );
  NAND2_X1 U12397 ( .A1(n10497), .A2(n13859), .ZN(n10500) );
  INV_X1 U12398 ( .A(n10497), .ZN(n10498) );
  NAND2_X1 U12399 ( .A1(n10498), .A2(n13884), .ZN(n10499) );
  NAND2_X1 U12400 ( .A1(n10500), .A2(n10499), .ZN(n13638) );
  INV_X1 U12401 ( .A(n10500), .ZN(n13612) );
  XNOR2_X1 U12402 ( .A(n14164), .B(n13236), .ZN(n10501) );
  NAND2_X1 U12403 ( .A1(n10501), .A2(n13838), .ZN(n10504) );
  INV_X1 U12404 ( .A(n10501), .ZN(n10502) );
  NAND2_X1 U12405 ( .A1(n10502), .A2(n13870), .ZN(n10503) );
  AND2_X1 U12406 ( .A1(n10504), .A2(n10503), .ZN(n13611) );
  XNOR2_X1 U12407 ( .A(n13686), .B(n10507), .ZN(n10505) );
  NOR2_X1 U12408 ( .A1(n10505), .A2(n13857), .ZN(n10506) );
  AOI21_X1 U12409 ( .B1(n10505), .B2(n13857), .A(n10506), .ZN(n13689) );
  INV_X1 U12410 ( .A(n10506), .ZN(n13232) );
  NAND2_X1 U12411 ( .A1(n13687), .A2(n13232), .ZN(n10509) );
  XNOR2_X1 U12412 ( .A(n8915), .B(n10507), .ZN(n10508) );
  NOR2_X1 U12413 ( .A1(n10508), .A2(n13702), .ZN(n13231) );
  AOI21_X1 U12414 ( .B1(n10508), .B2(n13702), .A(n13231), .ZN(n13234) );
  XNOR2_X1 U12415 ( .A(n10509), .B(n13234), .ZN(n10513) );
  NAND3_X1 U12416 ( .A1(n10525), .A2(n10510), .A3(n16609), .ZN(n10511) );
  OAI21_X1 U12417 ( .B1(n10521), .B2(n10519), .A(n10511), .ZN(n10512) );
  NAND2_X1 U12418 ( .A1(n10513), .A2(n13690), .ZN(n10537) );
  INV_X1 U12419 ( .A(n8915), .ZN(n13833) );
  NAND3_X1 U12420 ( .A1(n10525), .A2(n14105), .A3(n11722), .ZN(n10515) );
  INV_X1 U12421 ( .A(n16333), .ZN(n12397) );
  INV_X1 U12422 ( .A(n13673), .ZN(n13700) );
  INV_X1 U12423 ( .A(n11893), .ZN(n10516) );
  NAND2_X1 U12424 ( .A1(n11722), .A2(n10516), .ZN(n13543) );
  NOR2_X1 U12425 ( .A1(n13543), .A2(n10521), .ZN(n10530) );
  INV_X1 U12426 ( .A(n13671), .ZN(n13697) );
  INV_X1 U12427 ( .A(n13831), .ZN(n10532) );
  INV_X1 U12428 ( .A(n13543), .ZN(n10518) );
  OR2_X1 U12429 ( .A1(n11723), .A2(P3_U3151), .ZN(n13547) );
  INV_X1 U12430 ( .A(n13547), .ZN(n11721) );
  AOI21_X1 U12431 ( .B1(n10518), .B2(n10521), .A(n11721), .ZN(n10528) );
  INV_X1 U12432 ( .A(n10519), .ZN(n10520) );
  NAND2_X1 U12433 ( .A1(n10521), .A2(n10520), .ZN(n10523) );
  AND2_X1 U12434 ( .A1(n12398), .A2(n10955), .ZN(n10522) );
  OAI211_X1 U12435 ( .C1(n10525), .C2(n10524), .A(n10523), .B(n10522), .ZN(
        n10526) );
  NAND2_X1 U12436 ( .A1(n10526), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10527) );
  AOI22_X1 U12437 ( .A1(n13857), .A2(n13692), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10531) );
  OAI21_X1 U12438 ( .B1(n10532), .B2(n13694), .A(n10531), .ZN(n10533) );
  AOI21_X1 U12439 ( .B1(n13829), .B2(n13697), .A(n10533), .ZN(n10534) );
  NAND2_X1 U12440 ( .A1(n10537), .A2(n10536), .ZN(P3_U3154) );
  INV_X1 U12441 ( .A(n16349), .ZN(n10540) );
  NAND2_X1 U12442 ( .A1(n16350), .A2(n10540), .ZN(n10542) );
  NAND2_X1 U12443 ( .A1(n10542), .A2(n10541), .ZN(n12027) );
  NAND2_X1 U12444 ( .A1(n12027), .A2(n12036), .ZN(n10544) );
  NAND2_X1 U12445 ( .A1(n11992), .A2(n12178), .ZN(n10545) );
  INV_X1 U12446 ( .A(n12179), .ZN(n12176) );
  NAND2_X1 U12447 ( .A1(n12189), .A2(n12166), .ZN(n10546) );
  OR2_X1 U12448 ( .A1(n12236), .A2(n12570), .ZN(n10548) );
  NAND2_X1 U12449 ( .A1(n12165), .A2(n10548), .ZN(n12220) );
  INV_X1 U12450 ( .A(n12221), .ZN(n10549) );
  NAND2_X1 U12451 ( .A1(n12220), .A2(n10549), .ZN(n10551) );
  OR2_X1 U12452 ( .A1(n12573), .A2(n12888), .ZN(n10550) );
  INV_X1 U12453 ( .A(n12197), .ZN(n12195) );
  INV_X1 U12454 ( .A(n14935), .ZN(n12925) );
  INV_X1 U12455 ( .A(n14934), .ZN(n12887) );
  OR2_X1 U12456 ( .A1(n12928), .A2(n12887), .ZN(n10552) );
  NAND2_X1 U12457 ( .A1(n10554), .A2(n14933), .ZN(n10553) );
  NAND2_X1 U12458 ( .A1(n10553), .A2(n12614), .ZN(n10556) );
  INV_X1 U12459 ( .A(n14933), .ZN(n12924) );
  NAND2_X1 U12460 ( .A1(n12615), .A2(n12924), .ZN(n10555) );
  NAND2_X1 U12461 ( .A1(n10556), .A2(n10555), .ZN(n12552) );
  INV_X1 U12462 ( .A(n12552), .ZN(n10557) );
  OR2_X1 U12463 ( .A1(n12813), .A2(n13173), .ZN(n10558) );
  NAND2_X1 U12464 ( .A1(n13176), .A2(n16544), .ZN(n10559) );
  OR2_X1 U12465 ( .A1(n16561), .A2(n13172), .ZN(n10561) );
  NAND2_X1 U12466 ( .A1(n12965), .A2(n10561), .ZN(n16620) );
  INV_X1 U12467 ( .A(n14929), .ZN(n16541) );
  OR2_X1 U12468 ( .A1(n11055), .A2(n16541), .ZN(n10562) );
  INV_X1 U12469 ( .A(n14928), .ZN(n10564) );
  NAND2_X1 U12470 ( .A1(n15762), .A2(n10564), .ZN(n10565) );
  INV_X1 U12471 ( .A(n15232), .ZN(n14889) );
  OR2_X1 U12472 ( .A1(n15757), .A2(n14889), .ZN(n10566) );
  NAND2_X1 U12473 ( .A1(n15248), .A2(n10566), .ZN(n15231) );
  INV_X1 U12474 ( .A(n15227), .ZN(n15230) );
  OR2_X1 U12475 ( .A1(n15753), .A2(n15215), .ZN(n10567) );
  NAND2_X1 U12476 ( .A1(n15748), .A2(n14888), .ZN(n10568) );
  INV_X1 U12477 ( .A(n14926), .ZN(n15217) );
  OR2_X1 U12478 ( .A1(n15739), .A2(n15217), .ZN(n15174) );
  INV_X1 U12479 ( .A(n15194), .ZN(n15161) );
  OR2_X1 U12480 ( .A1(n15729), .A2(n15161), .ZN(n10569) );
  NAND2_X1 U12481 ( .A1(n15156), .A2(n10571), .ZN(n15141) );
  INV_X1 U12482 ( .A(n14924), .ZN(n15162) );
  AND2_X1 U12483 ( .A1(n15718), .A2(n15162), .ZN(n10572) );
  INV_X1 U12484 ( .A(n14923), .ZN(n14898) );
  NAND2_X1 U12485 ( .A1(n15123), .A2(n14898), .ZN(n10573) );
  NOR2_X1 U12486 ( .A1(n15696), .A2(n15112), .ZN(n13215) );
  NOR2_X1 U12487 ( .A1(n13214), .A2(n13215), .ZN(n10574) );
  INV_X1 U12488 ( .A(n15090), .ZN(n10575) );
  NAND2_X1 U12489 ( .A1(n10576), .A2(n10575), .ZN(n15072) );
  INV_X1 U12490 ( .A(n14921), .ZN(n14800) );
  NAND2_X1 U12491 ( .A1(n15686), .A2(n14800), .ZN(n10577) );
  NAND2_X1 U12492 ( .A1(n15072), .A2(n10577), .ZN(n10579) );
  INV_X1 U12493 ( .A(n10641), .ZN(n10578) );
  XNOR2_X1 U12494 ( .A(n10579), .B(n10578), .ZN(n10583) );
  INV_X1 U12495 ( .A(n10580), .ZN(n10581) );
  NAND2_X1 U12496 ( .A1(n15233), .A2(n14921), .ZN(n15677) );
  NAND2_X1 U12497 ( .A1(n15807), .A2(P1_B_REG_SCAN_IN), .ZN(n10584) );
  MUX2_X1 U12498 ( .A(P1_B_REG_SCAN_IN), .B(n10584), .S(n13205), .Z(n10585) );
  NAND2_X1 U12499 ( .A1(n10585), .A2(n15803), .ZN(n11235) );
  INV_X1 U12500 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10587) );
  INV_X1 U12501 ( .A(n13205), .ZN(n10586) );
  INV_X1 U12502 ( .A(n12157), .ZN(n11420) );
  INV_X1 U12503 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n11238) );
  INV_X1 U12504 ( .A(n15807), .ZN(n10588) );
  NOR2_X1 U12505 ( .A1(n15803), .A2(n10588), .ZN(n11236) );
  NOR4_X1 U12506 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10597) );
  NOR4_X1 U12507 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10596) );
  NOR4_X1 U12508 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10592) );
  NOR4_X1 U12509 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10591) );
  NOR4_X1 U12510 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10590) );
  NOR4_X1 U12511 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10589) );
  NAND4_X1 U12512 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .ZN(
        n10593) );
  NOR4_X1 U12513 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n10594), .A4(n10593), .ZN(n10595) );
  NAND3_X1 U12514 ( .A1(n10597), .A2(n10596), .A3(n10595), .ZN(n10598) );
  NAND2_X1 U12515 ( .A1(n10599), .A2(n10598), .ZN(n11416) );
  NAND4_X1 U12516 ( .A1(n11419), .A2(n11420), .A3(n11415), .A4(n11416), .ZN(
        n10655) );
  AOI21_X1 U12517 ( .B1(n15682), .B2(n15677), .A(n16398), .ZN(n10601) );
  NAND2_X1 U12518 ( .A1(n14943), .A2(n9115), .ZN(n16309) );
  NAND2_X1 U12519 ( .A1(n10602), .A2(n16309), .ZN(n10605) );
  OR2_X1 U12520 ( .A1(n10603), .A2(n9154), .ZN(n10604) );
  NAND2_X1 U12521 ( .A1(n16342), .A2(n16349), .ZN(n10607) );
  NAND2_X1 U12522 ( .A1(n9196), .A2(n16348), .ZN(n10606) );
  INV_X1 U12523 ( .A(n12036), .ZN(n10608) );
  NAND2_X1 U12524 ( .A1(n12037), .A2(n10608), .ZN(n10610) );
  OR2_X1 U12525 ( .A1(n16365), .A2(n14941), .ZN(n10609) );
  NAND2_X1 U12526 ( .A1(n10610), .A2(n10609), .ZN(n16376) );
  NAND2_X1 U12527 ( .A1(n16376), .A2(n16377), .ZN(n10612) );
  NAND2_X1 U12528 ( .A1(n9860), .A2(n11996), .ZN(n10611) );
  NAND2_X1 U12529 ( .A1(n10612), .A2(n10611), .ZN(n11991) );
  INV_X1 U12530 ( .A(n11994), .ZN(n10613) );
  NAND2_X1 U12531 ( .A1(n11991), .A2(n10613), .ZN(n10615) );
  NAND2_X1 U12532 ( .A1(n16401), .A2(n11845), .ZN(n10614) );
  NAND2_X1 U12533 ( .A1(n10615), .A2(n10614), .ZN(n12175) );
  OAI21_X1 U12534 ( .B1(n12175), .B2(n7550), .A(n7463), .ZN(n10616) );
  INV_X1 U12535 ( .A(n10616), .ZN(n12160) );
  NAND2_X1 U12536 ( .A1(n12160), .A2(n12163), .ZN(n12159) );
  OR2_X1 U12537 ( .A1(n12236), .A2(n14937), .ZN(n10617) );
  AND2_X2 U12538 ( .A1(n12159), .A2(n10617), .ZN(n12218) );
  NAND2_X1 U12539 ( .A1(n12573), .A2(n14936), .ZN(n10618) );
  NAND2_X1 U12540 ( .A1(n12217), .A2(n10618), .ZN(n12196) );
  INV_X1 U12541 ( .A(n10619), .ZN(n12366) );
  NAND2_X1 U12542 ( .A1(n12367), .A2(n12366), .ZN(n12365) );
  OR2_X1 U12543 ( .A1(n12928), .A2(n14934), .ZN(n10620) );
  AND2_X2 U12544 ( .A1(n12365), .A2(n10620), .ZN(n12610) );
  NAND2_X1 U12545 ( .A1(n12614), .A2(n14933), .ZN(n10622) );
  INV_X1 U12546 ( .A(n12553), .ZN(n10623) );
  OR2_X1 U12547 ( .A1(n12813), .A2(n14932), .ZN(n10624) );
  NAND2_X1 U12548 ( .A1(n12833), .A2(n8236), .ZN(n12832) );
  OR2_X1 U12549 ( .A1(n13176), .A2(n14931), .ZN(n10625) );
  NAND2_X1 U12550 ( .A1(n12832), .A2(n10625), .ZN(n12956) );
  INV_X1 U12551 ( .A(n12956), .ZN(n10626) );
  NAND2_X1 U12552 ( .A1(n16561), .A2(n14930), .ZN(n10627) );
  OR2_X1 U12553 ( .A1(n15762), .A2(n14928), .ZN(n10628) );
  NAND2_X2 U12554 ( .A1(n15258), .A2(n7696), .ZN(n15257) );
  NAND2_X1 U12555 ( .A1(n15757), .A2(n15232), .ZN(n10629) );
  AND2_X1 U12556 ( .A1(n15753), .A2(n14927), .ZN(n10630) );
  OR2_X1 U12557 ( .A1(n15753), .A2(n14927), .ZN(n10631) );
  INV_X1 U12558 ( .A(n15192), .ZN(n15200) );
  NAND2_X1 U12559 ( .A1(n15739), .A2(n14926), .ZN(n10632) );
  NAND2_X1 U12560 ( .A1(n15741), .A2(n10632), .ZN(n15181) );
  OR2_X1 U12561 ( .A1(n15729), .A2(n15194), .ZN(n10633) );
  NAND2_X1 U12562 ( .A1(n10645), .A2(n14830), .ZN(n10634) );
  NAND2_X1 U12563 ( .A1(n10635), .A2(n10634), .ZN(n15150) );
  INV_X1 U12564 ( .A(n15119), .ZN(n10637) );
  NAND2_X1 U12565 ( .A1(n15123), .A2(n14923), .ZN(n10638) );
  INV_X1 U12566 ( .A(n13214), .ZN(n13226) );
  OR2_X1 U12567 ( .A1(n15691), .A2(n15076), .ZN(n10639) );
  OR2_X1 U12568 ( .A1(n10958), .A2(n9825), .ZN(n10644) );
  NAND2_X1 U12569 ( .A1(n9824), .A2(n13032), .ZN(n10642) );
  INV_X1 U12570 ( .A(n15739), .ZN(n15199) );
  INV_X1 U12571 ( .A(n12891), .ZN(n12310) );
  INV_X1 U12572 ( .A(n12236), .ZN(n12162) );
  NAND2_X1 U12573 ( .A1(n16348), .A2(n16343), .ZN(n16344) );
  NAND2_X1 U12574 ( .A1(n12162), .A2(n12161), .ZN(n12227) );
  NOR2_X2 U12575 ( .A1(n12227), .A2(n12573), .ZN(n12226) );
  INV_X1 U12576 ( .A(n12614), .ZN(n16494) );
  INV_X1 U12577 ( .A(n12548), .ZN(n12837) );
  INV_X1 U12578 ( .A(n13176), .ZN(n16527) );
  NAND2_X1 U12579 ( .A1(n12837), .A2(n16527), .ZN(n12957) );
  NOR2_X2 U12580 ( .A1(n12957), .A2(n16561), .ZN(n16623) );
  NAND2_X1 U12581 ( .A1(n16641), .A2(n16623), .ZN(n16621) );
  NAND2_X1 U12582 ( .A1(n15199), .A2(n15221), .ZN(n15198) );
  NAND2_X1 U12583 ( .A1(n10645), .A2(n15163), .ZN(n15165) );
  OR2_X1 U12584 ( .A1(n15165), .A2(n15718), .ZN(n15142) );
  OR2_X2 U12585 ( .A1(n15711), .A2(n15142), .ZN(n15131) );
  INV_X1 U12586 ( .A(n15691), .ZN(n13224) );
  INV_X1 U12587 ( .A(n15686), .ZN(n15085) );
  NAND2_X1 U12588 ( .A1(n15083), .A2(n10658), .ZN(n15064) );
  INV_X1 U12589 ( .A(n15083), .ZN(n10648) );
  NAND2_X4 U12590 ( .A1(n10647), .A2(n7436), .ZN(n16566) );
  AOI21_X1 U12591 ( .B1(n10648), .B2(n15679), .A(n16566), .ZN(n10649) );
  NAND2_X1 U12592 ( .A1(n15064), .A2(n10649), .ZN(n15681) );
  INV_X1 U12593 ( .A(n15681), .ZN(n10660) );
  INV_X1 U12594 ( .A(n16640), .ZN(n16327) );
  INV_X1 U12595 ( .A(n9908), .ZN(n14957) );
  INV_X1 U12596 ( .A(P1_B_REG_SCAN_IN), .ZN(n10651) );
  NOR2_X1 U12597 ( .A1(n14954), .A2(n10651), .ZN(n15060) );
  NOR2_X1 U12598 ( .A1(n10652), .A2(n15060), .ZN(n10653) );
  NAND2_X1 U12599 ( .A1(n15234), .A2(n10653), .ZN(n15676) );
  OAI22_X1 U12600 ( .A1(n10655), .A2(n15676), .B1(n10654), .B2(n16653), .ZN(
        n10656) );
  AOI21_X1 U12601 ( .B1(n16398), .B2(P1_REG2_REG_29__SCAN_IN), .A(n10656), 
        .ZN(n10657) );
  OAI21_X1 U12602 ( .B1(n10658), .B2(n16493), .A(n10657), .ZN(n10659) );
  INV_X1 U12603 ( .A(n10661), .ZN(n10662) );
  NAND2_X1 U12604 ( .A1(n13208), .A2(n10871), .ZN(n10668) );
  OR2_X1 U12605 ( .A1(n10873), .A2(n14778), .ZN(n10667) );
  NAND2_X1 U12606 ( .A1(n10670), .A2(n10669), .ZN(n11509) );
  INV_X1 U12607 ( .A(n11509), .ZN(n10671) );
  NAND3_X1 U12608 ( .A1(n15822), .A2(n11499), .A3(n11512), .ZN(n10673) );
  INV_X1 U12609 ( .A(n11508), .ZN(n10672) );
  OR2_X1 U12610 ( .A1(n11852), .A2(n10331), .ZN(n10674) );
  OR2_X1 U12611 ( .A1(n16598), .A2(n14609), .ZN(n10675) );
  NAND2_X1 U12612 ( .A1(n10677), .A2(n10676), .ZN(n10679) );
  INV_X1 U12613 ( .A(P2_B_REG_SCAN_IN), .ZN(n10680) );
  NOR2_X1 U12614 ( .A1(n14784), .A2(n10680), .ZN(n10681) );
  NOR2_X1 U12615 ( .A1(n14604), .A2(n10681), .ZN(n14437) );
  INV_X1 U12616 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14444) );
  NAND2_X1 U12617 ( .A1(n10682), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U12618 ( .A1(n10683), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n10684) );
  OAI211_X1 U12619 ( .C1(n10877), .C2(n14444), .A(n10685), .B(n10684), .ZN(
        n14364) );
  NAND2_X1 U12620 ( .A1(n14437), .A2(n14364), .ZN(n10686) );
  INV_X2 U12621 ( .A(n14610), .ZN(n16598) );
  OR2_X1 U12622 ( .A1(n11491), .A2(n10329), .ZN(n11505) );
  INV_X1 U12623 ( .A(n14640), .ZN(n16596) );
  AOI22_X1 U12624 ( .A1(n10689), .A2(n16596), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n16598), .ZN(n10690) );
  OAI21_X1 U12625 ( .B1(n10891), .B2(n14621), .A(n10690), .ZN(n10691) );
  MUX2_X1 U12626 ( .A(n10697), .B(n14387), .S(n10702), .Z(n10701) );
  NAND2_X1 U12627 ( .A1(n10696), .A2(n10695), .ZN(n10698) );
  NAND2_X1 U12628 ( .A1(n10698), .A2(n10901), .ZN(n10700) );
  NAND2_X1 U12629 ( .A1(n11668), .A2(n10702), .ZN(n10703) );
  NAND2_X1 U12630 ( .A1(n10708), .A2(n10709), .ZN(n10707) );
  MUX2_X1 U12631 ( .A(n7435), .B(n11668), .S(n10714), .Z(n10706) );
  NAND2_X1 U12632 ( .A1(n10707), .A2(n10706), .ZN(n10713) );
  NAND2_X1 U12633 ( .A1(n10711), .A2(n10710), .ZN(n10712) );
  NAND2_X1 U12634 ( .A1(n10713), .A2(n10712), .ZN(n10717) );
  MUX2_X1 U12635 ( .A(n11679), .B(n14386), .S(n10919), .Z(n10718) );
  NAND2_X1 U12636 ( .A1(n10717), .A2(n10718), .ZN(n10716) );
  MUX2_X1 U12637 ( .A(n11679), .B(n14386), .S(n10899), .Z(n10715) );
  NAND2_X1 U12638 ( .A1(n10716), .A2(n10715), .ZN(n10722) );
  INV_X1 U12639 ( .A(n10717), .ZN(n10720) );
  NAND2_X1 U12640 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  MUX2_X1 U12641 ( .A(n14384), .B(n12045), .S(n10714), .Z(n10723) );
  INV_X1 U12642 ( .A(n11647), .ZN(n14383) );
  MUX2_X1 U12643 ( .A(n11612), .B(n14383), .S(n10919), .Z(n10728) );
  NAND2_X1 U12644 ( .A1(n10727), .A2(n10728), .ZN(n10726) );
  MUX2_X1 U12645 ( .A(n14383), .B(n11612), .S(n10919), .Z(n10725) );
  NAND2_X1 U12646 ( .A1(n10726), .A2(n10725), .ZN(n10732) );
  INV_X1 U12647 ( .A(n10727), .ZN(n10730) );
  INV_X1 U12648 ( .A(n10728), .ZN(n10729) );
  NAND2_X1 U12649 ( .A1(n10730), .A2(n10729), .ZN(n10731) );
  MUX2_X1 U12650 ( .A(n14382), .B(n11701), .S(n10919), .Z(n10734) );
  MUX2_X1 U12651 ( .A(n11701), .B(n14382), .S(n10919), .Z(n10733) );
  INV_X1 U12652 ( .A(n10734), .ZN(n10735) );
  MUX2_X1 U12653 ( .A(n16419), .B(n14381), .S(n10919), .Z(n10737) );
  MUX2_X1 U12654 ( .A(n16419), .B(n14381), .S(n10899), .Z(n10736) );
  INV_X1 U12655 ( .A(n10737), .ZN(n10738) );
  AND2_X1 U12656 ( .A1(n10739), .A2(n10738), .ZN(n10740) );
  NAND2_X1 U12657 ( .A1(n10741), .A2(n10740), .ZN(n10742) );
  MUX2_X1 U12658 ( .A(n12126), .B(n12088), .S(n10919), .Z(n10744) );
  MUX2_X1 U12659 ( .A(n12088), .B(n12126), .S(n10919), .Z(n10743) );
  INV_X1 U12660 ( .A(n10744), .ZN(n10745) );
  MUX2_X1 U12661 ( .A(n14380), .B(n12142), .S(n10899), .Z(n10748) );
  MUX2_X1 U12662 ( .A(n14380), .B(n12142), .S(n10919), .Z(n10746) );
  INV_X1 U12663 ( .A(n10748), .ZN(n10749) );
  MUX2_X1 U12664 ( .A(n14379), .B(n7849), .S(n10919), .Z(n10753) );
  MUX2_X1 U12665 ( .A(n14379), .B(n7849), .S(n10899), .Z(n10750) );
  NAND2_X1 U12666 ( .A1(n10751), .A2(n10750), .ZN(n10757) );
  INV_X1 U12667 ( .A(n10752), .ZN(n10755) );
  INV_X1 U12668 ( .A(n10753), .ZN(n10754) );
  NAND2_X1 U12669 ( .A1(n10755), .A2(n10754), .ZN(n10756) );
  MUX2_X1 U12670 ( .A(n12355), .B(n12463), .S(n10899), .Z(n10759) );
  MUX2_X1 U12671 ( .A(n12355), .B(n12463), .S(n10919), .Z(n10758) );
  MUX2_X1 U12672 ( .A(n14378), .B(n12644), .S(n10919), .Z(n10763) );
  MUX2_X1 U12673 ( .A(n14378), .B(n12644), .S(n10899), .Z(n10760) );
  NAND2_X1 U12674 ( .A1(n10761), .A2(n10760), .ZN(n10767) );
  INV_X1 U12675 ( .A(n10762), .ZN(n10765) );
  INV_X1 U12676 ( .A(n10763), .ZN(n10764) );
  NAND2_X1 U12677 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  NAND2_X1 U12678 ( .A1(n10767), .A2(n10766), .ZN(n10769) );
  MUX2_X1 U12679 ( .A(n12702), .B(n12770), .S(n10899), .Z(n10770) );
  MUX2_X1 U12680 ( .A(n12702), .B(n12770), .S(n10919), .Z(n10768) );
  INV_X1 U12681 ( .A(n10770), .ZN(n10771) );
  MUX2_X1 U12682 ( .A(n14377), .B(n12863), .S(n10919), .Z(n10775) );
  MUX2_X1 U12683 ( .A(n14377), .B(n12863), .S(n10899), .Z(n10772) );
  NAND2_X1 U12684 ( .A1(n10773), .A2(n10772), .ZN(n10779) );
  INV_X1 U12685 ( .A(n10774), .ZN(n10777) );
  INV_X1 U12686 ( .A(n10775), .ZN(n10776) );
  NAND2_X1 U12687 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  NAND2_X1 U12688 ( .A1(n10779), .A2(n10778), .ZN(n10782) );
  MUX2_X1 U12689 ( .A(n14376), .B(n16600), .S(n10899), .Z(n10783) );
  NAND2_X1 U12690 ( .A1(n10782), .A2(n10783), .ZN(n10781) );
  MUX2_X1 U12691 ( .A(n14376), .B(n16600), .S(n10919), .Z(n10780) );
  NAND2_X1 U12692 ( .A1(n10781), .A2(n10780), .ZN(n10790) );
  INV_X1 U12693 ( .A(n10782), .ZN(n10785) );
  INV_X1 U12694 ( .A(n10783), .ZN(n10784) );
  NAND2_X1 U12695 ( .A1(n10785), .A2(n10784), .ZN(n10788) );
  MUX2_X1 U12696 ( .A(n14375), .B(n13050), .S(n10919), .Z(n10787) );
  MUX2_X1 U12697 ( .A(n14375), .B(n13050), .S(n10714), .Z(n10786) );
  INV_X1 U12698 ( .A(n10787), .ZN(n10789) );
  MUX2_X1 U12699 ( .A(n14374), .B(n14720), .S(n10714), .Z(n10794) );
  NAND2_X1 U12700 ( .A1(n10793), .A2(n10794), .ZN(n10792) );
  MUX2_X1 U12701 ( .A(n14374), .B(n14720), .S(n10919), .Z(n10791) );
  NAND2_X1 U12702 ( .A1(n10792), .A2(n10791), .ZN(n10798) );
  INV_X1 U12703 ( .A(n10793), .ZN(n10796) );
  INV_X1 U12704 ( .A(n10794), .ZN(n10795) );
  NAND2_X1 U12705 ( .A1(n10796), .A2(n10795), .ZN(n10797) );
  MUX2_X1 U12706 ( .A(n14373), .B(n14716), .S(n10919), .Z(n10801) );
  MUX2_X1 U12707 ( .A(n14373), .B(n14716), .S(n10714), .Z(n10799) );
  INV_X1 U12708 ( .A(n10801), .ZN(n10802) );
  MUX2_X1 U12709 ( .A(n14372), .B(n14710), .S(n10714), .Z(n10805) );
  MUX2_X1 U12710 ( .A(n14372), .B(n14710), .S(n10919), .Z(n10803) );
  NAND2_X1 U12711 ( .A1(n10804), .A2(n10803), .ZN(n10808) );
  INV_X1 U12712 ( .A(n10805), .ZN(n10806) );
  NAND2_X1 U12713 ( .A1(n10808), .A2(n10807), .ZN(n10810) );
  MUX2_X1 U12714 ( .A(n14579), .B(n14594), .S(n10919), .Z(n10811) );
  MUX2_X1 U12715 ( .A(n14579), .B(n14594), .S(n10714), .Z(n10809) );
  MUX2_X1 U12716 ( .A(n14371), .B(n14698), .S(n10714), .Z(n10813) );
  MUX2_X1 U12717 ( .A(n14371), .B(n14698), .S(n10919), .Z(n10812) );
  MUX2_X1 U12718 ( .A(n14576), .B(n14566), .S(n10919), .Z(n10816) );
  MUX2_X1 U12719 ( .A(n14576), .B(n14566), .S(n10714), .Z(n10814) );
  INV_X1 U12720 ( .A(n10816), .ZN(n10817) );
  MUX2_X1 U12721 ( .A(n14551), .B(n14370), .S(n10919), .Z(n10820) );
  MUX2_X1 U12722 ( .A(n14551), .B(n14370), .S(n10714), .Z(n10818) );
  INV_X1 U12723 ( .A(n10820), .ZN(n10821) );
  MUX2_X1 U12724 ( .A(n14369), .B(n14527), .S(n10919), .Z(n10824) );
  MUX2_X1 U12725 ( .A(n14527), .B(n14369), .S(n10919), .Z(n10822) );
  INV_X1 U12726 ( .A(n10824), .ZN(n10825) );
  MUX2_X1 U12727 ( .A(n14492), .B(n14676), .S(n10714), .Z(n10828) );
  MUX2_X1 U12728 ( .A(n14492), .B(n14676), .S(n10919), .Z(n10826) );
  NAND2_X1 U12729 ( .A1(n10827), .A2(n10826), .ZN(n10831) );
  INV_X1 U12730 ( .A(n10828), .ZN(n10829) );
  NAND2_X1 U12731 ( .A1(n7517), .A2(n10829), .ZN(n10830) );
  MUX2_X1 U12732 ( .A(n14368), .B(n14498), .S(n10919), .Z(n10833) );
  MUX2_X1 U12733 ( .A(n14368), .B(n14498), .S(n10714), .Z(n10832) );
  MUX2_X1 U12734 ( .A(n14493), .B(n14480), .S(n10714), .Z(n10836) );
  MUX2_X1 U12735 ( .A(n14493), .B(n14480), .S(n10919), .Z(n10834) );
  INV_X1 U12736 ( .A(n10836), .ZN(n10837) );
  MUX2_X1 U12737 ( .A(n14367), .B(n14467), .S(n10702), .Z(n10841) );
  MUX2_X1 U12738 ( .A(n14367), .B(n14467), .S(n10714), .Z(n10838) );
  NAND2_X1 U12739 ( .A1(n10839), .A2(n10838), .ZN(n10843) );
  NAND2_X1 U12740 ( .A1(n10843), .A2(n10842), .ZN(n10952) );
  INV_X1 U12741 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13211) );
  OR2_X1 U12742 ( .A1(n10873), .A2(n13211), .ZN(n10844) );
  XNOR2_X1 U12743 ( .A(n14447), .B(n14364), .ZN(n10869) );
  NAND2_X1 U12744 ( .A1(n10847), .A2(n10846), .ZN(n14580) );
  XNOR2_X1 U12745 ( .A(n12770), .B(n12772), .ZN(n12595) );
  NAND2_X1 U12746 ( .A1(n11492), .A2(n14387), .ZN(n11535) );
  AND2_X1 U12747 ( .A1(n11665), .A2(n11535), .ZN(n11860) );
  NAND4_X1 U12748 ( .A1(n10849), .A2(n10848), .A3(n11860), .A4(n10333), .ZN(
        n10850) );
  NOR2_X1 U12749 ( .A1(n11614), .A2(n10850), .ZN(n10853) );
  NAND4_X1 U12750 ( .A1(n12245), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10854) );
  NOR3_X1 U12751 ( .A1(n10855), .A2(n12082), .A3(n10854), .ZN(n10856) );
  NAND4_X1 U12752 ( .A1(n12456), .A2(n12375), .A3(n10856), .A4(n12210), .ZN(
        n10857) );
  OR4_X1 U12753 ( .A1(n16581), .A2(n10858), .A3(n12595), .A4(n10857), .ZN(
        n10859) );
  NOR2_X1 U12754 ( .A1(n12912), .A2(n10859), .ZN(n10860) );
  NAND4_X1 U12755 ( .A1(n14626), .A2(n10860), .A3(n14632), .A4(n13085), .ZN(
        n10861) );
  NOR2_X1 U12756 ( .A1(n14580), .A2(n10861), .ZN(n10862) );
  NAND4_X1 U12757 ( .A1(n14549), .A2(n10862), .A3(n14570), .A4(n14600), .ZN(
        n10863) );
  OR2_X1 U12758 ( .A1(n14532), .A2(n10863), .ZN(n10864) );
  NOR2_X1 U12759 ( .A1(n10865), .A2(n10864), .ZN(n10868) );
  NAND2_X1 U12760 ( .A1(n14477), .A2(n14490), .ZN(n10870) );
  NAND2_X1 U12761 ( .A1(n10872), .A2(n10871), .ZN(n10875) );
  INV_X1 U12762 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14771) );
  OR2_X1 U12763 ( .A1(n10873), .A2(n14771), .ZN(n10874) );
  INV_X1 U12764 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14652) );
  OR2_X1 U12765 ( .A1(n10876), .A2(n14652), .ZN(n10881) );
  INV_X1 U12766 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14436) );
  OR2_X1 U12767 ( .A1(n10877), .A2(n14436), .ZN(n10880) );
  INV_X1 U12768 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14726) );
  OR2_X1 U12769 ( .A1(n10878), .A2(n14726), .ZN(n10879) );
  AND3_X1 U12770 ( .A1(n10881), .A2(n10880), .A3(n10879), .ZN(n14438) );
  NAND2_X1 U12771 ( .A1(n14434), .A2(n14438), .ZN(n10923) );
  XNOR2_X1 U12772 ( .A(n10882), .B(n10696), .ZN(n10883) );
  NAND2_X1 U12773 ( .A1(n10883), .A2(n10331), .ZN(n10915) );
  OR2_X1 U12774 ( .A1(n11852), .A2(n10695), .ZN(n10887) );
  NAND2_X1 U12775 ( .A1(n10696), .A2(n10884), .ZN(n10885) );
  AND2_X1 U12776 ( .A1(n10887), .A2(n10885), .ZN(n10886) );
  NAND2_X1 U12777 ( .A1(n10915), .A2(n10886), .ZN(n10918) );
  MUX2_X1 U12778 ( .A(n10905), .B(n10923), .S(n10714), .Z(n10896) );
  MUX2_X1 U12779 ( .A(n14447), .B(n14364), .S(n10714), .Z(n10898) );
  INV_X1 U12780 ( .A(n14438), .ZN(n14363) );
  NAND2_X1 U12781 ( .A1(n14363), .A2(n10919), .ZN(n10888) );
  NAND4_X1 U12782 ( .A1(n10902), .A2(n10888), .A3(n10946), .A4(n10887), .ZN(
        n10889) );
  AND2_X1 U12783 ( .A1(n10889), .A2(n14364), .ZN(n10890) );
  AOI21_X1 U12784 ( .B1(n14447), .B2(n10714), .A(n10890), .ZN(n10897) );
  INV_X1 U12785 ( .A(n10913), .ZN(n10894) );
  INV_X1 U12786 ( .A(n14365), .ZN(n10892) );
  MUX2_X1 U12787 ( .A(n10892), .B(n10891), .S(n10919), .Z(n10914) );
  INV_X1 U12788 ( .A(n10914), .ZN(n10893) );
  OAI22_X1 U12789 ( .A1(n10898), .A2(n10897), .B1(n10894), .B2(n10893), .ZN(
        n10895) );
  NAND2_X1 U12790 ( .A1(n10898), .A2(n10897), .ZN(n10911) );
  NAND2_X1 U12791 ( .A1(n10933), .A2(n10911), .ZN(n10908) );
  OR2_X1 U12792 ( .A1(n10923), .A2(n10714), .ZN(n10904) );
  NAND2_X1 U12793 ( .A1(n10908), .A2(n10904), .ZN(n10900) );
  NAND2_X1 U12794 ( .A1(n10918), .A2(n10900), .ZN(n10910) );
  NAND2_X1 U12795 ( .A1(n13114), .A2(n10902), .ZN(n10903) );
  OAI211_X1 U12796 ( .C1(n10948), .C2(n11485), .A(n10946), .B(n10903), .ZN(
        n10921) );
  OAI211_X1 U12797 ( .C1(n10905), .C2(n10919), .A(n10904), .B(n10921), .ZN(
        n10906) );
  INV_X1 U12798 ( .A(n10906), .ZN(n10907) );
  NAND2_X1 U12799 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  OAI211_X1 U12800 ( .C1(n10914), .C2(n10913), .A(n10912), .B(n10911), .ZN(
        n10917) );
  INV_X1 U12801 ( .A(n10915), .ZN(n10916) );
  OAI21_X1 U12802 ( .B1(n10933), .B2(n10917), .A(n10930), .ZN(n10929) );
  NOR2_X1 U12803 ( .A1(n10918), .A2(n10917), .ZN(n10941) );
  MUX2_X1 U12804 ( .A(n10920), .B(n14736), .S(n10702), .Z(n10935) );
  MUX2_X1 U12805 ( .A(n14366), .B(n14453), .S(n10714), .Z(n10931) );
  NAND3_X1 U12806 ( .A1(n10941), .A2(n10935), .A3(n10931), .ZN(n10928) );
  INV_X1 U12807 ( .A(n10921), .ZN(n10922) );
  AND2_X1 U12808 ( .A1(n10923), .A2(n10922), .ZN(n10934) );
  INV_X1 U12809 ( .A(n10931), .ZN(n10925) );
  INV_X1 U12810 ( .A(n10935), .ZN(n10924) );
  AND2_X1 U12811 ( .A1(n10925), .A2(n10924), .ZN(n10939) );
  INV_X1 U12812 ( .A(n10933), .ZN(n10926) );
  NAND4_X1 U12813 ( .A1(n10930), .A2(n10934), .A3(n10939), .A4(n10926), .ZN(
        n10927) );
  OAI211_X1 U12814 ( .C1(n10932), .C2(n10929), .A(n10928), .B(n10927), .ZN(
        n10945) );
  INV_X1 U12815 ( .A(n10934), .ZN(n10936) );
  INV_X1 U12816 ( .A(n11511), .ZN(n10938) );
  NAND2_X1 U12817 ( .A1(n10938), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13001) );
  INV_X1 U12818 ( .A(n10939), .ZN(n10940) );
  NAND2_X1 U12819 ( .A1(n10941), .A2(n10940), .ZN(n10943) );
  NAND2_X1 U12820 ( .A1(n10952), .A2(n8393), .ZN(n10950) );
  INV_X1 U12821 ( .A(n14784), .ZN(n11306) );
  INV_X1 U12822 ( .A(n10946), .ZN(n11503) );
  NAND4_X1 U12823 ( .A1(n14578), .A2(n11306), .A3(n11503), .A4(n15823), .ZN(
        n10947) );
  OAI211_X1 U12824 ( .C1(n10948), .C2(n13001), .A(n10947), .B(P2_B_REG_SCAN_IN), .ZN(n10949) );
  OAI211_X1 U12825 ( .C1(n10952), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        P2_U3328) );
  NOR2_X1 U12826 ( .A1(n10957), .A2(P1_U3086), .ZN(n10954) );
  NAND2_X2 U12827 ( .A1(n10958), .A2(n10957), .ZN(n10981) );
  INV_X2 U12828 ( .A(n10981), .ZN(n13302) );
  INV_X2 U12829 ( .A(n10968), .ZN(n13315) );
  AND2_X1 U12830 ( .A1(n14926), .A2(n13315), .ZN(n10959) );
  AOI21_X1 U12831 ( .B1(n15739), .B2(n13316), .A(n10959), .ZN(n13249) );
  NAND2_X1 U12832 ( .A1(n15739), .A2(n13313), .ZN(n10961) );
  NAND2_X1 U12833 ( .A1(n14926), .A2(n13316), .ZN(n10960) );
  NAND2_X1 U12834 ( .A1(n10961), .A2(n10960), .ZN(n10962) );
  XNOR2_X1 U12835 ( .A(n10962), .B(n10643), .ZN(n13251) );
  XOR2_X1 U12836 ( .A(n13249), .B(n13251), .Z(n11099) );
  NOR2_X1 U12837 ( .A1(n10968), .A2(n12166), .ZN(n10963) );
  AOI21_X1 U12838 ( .B1(n12189), .B2(n13316), .A(n10963), .ZN(n10997) );
  INV_X1 U12839 ( .A(n10997), .ZN(n11000) );
  AOI22_X1 U12840 ( .A1(n12189), .A2(n13313), .B1(n13316), .B2(n14938), .ZN(
        n10964) );
  XNOR2_X1 U12841 ( .A(n10964), .B(n10643), .ZN(n10998) );
  INV_X1 U12842 ( .A(n10998), .ZN(n10999) );
  OAI22_X1 U12843 ( .A1(n10968), .A2(n11602), .B1(n16314), .B2(n11059), .ZN(
        n10966) );
  OR2_X1 U12844 ( .A1(n10981), .A2(n16314), .ZN(n10965) );
  INV_X1 U12845 ( .A(n14943), .ZN(n11595) );
  NAND2_X1 U12846 ( .A1(n10969), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10972) );
  OR2_X1 U12847 ( .A1(n10981), .A2(n16310), .ZN(n10971) );
  OAI211_X1 U12848 ( .C1(n11059), .C2(n11595), .A(n10972), .B(n10971), .ZN(
        n11462) );
  OAI22_X1 U12849 ( .A1(n10968), .A2(n9196), .B1(n16348), .B2(n11059), .ZN(
        n10975) );
  OAI22_X1 U12850 ( .A1(n11059), .A2(n9196), .B1(n10981), .B2(n16348), .ZN(
        n10973) );
  XNOR2_X1 U12851 ( .A(n10973), .B(n10643), .ZN(n10974) );
  XOR2_X1 U12852 ( .A(n10975), .B(n10974), .Z(n11600) );
  NAND2_X1 U12853 ( .A1(n11599), .A2(n11600), .ZN(n11598) );
  NAND2_X1 U12854 ( .A1(n11598), .A2(n10976), .ZN(n11711) );
  AOI22_X1 U12855 ( .A1(n13316), .A2(n14941), .B1(n13313), .B2(n16365), .ZN(
        n10977) );
  XNOR2_X1 U12856 ( .A(n10977), .B(n10643), .ZN(n10979) );
  AOI22_X1 U12857 ( .A1(n13315), .A2(n14941), .B1(n13316), .B2(n16365), .ZN(
        n10978) );
  XNOR2_X1 U12858 ( .A(n10979), .B(n10978), .ZN(n11712) );
  NOR2_X1 U12859 ( .A1(n10979), .A2(n10978), .ZN(n10984) );
  NAND2_X1 U12860 ( .A1(n13315), .A2(n14940), .ZN(n10980) );
  OAI21_X1 U12861 ( .B1(n9860), .B2(n11059), .A(n10980), .ZN(n10983) );
  OAI22_X1 U12862 ( .A1(n9860), .A2(n10981), .B1(n11996), .B2(n11059), .ZN(
        n10982) );
  XNOR2_X1 U12863 ( .A(n10982), .B(n13305), .ZN(n11842) );
  NAND2_X1 U12864 ( .A1(n12003), .A2(n13302), .ZN(n10989) );
  NAND2_X1 U12865 ( .A1(n13316), .A2(n14939), .ZN(n10988) );
  NAND2_X1 U12866 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  XNOR2_X1 U12867 ( .A(n10990), .B(n10643), .ZN(n10996) );
  INV_X1 U12868 ( .A(n10996), .ZN(n10994) );
  NAND2_X1 U12869 ( .A1(n12003), .A2(n13316), .ZN(n10992) );
  NAND2_X1 U12870 ( .A1(n13315), .A2(n14939), .ZN(n10991) );
  NAND2_X1 U12871 ( .A1(n10992), .A2(n10991), .ZN(n10995) );
  INV_X1 U12872 ( .A(n10995), .ZN(n10993) );
  NAND2_X1 U12873 ( .A1(n10994), .A2(n10993), .ZN(n11883) );
  AND2_X1 U12874 ( .A1(n10996), .A2(n10995), .ZN(n11884) );
  XNOR2_X1 U12875 ( .A(n10998), .B(n10997), .ZN(n11114) );
  AOI22_X1 U12876 ( .A1(n12236), .A2(n13313), .B1(n13316), .B2(n14937), .ZN(
        n11001) );
  XNOR2_X1 U12877 ( .A(n11001), .B(n10643), .ZN(n11003) );
  NOR2_X1 U12878 ( .A1(n10968), .A2(n12570), .ZN(n11002) );
  AOI21_X1 U12879 ( .B1(n12236), .B2(n13316), .A(n11002), .ZN(n11004) );
  XNOR2_X1 U12880 ( .A(n11003), .B(n11004), .ZN(n11120) );
  INV_X1 U12881 ( .A(n11003), .ZN(n11006) );
  INV_X1 U12882 ( .A(n11004), .ZN(n11005) );
  AOI22_X1 U12883 ( .A1(n12573), .A2(n13316), .B1(n13315), .B2(n14936), .ZN(
        n11009) );
  AOI22_X1 U12884 ( .A1(n12573), .A2(n13313), .B1(n13316), .B2(n14936), .ZN(
        n11007) );
  XNOR2_X1 U12885 ( .A(n11007), .B(n10643), .ZN(n11008) );
  XOR2_X1 U12886 ( .A(n11009), .B(n11008), .Z(n12566) );
  NAND2_X1 U12887 ( .A1(n12565), .A2(n12566), .ZN(n12564) );
  NAND2_X1 U12888 ( .A1(n12564), .A2(n11010), .ZN(n11015) );
  NOR2_X1 U12889 ( .A1(n10968), .A2(n12925), .ZN(n11011) );
  AOI21_X1 U12890 ( .B1(n12891), .B2(n13316), .A(n11011), .ZN(n11014) );
  INV_X1 U12891 ( .A(n11014), .ZN(n11012) );
  AOI22_X1 U12892 ( .A1(n12891), .A2(n13313), .B1(n13316), .B2(n14935), .ZN(
        n11013) );
  XNOR2_X1 U12893 ( .A(n11013), .B(n10643), .ZN(n12884) );
  NAND2_X1 U12894 ( .A1(n12928), .A2(n13302), .ZN(n11018) );
  NAND2_X1 U12895 ( .A1(n13316), .A2(n14934), .ZN(n11017) );
  NAND2_X1 U12896 ( .A1(n11018), .A2(n11017), .ZN(n11019) );
  XNOR2_X1 U12897 ( .A(n11019), .B(n13305), .ZN(n11022) );
  NOR2_X1 U12898 ( .A1(n10968), .A2(n12887), .ZN(n11020) );
  AOI21_X1 U12899 ( .B1(n12928), .B2(n13316), .A(n11020), .ZN(n11021) );
  NOR2_X1 U12900 ( .A1(n11022), .A2(n11021), .ZN(n12920) );
  NAND2_X1 U12901 ( .A1(n12614), .A2(n13302), .ZN(n11024) );
  NAND2_X1 U12902 ( .A1(n13316), .A2(n14933), .ZN(n11023) );
  NAND2_X1 U12903 ( .A1(n11024), .A2(n11023), .ZN(n11025) );
  XNOR2_X1 U12904 ( .A(n11025), .B(n10643), .ZN(n11029) );
  NAND2_X1 U12905 ( .A1(n12614), .A2(n13316), .ZN(n11027) );
  NAND2_X1 U12906 ( .A1(n13315), .A2(n14933), .ZN(n11026) );
  NAND2_X1 U12907 ( .A1(n11027), .A2(n11026), .ZN(n11028) );
  NOR2_X1 U12908 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  AOI21_X1 U12909 ( .B1(n11029), .B2(n11028), .A(n11030), .ZN(n13042) );
  NAND2_X1 U12910 ( .A1(n12813), .A2(n13302), .ZN(n11032) );
  NAND2_X1 U12911 ( .A1(n13316), .A2(n14932), .ZN(n11031) );
  NAND2_X1 U12912 ( .A1(n11032), .A2(n11031), .ZN(n11033) );
  XNOR2_X1 U12913 ( .A(n11033), .B(n10643), .ZN(n11036) );
  AOI22_X1 U12914 ( .A1(n12813), .A2(n13316), .B1(n13315), .B2(n14932), .ZN(
        n11034) );
  XNOR2_X1 U12915 ( .A(n11036), .B(n11034), .ZN(n13142) );
  INV_X1 U12916 ( .A(n11034), .ZN(n11035) );
  NAND2_X1 U12917 ( .A1(n13176), .A2(n13302), .ZN(n11039) );
  NAND2_X1 U12918 ( .A1(n13316), .A2(n14931), .ZN(n11038) );
  NAND2_X1 U12919 ( .A1(n11039), .A2(n11038), .ZN(n11040) );
  XNOR2_X1 U12920 ( .A(n11040), .B(n13305), .ZN(n11046) );
  NOR2_X1 U12921 ( .A1(n10968), .A2(n16544), .ZN(n11041) );
  AOI21_X1 U12922 ( .B1(n13176), .B2(n13316), .A(n11041), .ZN(n11047) );
  NAND2_X1 U12923 ( .A1(n11046), .A2(n11047), .ZN(n13168) );
  NAND2_X1 U12924 ( .A1(n16561), .A2(n13302), .ZN(n11043) );
  NAND2_X1 U12925 ( .A1(n13316), .A2(n14930), .ZN(n11042) );
  NAND2_X1 U12926 ( .A1(n11043), .A2(n11042), .ZN(n11044) );
  XNOR2_X1 U12927 ( .A(n11044), .B(n10643), .ZN(n11053) );
  NOR2_X1 U12928 ( .A1(n10968), .A2(n13172), .ZN(n11045) );
  AOI21_X1 U12929 ( .B1(n16561), .B2(n13316), .A(n11045), .ZN(n11051) );
  XNOR2_X1 U12930 ( .A(n11053), .B(n11051), .ZN(n16545) );
  INV_X1 U12931 ( .A(n11046), .ZN(n11049) );
  INV_X1 U12932 ( .A(n11047), .ZN(n11048) );
  NAND2_X1 U12933 ( .A1(n11049), .A2(n11048), .ZN(n16546) );
  NAND2_X1 U12934 ( .A1(n16547), .A2(n11050), .ZN(n16550) );
  INV_X1 U12935 ( .A(n11051), .ZN(n11052) );
  OR2_X1 U12936 ( .A1(n11053), .A2(n11052), .ZN(n11054) );
  NAND2_X1 U12937 ( .A1(n11055), .A2(n13302), .ZN(n11057) );
  NAND2_X1 U12938 ( .A1(n13316), .A2(n14929), .ZN(n11056) );
  NAND2_X1 U12939 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  XNOR2_X1 U12940 ( .A(n11058), .B(n10643), .ZN(n11060) );
  OAI22_X1 U12941 ( .A1(n16641), .A2(n11059), .B1(n16541), .B2(n10968), .ZN(
        n14907) );
  AOI22_X1 U12942 ( .A1(n15762), .A2(n13313), .B1(n13316), .B2(n14928), .ZN(
        n11062) );
  XNOR2_X1 U12943 ( .A(n11062), .B(n10643), .ZN(n11064) );
  AOI22_X1 U12944 ( .A1(n15762), .A2(n13316), .B1(n13315), .B2(n14928), .ZN(
        n11063) );
  XNOR2_X1 U12945 ( .A(n11064), .B(n11063), .ZN(n14851) );
  NAND2_X1 U12946 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U12947 ( .A1(n14849), .A2(n11065), .ZN(n14857) );
  NAND2_X1 U12948 ( .A1(n15757), .A2(n13313), .ZN(n11067) );
  NAND2_X1 U12949 ( .A1(n15232), .A2(n13316), .ZN(n11066) );
  NAND2_X1 U12950 ( .A1(n11067), .A2(n11066), .ZN(n11068) );
  XNOR2_X1 U12951 ( .A(n11068), .B(n10643), .ZN(n11069) );
  AOI22_X1 U12952 ( .A1(n15757), .A2(n13316), .B1(n13315), .B2(n15232), .ZN(
        n11070) );
  XNOR2_X1 U12953 ( .A(n11069), .B(n11070), .ZN(n14859) );
  INV_X1 U12954 ( .A(n11069), .ZN(n11071) );
  NAND2_X1 U12955 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  NAND2_X1 U12956 ( .A1(n15753), .A2(n13313), .ZN(n11074) );
  NAND2_X1 U12957 ( .A1(n14927), .A2(n13316), .ZN(n11073) );
  NAND2_X1 U12958 ( .A1(n11074), .A2(n11073), .ZN(n11075) );
  XNOR2_X1 U12959 ( .A(n11075), .B(n10643), .ZN(n11085) );
  AOI22_X1 U12960 ( .A1(n15753), .A2(n13316), .B1(n13315), .B2(n14927), .ZN(
        n11086) );
  XNOR2_X1 U12961 ( .A(n11085), .B(n11086), .ZN(n14886) );
  NAND2_X1 U12962 ( .A1(n15748), .A2(n13313), .ZN(n11077) );
  NAND2_X1 U12963 ( .A1(n15235), .A2(n13316), .ZN(n11076) );
  NAND2_X1 U12964 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  XNOR2_X1 U12965 ( .A(n11078), .B(n10643), .ZN(n11081) );
  INV_X1 U12966 ( .A(n11081), .ZN(n11079) );
  AOI22_X1 U12967 ( .A1(n15748), .A2(n13316), .B1(n13315), .B2(n15235), .ZN(
        n11080) );
  NAND2_X1 U12968 ( .A1(n11079), .A2(n11080), .ZN(n11088) );
  INV_X1 U12969 ( .A(n11088), .ZN(n11082) );
  XNOR2_X1 U12970 ( .A(n11081), .B(n11080), .ZN(n14820) );
  OR2_X1 U12971 ( .A1(n11082), .A2(n14820), .ZN(n11084) );
  AND2_X1 U12972 ( .A1(n14886), .A2(n11084), .ZN(n11083) );
  INV_X1 U12973 ( .A(n11084), .ZN(n11090) );
  INV_X1 U12974 ( .A(n11085), .ZN(n11087) );
  NAND2_X1 U12975 ( .A1(n11087), .A2(n11086), .ZN(n14817) );
  AND2_X1 U12976 ( .A1(n14817), .A2(n11088), .ZN(n11089) );
  NAND3_X1 U12977 ( .A1(n12157), .A2(n11415), .A3(n11416), .ZN(n11101) );
  INV_X1 U12978 ( .A(n11237), .ZN(n11091) );
  OR2_X1 U12979 ( .A1(n11101), .A2(n11091), .ZN(n11108) );
  INV_X1 U12980 ( .A(n11108), .ZN(n11095) );
  INV_X1 U12981 ( .A(n11093), .ZN(n11145) );
  NOR2_X1 U12982 ( .A1(n16560), .A2(n11145), .ZN(n11094) );
  INV_X1 U12983 ( .A(n11099), .ZN(n11097) );
  INV_X1 U12984 ( .A(n13253), .ZN(n11098) );
  AOI211_X1 U12985 ( .C1(n11099), .C2(n11096), .A(n16549), .B(n11098), .ZN(
        n11112) );
  OAI21_X2 U12986 ( .B1(n11108), .B2(n16640), .A(n16653), .ZN(n16554) );
  INV_X1 U12987 ( .A(n16554), .ZN(n14918) );
  NOR2_X1 U12988 ( .A1(n15199), .A2(n14918), .ZN(n11111) );
  INV_X1 U12989 ( .A(n11100), .ZN(n11417) );
  NAND2_X1 U12990 ( .A1(n11101), .A2(n11417), .ZN(n11104) );
  INV_X1 U12991 ( .A(n11102), .ZN(n11103) );
  NAND2_X1 U12992 ( .A1(n11104), .A2(n11103), .ZN(n11464) );
  OAI22_X1 U12993 ( .A1(n16558), .A2(n15202), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11105), .ZN(n11110) );
  INV_X1 U12994 ( .A(n11106), .ZN(n11107) );
  NAND2_X1 U12995 ( .A1(n14899), .A2(n15234), .ZN(n16542) );
  NAND2_X1 U12996 ( .A1(n14899), .A2(n15233), .ZN(n16543) );
  OAI22_X1 U12997 ( .A1(n15161), .A2(n16542), .B1(n14888), .B2(n16543), .ZN(
        n11109) );
  AOI211_X1 U12998 ( .C1(n11115), .C2(n11114), .A(n16549), .B(n11113), .ZN(
        n11119) );
  NOR2_X1 U12999 ( .A1(n16543), .A2(n11845), .ZN(n11118) );
  OAI22_X1 U13000 ( .A1(n7943), .A2(n14918), .B1(n16542), .B2(n12570), .ZN(
        n11117) );
  NAND2_X1 U13001 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n15002) );
  OAI21_X1 U13002 ( .B1(n16558), .B2(n12184), .A(n15002), .ZN(n11116) );
  OR4_X1 U13003 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        P1_U3239) );
  AOI211_X1 U13004 ( .C1(n11121), .C2(n11120), .A(n16549), .B(n8205), .ZN(
        n11125) );
  NOR2_X1 U13005 ( .A1(n14918), .A2(n12162), .ZN(n11124) );
  NAND2_X1 U13006 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n15014) );
  OAI21_X1 U13007 ( .B1(n16558), .B2(n12234), .A(n15014), .ZN(n11123) );
  OAI22_X1 U13008 ( .A1(n12166), .A2(n16543), .B1(n16542), .B2(n12888), .ZN(
        n11122) );
  OR4_X1 U13009 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        P1_U3213) );
  INV_X1 U13010 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n11126) );
  MUX2_X1 U13011 ( .A(n11126), .B(P1_REG1_REG_1__SCAN_IN), .S(n11190), .Z(
        n14947) );
  AND2_X1 U13012 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14948) );
  NAND2_X1 U13013 ( .A1(n14947), .A2(n14948), .ZN(n14946) );
  NAND2_X1 U13014 ( .A1(n14949), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U13015 ( .A1(n14946), .A2(n11127), .ZN(n14968) );
  INV_X1 U13016 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n11128) );
  MUX2_X1 U13017 ( .A(n11128), .B(P1_REG1_REG_2__SCAN_IN), .S(n11185), .Z(
        n14969) );
  NAND2_X1 U13018 ( .A1(n14968), .A2(n14969), .ZN(n14982) );
  NAND2_X1 U13019 ( .A1(n14965), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14981) );
  NAND2_X1 U13020 ( .A1(n14982), .A2(n14981), .ZN(n11131) );
  MUX2_X1 U13021 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n11129), .S(n14979), .Z(
        n11130) );
  NAND2_X1 U13022 ( .A1(n11131), .A2(n11130), .ZN(n16280) );
  NAND2_X1 U13023 ( .A1(n14979), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n16279) );
  NAND2_X1 U13024 ( .A1(n16280), .A2(n16279), .ZN(n11134) );
  MUX2_X1 U13025 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n11132), .S(n16284), .Z(
        n11133) );
  NAND2_X1 U13026 ( .A1(n11134), .A2(n11133), .ZN(n16282) );
  NAND2_X1 U13027 ( .A1(n16284), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n11135) );
  AND2_X1 U13028 ( .A1(n16282), .A2(n11135), .ZN(n14991) );
  MUX2_X1 U13029 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9250), .S(n14994), .Z(
        n14992) );
  NAND2_X1 U13030 ( .A1(n14991), .A2(n14992), .ZN(n14990) );
  OR2_X1 U13031 ( .A1(n14994), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11136) );
  AND2_X1 U13032 ( .A1(n14990), .A2(n11136), .ZN(n15005) );
  INV_X1 U13033 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11137) );
  MUX2_X1 U13034 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n11137), .S(n15006), .Z(
        n15004) );
  NAND2_X1 U13035 ( .A1(n15005), .A2(n15004), .ZN(n15025) );
  NAND2_X1 U13036 ( .A1(n15006), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n15024) );
  NAND2_X1 U13037 ( .A1(n15025), .A2(n15024), .ZN(n11139) );
  MUX2_X1 U13038 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15022), .S(n15021), .Z(
        n11138) );
  NAND2_X1 U13039 ( .A1(n11139), .A2(n11138), .ZN(n15027) );
  NAND2_X1 U13040 ( .A1(n15021), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U13041 ( .A1(n15027), .A2(n11140), .ZN(n11256) );
  MUX2_X1 U13042 ( .A(n11141), .B(P1_REG1_REG_8__SCAN_IN), .S(n11260), .Z(
        n11257) );
  OR2_X1 U13043 ( .A1(n11256), .A2(n11257), .ZN(n11270) );
  OR2_X1 U13044 ( .A1(n11260), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U13045 ( .A1(n11270), .A2(n11268), .ZN(n11142) );
  INV_X1 U13046 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n12316) );
  MUX2_X1 U13047 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n12316), .S(n11275), .Z(
        n11267) );
  NAND2_X1 U13048 ( .A1(n11142), .A2(n11267), .ZN(n11272) );
  INV_X1 U13049 ( .A(n11275), .ZN(n11245) );
  NAND2_X1 U13050 ( .A1(n11245), .A2(n12316), .ZN(n11143) );
  NAND2_X1 U13051 ( .A1(n11272), .A2(n11143), .ZN(n11149) );
  INV_X1 U13052 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n12509) );
  MUX2_X1 U13053 ( .A(n12509), .B(P1_REG1_REG_10__SCAN_IN), .S(n11353), .Z(
        n11148) );
  AOI21_X1 U13054 ( .B1(n11145), .B2(n11146), .A(n7442), .ZN(n11175) );
  AOI21_X1 U13055 ( .B1(n11146), .B2(n10969), .A(P1_U3086), .ZN(n11176) );
  AND2_X1 U13056 ( .A1(n11175), .A2(n11176), .ZN(n13023) );
  NAND2_X1 U13057 ( .A1(n13023), .A2(n14954), .ZN(n13030) );
  OR2_X1 U13058 ( .A1(n11149), .A2(n11148), .ZN(n11355) );
  INV_X1 U13059 ( .A(n11355), .ZN(n11147) );
  AOI211_X1 U13060 ( .C1(n11149), .C2(n11148), .A(n13030), .B(n11147), .ZN(
        n11182) );
  MUX2_X1 U13061 ( .A(n11150), .B(P1_REG2_REG_1__SCAN_IN), .S(n11190), .Z(
        n14945) );
  AND2_X1 U13062 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14956) );
  NAND2_X1 U13063 ( .A1(n14945), .A2(n14956), .ZN(n14944) );
  NAND2_X1 U13064 ( .A1(n14949), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U13065 ( .A1(n14944), .A2(n11151), .ZN(n14966) );
  MUX2_X1 U13066 ( .A(n11152), .B(P1_REG2_REG_2__SCAN_IN), .S(n11185), .Z(
        n14967) );
  NAND2_X1 U13067 ( .A1(n14966), .A2(n14967), .ZN(n14977) );
  NAND2_X1 U13068 ( .A1(n14965), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14976) );
  NAND2_X1 U13069 ( .A1(n14977), .A2(n14976), .ZN(n11155) );
  MUX2_X1 U13070 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11153), .S(n14979), .Z(
        n11154) );
  NAND2_X1 U13071 ( .A1(n11155), .A2(n11154), .ZN(n16274) );
  NAND2_X1 U13072 ( .A1(n14979), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n16273) );
  NAND2_X1 U13073 ( .A1(n16274), .A2(n16273), .ZN(n11158) );
  MUX2_X1 U13074 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11156), .S(n16284), .Z(
        n11157) );
  NAND2_X1 U13075 ( .A1(n11158), .A2(n11157), .ZN(n16276) );
  NAND2_X1 U13076 ( .A1(n16284), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U13077 ( .A1(n16276), .A2(n14997), .ZN(n11160) );
  INV_X1 U13078 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n14995) );
  MUX2_X1 U13079 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n14995), .S(n14994), .Z(
        n11159) );
  NAND2_X1 U13080 ( .A1(n11160), .A2(n11159), .ZN(n15009) );
  NAND2_X1 U13081 ( .A1(n14994), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n15008) );
  NAND2_X1 U13082 ( .A1(n15009), .A2(n15008), .ZN(n11163) );
  MUX2_X1 U13083 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11161), .S(n15006), .Z(
        n11162) );
  NAND2_X1 U13084 ( .A1(n11163), .A2(n11162), .ZN(n15018) );
  NAND2_X1 U13085 ( .A1(n15006), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n15017) );
  NAND2_X1 U13086 ( .A1(n15018), .A2(n15017), .ZN(n11166) );
  MUX2_X1 U13087 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11164), .S(n15021), .Z(
        n11165) );
  NAND2_X1 U13088 ( .A1(n11166), .A2(n11165), .ZN(n15020) );
  NAND2_X1 U13089 ( .A1(n15021), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U13090 ( .A1(n15020), .A2(n11262), .ZN(n11169) );
  MUX2_X1 U13091 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11167), .S(n11260), .Z(
        n11168) );
  NAND2_X1 U13092 ( .A1(n11169), .A2(n11168), .ZN(n11279) );
  NAND2_X1 U13093 ( .A1(n11260), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11278) );
  MUX2_X1 U13094 ( .A(n12199), .B(P1_REG2_REG_9__SCAN_IN), .S(n11275), .Z(
        n11277) );
  AOI21_X1 U13095 ( .B1(n11279), .B2(n11278), .A(n11277), .ZN(n11276) );
  NOR2_X1 U13096 ( .A1(n11245), .A2(n12199), .ZN(n11172) );
  MUX2_X1 U13097 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12362), .S(n11353), .Z(
        n11171) );
  OAI21_X1 U13098 ( .B1(n11276), .B2(n11172), .A(n11171), .ZN(n11351) );
  INV_X1 U13099 ( .A(n11351), .ZN(n11174) );
  NOR2_X1 U13100 ( .A1(n9908), .A2(n14954), .ZN(n11170) );
  NAND2_X1 U13101 ( .A1(n13023), .A2(n11170), .ZN(n13028) );
  NOR3_X1 U13102 ( .A1(n11276), .A2(n11172), .A3(n11171), .ZN(n11173) );
  NOR3_X1 U13103 ( .A1(n11174), .A2(n13028), .A3(n11173), .ZN(n11181) );
  NAND2_X1 U13104 ( .A1(n13023), .A2(n9908), .ZN(n13026) );
  INV_X1 U13105 ( .A(n11353), .ZN(n11286) );
  NOR2_X1 U13106 ( .A1(n13026), .A2(n11286), .ZN(n11180) );
  INV_X1 U13107 ( .A(n11175), .ZN(n11177) );
  INV_X1 U13108 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U13109 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12922)
         );
  OAI21_X1 U13110 ( .B1(n15046), .B2(n11178), .A(n12922), .ZN(n11179) );
  OR4_X1 U13111 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(
        P1_U3253) );
  MUX2_X1 U13112 ( .A(P2_RD_REG_SCAN_IN), .B(n8433), .S(P1_RD_REG_SCAN_IN), 
        .Z(n11184) );
  INV_X1 U13113 ( .A(P3_RD_REG_SCAN_IN), .ZN(n11183) );
  NAND2_X1 U13114 ( .A1(n11184), .A2(n11183), .ZN(U29) );
  NAND2_X2 U13115 ( .A1(n11209), .A2(P1_U3086), .ZN(n15810) );
  INV_X1 U13116 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n11186) );
  OAI222_X1 U13117 ( .A1(n15810), .A2(n11186), .B1(n15805), .B2(n11216), .C1(
        n11185), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U13118 ( .A(n11187), .ZN(n11214) );
  INV_X1 U13119 ( .A(n14979), .ZN(n11188) );
  OAI222_X1 U13120 ( .A1(n15810), .A2(n7593), .B1(n15805), .B2(n11214), .C1(
        P1_U3086), .C2(n11188), .ZN(P1_U3352) );
  OAI222_X1 U13121 ( .A1(n15810), .A2(n9137), .B1(n15805), .B2(n9974), .C1(
        n11190), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U13122 ( .A(n16284), .ZN(n11192) );
  OAI222_X1 U13123 ( .A1(P1_U3086), .A2(n11192), .B1(n15805), .B2(n8178), .C1(
        n9207), .C2(n15810), .ZN(P1_U3351) );
  INV_X1 U13124 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n11194) );
  INV_X1 U13125 ( .A(n14994), .ZN(n11193) );
  OAI222_X1 U13126 ( .A1(n15810), .A2(n11194), .B1(n15805), .B2(n11210), .C1(
        n11193), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X2 U13127 ( .A(n14212), .ZN(n14221) );
  NAND2_X2 U13128 ( .A1(n11209), .A2(P3_U3151), .ZN(n14223) );
  OAI222_X1 U13129 ( .A1(n11738), .A2(P3_U3151), .B1(n14221), .B2(n11195), 
        .C1(n15502), .C2(n14223), .ZN(P3_U3294) );
  OAI222_X1 U13130 ( .A1(P3_U3151), .A2(n16108), .B1(n14221), .B2(n11197), 
        .C1(n11196), .C2(n14223), .ZN(P3_U3289) );
  INV_X1 U13131 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n11199) );
  INV_X1 U13132 ( .A(n15006), .ZN(n11198) );
  OAI222_X1 U13133 ( .A1(n15810), .A2(n11199), .B1(n15805), .B2(n11253), .C1(
        n11198), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U13134 ( .A(n15021), .ZN(n11200) );
  OAI222_X1 U13135 ( .A1(n15810), .A2(n11288), .B1(n15805), .B2(n11212), .C1(
        n11200), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U13136 ( .A(n11201), .ZN(n11202) );
  OAI222_X1 U13137 ( .A1(P3_U3151), .A2(n12101), .B1(n14223), .B2(n15306), 
        .C1(n14221), .C2(n11202), .ZN(P3_U3288) );
  INV_X1 U13138 ( .A(SI_9_), .ZN(n11205) );
  INV_X1 U13139 ( .A(n11203), .ZN(n11204) );
  OAI222_X1 U13140 ( .A1(P3_U3151), .A2(n12681), .B1(n14223), .B2(n11205), 
        .C1(n14221), .C2(n11204), .ZN(P3_U3286) );
  OAI222_X1 U13141 ( .A1(n14221), .A2(n11207), .B1(n14223), .B2(n11206), .C1(
        P3_U3151), .C2(n12283), .ZN(P3_U3287) );
  NAND2_X2 U13142 ( .A1(n11209), .A2(P2_U3088), .ZN(n14775) );
  INV_X1 U13143 ( .A(n14424), .ZN(n14417) );
  OAI222_X1 U13144 ( .A1(n14792), .A2(n11211), .B1(n14775), .B2(n11210), .C1(
        n14417), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U13145 ( .A(n11366), .ZN(n11337) );
  OAI222_X1 U13146 ( .A1(n14792), .A2(n11213), .B1(n14775), .B2(n11212), .C1(
        n11337), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U13147 ( .A(n14391), .ZN(n11317) );
  OAI222_X1 U13148 ( .A1(n14792), .A2(n11215), .B1(n14775), .B2(n11214), .C1(
        P2_U3088), .C2(n11317), .ZN(P2_U3324) );
  OAI222_X1 U13149 ( .A1(n14792), .A2(n11217), .B1(n14775), .B2(n11216), .C1(
        n11316), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U13150 ( .A(n11218), .ZN(n11220) );
  INV_X1 U13151 ( .A(SI_5_), .ZN(n11219) );
  OAI222_X1 U13152 ( .A1(n11942), .A2(P3_U3151), .B1(n14221), .B2(n11220), 
        .C1(n11219), .C2(n14223), .ZN(P3_U3290) );
  INV_X1 U13153 ( .A(n11792), .ZN(n11801) );
  INV_X1 U13154 ( .A(n11221), .ZN(n11223) );
  INV_X1 U13155 ( .A(SI_4_), .ZN(n11222) );
  OAI222_X1 U13156 ( .A1(n11801), .A2(P3_U3151), .B1(n14221), .B2(n11223), 
        .C1(n11222), .C2(n14223), .ZN(P3_U3291) );
  INV_X1 U13157 ( .A(n11224), .ZN(n11225) );
  OAI222_X1 U13158 ( .A1(n11771), .A2(P3_U3151), .B1(n14221), .B2(n11225), 
        .C1(n15308), .C2(n14223), .ZN(P3_U3293) );
  INV_X1 U13159 ( .A(n11838), .ZN(n11777) );
  INV_X1 U13160 ( .A(n11226), .ZN(n11227) );
  INV_X1 U13161 ( .A(SI_3_), .ZN(n15309) );
  OAI222_X1 U13162 ( .A1(n11777), .A2(P3_U3151), .B1(n14221), .B2(n11227), 
        .C1(n15309), .C2(n14223), .ZN(P3_U3292) );
  INV_X1 U13163 ( .A(n13762), .ZN(n13717) );
  INV_X1 U13164 ( .A(SI_10_), .ZN(n11230) );
  INV_X1 U13165 ( .A(n11228), .ZN(n11229) );
  OAI222_X1 U13166 ( .A1(P3_U3151), .A2(n13717), .B1(n14223), .B2(n11230), 
        .C1(n14221), .C2(n11229), .ZN(P3_U3285) );
  INV_X1 U13167 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11231) );
  AOI21_X1 U13168 ( .B1(n13024), .B2(n11231), .A(n9908), .ZN(n14961) );
  OAI21_X1 U13169 ( .B1(n13024), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14961), .ZN(
        n11232) );
  XNOR2_X1 U13170 ( .A(n11232), .B(P1_IR_REG_0__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U13171 ( .A1(n13023), .A2(n11233), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11234) );
  OAI21_X1 U13172 ( .B1(n15046), .B2(n7668), .A(n11234), .ZN(P1_U3243) );
  NAND2_X2 U13173 ( .A1(n11237), .A2(n11235), .ZN(n15814) );
  AOI22_X1 U13174 ( .A1(n15814), .A2(n11238), .B1(n11237), .B2(n11236), .ZN(
        P1_U3446) );
  INV_X1 U13175 ( .A(n11260), .ZN(n11240) );
  INV_X1 U13176 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n11239) );
  OAI222_X1 U13177 ( .A1(P1_U3086), .A2(n11240), .B1(n15805), .B2(n11248), 
        .C1(n11239), .C2(n15810), .ZN(P1_U3347) );
  NAND2_X1 U13178 ( .A1(n15814), .A2(P1_D_REG_0__SCAN_IN), .ZN(n11241) );
  OAI21_X1 U13179 ( .B1(n15814), .B2(n11242), .A(n11241), .ZN(P1_U3445) );
  OAI222_X1 U13180 ( .A1(n14792), .A2(n8454), .B1(n14775), .B2(n9974), .C1(
        n11313), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U13181 ( .A(n11243), .ZN(n11244) );
  OAI222_X1 U13182 ( .A1(P3_U3151), .A2(n16134), .B1(n14223), .B2(n15493), 
        .C1(n14221), .C2(n11244), .ZN(P3_U3284) );
  OAI222_X1 U13183 ( .A1(n15810), .A2(n11246), .B1(n15805), .B2(n11251), .C1(
        n11245), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U13184 ( .A(n11423), .ZN(n11430) );
  OAI222_X1 U13185 ( .A1(P2_U3088), .A2(n11430), .B1(n14775), .B2(n11248), 
        .C1(n11247), .C2(n14792), .ZN(P2_U3319) );
  OAI222_X1 U13186 ( .A1(P2_U3088), .A2(n11319), .B1(n14775), .B2(n8178), .C1(
        n11249), .C2(n14792), .ZN(P2_U3323) );
  INV_X1 U13187 ( .A(n15923), .ZN(n11431) );
  OAI222_X1 U13188 ( .A1(P2_U3088), .A2(n11431), .B1(n14775), .B2(n11251), 
        .C1(n11250), .C2(n14792), .ZN(P2_U3318) );
  INV_X1 U13189 ( .A(n11297), .ZN(n11330) );
  OAI222_X1 U13190 ( .A1(P2_U3088), .A2(n11330), .B1(n14775), .B2(n11253), 
        .C1(n11252), .C2(n14792), .ZN(P2_U3321) );
  INV_X1 U13191 ( .A(n13741), .ZN(n16152) );
  OAI222_X1 U13192 ( .A1(P3_U3151), .A2(n16152), .B1(n14223), .B2(n15487), 
        .C1(n14221), .C2(n11254), .ZN(P3_U3283) );
  INV_X1 U13193 ( .A(n11270), .ZN(n11255) );
  AOI21_X1 U13194 ( .B1(n11257), .B2(n11256), .A(n11255), .ZN(n11266) );
  NAND2_X1 U13195 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11258) );
  OAI21_X1 U13196 ( .B1(n15046), .B2(n15992), .A(n11258), .ZN(n11259) );
  AOI21_X1 U13197 ( .B1(n16285), .B2(n11260), .A(n11259), .ZN(n11265) );
  MUX2_X1 U13198 ( .A(n11167), .B(P1_REG2_REG_8__SCAN_IN), .S(n11260), .Z(
        n11261) );
  NAND3_X1 U13199 ( .A1(n15020), .A2(n11262), .A3(n11261), .ZN(n11263) );
  NAND3_X1 U13200 ( .A1(n16277), .A2(n11279), .A3(n11263), .ZN(n11264) );
  OAI211_X1 U13201 ( .C1(n11266), .C2(n13030), .A(n11265), .B(n11264), .ZN(
        P1_U3251) );
  INV_X1 U13202 ( .A(n11267), .ZN(n11269) );
  NAND3_X1 U13203 ( .A1(n11270), .A2(n11269), .A3(n11268), .ZN(n11271) );
  AND2_X1 U13204 ( .A1(n11272), .A2(n11271), .ZN(n11284) );
  INV_X1 U13205 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11273) );
  NAND2_X1 U13206 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n12885) );
  OAI21_X1 U13207 ( .B1(n15046), .B2(n11273), .A(n12885), .ZN(n11274) );
  AOI21_X1 U13208 ( .B1(n16285), .B2(n11275), .A(n11274), .ZN(n11283) );
  INV_X1 U13209 ( .A(n11276), .ZN(n11281) );
  NAND3_X1 U13210 ( .A1(n11279), .A2(n11278), .A3(n11277), .ZN(n11280) );
  NAND3_X1 U13211 ( .A1(n16277), .A2(n11281), .A3(n11280), .ZN(n11282) );
  OAI211_X1 U13212 ( .C1(n11284), .C2(n13030), .A(n11283), .B(n11282), .ZN(
        P1_U3252) );
  INV_X1 U13213 ( .A(n11474), .ZN(n11470) );
  OAI222_X1 U13214 ( .A1(n14792), .A2(n11285), .B1(n14775), .B2(n11287), .C1(
        n11470), .C2(P2_U3088), .ZN(P2_U3317) );
  OAI222_X1 U13215 ( .A1(n15810), .A2(n11291), .B1(n15805), .B2(n11287), .C1(
        n11286), .C2(P1_U3086), .ZN(P1_U3345) );
  MUX2_X1 U13216 ( .A(n11288), .B(n12247), .S(P2_U3947), .Z(n11289) );
  INV_X1 U13217 ( .A(n11289), .ZN(P2_U3538) );
  MUX2_X1 U13218 ( .A(n11438), .B(n12772), .S(P2_U3947), .Z(n11290) );
  INV_X1 U13219 ( .A(n11290), .ZN(P2_U3543) );
  MUX2_X1 U13220 ( .A(n11291), .B(n12634), .S(P2_U3947), .Z(n11292) );
  INV_X1 U13221 ( .A(n11292), .ZN(P2_U3541) );
  INV_X1 U13222 ( .A(n11313), .ZN(n15832) );
  MUX2_X1 U13223 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9969), .S(n11313), .Z(
        n15839) );
  NAND2_X1 U13224 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15838) );
  NOR2_X1 U13225 ( .A1(n15839), .A2(n15838), .ZN(n15837) );
  AOI21_X1 U13226 ( .B1(n15832), .B2(P2_REG1_REG_1__SCAN_IN), .A(n15837), .ZN(
        n15852) );
  MUX2_X1 U13227 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9986), .S(n11316), .Z(
        n15851) );
  NOR2_X1 U13228 ( .A1(n15852), .A2(n15851), .ZN(n15850) );
  NOR2_X1 U13229 ( .A1(n11316), .A2(n9986), .ZN(n14396) );
  MUX2_X1 U13230 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n11293), .S(n14391), .Z(
        n14395) );
  OAI21_X1 U13231 ( .B1(n15850), .B2(n14396), .A(n14395), .ZN(n14410) );
  NAND2_X1 U13232 ( .A1(n14391), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n14409) );
  MUX2_X1 U13233 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n11294), .S(n11319), .Z(
        n14408) );
  AOI21_X1 U13234 ( .B1(n14410), .B2(n14409), .A(n14408), .ZN(n14430) );
  NOR2_X1 U13235 ( .A1(n11319), .A2(n11294), .ZN(n14425) );
  MUX2_X1 U13236 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n11295), .S(n14424), .Z(
        n11296) );
  OAI21_X1 U13237 ( .B1(n14430), .B2(n14425), .A(n11296), .ZN(n14428) );
  NAND2_X1 U13238 ( .A1(n14424), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11299) );
  INV_X1 U13239 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n16426) );
  MUX2_X1 U13240 ( .A(n16426), .B(P2_REG1_REG_6__SCAN_IN), .S(n11297), .Z(
        n11298) );
  AOI21_X1 U13241 ( .B1(n14428), .B2(n11299), .A(n11298), .ZN(n11336) );
  NAND3_X1 U13242 ( .A1(n14428), .A2(n11299), .A3(n11298), .ZN(n11307) );
  NAND2_X1 U13243 ( .A1(n11501), .A2(n11511), .ZN(n11301) );
  NAND2_X1 U13244 ( .A1(n11301), .A2(n11300), .ZN(n11304) );
  INV_X1 U13245 ( .A(n11302), .ZN(n11303) );
  NAND2_X1 U13246 ( .A1(n11304), .A2(n11303), .ZN(n11310) );
  OR2_X1 U13247 ( .A1(n11308), .A2(P2_U3088), .ZN(n14780) );
  INV_X1 U13248 ( .A(n14780), .ZN(n11305) );
  NAND2_X1 U13249 ( .A1(n11310), .A2(n11305), .ZN(n11321) );
  NOR2_X2 U13250 ( .A1(n11321), .A2(n11306), .ZN(n15920) );
  NAND2_X1 U13251 ( .A1(n11307), .A2(n15920), .ZN(n11326) );
  INV_X1 U13252 ( .A(n15928), .ZN(n15880) );
  NAND2_X1 U13253 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n11655) );
  INV_X1 U13254 ( .A(n11655), .ZN(n11312) );
  AND2_X1 U13255 ( .A1(n11308), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11309) );
  NOR2_X1 U13256 ( .A1(n14418), .A2(n11330), .ZN(n11311) );
  AOI211_X1 U13257 ( .C1(n15880), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n11312), .B(
        n11311), .ZN(n11325) );
  XNOR2_X1 U13258 ( .A(n11330), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n11323) );
  MUX2_X1 U13259 ( .A(n12058), .B(P2_REG2_REG_1__SCAN_IN), .S(n11313), .Z(
        n15830) );
  AND2_X1 U13260 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15829) );
  NAND2_X1 U13261 ( .A1(n15830), .A2(n15829), .ZN(n15828) );
  NAND2_X1 U13262 ( .A1(n15832), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U13263 ( .A1(n15828), .A2(n11314), .ZN(n15844) );
  MUX2_X1 U13264 ( .A(n11315), .B(P2_REG2_REG_2__SCAN_IN), .S(n11316), .Z(
        n15845) );
  NAND2_X1 U13265 ( .A1(n15844), .A2(n15845), .ZN(n15843) );
  OAI21_X1 U13266 ( .B1(n11316), .B2(n11315), .A(n15843), .ZN(n14393) );
  MUX2_X1 U13267 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n12044), .S(n14391), .Z(
        n14394) );
  NAND2_X1 U13268 ( .A1(n14393), .A2(n14394), .ZN(n14392) );
  OAI21_X1 U13269 ( .B1(n12044), .B2(n11317), .A(n14392), .ZN(n14406) );
  XNOR2_X1 U13270 ( .A(n11319), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U13271 ( .A1(n14406), .A2(n14407), .ZN(n14405) );
  OAI21_X1 U13272 ( .B1(n11319), .B2(n11318), .A(n14405), .ZN(n14422) );
  MUX2_X1 U13273 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11320), .S(n14424), .Z(
        n14423) );
  NAND2_X1 U13274 ( .A1(n14422), .A2(n14423), .ZN(n14421) );
  OAI21_X1 U13275 ( .B1(n11320), .B2(n14417), .A(n14421), .ZN(n11322) );
  INV_X1 U13276 ( .A(n15897), .ZN(n15924) );
  NAND2_X1 U13277 ( .A1(n11322), .A2(n11323), .ZN(n11327) );
  OAI211_X1 U13278 ( .C1(n11323), .C2(n11322), .A(n15924), .B(n11327), .ZN(
        n11324) );
  OAI211_X1 U13279 ( .C1(n11336), .C2(n11326), .A(n11325), .B(n11324), .ZN(
        P2_U3220) );
  OAI21_X1 U13280 ( .B1(n11330), .B2(n12260), .A(n11327), .ZN(n11329) );
  MUX2_X1 U13281 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n12086), .S(n11366), .Z(
        n11328) );
  AND2_X1 U13282 ( .A1(n11329), .A2(n11328), .ZN(n11363) );
  OAI21_X1 U13283 ( .B1(n11329), .B2(n11328), .A(n15924), .ZN(n11342) );
  NOR2_X1 U13284 ( .A1(n11330), .A2(n16426), .ZN(n11334) );
  INV_X1 U13285 ( .A(n11334), .ZN(n11332) );
  INV_X1 U13286 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n12150) );
  MUX2_X1 U13287 ( .A(n12150), .B(P2_REG1_REG_7__SCAN_IN), .S(n11366), .Z(
        n11331) );
  NAND2_X1 U13288 ( .A1(n11332), .A2(n11331), .ZN(n11335) );
  MUX2_X1 U13289 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n12150), .S(n11366), .Z(
        n11333) );
  OAI21_X1 U13290 ( .B1(n11336), .B2(n11334), .A(n11333), .ZN(n11369) );
  OAI211_X1 U13291 ( .C1(n11336), .C2(n11335), .A(n11369), .B(n15920), .ZN(
        n11341) );
  NAND2_X1 U13292 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11971) );
  INV_X1 U13293 ( .A(n11971), .ZN(n11339) );
  NOR2_X1 U13294 ( .A1(n14418), .A2(n11337), .ZN(n11338) );
  AOI211_X1 U13295 ( .C1(n15880), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n11339), .B(
        n11338), .ZN(n11340) );
  OAI211_X1 U13296 ( .C1(n11363), .C2(n11342), .A(n11341), .B(n11340), .ZN(
        P2_U3221) );
  OAI222_X1 U13297 ( .A1(P3_U3151), .A2(n13776), .B1(n14223), .B2(n15488), 
        .C1(n14221), .C2(n11343), .ZN(P3_U3282) );
  INV_X1 U13298 ( .A(n11344), .ZN(n11347) );
  INV_X1 U13299 ( .A(n11450), .ZN(n11345) );
  OAI222_X1 U13300 ( .A1(n15810), .A2(n11346), .B1(n15805), .B2(n11347), .C1(
        P1_U3086), .C2(n11345), .ZN(P1_U3344) );
  INV_X1 U13301 ( .A(n11874), .ZN(n11862) );
  OAI222_X1 U13302 ( .A1(n14792), .A2(n11348), .B1(n14775), .B2(n11347), .C1(
        P2_U3088), .C2(n11862), .ZN(P2_U3316) );
  INV_X1 U13303 ( .A(n15046), .ZN(n16287) );
  NOR2_X1 U13304 ( .A1(n16287), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U13305 ( .A1(n11353), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11350) );
  MUX2_X1 U13306 ( .A(n9389), .B(P1_REG2_REG_11__SCAN_IN), .S(n11450), .Z(
        n11349) );
  AOI21_X1 U13307 ( .B1(n11351), .B2(n11350), .A(n11349), .ZN(n11446) );
  NAND3_X1 U13308 ( .A1(n11351), .A2(n11350), .A3(n11349), .ZN(n11352) );
  NAND2_X1 U13309 ( .A1(n16277), .A2(n11352), .ZN(n11362) );
  MUX2_X1 U13310 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9388), .S(n11450), .Z(
        n11357) );
  NAND2_X1 U13311 ( .A1(n11353), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11354) );
  AND2_X1 U13312 ( .A1(n11355), .A2(n11354), .ZN(n11356) );
  NAND2_X1 U13313 ( .A1(n11356), .A2(n11357), .ZN(n11455) );
  OAI21_X1 U13314 ( .B1(n11357), .B2(n11356), .A(n11455), .ZN(n11358) );
  INV_X1 U13315 ( .A(n13030), .ZN(n16283) );
  NAND2_X1 U13316 ( .A1(n11358), .A2(n16283), .ZN(n11361) );
  NAND2_X1 U13317 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n13045)
         );
  OAI21_X1 U13318 ( .B1(n15046), .B2(n16017), .A(n13045), .ZN(n11359) );
  AOI21_X1 U13319 ( .B1(n16285), .B2(n11450), .A(n11359), .ZN(n11360) );
  OAI211_X1 U13320 ( .C1(n11446), .C2(n11362), .A(n11361), .B(n11360), .ZN(
        P1_U3254) );
  AOI21_X1 U13321 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n11366), .A(n11363), .ZN(
        n11365) );
  XNOR2_X1 U13322 ( .A(n11423), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n11364) );
  NOR2_X1 U13323 ( .A1(n11365), .A2(n11364), .ZN(n15914) );
  AOI211_X1 U13324 ( .C1(n11365), .C2(n11364), .A(n15897), .B(n15914), .ZN(
        n11375) );
  NAND2_X1 U13325 ( .A1(n11366), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11368) );
  MUX2_X1 U13326 ( .A(n10068), .B(P2_REG1_REG_8__SCAN_IN), .S(n11423), .Z(
        n11367) );
  AOI21_X1 U13327 ( .B1(n11369), .B2(n11368), .A(n11367), .ZN(n11422) );
  AND3_X1 U13328 ( .A1(n11369), .A2(n11368), .A3(n11367), .ZN(n11370) );
  INV_X1 U13329 ( .A(n15920), .ZN(n15903) );
  NOR3_X1 U13330 ( .A1(n11422), .A2(n11370), .A3(n15903), .ZN(n11374) );
  NAND2_X1 U13331 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11982) );
  INV_X1 U13332 ( .A(n11982), .ZN(n11371) );
  AOI21_X1 U13333 ( .B1(n15880), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n11371), .ZN(
        n11372) );
  OAI21_X1 U13334 ( .B1(n11430), .B2(n14418), .A(n11372), .ZN(n11373) );
  OR3_X1 U13335 ( .A1(n11375), .A2(n11374), .A3(n11373), .ZN(P2_U3222) );
  INV_X1 U13336 ( .A(n14210), .ZN(n11377) );
  CLKBUF_X1 U13337 ( .A(n11382), .Z(n11408) );
  INV_X1 U13338 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n11378) );
  NOR2_X1 U13339 ( .A1(n11408), .A2(n11378), .ZN(P3_U3248) );
  INV_X1 U13340 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n11379) );
  NOR2_X1 U13341 ( .A1(n11408), .A2(n11379), .ZN(P3_U3252) );
  INV_X1 U13342 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n11380) );
  NOR2_X1 U13343 ( .A1(n11408), .A2(n11380), .ZN(P3_U3253) );
  INV_X1 U13344 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n11381) );
  NOR2_X1 U13345 ( .A1(n11408), .A2(n11381), .ZN(P3_U3254) );
  INV_X1 U13346 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n11383) );
  NOR2_X1 U13347 ( .A1(n11408), .A2(n11383), .ZN(P3_U3234) );
  INV_X1 U13348 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n11384) );
  NOR2_X1 U13349 ( .A1(n11382), .A2(n11384), .ZN(P3_U3235) );
  INV_X1 U13350 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n11385) );
  NOR2_X1 U13351 ( .A1(n11382), .A2(n11385), .ZN(P3_U3236) );
  INV_X1 U13352 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n11386) );
  NOR2_X1 U13353 ( .A1(n11382), .A2(n11386), .ZN(P3_U3237) );
  INV_X1 U13354 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n11387) );
  NOR2_X1 U13355 ( .A1(n11382), .A2(n11387), .ZN(P3_U3238) );
  INV_X1 U13356 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n11388) );
  NOR2_X1 U13357 ( .A1(n11382), .A2(n11388), .ZN(P3_U3239) );
  INV_X1 U13358 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n11389) );
  NOR2_X1 U13359 ( .A1(n11382), .A2(n11389), .ZN(P3_U3240) );
  INV_X1 U13360 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n11390) );
  NOR2_X1 U13361 ( .A1(n11382), .A2(n11390), .ZN(P3_U3241) );
  INV_X1 U13362 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n11391) );
  NOR2_X1 U13363 ( .A1(n11382), .A2(n11391), .ZN(P3_U3242) );
  INV_X1 U13364 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n11392) );
  NOR2_X1 U13365 ( .A1(n11382), .A2(n11392), .ZN(P3_U3243) );
  INV_X1 U13366 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n11393) );
  NOR2_X1 U13367 ( .A1(n11382), .A2(n11393), .ZN(P3_U3244) );
  INV_X1 U13368 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n11394) );
  NOR2_X1 U13369 ( .A1(n11382), .A2(n11394), .ZN(P3_U3245) );
  INV_X1 U13370 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n11395) );
  NOR2_X1 U13371 ( .A1(n11408), .A2(n11395), .ZN(P3_U3246) );
  INV_X1 U13372 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n11396) );
  NOR2_X1 U13373 ( .A1(n11408), .A2(n11396), .ZN(P3_U3247) );
  INV_X1 U13374 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n11397) );
  NOR2_X1 U13375 ( .A1(n11408), .A2(n11397), .ZN(P3_U3257) );
  INV_X1 U13376 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n11398) );
  NOR2_X1 U13377 ( .A1(n11408), .A2(n11398), .ZN(P3_U3249) );
  INV_X1 U13378 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n11399) );
  NOR2_X1 U13379 ( .A1(n11408), .A2(n11399), .ZN(P3_U3250) );
  INV_X1 U13380 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n11400) );
  NOR2_X1 U13381 ( .A1(n11408), .A2(n11400), .ZN(P3_U3251) );
  INV_X1 U13382 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n11401) );
  NOR2_X1 U13383 ( .A1(n11408), .A2(n11401), .ZN(P3_U3261) );
  INV_X1 U13384 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n11402) );
  NOR2_X1 U13385 ( .A1(n11408), .A2(n11402), .ZN(P3_U3262) );
  INV_X1 U13386 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n11403) );
  NOR2_X1 U13387 ( .A1(n11408), .A2(n11403), .ZN(P3_U3263) );
  INV_X1 U13388 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n11404) );
  NOR2_X1 U13389 ( .A1(n11408), .A2(n11404), .ZN(P3_U3255) );
  INV_X1 U13390 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n11405) );
  NOR2_X1 U13391 ( .A1(n11408), .A2(n11405), .ZN(P3_U3256) );
  INV_X1 U13392 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n11406) );
  NOR2_X1 U13393 ( .A1(n11408), .A2(n11406), .ZN(P3_U3258) );
  INV_X1 U13394 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n11407) );
  NOR2_X1 U13395 ( .A1(n11408), .A2(n11407), .ZN(P3_U3259) );
  INV_X1 U13396 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n11409) );
  NOR2_X1 U13397 ( .A1(n11408), .A2(n11409), .ZN(P3_U3260) );
  OAI222_X1 U13398 ( .A1(P3_U3151), .A2(n16185), .B1(n14223), .B2(n11411), 
        .C1(n14221), .C2(n11410), .ZN(P3_U3281) );
  NOR2_X1 U13399 ( .A1(n11092), .A2(n16310), .ZN(n16299) );
  NAND2_X1 U13400 ( .A1(n16324), .A2(n16351), .ZN(n11413) );
  AOI22_X1 U13401 ( .A1(n11413), .A2(n16296), .B1(n15234), .B2(n10603), .ZN(
        n16302) );
  INV_X1 U13402 ( .A(n16302), .ZN(n11414) );
  AOI211_X1 U13403 ( .C1(n16452), .C2(n16296), .A(n16299), .B(n11414), .ZN(
        n16294) );
  INV_X1 U13404 ( .A(n11415), .ZN(n11418) );
  NAND4_X1 U13405 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n12158) );
  NAND2_X1 U13406 ( .A1(n16633), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11421) );
  OAI21_X1 U13407 ( .B1(n16294), .B2(n16633), .A(n11421), .ZN(P1_U3528) );
  AOI21_X1 U13408 ( .B1(n11423), .B2(P2_REG1_REG_8__SCAN_IN), .A(n11422), .ZN(
        n15919) );
  INV_X1 U13409 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11424) );
  MUX2_X1 U13410 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11424), .S(n15923), .Z(
        n15918) );
  NAND2_X1 U13411 ( .A1(n15919), .A2(n15918), .ZN(n15917) );
  OAI21_X1 U13412 ( .B1(n15923), .B2(P2_REG1_REG_9__SCAN_IN), .A(n15917), .ZN(
        n11426) );
  INV_X1 U13413 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n16480) );
  MUX2_X1 U13414 ( .A(n16480), .B(P2_REG1_REG_10__SCAN_IN), .S(n11474), .Z(
        n11425) );
  OR2_X1 U13415 ( .A1(n11426), .A2(n11425), .ZN(n11477) );
  INV_X1 U13416 ( .A(n11477), .ZN(n11481) );
  AOI211_X1 U13417 ( .C1(n11426), .C2(n11425), .A(n15903), .B(n11481), .ZN(
        n11429) );
  AND2_X1 U13418 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n12477) );
  AOI21_X1 U13419 ( .B1(n15880), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n12477), 
        .ZN(n11427) );
  OAI21_X1 U13420 ( .B1(n11470), .B2(n14418), .A(n11427), .ZN(n11428) );
  NOR2_X1 U13421 ( .A1(n11429), .A2(n11428), .ZN(n11435) );
  NOR2_X1 U13422 ( .A1(n11430), .A2(n12137), .ZN(n15913) );
  XNOR2_X1 U13423 ( .A(n15923), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n15912) );
  NOR3_X1 U13424 ( .A1(n15914), .A2(n15913), .A3(n15912), .ZN(n15911) );
  AOI21_X1 U13425 ( .B1(n11431), .B2(n12207), .A(n15911), .ZN(n11433) );
  MUX2_X1 U13426 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n12379), .S(n11474), .Z(
        n11432) );
  NAND2_X1 U13427 ( .A1(n11433), .A2(n11432), .ZN(n11469) );
  OAI211_X1 U13428 ( .C1(n11433), .C2(n11432), .A(n11469), .B(n15924), .ZN(
        n11434) );
  NAND2_X1 U13429 ( .A1(n11435), .A2(n11434), .ZN(P2_U3224) );
  INV_X1 U13430 ( .A(n11436), .ZN(n11439) );
  INV_X1 U13431 ( .A(n11558), .ZN(n11437) );
  OAI222_X1 U13432 ( .A1(n15810), .A2(n11438), .B1(n15805), .B2(n11439), .C1(
        n11437), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U13433 ( .A1(n14792), .A2(n11440), .B1(n14775), .B2(n11439), .C1(
        n15896), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13434 ( .A(n16197), .ZN(n13785) );
  OAI222_X1 U13435 ( .A1(n14223), .A2(n11442), .B1(n14221), .B2(n11441), .C1(
        n13785), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U13436 ( .A(n11627), .ZN(n11443) );
  OAI222_X1 U13437 ( .A1(n15810), .A2(n11444), .B1(n15805), .B2(n11445), .C1(
        n11443), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13438 ( .A(n12583), .ZN(n12577) );
  OAI222_X1 U13439 ( .A1(n14792), .A2(n8077), .B1(n14775), .B2(n11445), .C1(
        n12577), .C2(P2_U3088), .ZN(P2_U3314) );
  MUX2_X1 U13440 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12546), .S(n11558), .Z(
        n11448) );
  AOI21_X1 U13441 ( .B1(n11450), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11446), 
        .ZN(n11447) );
  NAND2_X1 U13442 ( .A1(n11447), .A2(n11448), .ZN(n11552) );
  OAI21_X1 U13443 ( .B1(n11448), .B2(n11447), .A(n11552), .ZN(n11459) );
  NAND2_X1 U13444 ( .A1(n16285), .A2(n11558), .ZN(n11449) );
  NAND2_X1 U13445 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n13144)
         );
  OAI211_X1 U13446 ( .C1(n16032), .C2(n15046), .A(n11449), .B(n13144), .ZN(
        n11458) );
  OR2_X1 U13447 ( .A1(n11450), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U13448 ( .A1(n11455), .A2(n11453), .ZN(n11451) );
  MUX2_X1 U13449 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9408), .S(n11558), .Z(
        n11452) );
  NAND2_X1 U13450 ( .A1(n11451), .A2(n11452), .ZN(n11560) );
  INV_X1 U13451 ( .A(n11452), .ZN(n11454) );
  NAND3_X1 U13452 ( .A1(n11455), .A2(n11454), .A3(n11453), .ZN(n11456) );
  AOI21_X1 U13453 ( .B1(n11560), .B2(n11456), .A(n13030), .ZN(n11457) );
  AOI211_X1 U13454 ( .C1(n16277), .C2(n11459), .A(n11458), .B(n11457), .ZN(
        n11460) );
  INV_X1 U13455 ( .A(n11460), .ZN(P1_U3255) );
  XOR2_X1 U13456 ( .A(n11462), .B(n11461), .Z(n14955) );
  INV_X1 U13457 ( .A(n16542), .ZN(n11463) );
  AOI22_X1 U13458 ( .A1(n11463), .A2(n10603), .B1(n9115), .B2(n16554), .ZN(
        n11466) );
  OR2_X1 U13459 ( .A1(n11464), .A2(P1_U3086), .ZN(n11603) );
  NAND2_X1 U13460 ( .A1(n11603), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n11465) );
  OAI211_X1 U13461 ( .C1(n14955), .C2(n16549), .A(n11466), .B(n11465), .ZN(
        P1_U3232) );
  INV_X1 U13462 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U13463 ( .A1(n13585), .A2(P3_U3897), .ZN(n11467) );
  OAI21_X1 U13464 ( .B1(P3_U3897), .B2(n11468), .A(n11467), .ZN(P3_U3491) );
  MUX2_X1 U13465 ( .A(n12452), .B(P2_REG2_REG_11__SCAN_IN), .S(n11874), .Z(
        n11472) );
  OAI21_X1 U13466 ( .B1(n11470), .B2(n12379), .A(n11469), .ZN(n11471) );
  NOR2_X1 U13467 ( .A1(n11471), .A2(n11472), .ZN(n15892) );
  AOI21_X1 U13468 ( .B1(n11472), .B2(n11471), .A(n15892), .ZN(n11484) );
  NAND2_X1 U13469 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n12632)
         );
  OAI21_X1 U13470 ( .B1(n14418), .B2(n11862), .A(n12632), .ZN(n11473) );
  AOI21_X1 U13471 ( .B1(n15880), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n11473), 
        .ZN(n11483) );
  NAND2_X1 U13472 ( .A1(n11474), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11476) );
  INV_X1 U13473 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11863) );
  OR2_X1 U13474 ( .A1(n11874), .A2(n11863), .ZN(n11475) );
  OAI211_X1 U13475 ( .C1(n11862), .C2(P2_REG1_REG_11__SCAN_IN), .A(n11476), 
        .B(n11475), .ZN(n11480) );
  NAND2_X1 U13476 ( .A1(n11477), .A2(n11476), .ZN(n11479) );
  NAND2_X1 U13477 ( .A1(n11874), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11478) );
  OAI211_X1 U13478 ( .C1(n11874), .C2(P2_REG1_REG_11__SCAN_IN), .A(n11479), 
        .B(n11478), .ZN(n11861) );
  OAI211_X1 U13479 ( .C1(n11481), .C2(n11480), .A(n11861), .B(n15920), .ZN(
        n11482) );
  OAI211_X1 U13480 ( .C1(n11484), .C2(n15897), .A(n11483), .B(n11482), .ZN(
        P2_U3225) );
  NAND2_X1 U13481 ( .A1(n14386), .A2(n11533), .ZN(n11487) );
  NAND2_X1 U13482 ( .A1(n11486), .A2(n11487), .ZN(n11498) );
  INV_X1 U13483 ( .A(n11487), .ZN(n11488) );
  XNOR2_X1 U13484 ( .A(n11490), .B(n11668), .ZN(n11494) );
  NAND2_X1 U13485 ( .A1(n7435), .A2(n11533), .ZN(n11495) );
  XNOR2_X1 U13486 ( .A(n11494), .B(n11495), .ZN(n11522) );
  NAND2_X1 U13487 ( .A1(n11490), .A2(n11492), .ZN(n11493) );
  OR2_X1 U13488 ( .A1(n11492), .A2(n11491), .ZN(n11853) );
  AND2_X1 U13489 ( .A1(n11665), .A2(n11853), .ZN(n11534) );
  NAND2_X1 U13490 ( .A1(n11493), .A2(n11534), .ZN(n11521) );
  NAND2_X1 U13491 ( .A1(n11522), .A2(n11521), .ZN(n11520) );
  INV_X1 U13492 ( .A(n11494), .ZN(n11496) );
  NAND2_X1 U13493 ( .A1(n11496), .A2(n11495), .ZN(n11497) );
  NAND2_X1 U13494 ( .A1(n14384), .A2(n11533), .ZN(n11573) );
  XNOR2_X1 U13495 ( .A(n11572), .B(n11573), .ZN(n11577) );
  XNOR2_X1 U13496 ( .A(n11577), .B(n11578), .ZN(n11517) );
  INV_X1 U13497 ( .A(n11499), .ZN(n11500) );
  NOR2_X1 U13498 ( .A1(n16418), .A2(n11501), .ZN(n11502) );
  INV_X1 U13499 ( .A(n14297), .ZN(n14358) );
  AOI22_X1 U13500 ( .A1(n14383), .A2(n14575), .B1(n14578), .B2(n14386), .ZN(
        n11687) );
  INV_X1 U13501 ( .A(n11687), .ZN(n11507) );
  AOI22_X1 U13502 ( .A1(n14358), .A2(n11507), .B1(n14324), .B2(n12045), .ZN(
        n11516) );
  OAI21_X1 U13503 ( .B1(n15822), .B2(n11509), .A(n11508), .ZN(n11514) );
  AND3_X1 U13504 ( .A1(n11512), .A2(n11511), .A3(n11510), .ZN(n11513) );
  NAND2_X1 U13505 ( .A1(n11514), .A2(n11513), .ZN(n11518) );
  MUX2_X1 U13506 ( .A(n14355), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n11515) );
  OAI211_X1 U13507 ( .C1(n11517), .C2(n14326), .A(n11516), .B(n11515), .ZN(
        P2_U3190) );
  NOR2_X1 U13508 ( .A1(n11518), .A2(P2_U3088), .ZN(n11539) );
  AOI22_X1 U13509 ( .A1(n14386), .A2(n14575), .B1(n14578), .B2(n14387), .ZN(
        n11666) );
  INV_X1 U13510 ( .A(n11666), .ZN(n11519) );
  AOI22_X1 U13511 ( .A1(n14358), .A2(n11519), .B1(n14324), .B2(n11668), .ZN(
        n11525) );
  OAI21_X1 U13512 ( .B1(n11522), .B2(n11521), .A(n11520), .ZN(n11523) );
  NAND2_X1 U13513 ( .A1(n14352), .A2(n11523), .ZN(n11524) );
  OAI211_X1 U13514 ( .C1(n11539), .C2(n12053), .A(n11525), .B(n11524), .ZN(
        P2_U3194) );
  AOI22_X1 U13515 ( .A1(n14578), .A2(n7435), .B1(n14384), .B2(n14575), .ZN(
        n11677) );
  INV_X1 U13516 ( .A(n11677), .ZN(n11526) );
  AOI22_X1 U13517 ( .A1(n14358), .A2(n11526), .B1(n14324), .B2(n11679), .ZN(
        n11532) );
  OAI21_X1 U13518 ( .B1(n11529), .B2(n11528), .A(n11527), .ZN(n11530) );
  NAND2_X1 U13519 ( .A1(n11530), .A2(n14352), .ZN(n11531) );
  OAI211_X1 U13520 ( .C1(n11539), .C2(n9985), .A(n11532), .B(n11531), .ZN(
        P2_U3209) );
  INV_X1 U13521 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11855) );
  OAI21_X1 U13522 ( .B1(n12771), .B2(n11535), .A(n11534), .ZN(n11536) );
  AOI22_X1 U13523 ( .A1(n14352), .A2(n11536), .B1(n14324), .B2(n10697), .ZN(
        n11538) );
  NAND2_X1 U13524 ( .A1(n14331), .A2(n7435), .ZN(n11537) );
  OAI211_X1 U13525 ( .C1(n11539), .C2(n11855), .A(n11538), .B(n11537), .ZN(
        P2_U3204) );
  INV_X1 U13526 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U13527 ( .A1(n11540), .A2(P3_U3897), .ZN(n11541) );
  OAI21_X1 U13528 ( .B1(P3_U3897), .B2(n11542), .A(n11541), .ZN(P3_U3500) );
  INV_X1 U13529 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15594) );
  NAND2_X1 U13530 ( .A1(n13655), .A2(P3_U3897), .ZN(n11543) );
  OAI21_X1 U13531 ( .B1(P3_U3897), .B2(n15594), .A(n11543), .ZN(P3_U3505) );
  INV_X1 U13532 ( .A(n11544), .ZN(n11546) );
  INV_X1 U13533 ( .A(n11904), .ZN(n11908) );
  OAI222_X1 U13534 ( .A1(n15810), .A2(n11545), .B1(n15805), .B2(n11546), .C1(
        P1_U3086), .C2(n11908), .ZN(P1_U3341) );
  INV_X1 U13535 ( .A(n15859), .ZN(n12579) );
  OAI222_X1 U13536 ( .A1(n14792), .A2(n11547), .B1(n14775), .B2(n11546), .C1(
        P2_U3088), .C2(n12579), .ZN(P2_U3313) );
  INV_X1 U13537 ( .A(n11548), .ZN(n11549) );
  INV_X1 U13538 ( .A(n16213), .ZN(n13758) );
  OAI222_X1 U13539 ( .A1(n14223), .A2(n15479), .B1(n14221), .B2(n11549), .C1(
        n13758), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U13540 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U13541 ( .A1(n13625), .A2(P3_U3897), .ZN(n11550) );
  OAI21_X1 U13542 ( .B1(P3_U3897), .B2(n15596), .A(n11550), .ZN(P3_U3506) );
  INV_X1 U13543 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U13544 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13170)
         );
  OAI21_X1 U13545 ( .B1(n15046), .B2(n11551), .A(n13170), .ZN(n11557) );
  OAI21_X1 U13546 ( .B1(n11558), .B2(P1_REG2_REG_12__SCAN_IN), .A(n11552), 
        .ZN(n11555) );
  INV_X1 U13547 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11553) );
  MUX2_X1 U13548 ( .A(n11553), .B(P1_REG2_REG_13__SCAN_IN), .S(n11627), .Z(
        n11554) );
  NOR2_X1 U13549 ( .A1(n11555), .A2(n11554), .ZN(n11626) );
  AOI211_X1 U13550 ( .C1(n11555), .C2(n11554), .A(n13028), .B(n11626), .ZN(
        n11556) );
  AOI211_X1 U13551 ( .C1(n16285), .C2(n11627), .A(n11557), .B(n11556), .ZN(
        n11567) );
  OR2_X1 U13552 ( .A1(n11558), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U13553 ( .A1(n11560), .A2(n11559), .ZN(n11563) );
  INV_X1 U13554 ( .A(n11563), .ZN(n11565) );
  MUX2_X1 U13555 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11561), .S(n11627), .Z(
        n11564) );
  MUX2_X1 U13556 ( .A(n11561), .B(P1_REG1_REG_13__SCAN_IN), .S(n11627), .Z(
        n11562) );
  OR2_X1 U13557 ( .A1(n11563), .A2(n11562), .ZN(n11629) );
  OAI211_X1 U13558 ( .C1(n11565), .C2(n11564), .A(n16283), .B(n11629), .ZN(
        n11566) );
  NAND2_X1 U13559 ( .A1(n11567), .A2(n11566), .ZN(P1_U3256) );
  INV_X1 U13560 ( .A(n11568), .ZN(n12300) );
  NAND2_X1 U13561 ( .A1(n14382), .A2(n14575), .ZN(n11570) );
  NAND2_X1 U13562 ( .A1(n14384), .A2(n14578), .ZN(n11569) );
  AND2_X1 U13563 ( .A1(n11570), .A2(n11569), .ZN(n11615) );
  NAND2_X1 U13564 ( .A1(n14324), .A2(n11612), .ZN(n11571) );
  NAND2_X1 U13565 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14401) );
  OAI211_X1 U13566 ( .C1(n11615), .C2(n14297), .A(n11571), .B(n14401), .ZN(
        n11588) );
  INV_X1 U13567 ( .A(n11572), .ZN(n11575) );
  INV_X1 U13568 ( .A(n11573), .ZN(n11574) );
  NAND2_X1 U13569 ( .A1(n11575), .A2(n11574), .ZN(n11576) );
  XNOR2_X1 U13570 ( .A(n11612), .B(n14244), .ZN(n11579) );
  OR2_X1 U13571 ( .A1(n11647), .A2(n12771), .ZN(n11580) );
  NAND2_X1 U13572 ( .A1(n11579), .A2(n11580), .ZN(n11643) );
  INV_X1 U13573 ( .A(n11579), .ZN(n11582) );
  INV_X1 U13574 ( .A(n11580), .ZN(n11581) );
  NAND2_X1 U13575 ( .A1(n11582), .A2(n11581), .ZN(n11583) );
  NAND2_X1 U13576 ( .A1(n11643), .A2(n11583), .ZN(n11584) );
  NAND2_X1 U13577 ( .A1(n11585), .A2(n11584), .ZN(n11586) );
  AOI21_X1 U13578 ( .B1(n11644), .B2(n11586), .A(n14326), .ZN(n11587) );
  AOI211_X1 U13579 ( .C1(n14332), .C2(n12300), .A(n11588), .B(n11587), .ZN(
        n11589) );
  INV_X1 U13580 ( .A(n11589), .ZN(P2_U3202) );
  INV_X1 U13581 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15593) );
  NAND2_X1 U13582 ( .A1(n13656), .A2(P3_U3897), .ZN(n11590) );
  OAI21_X1 U13583 ( .B1(P3_U3897), .B2(n15593), .A(n11590), .ZN(P3_U3503) );
  OAI21_X1 U13584 ( .B1(n11591), .B2(n11593), .A(n11592), .ZN(n11594) );
  NAND2_X1 U13585 ( .A1(n11594), .A2(n14905), .ZN(n11597) );
  OAI22_X1 U13586 ( .A1(n11595), .A2(n15216), .B1(n15218), .B2(n9196), .ZN(
        n16316) );
  AOI22_X1 U13587 ( .A1(n14899), .A2(n16316), .B1(n11603), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n11596) );
  OAI211_X1 U13588 ( .C1(n16314), .C2(n14918), .A(n11597), .B(n11596), .ZN(
        P1_U3222) );
  OAI21_X1 U13589 ( .B1(n11600), .B2(n11599), .A(n11598), .ZN(n11601) );
  NAND2_X1 U13590 ( .A1(n11601), .A2(n14905), .ZN(n11605) );
  OAI22_X1 U13591 ( .A1(n11602), .A2(n15216), .B1(n15218), .B2(n11846), .ZN(
        n16354) );
  AOI22_X1 U13592 ( .A1(n14899), .A2(n16354), .B1(n11603), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n11604) );
  OAI211_X1 U13593 ( .C1(n16348), .C2(n14918), .A(n11605), .B(n11604), .ZN(
        P1_U3237) );
  NAND2_X1 U13594 ( .A1(n13694), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13584) );
  INV_X1 U13595 ( .A(n13584), .ZN(n11609) );
  INV_X1 U13596 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11608) );
  INV_X1 U13597 ( .A(n12443), .ZN(n11988) );
  AND2_X1 U13598 ( .A1(n13585), .A2(n11988), .ZN(n13365) );
  INV_X1 U13599 ( .A(n13365), .ZN(n13520) );
  NAND2_X1 U13600 ( .A1(n13520), .A2(n12404), .ZN(n11894) );
  OAI22_X1 U13601 ( .A1(n12330), .A2(n13671), .B1(n11988), .B2(n13700), .ZN(
        n11606) );
  AOI21_X1 U13602 ( .B1(n11894), .B2(n13690), .A(n11606), .ZN(n11607) );
  OAI21_X1 U13603 ( .B1(n11609), .B2(n11608), .A(n11607), .ZN(P3_U3172) );
  OAI21_X1 U13604 ( .B1(n11611), .B2(n11614), .A(n11610), .ZN(n12305) );
  AOI211_X1 U13605 ( .C1(n11612), .C2(n11684), .A(n11533), .B(n11698), .ZN(
        n12299) );
  XNOR2_X1 U13606 ( .A(n11613), .B(n11614), .ZN(n11616) );
  OAI21_X1 U13607 ( .B1(n11616), .B2(n14510), .A(n11615), .ZN(n12298) );
  AOI211_X1 U13608 ( .C1(n16588), .C2(n12305), .A(n12299), .B(n12298), .ZN(
        n12026) );
  OAI22_X1 U13609 ( .A1(n14708), .A2(n12303), .B1(n16591), .B2(n11294), .ZN(
        n11617) );
  INV_X1 U13610 ( .A(n11617), .ZN(n11618) );
  OAI21_X1 U13611 ( .B1(n12026), .B2(n16589), .A(n11618), .ZN(P2_U3503) );
  INV_X1 U13612 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U13613 ( .A1(n11619), .A2(P3_U3897), .ZN(n11620) );
  OAI21_X1 U13614 ( .B1(P3_U3897), .B2(n15389), .A(n11620), .ZN(P3_U3501) );
  INV_X1 U13615 ( .A(n11626), .ZN(n11622) );
  NAND2_X1 U13616 ( .A1(n11627), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11623) );
  INV_X1 U13617 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11621) );
  MUX2_X1 U13618 ( .A(n11621), .B(P1_REG2_REG_14__SCAN_IN), .S(n11904), .Z(
        n11624) );
  AOI21_X1 U13619 ( .B1(n11622), .B2(n11623), .A(n11624), .ZN(n11906) );
  NAND2_X1 U13620 ( .A1(n11624), .A2(n11623), .ZN(n11625) );
  OAI21_X1 U13621 ( .B1(n11626), .B2(n11625), .A(n16277), .ZN(n11636) );
  INV_X1 U13622 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n16570) );
  MUX2_X1 U13623 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n16570), .S(n11904), .Z(
        n11631) );
  NAND2_X1 U13624 ( .A1(n11627), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11628) );
  AND2_X1 U13625 ( .A1(n11629), .A2(n11628), .ZN(n11630) );
  NAND2_X1 U13626 ( .A1(n11630), .A2(n11631), .ZN(n11903) );
  OAI21_X1 U13627 ( .B1(n11631), .B2(n11630), .A(n11903), .ZN(n11632) );
  NAND2_X1 U13628 ( .A1(n11632), .A2(n16283), .ZN(n11635) );
  INV_X1 U13629 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n16047) );
  NAND2_X1 U13630 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n16555)
         );
  OAI21_X1 U13631 ( .B1(n15046), .B2(n16047), .A(n16555), .ZN(n11633) );
  AOI21_X1 U13632 ( .B1(n16285), .B2(n11904), .A(n11633), .ZN(n11634) );
  OAI211_X1 U13633 ( .C1(n11906), .C2(n11636), .A(n11635), .B(n11634), .ZN(
        P1_U3257) );
  INV_X1 U13634 ( .A(n13756), .ZN(n16243) );
  OAI222_X1 U13635 ( .A1(n14223), .A2(n15480), .B1(n14221), .B2(n11637), .C1(
        n16243), .C2(P3_U3151), .ZN(P3_U3278) );
  XNOR2_X1 U13636 ( .A(n11701), .B(n14244), .ZN(n11638) );
  NAND2_X1 U13637 ( .A1(n14382), .A2(n11533), .ZN(n11639) );
  NAND2_X1 U13638 ( .A1(n11638), .A2(n11639), .ZN(n11653) );
  INV_X1 U13639 ( .A(n11638), .ZN(n11641) );
  INV_X1 U13640 ( .A(n11639), .ZN(n11640) );
  NAND2_X1 U13641 ( .A1(n11641), .A2(n11640), .ZN(n11642) );
  AND2_X1 U13642 ( .A1(n11653), .A2(n11642), .ZN(n11646) );
  OAI21_X1 U13643 ( .B1(n11646), .B2(n11645), .A(n11654), .ZN(n11651) );
  NOR2_X1 U13644 ( .A1(n14297), .A2(n14602), .ZN(n14333) );
  OAI22_X1 U13645 ( .A1(n14281), .A2(n11647), .B1(n12070), .B2(n14355), .ZN(
        n11650) );
  NAND2_X1 U13646 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14416) );
  NAND2_X1 U13647 ( .A1(n14324), .A2(n11701), .ZN(n11648) );
  OAI211_X1 U13648 ( .C1(n14320), .C2(n12079), .A(n14416), .B(n11648), .ZN(
        n11649) );
  AOI211_X1 U13649 ( .C1(n11651), .C2(n14352), .A(n11650), .B(n11649), .ZN(
        n11652) );
  INV_X1 U13650 ( .A(n11652), .ZN(P2_U3199) );
  XNOR2_X1 U13651 ( .A(n16419), .B(n14244), .ZN(n11961) );
  NAND2_X1 U13652 ( .A1(n14381), .A2(n11533), .ZN(n11960) );
  XNOR2_X1 U13653 ( .A(n11961), .B(n11960), .ZN(n11962) );
  XNOR2_X1 U13654 ( .A(n11963), .B(n11962), .ZN(n11660) );
  OAI21_X1 U13655 ( .B1(n14320), .B2(n12247), .A(n11655), .ZN(n11658) );
  OAI22_X1 U13656 ( .A1(n14281), .A2(n11656), .B1(n12259), .B2(n14355), .ZN(
        n11657) );
  AOI211_X1 U13657 ( .C1(n16419), .C2(n14324), .A(n11658), .B(n11657), .ZN(
        n11659) );
  OAI21_X1 U13658 ( .B1(n11660), .B2(n14326), .A(n11659), .ZN(P2_U3211) );
  OAI21_X1 U13659 ( .B1(n11662), .B2(n7506), .A(n11661), .ZN(n12052) );
  NAND2_X1 U13660 ( .A1(n10697), .A2(n11668), .ZN(n11663) );
  NAND2_X1 U13661 ( .A1(n11663), .A2(n12771), .ZN(n11664) );
  NOR2_X1 U13662 ( .A1(n11672), .A2(n11664), .ZN(n12056) );
  XNOR2_X1 U13663 ( .A(n10333), .B(n11665), .ZN(n11667) );
  OAI21_X1 U13664 ( .B1(n11667), .B2(n14510), .A(n11666), .ZN(n12057) );
  AOI211_X1 U13665 ( .C1(n16588), .C2(n12052), .A(n12056), .B(n12057), .ZN(
        n12018) );
  INV_X1 U13666 ( .A(n14708), .ZN(n12643) );
  AOI22_X1 U13667 ( .A1(n12643), .A2(n11668), .B1(n16589), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n11669) );
  OAI21_X1 U13668 ( .B1(n12018), .B2(n16589), .A(n11669), .ZN(P2_U3500) );
  OAI21_X1 U13669 ( .B1(n11671), .B2(n11675), .A(n11670), .ZN(n12273) );
  INV_X1 U13670 ( .A(n11672), .ZN(n11673) );
  AOI21_X1 U13671 ( .B1(n11673), .B2(n11679), .A(n11533), .ZN(n11674) );
  AND2_X1 U13672 ( .A1(n11674), .A2(n11683), .ZN(n12267) );
  XNOR2_X1 U13673 ( .A(n11676), .B(n11675), .ZN(n11678) );
  OAI21_X1 U13674 ( .B1(n11678), .B2(n14510), .A(n11677), .ZN(n12266) );
  AOI211_X1 U13675 ( .C1(n16588), .C2(n12273), .A(n12267), .B(n12266), .ZN(
        n12022) );
  AOI22_X1 U13676 ( .A1(n12643), .A2(n11679), .B1(n16589), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n11680) );
  OAI21_X1 U13677 ( .B1(n12022), .B2(n16589), .A(n11680), .ZN(P2_U3501) );
  OAI21_X1 U13678 ( .B1(n11682), .B2(n11686), .A(n11681), .ZN(n12041) );
  AOI21_X1 U13679 ( .B1(n12045), .B2(n11683), .A(n11533), .ZN(n11685) );
  AND2_X1 U13680 ( .A1(n11685), .A2(n11684), .ZN(n12048) );
  OAI21_X1 U13681 ( .B1(n11688), .B2(n14510), .A(n11687), .ZN(n12042) );
  AOI211_X1 U13682 ( .C1(n16588), .C2(n12041), .A(n12048), .B(n12042), .ZN(
        n11959) );
  AOI22_X1 U13683 ( .A1(n12643), .A2(n12045), .B1(n16589), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n11689) );
  OAI21_X1 U13684 ( .B1(n11959), .B2(n16589), .A(n11689), .ZN(P2_U3502) );
  AOI21_X1 U13685 ( .B1(n14510), .B2(n14609), .A(n11860), .ZN(n11691) );
  AOI21_X1 U13686 ( .B1(n14575), .B2(n7435), .A(n11691), .ZN(n11851) );
  OAI211_X1 U13687 ( .C1(n11860), .C2(n12148), .A(n11851), .B(n11853), .ZN(
        n14725) );
  NAND2_X1 U13688 ( .A1(n16595), .A2(n14725), .ZN(n11692) );
  OAI21_X1 U13689 ( .B1(n16595), .B2(n9953), .A(n11692), .ZN(P2_U3430) );
  INV_X1 U13690 ( .A(n16253), .ZN(n13793) );
  OAI222_X1 U13691 ( .A1(P3_U3151), .A2(n13793), .B1(n14223), .B2(n11694), 
        .C1(n14221), .C2(n11693), .ZN(P3_U3277) );
  OR2_X1 U13692 ( .A1(n11695), .A2(n11703), .ZN(n11696) );
  NAND2_X1 U13693 ( .A1(n11697), .A2(n11696), .ZN(n12067) );
  INV_X1 U13694 ( .A(n11698), .ZN(n11700) );
  INV_X1 U13695 ( .A(n12257), .ZN(n11699) );
  AOI211_X1 U13696 ( .C1(n11701), .C2(n11700), .A(n11533), .B(n11699), .ZN(
        n12073) );
  XNOR2_X1 U13697 ( .A(n11702), .B(n11703), .ZN(n11706) );
  INV_X1 U13698 ( .A(n14609), .ZN(n12254) );
  NAND2_X1 U13699 ( .A1(n12067), .A2(n12254), .ZN(n11705) );
  AOI22_X1 U13700 ( .A1(n14383), .A2(n14578), .B1(n14575), .B2(n14381), .ZN(
        n11704) );
  OAI211_X1 U13701 ( .C1(n14510), .C2(n11706), .A(n11705), .B(n11704), .ZN(
        n12068) );
  AOI211_X1 U13702 ( .C1(n16514), .C2(n12067), .A(n12073), .B(n12068), .ZN(
        n12014) );
  OAI22_X1 U13703 ( .A1(n14708), .A2(n12071), .B1(n16591), .B2(n11295), .ZN(
        n11707) );
  INV_X1 U13704 ( .A(n11707), .ZN(n11708) );
  OAI21_X1 U13705 ( .B1(n12014), .B2(n16589), .A(n11708), .ZN(P2_U3504) );
  INV_X1 U13706 ( .A(n16558), .ZN(n14914) );
  INV_X1 U13707 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14973) );
  INV_X1 U13708 ( .A(n16365), .ZN(n12034) );
  OAI22_X1 U13709 ( .A1(n9196), .A2(n15216), .B1(n15218), .B2(n11996), .ZN(
        n12028) );
  AOI22_X1 U13710 ( .A1(n14899), .A2(n12028), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11709) );
  OAI21_X1 U13711 ( .B1(n14918), .B2(n12034), .A(n11709), .ZN(n11714) );
  AOI211_X1 U13712 ( .C1(n11712), .C2(n11711), .A(n16549), .B(n11710), .ZN(
        n11713) );
  AOI211_X1 U13713 ( .C1(n14914), .C2(n14973), .A(n11714), .B(n11713), .ZN(
        n11715) );
  INV_X1 U13714 ( .A(n11715), .ZN(P1_U3218) );
  INV_X1 U13715 ( .A(n11716), .ZN(n11718) );
  INV_X1 U13716 ( .A(n12758), .ZN(n12750) );
  OAI222_X1 U13717 ( .A1(n15810), .A2(n11717), .B1(n15805), .B2(n11718), .C1(
        n12750), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13718 ( .A(n12718), .ZN(n12725) );
  OAI222_X1 U13719 ( .A1(n14792), .A2(n11719), .B1(n14775), .B2(n11718), .C1(
        n12725), .C2(P2_U3088), .ZN(P2_U3312) );
  MUX2_X1 U13720 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n7414), .Z(n11750) );
  INV_X1 U13721 ( .A(n11738), .ZN(n11751) );
  XNOR2_X1 U13722 ( .A(n11750), .B(n11751), .ZN(n11749) );
  INV_X1 U13723 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11720) );
  INV_X1 U13724 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11987) );
  MUX2_X1 U13725 ( .A(n11720), .B(n11987), .S(n7414), .Z(n16100) );
  NAND2_X1 U13726 ( .A1(n16100), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n16099) );
  XNOR2_X1 U13727 ( .A(n11749), .B(n16099), .ZN(n11747) );
  NAND2_X1 U13728 ( .A1(n13466), .A2(n11723), .ZN(n11725) );
  AND2_X1 U13729 ( .A1(n11725), .A2(n11724), .ZN(n11730) );
  INV_X1 U13730 ( .A(n11742), .ZN(n11726) );
  MUX2_X1 U13731 ( .A(n13711), .B(n11726), .S(n8956), .Z(n16244) );
  INV_X1 U13732 ( .A(n16262), .ZN(n16116) );
  NAND2_X1 U13733 ( .A1(n11736), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U13734 ( .A1(n11738), .A2(n11764), .ZN(n11729) );
  NAND2_X1 U13735 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n11735), .ZN(n11727) );
  OR2_X1 U13736 ( .A1(n11727), .A2(n11736), .ZN(n11728) );
  NAND2_X1 U13737 ( .A1(n11729), .A2(n11728), .ZN(n11763) );
  XOR2_X1 U13738 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n11763), .Z(n11734) );
  INV_X1 U13739 ( .A(n11730), .ZN(n11731) );
  AOI22_X1 U13740 ( .A1(n16252), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11733) );
  OAI21_X1 U13741 ( .B1(n16116), .B2(n11734), .A(n11733), .ZN(n11745) );
  AND2_X1 U13742 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n11735), .ZN(n11737) );
  NAND2_X1 U13743 ( .A1(n11736), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11773) );
  OAI21_X1 U13744 ( .B1(n11738), .B2(n11737), .A(n11773), .ZN(n11739) );
  INV_X1 U13745 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U13746 ( .A1(n11739), .A2(n12409), .ZN(n11743) );
  INV_X1 U13747 ( .A(n11740), .ZN(n11741) );
  AOI21_X1 U13748 ( .B1(n11774), .B2(n11743), .A(n16250), .ZN(n11744) );
  AOI211_X1 U13749 ( .C1(n16254), .C2(n11751), .A(n11745), .B(n11744), .ZN(
        n11746) );
  OAI21_X1 U13750 ( .B1(n16190), .B2(n11747), .A(n11746), .ZN(P3_U3183) );
  MUX2_X1 U13751 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13791), .Z(n11791) );
  XNOR2_X1 U13752 ( .A(n11791), .B(n11792), .ZN(n11789) );
  INV_X1 U13753 ( .A(n16099), .ZN(n11748) );
  NAND2_X1 U13754 ( .A1(n11749), .A2(n11748), .ZN(n11754) );
  INV_X1 U13755 ( .A(n11750), .ZN(n11752) );
  NAND2_X1 U13756 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U13757 ( .A1(n11754), .A2(n11753), .ZN(n11811) );
  MUX2_X1 U13758 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n7414), .Z(n11755) );
  XNOR2_X1 U13759 ( .A(n11755), .B(n11772), .ZN(n11812) );
  NAND2_X1 U13760 ( .A1(n11811), .A2(n11812), .ZN(n11758) );
  INV_X1 U13761 ( .A(n11755), .ZN(n11756) );
  NAND2_X1 U13762 ( .A1(n11758), .A2(n11757), .ZN(n11827) );
  MUX2_X1 U13763 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13791), .Z(n11759) );
  XNOR2_X1 U13764 ( .A(n11759), .B(n11838), .ZN(n11828) );
  NAND2_X1 U13765 ( .A1(n11827), .A2(n11828), .ZN(n11762) );
  INV_X1 U13766 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U13767 ( .A1(n11760), .A2(n11838), .ZN(n11761) );
  NAND2_X1 U13768 ( .A1(n11762), .A2(n11761), .ZN(n11790) );
  XOR2_X1 U13769 ( .A(n11789), .B(n11790), .Z(n11788) );
  INV_X1 U13770 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n12487) );
  MUX2_X1 U13771 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n12487), .S(n11792), .Z(
        n11770) );
  INV_X1 U13772 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U13773 ( .A1(n11763), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11765) );
  NAND2_X1 U13774 ( .A1(n11765), .A2(n11764), .ZN(n11818) );
  NAND2_X1 U13775 ( .A1(n11819), .A2(n11818), .ZN(n11817) );
  OR2_X1 U13776 ( .A1(n11772), .A2(n11766), .ZN(n11767) );
  NAND2_X1 U13777 ( .A1(n11817), .A2(n11767), .ZN(n11768) );
  XNOR2_X1 U13778 ( .A(n11768), .B(n11838), .ZN(n11832) );
  AOI22_X1 U13779 ( .A1(n11832), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n11777), 
        .B2(n11768), .ZN(n11769) );
  AOI21_X1 U13780 ( .B1(n11770), .B2(n11769), .A(n11800), .ZN(n11785) );
  NOR2_X1 U13781 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15542), .ZN(n12389) );
  AOI21_X1 U13782 ( .B1(n16252), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n12389), .ZN(
        n11784) );
  XNOR2_X1 U13783 ( .A(n11792), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11781) );
  XNOR2_X1 U13784 ( .A(n11772), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n11815) );
  INV_X1 U13785 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11775) );
  OR2_X1 U13786 ( .A1(n11772), .A2(n11775), .ZN(n11776) );
  XNOR2_X1 U13787 ( .A(n11778), .B(n11777), .ZN(n11830) );
  INV_X1 U13788 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11829) );
  INV_X1 U13789 ( .A(n11778), .ZN(n11779) );
  OAI22_X1 U13790 ( .A1(n11830), .A2(n11829), .B1(n11838), .B2(n11779), .ZN(
        n11780) );
  OAI21_X1 U13791 ( .B1(n11781), .B2(n11780), .A(n11797), .ZN(n11782) );
  NAND2_X1 U13792 ( .A1(n16265), .A2(n11782), .ZN(n11783) );
  OAI211_X1 U13793 ( .C1(n16116), .C2(n11785), .A(n11784), .B(n11783), .ZN(
        n11786) );
  AOI21_X1 U13794 ( .B1(n11792), .B2(n16254), .A(n11786), .ZN(n11787) );
  OAI21_X1 U13795 ( .B1(n11788), .B2(n16190), .A(n11787), .ZN(P3_U3186) );
  MUX2_X1 U13796 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13791), .Z(n11926) );
  XNOR2_X1 U13797 ( .A(n11926), .B(n11927), .ZN(n11924) );
  NAND2_X1 U13798 ( .A1(n11790), .A2(n11789), .ZN(n11795) );
  INV_X1 U13799 ( .A(n11791), .ZN(n11793) );
  NAND2_X1 U13800 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  NAND2_X1 U13801 ( .A1(n11795), .A2(n11794), .ZN(n11925) );
  XOR2_X1 U13802 ( .A(n11924), .B(n11925), .Z(n11810) );
  INV_X1 U13803 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11798) );
  AOI21_X1 U13804 ( .B1(n11799), .B2(n11798), .A(n11936), .ZN(n11807) );
  NAND2_X1 U13805 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n11802), .ZN(n11943) );
  OAI21_X1 U13806 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11802), .A(n11943), .ZN(
        n11805) );
  NOR2_X1 U13807 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11803), .ZN(n12533) );
  INV_X1 U13808 ( .A(n16252), .ZN(n16241) );
  NOR2_X1 U13809 ( .A1(n16241), .A2(n15971), .ZN(n11804) );
  AOI211_X1 U13810 ( .C1(n16262), .C2(n11805), .A(n12533), .B(n11804), .ZN(
        n11806) );
  OAI21_X1 U13811 ( .B1(n11807), .B2(n16250), .A(n11806), .ZN(n11808) );
  AOI21_X1 U13812 ( .B1(n11927), .B2(n16254), .A(n11808), .ZN(n11809) );
  OAI21_X1 U13813 ( .B1(n11810), .B2(n16190), .A(n11809), .ZN(P3_U3187) );
  XOR2_X1 U13814 ( .A(n11812), .B(n11811), .Z(n11826) );
  OAI21_X1 U13815 ( .B1(n11815), .B2(n11814), .A(n11813), .ZN(n11816) );
  NAND2_X1 U13816 ( .A1(n16265), .A2(n11816), .ZN(n11823) );
  OAI21_X1 U13817 ( .B1(n11819), .B2(n11818), .A(n11817), .ZN(n11820) );
  NAND2_X1 U13818 ( .A1(n16262), .A2(n11820), .ZN(n11822) );
  AOI22_X1 U13819 ( .A1(n16252), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11821) );
  NAND3_X1 U13820 ( .A1(n11823), .A2(n11822), .A3(n11821), .ZN(n11824) );
  AOI21_X1 U13821 ( .B1(n16254), .B2(n11772), .A(n11824), .ZN(n11825) );
  OAI21_X1 U13822 ( .B1(n11826), .B2(n16190), .A(n11825), .ZN(P3_U3184) );
  XOR2_X1 U13823 ( .A(n11828), .B(n11827), .Z(n11840) );
  XNOR2_X1 U13824 ( .A(n11830), .B(n11829), .ZN(n11831) );
  NAND2_X1 U13825 ( .A1(n16265), .A2(n11831), .ZN(n11836) );
  XNOR2_X1 U13826 ( .A(n11832), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n11833) );
  NAND2_X1 U13827 ( .A1(n16262), .A2(n11833), .ZN(n11835) );
  AOI22_X1 U13828 ( .A1(n16252), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11834) );
  NAND3_X1 U13829 ( .A1(n11836), .A2(n11835), .A3(n11834), .ZN(n11837) );
  AOI21_X1 U13830 ( .B1(n16254), .B2(n11838), .A(n11837), .ZN(n11839) );
  OAI21_X1 U13831 ( .B1(n11840), .B2(n16190), .A(n11839), .ZN(P3_U3185) );
  NAND2_X1 U13832 ( .A1(n7573), .A2(n11841), .ZN(n11843) );
  XNOR2_X1 U13833 ( .A(n11843), .B(n11842), .ZN(n11850) );
  INV_X1 U13834 ( .A(n11844), .ZN(n16388) );
  OAI22_X1 U13835 ( .A1(n11846), .A2(n15216), .B1(n15218), .B2(n11845), .ZN(
        n16382) );
  AOI22_X1 U13836 ( .A1(n14899), .A2(n16382), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11847) );
  OAI21_X1 U13837 ( .B1(n14918), .B2(n9860), .A(n11847), .ZN(n11848) );
  AOI21_X1 U13838 ( .B1(n16388), .B2(n14914), .A(n11848), .ZN(n11849) );
  OAI21_X1 U13839 ( .B1(n11850), .B2(n16549), .A(n11849), .ZN(P1_U3230) );
  INV_X1 U13840 ( .A(n11851), .ZN(n11857) );
  INV_X1 U13841 ( .A(n11852), .ZN(n11854) );
  OAI22_X1 U13842 ( .A1(n14640), .A2(n11855), .B1(n11854), .B2(n11853), .ZN(
        n11856) );
  OAI21_X1 U13843 ( .B1(n11857), .B2(n11856), .A(n14610), .ZN(n11859) );
  NAND2_X1 U13844 ( .A1(n16598), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n11858) );
  OAI211_X1 U13845 ( .C1(n14613), .C2(n11860), .A(n11859), .B(n11858), .ZN(
        P2_U3265) );
  INV_X1 U13846 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n16515) );
  NOR2_X1 U13847 ( .A1(n15896), .A2(n16515), .ZN(n11864) );
  OAI21_X1 U13848 ( .B1(n11863), .B2(n11862), .A(n11861), .ZN(n15902) );
  AOI211_X1 U13849 ( .C1(n16515), .C2(n15896), .A(n11864), .B(n15902), .ZN(
        n15900) );
  AOI21_X1 U13850 ( .B1(n16515), .B2(n15896), .A(n15900), .ZN(n11868) );
  INV_X1 U13851 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12805) );
  OR2_X1 U13852 ( .A1(n12583), .A2(n12805), .ZN(n11865) );
  OAI21_X1 U13853 ( .B1(n12577), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11865), 
        .ZN(n11867) );
  NAND2_X1 U13854 ( .A1(n12583), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11866) );
  OAI211_X1 U13855 ( .C1(n12583), .C2(P2_REG1_REG_13__SCAN_IN), .A(n11868), 
        .B(n11866), .ZN(n12576) );
  OAI211_X1 U13856 ( .C1(n11868), .C2(n11867), .A(n12576), .B(n15920), .ZN(
        n11871) );
  NOR2_X1 U13857 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12876), .ZN(n11869) );
  AOI21_X1 U13858 ( .B1(n15880), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11869), 
        .ZN(n11870) );
  OAI211_X1 U13859 ( .C1(n14418), .C2(n12577), .A(n11871), .B(n11870), .ZN(
        n11880) );
  NOR2_X1 U13860 ( .A1(n12583), .A2(n11872), .ZN(n11873) );
  AOI21_X1 U13861 ( .B1(n12583), .B2(n11872), .A(n11873), .ZN(n11878) );
  INV_X1 U13862 ( .A(n15896), .ZN(n15908) );
  NOR2_X1 U13863 ( .A1(n11874), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15893) );
  NAND2_X1 U13864 ( .A1(n15908), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U13865 ( .A1(n15896), .A2(n12599), .ZN(n11875) );
  OAI211_X1 U13866 ( .C1(n15892), .C2(n15893), .A(n11876), .B(n11875), .ZN(
        n15899) );
  OAI21_X1 U13867 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n15908), .A(n15899), 
        .ZN(n11877) );
  NOR2_X1 U13868 ( .A1(n11877), .A2(n11878), .ZN(n12582) );
  AOI211_X1 U13869 ( .C1(n11878), .C2(n11877), .A(n15897), .B(n12582), .ZN(
        n11879) );
  OR2_X1 U13870 ( .A1(n11880), .A2(n11879), .ZN(P2_U3227) );
  OAI222_X1 U13871 ( .A1(n14223), .A2(n15474), .B1(P3_U3151), .B2(n13799), 
        .C1(n14221), .C2(n11881), .ZN(P3_U3276) );
  INV_X1 U13872 ( .A(n11883), .ZN(n11885) );
  NOR2_X1 U13873 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  XNOR2_X1 U13874 ( .A(n11887), .B(n11886), .ZN(n11892) );
  INV_X1 U13875 ( .A(n16543), .ZN(n11890) );
  OAI22_X1 U13876 ( .A1(n16542), .A2(n12166), .B1(n16558), .B2(n12007), .ZN(
        n11889) );
  NAND2_X1 U13877 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14987) );
  OAI21_X1 U13878 ( .B1(n14918), .B2(n16401), .A(n14987), .ZN(n11888) );
  AOI211_X1 U13879 ( .C1(n11890), .C2(n14940), .A(n11889), .B(n11888), .ZN(
        n11891) );
  OAI21_X1 U13880 ( .B1(n11892), .B2(n16549), .A(n11891), .ZN(P1_U3227) );
  NAND3_X1 U13881 ( .A1(n11894), .A2(n16609), .A3(n11893), .ZN(n11895) );
  OAI21_X1 U13882 ( .B1(n12330), .B2(n14089), .A(n11895), .ZN(n12439) );
  INV_X1 U13883 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11896) );
  OAI22_X1 U13884 ( .A1(n14207), .A2(n11988), .B1(n16618), .B2(n11896), .ZN(
        n11897) );
  AOI21_X1 U13885 ( .B1(n12439), .B2(n16618), .A(n11897), .ZN(n11898) );
  INV_X1 U13886 ( .A(n11898), .ZN(P3_U3390) );
  INV_X1 U13887 ( .A(n11899), .ZN(n11901) );
  INV_X1 U13888 ( .A(n15037), .ZN(n12762) );
  OAI222_X1 U13889 ( .A1(n15810), .A2(n11900), .B1(n15805), .B2(n11901), .C1(
        n12762), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13890 ( .A(n15874), .ZN(n12730) );
  OAI222_X1 U13891 ( .A1(n14792), .A2(n11902), .B1(n14775), .B2(n11901), .C1(
        n12730), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI21_X1 U13892 ( .B1(n11904), .B2(P1_REG1_REG_14__SCAN_IN), .A(n11903), 
        .ZN(n12751) );
  XNOR2_X1 U13893 ( .A(n12751), .B(n12750), .ZN(n11905) );
  NOR2_X1 U13894 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11905), .ZN(n12749) );
  AOI21_X1 U13895 ( .B1(n11905), .B2(P1_REG1_REG_15__SCAN_IN), .A(n12749), 
        .ZN(n11916) );
  INV_X1 U13896 ( .A(n11906), .ZN(n11907) );
  OAI21_X1 U13897 ( .B1(n11621), .B2(n11908), .A(n11907), .ZN(n12757) );
  XNOR2_X1 U13898 ( .A(n12757), .B(n12758), .ZN(n11909) );
  NOR2_X1 U13899 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11909), .ZN(n12759) );
  AOI21_X1 U13900 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11909), .A(n12759), 
        .ZN(n11910) );
  NOR2_X1 U13901 ( .A1(n11910), .A2(n13028), .ZN(n11914) );
  NOR2_X1 U13902 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14911), .ZN(n11911) );
  AOI21_X1 U13903 ( .B1(n16287), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n11911), 
        .ZN(n11912) );
  OAI21_X1 U13904 ( .B1(n13026), .B2(n12750), .A(n11912), .ZN(n11913) );
  NOR2_X1 U13905 ( .A1(n11914), .A2(n11913), .ZN(n11915) );
  OAI21_X1 U13906 ( .B1(n11916), .B2(n13030), .A(n11915), .ZN(P1_U3258) );
  XOR2_X1 U13907 ( .A(n11917), .B(n11918), .Z(n11923) );
  AOI22_X1 U13908 ( .A1(n13713), .A2(n13697), .B1(n11919), .B2(n13673), .ZN(
        n11920) );
  OAI21_X1 U13909 ( .B1(n12330), .B2(n13681), .A(n11920), .ZN(n11921) );
  AOI21_X1 U13910 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n13584), .A(n11921), .ZN(
        n11922) );
  OAI21_X1 U13911 ( .B1(n11923), .B2(n13675), .A(n11922), .ZN(P3_U3177) );
  MUX2_X1 U13912 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n7414), .Z(n12096) );
  XNOR2_X1 U13913 ( .A(n12096), .B(n12111), .ZN(n12094) );
  NAND2_X1 U13914 ( .A1(n11925), .A2(n11924), .ZN(n11930) );
  INV_X1 U13915 ( .A(n11926), .ZN(n11928) );
  NAND2_X1 U13916 ( .A1(n11928), .A2(n11927), .ZN(n11929) );
  NAND2_X1 U13917 ( .A1(n11930), .A2(n11929), .ZN(n16107) );
  MUX2_X1 U13918 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13791), .Z(n11931) );
  INV_X1 U13919 ( .A(n16108), .ZN(n11932) );
  XNOR2_X1 U13920 ( .A(n11931), .B(n11932), .ZN(n16106) );
  NAND2_X1 U13921 ( .A1(n16107), .A2(n16106), .ZN(n11935) );
  INV_X1 U13922 ( .A(n11931), .ZN(n11933) );
  NAND2_X1 U13923 ( .A1(n11933), .A2(n11932), .ZN(n11934) );
  NAND2_X1 U13924 ( .A1(n11935), .A2(n11934), .ZN(n12095) );
  XOR2_X1 U13925 ( .A(n12094), .B(n12095), .Z(n11954) );
  INV_X1 U13926 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U13927 ( .A1(n16108), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11939) );
  OR2_X1 U13928 ( .A1(n16108), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U13929 ( .A1(n11939), .A2(n11938), .ZN(n16111) );
  XOR2_X1 U13930 ( .A(n12110), .B(n12101), .Z(n12109) );
  XNOR2_X1 U13931 ( .A(n12744), .B(n12109), .ZN(n11952) );
  NOR2_X1 U13932 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15512), .ZN(n12662) );
  AOI21_X1 U13933 ( .B1(n16252), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12662), .ZN(
        n11950) );
  NAND2_X1 U13934 ( .A1(n16108), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11946) );
  INV_X1 U13935 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11940) );
  MUX2_X1 U13936 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n11940), .S(n16108), .Z(
        n16114) );
  NAND2_X1 U13937 ( .A1(n11942), .A2(n11941), .ZN(n11944) );
  NAND2_X1 U13938 ( .A1(n11944), .A2(n11943), .ZN(n16113) );
  NAND2_X1 U13939 ( .A1(n16114), .A2(n16113), .ZN(n11945) );
  NAND2_X1 U13940 ( .A1(n11946), .A2(n11945), .ZN(n12100) );
  XNOR2_X1 U13941 ( .A(n12100), .B(n12111), .ZN(n11947) );
  NAND2_X1 U13942 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n11947), .ZN(n12102) );
  OAI21_X1 U13943 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11947), .A(n12102), .ZN(
        n11948) );
  NAND2_X1 U13944 ( .A1(n11948), .A2(n16262), .ZN(n11949) );
  OAI211_X1 U13945 ( .C1(n16244), .C2(n12101), .A(n11950), .B(n11949), .ZN(
        n11951) );
  AOI21_X1 U13946 ( .B1(n16265), .B2(n11952), .A(n11951), .ZN(n11953) );
  OAI21_X1 U13947 ( .B1(n11954), .B2(n16190), .A(n11953), .ZN(P3_U3189) );
  INV_X1 U13948 ( .A(n14764), .ZN(n11957) );
  INV_X1 U13949 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11955) );
  NOR2_X1 U13950 ( .A1(n16595), .A2(n11955), .ZN(n11956) );
  AOI21_X1 U13951 ( .B1(n11957), .B2(n12045), .A(n11956), .ZN(n11958) );
  OAI21_X1 U13952 ( .B1(n11959), .B2(n16592), .A(n11958), .ZN(P2_U3439) );
  XNOR2_X1 U13953 ( .A(n12088), .B(n14244), .ZN(n11964) );
  OR2_X1 U13954 ( .A1(n12247), .A2(n12771), .ZN(n11965) );
  NAND2_X1 U13955 ( .A1(n11964), .A2(n11965), .ZN(n11976) );
  INV_X1 U13956 ( .A(n11964), .ZN(n11967) );
  INV_X1 U13957 ( .A(n11965), .ZN(n11966) );
  NAND2_X1 U13958 ( .A1(n11967), .A2(n11966), .ZN(n11968) );
  NAND2_X1 U13959 ( .A1(n11976), .A2(n11968), .ZN(n11969) );
  AOI21_X1 U13960 ( .B1(n11970), .B2(n11969), .A(n7572), .ZN(n11975) );
  OAI21_X1 U13961 ( .B1(n14320), .B2(n12352), .A(n11971), .ZN(n11973) );
  OAI22_X1 U13962 ( .A1(n14281), .A2(n12079), .B1(n12090), .B2(n14355), .ZN(
        n11972) );
  AOI211_X1 U13963 ( .C1(n12088), .C2(n14324), .A(n11973), .B(n11972), .ZN(
        n11974) );
  OAI21_X1 U13964 ( .B1(n11975), .B2(n14326), .A(n11974), .ZN(P2_U3185) );
  XNOR2_X1 U13965 ( .A(n12142), .B(n14244), .ZN(n11977) );
  OR2_X1 U13966 ( .A1(n12352), .A2(n12771), .ZN(n11978) );
  INV_X1 U13967 ( .A(n11977), .ZN(n11980) );
  INV_X1 U13968 ( .A(n11978), .ZN(n11979) );
  NAND2_X1 U13969 ( .A1(n11980), .A2(n11979), .ZN(n12348) );
  NAND2_X1 U13970 ( .A1(n7470), .A2(n12348), .ZN(n11981) );
  XNOR2_X1 U13971 ( .A(n12347), .B(n11981), .ZN(n11986) );
  OAI21_X1 U13972 ( .B1(n14320), .B2(n12475), .A(n11982), .ZN(n11984) );
  OAI22_X1 U13973 ( .A1(n14281), .A2(n12247), .B1(n12136), .B2(n14355), .ZN(
        n11983) );
  AOI211_X1 U13974 ( .C1(n12142), .C2(n14324), .A(n11984), .B(n11983), .ZN(
        n11985) );
  OAI21_X1 U13975 ( .B1(n11986), .B2(n14326), .A(n11985), .ZN(P2_U3193) );
  OAI22_X1 U13976 ( .A1(n14149), .A2(n11988), .B1(n16615), .B2(n11987), .ZN(
        n11989) );
  AOI21_X1 U13977 ( .B1(n12439), .B2(n16615), .A(n11989), .ZN(n11990) );
  INV_X1 U13978 ( .A(n11990), .ZN(P3_U3459) );
  XNOR2_X1 U13979 ( .A(n11991), .B(n11994), .ZN(n12001) );
  OAI21_X1 U13980 ( .B1(n11994), .B2(n11993), .A(n11992), .ZN(n11995) );
  NAND2_X1 U13981 ( .A1(n11995), .A2(n16631), .ZN(n11999) );
  OAI22_X1 U13982 ( .A1(n11996), .A2(n15216), .B1(n15218), .B2(n12166), .ZN(
        n11997) );
  INV_X1 U13983 ( .A(n11997), .ZN(n11998) );
  OAI211_X1 U13984 ( .C1(n12001), .C2(n16324), .A(n11999), .B(n11998), .ZN(
        n16402) );
  MUX2_X1 U13985 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n16402), .S(n7416), .Z(
        n12000) );
  INV_X1 U13986 ( .A(n12000), .ZN(n12010) );
  INV_X1 U13987 ( .A(n16323), .ZN(n16297) );
  NAND2_X1 U13988 ( .A1(n7416), .A2(n16297), .ZN(n12233) );
  INV_X1 U13989 ( .A(n12233), .ZN(n16361) );
  INV_X1 U13990 ( .A(n12001), .ZN(n16404) );
  INV_X1 U13991 ( .A(n12002), .ZN(n16378) );
  NAND2_X1 U13992 ( .A1(n16378), .A2(n12003), .ZN(n12004) );
  AND3_X1 U13993 ( .A1(n12004), .A2(n16622), .A3(n12185), .ZN(n16399) );
  NAND2_X1 U13994 ( .A1(n16498), .A2(n16399), .ZN(n12006) );
  OR2_X1 U13995 ( .A1(n16493), .A2(n16401), .ZN(n12005) );
  OAI211_X1 U13996 ( .C1(n16653), .C2(n12007), .A(n12006), .B(n12005), .ZN(
        n12008) );
  AOI21_X1 U13997 ( .B1(n16361), .B2(n16404), .A(n12008), .ZN(n12009) );
  NAND2_X1 U13998 ( .A1(n12010), .A2(n12009), .ZN(P1_U3288) );
  INV_X1 U13999 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n12011) );
  OAI22_X1 U14000 ( .A1(n14764), .A2(n12071), .B1(n16595), .B2(n12011), .ZN(
        n12012) );
  INV_X1 U14001 ( .A(n12012), .ZN(n12013) );
  OAI21_X1 U14002 ( .B1(n12014), .B2(n16592), .A(n12013), .ZN(P2_U3445) );
  INV_X1 U14003 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n12015) );
  OAI22_X1 U14004 ( .A1(n14764), .A2(n12054), .B1(n16595), .B2(n12015), .ZN(
        n12016) );
  INV_X1 U14005 ( .A(n12016), .ZN(n12017) );
  OAI21_X1 U14006 ( .B1(n12018), .B2(n16592), .A(n12017), .ZN(P2_U3433) );
  INV_X1 U14007 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n12019) );
  OAI22_X1 U14008 ( .A1(n14764), .A2(n12271), .B1(n16595), .B2(n12019), .ZN(
        n12020) );
  INV_X1 U14009 ( .A(n12020), .ZN(n12021) );
  OAI21_X1 U14010 ( .B1(n12022), .B2(n16592), .A(n12021), .ZN(P2_U3436) );
  INV_X1 U14011 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n12023) );
  OAI22_X1 U14012 ( .A1(n14764), .A2(n12303), .B1(n16595), .B2(n12023), .ZN(
        n12024) );
  INV_X1 U14013 ( .A(n12024), .ZN(n12025) );
  OAI21_X1 U14014 ( .B1(n12026), .B2(n16592), .A(n12025), .ZN(P2_U3442) );
  XNOR2_X1 U14015 ( .A(n12027), .B(n12036), .ZN(n12029) );
  AOI21_X1 U14016 ( .B1(n12029), .B2(n16631), .A(n12028), .ZN(n16373) );
  INV_X1 U14017 ( .A(n16379), .ZN(n12032) );
  AND2_X1 U14018 ( .A1(n16365), .A2(n16344), .ZN(n12030) );
  NOR2_X1 U14019 ( .A1(n12030), .A2(n16566), .ZN(n12031) );
  AND2_X1 U14020 ( .A1(n12032), .A2(n12031), .ZN(n16367) );
  INV_X1 U14021 ( .A(n16653), .ZN(n16490) );
  AOI22_X1 U14022 ( .A1(n16398), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n16490), 
        .B2(n14973), .ZN(n12033) );
  OAI21_X1 U14023 ( .B1(n12034), .B2(n16493), .A(n12033), .ZN(n12039) );
  INV_X1 U14024 ( .A(n16324), .ZN(n16370) );
  NAND2_X1 U14025 ( .A1(n7416), .A2(n16370), .ZN(n12035) );
  XNOR2_X1 U14026 ( .A(n12037), .B(n12036), .ZN(n16368) );
  NOR2_X1 U14027 ( .A1(n15247), .A2(n16368), .ZN(n12038) );
  AOI211_X1 U14028 ( .C1(n16367), .C2(n16498), .A(n12039), .B(n12038), .ZN(
        n12040) );
  OAI21_X1 U14029 ( .B1(n16398), .B2(n16373), .A(n12040), .ZN(P1_U3290) );
  INV_X1 U14030 ( .A(n12041), .ZN(n12051) );
  INV_X1 U14031 ( .A(n12042), .ZN(n12043) );
  MUX2_X1 U14032 ( .A(n12044), .B(n12043), .S(n14610), .Z(n12050) );
  INV_X1 U14033 ( .A(n12045), .ZN(n12046) );
  OAI22_X1 U14034 ( .A1(n14621), .A2(n12046), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14640), .ZN(n12047) );
  AOI21_X1 U14035 ( .B1(n14645), .B2(n12048), .A(n12047), .ZN(n12049) );
  OAI211_X1 U14036 ( .C1(n14648), .C2(n12051), .A(n12050), .B(n12049), .ZN(
        P2_U3262) );
  INV_X1 U14037 ( .A(n12052), .ZN(n12062) );
  OAI22_X1 U14038 ( .A1(n14621), .A2(n12054), .B1(n14640), .B2(n12053), .ZN(
        n12055) );
  AOI21_X1 U14039 ( .B1(n14645), .B2(n12056), .A(n12055), .ZN(n12061) );
  INV_X1 U14040 ( .A(n12057), .ZN(n12059) );
  MUX2_X1 U14041 ( .A(n12059), .B(n12058), .S(n16598), .Z(n12060) );
  OAI211_X1 U14042 ( .C1(n14648), .C2(n12062), .A(n12061), .B(n12060), .ZN(
        P2_U3264) );
  INV_X1 U14043 ( .A(n12063), .ZN(n12065) );
  OAI222_X1 U14044 ( .A1(n15810), .A2(n12064), .B1(n15805), .B2(n12065), .C1(
        n15044), .C2(P1_U3086), .ZN(P1_U3338) );
  OAI222_X1 U14045 ( .A1(n14792), .A2(n12066), .B1(n14775), .B2(n12065), .C1(
        n13105), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U14046 ( .A(n12067), .ZN(n12076) );
  MUX2_X1 U14047 ( .A(n12068), .B(P2_REG2_REG_5__SCAN_IN), .S(n16598), .Z(
        n12069) );
  INV_X1 U14048 ( .A(n12069), .ZN(n12075) );
  OAI22_X1 U14049 ( .A1(n14621), .A2(n12071), .B1(n14640), .B2(n12070), .ZN(
        n12072) );
  AOI21_X1 U14050 ( .B1(n12073), .B2(n14645), .A(n12072), .ZN(n12074) );
  OAI211_X1 U14051 ( .C1(n12076), .C2(n14613), .A(n12075), .B(n12074), .ZN(
        P2_U3260) );
  OAI21_X1 U14052 ( .B1(n12078), .B2(n12082), .A(n12077), .ZN(n12085) );
  INV_X1 U14053 ( .A(n12085), .ZN(n12149) );
  OAI22_X1 U14054 ( .A1(n12079), .A2(n14602), .B1(n12352), .B2(n14604), .ZN(
        n12084) );
  INV_X1 U14055 ( .A(n12130), .ZN(n12080) );
  AOI211_X1 U14056 ( .C1(n12082), .C2(n12081), .A(n14510), .B(n12080), .ZN(
        n12083) );
  AOI211_X1 U14057 ( .C1(n12254), .C2(n12085), .A(n12084), .B(n12083), .ZN(
        n12147) );
  MUX2_X1 U14058 ( .A(n12086), .B(n12147), .S(n14610), .Z(n12093) );
  AOI21_X1 U14059 ( .B1(n12088), .B2(n7850), .A(n11533), .ZN(n12089) );
  AND2_X1 U14060 ( .A1(n12138), .A2(n12089), .ZN(n12145) );
  OAI22_X1 U14061 ( .A1(n12153), .A2(n14621), .B1(n14640), .B2(n12090), .ZN(
        n12091) );
  AOI21_X1 U14062 ( .B1(n12145), .B2(n14645), .A(n12091), .ZN(n12092) );
  OAI211_X1 U14063 ( .C1(n12149), .C2(n14613), .A(n12093), .B(n12092), .ZN(
        P2_U3258) );
  MUX2_X1 U14064 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n7414), .Z(n12278) );
  INV_X1 U14065 ( .A(n12283), .ZN(n12279) );
  XNOR2_X1 U14066 ( .A(n12278), .B(n12279), .ZN(n12276) );
  NAND2_X1 U14067 ( .A1(n12095), .A2(n12094), .ZN(n12099) );
  INV_X1 U14068 ( .A(n12096), .ZN(n12097) );
  NAND2_X1 U14069 ( .A1(n12097), .A2(n12111), .ZN(n12098) );
  NAND2_X1 U14070 ( .A1(n12099), .A2(n12098), .ZN(n12277) );
  XOR2_X1 U14071 ( .A(n12277), .B(n12276), .Z(n12122) );
  NAND2_X1 U14072 ( .A1(n12101), .A2(n12100), .ZN(n12103) );
  INV_X1 U14073 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12104) );
  MUX2_X1 U14074 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n12104), .S(n12283), .Z(
        n12105) );
  OAI21_X1 U14075 ( .B1(n12106), .B2(n12105), .A(n12284), .ZN(n12120) );
  INV_X1 U14076 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12107) );
  NOR2_X1 U14077 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12107), .ZN(n12796) );
  AOI21_X1 U14078 ( .B1(n16252), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12796), .ZN(
        n12108) );
  OAI21_X1 U14079 ( .B1(n16244), .B2(n12283), .A(n12108), .ZN(n12119) );
  NAND2_X1 U14080 ( .A1(n12283), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12288) );
  OR2_X1 U14081 ( .A1(n12283), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12112) );
  NAND2_X1 U14082 ( .A1(n12288), .A2(n12112), .ZN(n12115) );
  INV_X1 U14083 ( .A(n12114), .ZN(n12116) );
  NAND2_X1 U14084 ( .A1(n12116), .A2(n12115), .ZN(n12117) );
  AOI21_X1 U14085 ( .B1(n12289), .B2(n12117), .A(n16250), .ZN(n12118) );
  AOI211_X1 U14086 ( .C1(n16262), .C2(n12120), .A(n12119), .B(n12118), .ZN(
        n12121) );
  OAI21_X1 U14087 ( .B1(n12122), .B2(n16190), .A(n12121), .ZN(P3_U3190) );
  NAND2_X1 U14088 ( .A1(n12123), .A2(n12128), .ZN(n12124) );
  NAND2_X1 U14089 ( .A1(n12125), .A2(n12124), .ZN(n16455) );
  AOI22_X1 U14090 ( .A1(n12126), .A2(n14578), .B1(n14575), .B2(n14379), .ZN(
        n12135) );
  INV_X1 U14091 ( .A(n12127), .ZN(n12129) );
  AOI21_X1 U14092 ( .B1(n12130), .B2(n12129), .A(n12128), .ZN(n12133) );
  INV_X1 U14093 ( .A(n12131), .ZN(n12132) );
  OAI21_X1 U14094 ( .B1(n12133), .B2(n12132), .A(n16584), .ZN(n12134) );
  OAI211_X1 U14095 ( .C1(n16455), .C2(n14609), .A(n12135), .B(n12134), .ZN(
        n16457) );
  NAND2_X1 U14096 ( .A1(n16457), .A2(n14610), .ZN(n12144) );
  OAI22_X1 U14097 ( .A1(n14610), .A2(n12137), .B1(n12136), .B2(n14640), .ZN(
        n12141) );
  INV_X1 U14098 ( .A(n12138), .ZN(n12139) );
  OAI211_X1 U14099 ( .C1(n8299), .C2(n12139), .A(n12206), .B(n12771), .ZN(
        n16456) );
  NOR2_X1 U14100 ( .A1(n16456), .A2(n16601), .ZN(n12140) );
  AOI211_X1 U14101 ( .C1(n16599), .C2(n12142), .A(n12141), .B(n12140), .ZN(
        n12143) );
  OAI211_X1 U14102 ( .C1(n16455), .C2(n14613), .A(n12144), .B(n12143), .ZN(
        P2_U3257) );
  INV_X1 U14103 ( .A(n12145), .ZN(n12146) );
  OAI211_X1 U14104 ( .C1(n12149), .C2(n12148), .A(n12147), .B(n12146), .ZN(
        n12155) );
  OAI22_X1 U14105 ( .A1(n14708), .A2(n12153), .B1(n16591), .B2(n12150), .ZN(
        n12151) );
  AOI21_X1 U14106 ( .B1(n12155), .B2(n16591), .A(n12151), .ZN(n12152) );
  INV_X1 U14107 ( .A(n12152), .ZN(P2_U3506) );
  OAI22_X1 U14108 ( .A1(n14764), .A2(n12153), .B1(n16595), .B2(n10050), .ZN(
        n12154) );
  AOI21_X1 U14109 ( .B1(n12155), .B2(n16595), .A(n12154), .ZN(n12156) );
  INV_X1 U14110 ( .A(n12156), .ZN(P2_U3451) );
  OAI21_X1 U14111 ( .B1(n12160), .B2(n12163), .A(n12159), .ZN(n12242) );
  OAI211_X1 U14112 ( .C1(n12162), .C2(n12161), .A(n16622), .B(n12227), .ZN(
        n12238) );
  OAI21_X1 U14113 ( .B1(n12162), .B2(n16624), .A(n12238), .ZN(n12171) );
  AOI21_X1 U14114 ( .B1(n12164), .B2(n12163), .A(n16351), .ZN(n12168) );
  OAI22_X1 U14115 ( .A1(n12166), .A2(n15216), .B1(n15218), .B2(n12888), .ZN(
        n12167) );
  AOI21_X1 U14116 ( .B1(n12168), .B2(n12165), .A(n12167), .ZN(n12170) );
  NAND2_X1 U14117 ( .A1(n12242), .A2(n16370), .ZN(n12169) );
  NAND2_X1 U14118 ( .A1(n12170), .A2(n12169), .ZN(n12239) );
  AOI211_X1 U14119 ( .C1(n16452), .C2(n12242), .A(n12171), .B(n12239), .ZN(
        n12173) );
  OR2_X1 U14120 ( .A1(n12173), .A2(n16636), .ZN(n12172) );
  OAI21_X1 U14121 ( .B1(n16638), .B2(n9293), .A(n12172), .ZN(P1_U3480) );
  INV_X1 U14122 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15022) );
  OR2_X1 U14123 ( .A1(n12173), .A2(n16633), .ZN(n12174) );
  OAI21_X1 U14124 ( .B1(n16635), .B2(n15022), .A(n12174), .ZN(P1_U3535) );
  XNOR2_X1 U14125 ( .A(n12175), .B(n12176), .ZN(n16412) );
  INV_X1 U14126 ( .A(n12177), .ZN(n12181) );
  AND3_X1 U14127 ( .A1(n11992), .A2(n12179), .A3(n12178), .ZN(n12180) );
  OAI21_X1 U14128 ( .B1(n12181), .B2(n12180), .A(n16631), .ZN(n12183) );
  AOI22_X1 U14129 ( .A1(n15233), .A2(n14939), .B1(n15234), .B2(n14937), .ZN(
        n12182) );
  OAI211_X1 U14130 ( .C1(n16412), .C2(n16324), .A(n12183), .B(n12182), .ZN(
        n16414) );
  NAND2_X1 U14131 ( .A1(n16414), .A2(n7416), .ZN(n12191) );
  OAI22_X1 U14132 ( .A1(n7416), .A2(n11161), .B1(n12184), .B2(n16653), .ZN(
        n12188) );
  OAI211_X1 U14133 ( .C1(n7943), .C2(n7944), .A(n16622), .B(n12186), .ZN(
        n16413) );
  NOR2_X1 U14134 ( .A1(n16413), .A2(n16644), .ZN(n12187) );
  AOI211_X1 U14135 ( .C1(n16389), .C2(n12189), .A(n12188), .B(n12187), .ZN(
        n12190) );
  OAI211_X1 U14136 ( .C1(n16412), .C2(n12233), .A(n12191), .B(n12190), .ZN(
        P1_U3287) );
  OAI222_X1 U14137 ( .A1(n14221), .A2(n12194), .B1(n14223), .B2(n12193), .C1(
        P3_U3151), .C2(n12192), .ZN(P3_U3275) );
  XNOR2_X1 U14138 ( .A(n12196), .B(n12195), .ZN(n12314) );
  NAND2_X1 U14139 ( .A1(n7416), .A2(n16631), .ZN(n16647) );
  INV_X1 U14140 ( .A(n16647), .ZN(n12966) );
  OAI21_X1 U14141 ( .B1(n7469), .B2(n12197), .A(n8247), .ZN(n12312) );
  XNOR2_X1 U14142 ( .A(n12226), .B(n12891), .ZN(n12198) );
  AOI222_X1 U14143 ( .A1(n14934), .A2(n15234), .B1(n12198), .B2(n16622), .C1(
        n14936), .C2(n15233), .ZN(n12309) );
  OAI22_X1 U14144 ( .A1(n7416), .A2(n12199), .B1(n12886), .B2(n16653), .ZN(
        n12200) );
  AOI21_X1 U14145 ( .B1(n12891), .B2(n16389), .A(n12200), .ZN(n12201) );
  OAI21_X1 U14146 ( .B1(n12309), .B2(n16644), .A(n12201), .ZN(n12202) );
  AOI21_X1 U14147 ( .B1(n12966), .B2(n12312), .A(n12202), .ZN(n12203) );
  OAI21_X1 U14148 ( .B1(n12314), .B2(n16646), .A(n12203), .ZN(P1_U3284) );
  XNOR2_X1 U14149 ( .A(n12204), .B(n12205), .ZN(n12416) );
  AOI211_X1 U14150 ( .C1(n7849), .C2(n12206), .A(n11533), .B(n7570), .ZN(
        n12418) );
  NOR2_X1 U14151 ( .A1(n12421), .A2(n14621), .ZN(n12209) );
  OAI22_X1 U14152 ( .A1(n14610), .A2(n12207), .B1(n12351), .B2(n14640), .ZN(
        n12208) );
  AOI211_X1 U14153 ( .C1(n12418), .C2(n14645), .A(n12209), .B(n12208), .ZN(
        n12216) );
  OAI21_X1 U14154 ( .B1(n12211), .B2(n12210), .A(n12373), .ZN(n12213) );
  OAI22_X1 U14155 ( .A1(n12352), .A2(n14602), .B1(n12634), .B2(n14604), .ZN(
        n12212) );
  AOI21_X1 U14156 ( .B1(n12213), .B2(n16584), .A(n12212), .ZN(n12214) );
  OAI21_X1 U14157 ( .B1(n12416), .B2(n14609), .A(n12214), .ZN(n12417) );
  NAND2_X1 U14158 ( .A1(n12417), .A2(n14610), .ZN(n12215) );
  OAI211_X1 U14159 ( .C1(n12416), .C2(n14613), .A(n12216), .B(n12215), .ZN(
        P2_U3256) );
  OAI21_X1 U14160 ( .B1(n12218), .B2(n12221), .A(n12217), .ZN(n16445) );
  OAI22_X1 U14161 ( .A1(n12570), .A2(n15216), .B1(n15218), .B2(n12925), .ZN(
        n12219) );
  INV_X1 U14162 ( .A(n12219), .ZN(n12224) );
  XNOR2_X1 U14163 ( .A(n12220), .B(n12221), .ZN(n12222) );
  NAND2_X1 U14164 ( .A1(n12222), .A2(n16631), .ZN(n12223) );
  OAI211_X1 U14165 ( .C1(n16445), .C2(n16324), .A(n12224), .B(n12223), .ZN(
        n16449) );
  MUX2_X1 U14166 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n16449), .S(n7416), .Z(
        n12225) );
  INV_X1 U14167 ( .A(n12225), .ZN(n12232) );
  INV_X1 U14168 ( .A(n12226), .ZN(n12229) );
  NAND2_X1 U14169 ( .A1(n12227), .A2(n12573), .ZN(n12228) );
  AND3_X1 U14170 ( .A1(n12229), .A2(n16622), .A3(n12228), .ZN(n16446) );
  INV_X1 U14171 ( .A(n12573), .ZN(n16448) );
  OAI22_X1 U14172 ( .A1(n16448), .A2(n16493), .B1(n16653), .B2(n12569), .ZN(
        n12230) );
  AOI21_X1 U14173 ( .B1(n16446), .B2(n16498), .A(n12230), .ZN(n12231) );
  OAI211_X1 U14174 ( .C1(n16445), .C2(n12233), .A(n12232), .B(n12231), .ZN(
        P1_U3285) );
  INV_X1 U14175 ( .A(n12234), .ZN(n12235) );
  AOI22_X1 U14176 ( .A1(n16389), .A2(n12236), .B1(n12235), .B2(n16490), .ZN(
        n12237) );
  OAI21_X1 U14177 ( .B1(n12238), .B2(n16644), .A(n12237), .ZN(n12241) );
  MUX2_X1 U14178 ( .A(n12239), .B(P1_REG2_REG_7__SCAN_IN), .S(n16398), .Z(
        n12240) );
  AOI211_X1 U14179 ( .C1(n16361), .C2(n12242), .A(n12241), .B(n12240), .ZN(
        n12243) );
  INV_X1 U14180 ( .A(n12243), .ZN(P1_U3286) );
  OAI21_X1 U14181 ( .B1(n7579), .B2(n12245), .A(n12244), .ZN(n12249) );
  NAND2_X1 U14182 ( .A1(n14382), .A2(n14578), .ZN(n12246) );
  OAI21_X1 U14183 ( .B1(n12247), .B2(n14604), .A(n12246), .ZN(n12248) );
  AOI21_X1 U14184 ( .B1(n12249), .B2(n16584), .A(n12248), .ZN(n12256) );
  OR2_X1 U14185 ( .A1(n12251), .A2(n12250), .ZN(n12252) );
  NAND2_X1 U14186 ( .A1(n12253), .A2(n12252), .ZN(n16423) );
  NAND2_X1 U14187 ( .A1(n16423), .A2(n12254), .ZN(n12255) );
  INV_X1 U14188 ( .A(n14613), .ZN(n12264) );
  AOI21_X1 U14189 ( .B1(n16419), .B2(n12257), .A(n11533), .ZN(n12258) );
  NAND2_X1 U14190 ( .A1(n12258), .A2(n7850), .ZN(n16421) );
  OAI22_X1 U14191 ( .A1(n14610), .A2(n12260), .B1(n12259), .B2(n14640), .ZN(
        n12261) );
  AOI21_X1 U14192 ( .B1(n16599), .B2(n16419), .A(n12261), .ZN(n12262) );
  OAI21_X1 U14193 ( .B1(n16421), .B2(n16601), .A(n12262), .ZN(n12263) );
  AOI21_X1 U14194 ( .B1(n16423), .B2(n12264), .A(n12263), .ZN(n12265) );
  OAI21_X1 U14195 ( .B1(n16425), .B2(n16598), .A(n12265), .ZN(P2_U3259) );
  INV_X1 U14196 ( .A(n12266), .ZN(n12275) );
  NAND2_X1 U14197 ( .A1(n14645), .A2(n12267), .ZN(n12270) );
  NOR2_X1 U14198 ( .A1(n14640), .A2(n9985), .ZN(n12268) );
  AOI21_X1 U14199 ( .B1(n16598), .B2(P2_REG2_REG_2__SCAN_IN), .A(n12268), .ZN(
        n12269) );
  OAI211_X1 U14200 ( .C1(n12271), .C2(n14621), .A(n12270), .B(n12269), .ZN(
        n12272) );
  AOI21_X1 U14201 ( .B1(n16604), .B2(n12273), .A(n12272), .ZN(n12274) );
  OAI21_X1 U14202 ( .B1(n16598), .B2(n12275), .A(n12274), .ZN(P2_U3263) );
  MUX2_X1 U14203 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13791), .Z(n12676) );
  XNOR2_X1 U14204 ( .A(n12676), .B(n12688), .ZN(n12674) );
  NAND2_X1 U14205 ( .A1(n12277), .A2(n12276), .ZN(n12282) );
  INV_X1 U14206 ( .A(n12278), .ZN(n12280) );
  NAND2_X1 U14207 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  NAND2_X1 U14208 ( .A1(n12282), .A2(n12281), .ZN(n12675) );
  XOR2_X1 U14209 ( .A(n12674), .B(n12675), .Z(n12297) );
  NAND2_X1 U14210 ( .A1(n12283), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U14211 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n12286), .ZN(n12682) );
  OAI21_X1 U14212 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n12286), .A(n12682), .ZN(
        n12295) );
  AND2_X1 U14213 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12827) );
  AOI21_X1 U14214 ( .B1(n16252), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12827), .ZN(
        n12287) );
  OAI21_X1 U14215 ( .B1(n16244), .B2(n12681), .A(n12287), .ZN(n12294) );
  INV_X1 U14216 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12290) );
  AOI21_X1 U14217 ( .B1(n12291), .B2(n12290), .A(n12689), .ZN(n12292) );
  NOR2_X1 U14218 ( .A1(n12292), .A2(n16250), .ZN(n12293) );
  AOI211_X1 U14219 ( .C1(n16262), .C2(n12295), .A(n12294), .B(n12293), .ZN(
        n12296) );
  OAI21_X1 U14220 ( .B1(n12297), .B2(n16190), .A(n12296), .ZN(P3_U3191) );
  INV_X1 U14221 ( .A(n12298), .ZN(n12307) );
  NAND2_X1 U14222 ( .A1(n12299), .A2(n14645), .ZN(n12302) );
  AOI22_X1 U14223 ( .A1(n16598), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n12300), 
        .B2(n16596), .ZN(n12301) );
  OAI211_X1 U14224 ( .C1(n12303), .C2(n14621), .A(n12302), .B(n12301), .ZN(
        n12304) );
  AOI21_X1 U14225 ( .B1(n16604), .B2(n12305), .A(n12304), .ZN(n12306) );
  OAI21_X1 U14226 ( .B1(n16598), .B2(n12307), .A(n12306), .ZN(P2_U3261) );
  INV_X1 U14227 ( .A(n16452), .ZN(n12308) );
  OAI21_X1 U14228 ( .B1(n12310), .B2(n16624), .A(n12309), .ZN(n12311) );
  AOI21_X1 U14229 ( .B1(n16631), .B2(n12312), .A(n12311), .ZN(n12313) );
  OAI21_X1 U14230 ( .B1(n16628), .B2(n12314), .A(n12313), .ZN(n12317) );
  NAND2_X1 U14231 ( .A1(n12317), .A2(n16635), .ZN(n12315) );
  OAI21_X1 U14232 ( .B1(n16635), .B2(n12316), .A(n12315), .ZN(P1_U3537) );
  INV_X1 U14233 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U14234 ( .A1(n12317), .A2(n16638), .ZN(n12318) );
  OAI21_X1 U14235 ( .B1(n16638), .B2(n12319), .A(n12318), .ZN(P1_U3486) );
  INV_X1 U14236 ( .A(n12320), .ZN(n12321) );
  AOI211_X1 U14237 ( .C1(n12323), .C2(n12322), .A(n13675), .B(n12321), .ZN(
        n12327) );
  MUX2_X1 U14238 ( .A(n13694), .B(P3_STATE_REG_SCAN_IN), .S(
        P3_REG3_REG_3__SCAN_IN), .Z(n12325) );
  AOI22_X1 U14239 ( .A1(n13697), .A2(n13712), .B1(n12560), .B2(n13673), .ZN(
        n12324) );
  OAI211_X1 U14240 ( .C1(n13582), .C2(n13681), .A(n12325), .B(n12324), .ZN(
        n12326) );
  OR2_X1 U14241 ( .A1(n12327), .A2(n12326), .ZN(P3_U3158) );
  OAI21_X1 U14242 ( .B1(n8388), .B2(n8970), .A(n12329), .ZN(n16336) );
  OAI22_X1 U14243 ( .A1(n12330), .A2(n14087), .B1(n10438), .B2(n14089), .ZN(
        n12334) );
  XNOR2_X1 U14244 ( .A(n12331), .B(n8970), .ZN(n12332) );
  NOR2_X1 U14245 ( .A1(n12332), .A2(n14084), .ZN(n12333) );
  AOI211_X1 U14246 ( .C1(n16428), .C2(n16336), .A(n12334), .B(n12333), .ZN(
        n16334) );
  OAI21_X1 U14247 ( .B1(n16609), .B2(n12335), .A(n16334), .ZN(n16338) );
  INV_X1 U14248 ( .A(n16338), .ZN(n12337) );
  NAND2_X1 U14249 ( .A1(n16618), .A2(n16521), .ZN(n14188) );
  INV_X1 U14250 ( .A(n14188), .ZN(n12515) );
  AOI22_X1 U14251 ( .A1(n16336), .A2(n12515), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n9044), .ZN(n12336) );
  OAI21_X1 U14252 ( .B1(n12337), .B2(n9044), .A(n12336), .ZN(P3_U3396) );
  INV_X1 U14253 ( .A(n15885), .ZN(n12339) );
  OAI222_X1 U14254 ( .A1(P2_U3088), .A2(n12339), .B1(n14775), .B2(n12341), 
        .C1(n12338), .C2(n14792), .ZN(P2_U3309) );
  INV_X1 U14255 ( .A(n13019), .ZN(n12763) );
  OAI222_X1 U14256 ( .A1(P1_U3086), .A2(n12763), .B1(n15805), .B2(n12341), 
        .C1(n12340), .C2(n15810), .ZN(P1_U3337) );
  INV_X1 U14257 ( .A(n14324), .ZN(n14362) );
  XNOR2_X1 U14258 ( .A(n7849), .B(n14244), .ZN(n12342) );
  NAND2_X1 U14259 ( .A1(n14379), .A2(n11533), .ZN(n12343) );
  NAND2_X1 U14260 ( .A1(n12342), .A2(n12343), .ZN(n12469) );
  INV_X1 U14261 ( .A(n12342), .ZN(n12345) );
  INV_X1 U14262 ( .A(n12343), .ZN(n12344) );
  NAND2_X1 U14263 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  AND2_X1 U14264 ( .A1(n12469), .A2(n12346), .ZN(n12349) );
  OAI21_X1 U14265 ( .B1(n12349), .B2(n7580), .A(n12470), .ZN(n12350) );
  NAND2_X1 U14266 ( .A1(n12350), .A2(n14352), .ZN(n12357) );
  NAND2_X1 U14267 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15926) );
  INV_X1 U14268 ( .A(n15926), .ZN(n12354) );
  OAI22_X1 U14269 ( .A1(n14281), .A2(n12352), .B1(n12351), .B2(n14355), .ZN(
        n12353) );
  AOI211_X1 U14270 ( .C1(n14331), .C2(n12355), .A(n12354), .B(n12353), .ZN(
        n12356) );
  OAI211_X1 U14271 ( .C1(n12421), .C2(n14362), .A(n12357), .B(n12356), .ZN(
        P2_U3203) );
  AOI21_X1 U14272 ( .B1(n7575), .B2(n12366), .A(n16351), .ZN(n12359) );
  AOI22_X1 U14273 ( .A1(n12359), .A2(n12358), .B1(n15233), .B2(n14935), .ZN(
        n12506) );
  OAI211_X1 U14274 ( .C1(n7947), .C2(n7577), .A(n16622), .B(n12613), .ZN(
        n12361) );
  OAI21_X1 U14275 ( .B1(n12924), .B2(n15218), .A(n12361), .ZN(n12504) );
  OAI22_X1 U14276 ( .A1(n7416), .A2(n12362), .B1(n12923), .B2(n16653), .ZN(
        n12364) );
  NOR2_X1 U14277 ( .A1(n7947), .A2(n16493), .ZN(n12363) );
  AOI211_X1 U14278 ( .C1(n12504), .C2(n16498), .A(n12364), .B(n12363), .ZN(
        n12369) );
  OAI21_X1 U14279 ( .B1(n12367), .B2(n12366), .A(n12365), .ZN(n12503) );
  NAND2_X1 U14280 ( .A1(n12503), .A2(n16394), .ZN(n12368) );
  OAI211_X1 U14281 ( .C1(n12506), .C2(n16398), .A(n12369), .B(n12368), .ZN(
        P1_U3283) );
  XNOR2_X1 U14282 ( .A(n12370), .B(n12371), .ZN(n16475) );
  AOI22_X1 U14283 ( .A1(n14578), .A2(n14379), .B1(n14378), .B2(n14575), .ZN(
        n12378) );
  AND2_X1 U14284 ( .A1(n12373), .A2(n12372), .ZN(n12376) );
  OAI211_X1 U14285 ( .C1(n12376), .C2(n12375), .A(n16584), .B(n12374), .ZN(
        n12377) );
  OAI211_X1 U14286 ( .C1(n16475), .C2(n14609), .A(n12378), .B(n12377), .ZN(
        n16477) );
  NAND2_X1 U14287 ( .A1(n16477), .A2(n14610), .ZN(n12383) );
  OAI22_X1 U14288 ( .A1(n14610), .A2(n12379), .B1(n12474), .B2(n14640), .ZN(
        n12381) );
  OAI211_X1 U14289 ( .C1(n7847), .C2(n7570), .A(n12771), .B(n12451), .ZN(
        n16476) );
  NOR2_X1 U14290 ( .A1(n16476), .A2(n16601), .ZN(n12380) );
  AOI211_X1 U14291 ( .C1(n16599), .C2(n12463), .A(n12381), .B(n12380), .ZN(
        n12382) );
  OAI211_X1 U14292 ( .C1(n16475), .C2(n14613), .A(n12383), .B(n12382), .ZN(
        P2_U3255) );
  INV_X1 U14293 ( .A(n12384), .ZN(n12385) );
  AOI21_X1 U14294 ( .B1(n12387), .B2(n12386), .A(n12385), .ZN(n12392) );
  OAI22_X1 U14295 ( .A1(n10438), .A2(n13681), .B1(n12850), .B2(n13671), .ZN(
        n12388) );
  AOI211_X1 U14296 ( .C1(n12654), .C2(n13673), .A(n12389), .B(n12388), .ZN(
        n12391) );
  NAND2_X1 U14297 ( .A1(n13683), .A2(n12653), .ZN(n12390) );
  OAI211_X1 U14298 ( .C1(n12392), .C2(n13675), .A(n12391), .B(n12390), .ZN(
        P3_U3170) );
  NOR2_X1 U14299 ( .A1(n8448), .A2(n16609), .ZN(n16304) );
  XNOR2_X1 U14300 ( .A(n12405), .B(n12393), .ZN(n12394) );
  NAND2_X1 U14301 ( .A1(n12394), .A2(n13979), .ZN(n12396) );
  AOI22_X1 U14302 ( .A1(n13714), .A2(n13986), .B1(n13987), .B2(n13585), .ZN(
        n12395) );
  NAND2_X1 U14303 ( .A1(n12396), .A2(n12395), .ZN(n16303) );
  AOI21_X1 U14304 ( .B1(n16304), .B2(n12397), .A(n16303), .ZN(n12412) );
  NAND2_X1 U14305 ( .A1(n12399), .A2(n12398), .ZN(n12400) );
  NAND2_X1 U14306 ( .A1(n12403), .A2(n12400), .ZN(n12401) );
  INV_X1 U14307 ( .A(n12404), .ZN(n12406) );
  INV_X1 U14308 ( .A(n13367), .ZN(n13361) );
  NOR2_X1 U14309 ( .A1(n13364), .A2(n13361), .ZN(n13522) );
  AOI21_X1 U14310 ( .B1(n12406), .B2(n12405), .A(n13522), .ZN(n16305) );
  AND2_X1 U14311 ( .A1(n13363), .A2(n16333), .ZN(n16335) );
  OR2_X1 U14312 ( .A1(n16428), .A2(n16335), .ZN(n12407) );
  NAND2_X1 U14313 ( .A1(n16340), .A2(n12407), .ZN(n13892) );
  INV_X1 U14314 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n12408) );
  OAI22_X1 U14315 ( .A1(n16340), .A2(n12409), .B1(n12408), .B2(n14073), .ZN(
        n12410) );
  AOI21_X1 U14316 ( .B1(n16305), .B2(n14098), .A(n12410), .ZN(n12411) );
  OAI21_X1 U14317 ( .B1(n12412), .B2(n14100), .A(n12411), .ZN(P3_U3232) );
  OAI222_X1 U14318 ( .A1(n14221), .A2(n12415), .B1(n14223), .B2(n12414), .C1(
        P3_U3151), .C2(n12413), .ZN(P3_U3274) );
  INV_X1 U14319 ( .A(n12416), .ZN(n12419) );
  AOI211_X1 U14320 ( .C1(n16514), .C2(n12419), .A(n12418), .B(n12417), .ZN(
        n12424) );
  AOI22_X1 U14321 ( .A1(n7849), .A2(n12643), .B1(n16589), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n12420) );
  OAI21_X1 U14322 ( .B1(n12424), .B2(n16589), .A(n12420), .ZN(P2_U3508) );
  OAI22_X1 U14323 ( .A1(n12421), .A2(n14764), .B1(n16595), .B2(n10082), .ZN(
        n12422) );
  INV_X1 U14324 ( .A(n12422), .ZN(n12423) );
  OAI21_X1 U14325 ( .B1(n12424), .B2(n16592), .A(n12423), .ZN(P2_U3457) );
  XNOR2_X1 U14326 ( .A(n12425), .B(n12429), .ZN(n12557) );
  OAI22_X1 U14327 ( .A1(n12531), .A2(n14089), .B1(n13582), .B2(n14087), .ZN(
        n12431) );
  INV_X1 U14328 ( .A(n12426), .ZN(n12427) );
  AOI211_X1 U14329 ( .C1(n12429), .C2(n12428), .A(n14084), .B(n12427), .ZN(
        n12430) );
  AOI211_X1 U14330 ( .C1(n12557), .C2(n16428), .A(n12431), .B(n12430), .ZN(
        n12558) );
  INV_X1 U14331 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n12432) );
  OAI22_X1 U14332 ( .A1(n14207), .A2(n12436), .B1(n16618), .B2(n12432), .ZN(
        n12433) );
  AOI21_X1 U14333 ( .B1(n12557), .B2(n12515), .A(n12433), .ZN(n12434) );
  OAI21_X1 U14334 ( .B1(n12558), .B2(n9044), .A(n12434), .ZN(P3_U3399) );
  NAND2_X1 U14335 ( .A1(n16615), .A2(n16521), .ZN(n14130) );
  INV_X1 U14336 ( .A(n14130), .ZN(n16331) );
  INV_X1 U14337 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n12435) );
  OAI22_X1 U14338 ( .A1(n14149), .A2(n12436), .B1(n16615), .B2(n12435), .ZN(
        n12437) );
  AOI21_X1 U14339 ( .B1(n12557), .B2(n16331), .A(n12437), .ZN(n12438) );
  OAI21_X1 U14340 ( .B1(n12558), .B2(n9060), .A(n12438), .ZN(P3_U3462) );
  AOI21_X1 U14341 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n16337), .A(n12439), .ZN(
        n12445) );
  INV_X1 U14342 ( .A(n12440), .ZN(n12442) );
  NOR2_X1 U14343 ( .A1(n16609), .A2(n16333), .ZN(n12441) );
  AOI22_X1 U14344 ( .A1(n14095), .A2(n12443), .B1(n14100), .B2(
        P3_REG2_REG_0__SCAN_IN), .ZN(n12444) );
  OAI21_X1 U14345 ( .B1(n12445), .B2(n14100), .A(n12444), .ZN(P3_U3233) );
  OAI22_X1 U14346 ( .A1(n13544), .A2(P3_U3151), .B1(SI_22_), .B2(n14223), .ZN(
        n12446) );
  AOI21_X1 U14347 ( .B1(n12447), .B2(n14212), .A(n12446), .ZN(P3_U3273) );
  XNOR2_X1 U14348 ( .A(n12448), .B(n12449), .ZN(n12639) );
  INV_X1 U14349 ( .A(n12450), .ZN(n12601) );
  AOI211_X1 U14350 ( .C1(n12644), .C2(n12451), .A(n11533), .B(n12601), .ZN(
        n12641) );
  NOR2_X1 U14351 ( .A1(n12646), .A2(n14621), .ZN(n12454) );
  OAI22_X1 U14352 ( .A1(n14610), .A2(n12452), .B1(n12633), .B2(n14640), .ZN(
        n12453) );
  AOI211_X1 U14353 ( .C1(n12641), .C2(n14645), .A(n12454), .B(n12453), .ZN(
        n12462) );
  OAI21_X1 U14354 ( .B1(n12457), .B2(n12456), .A(n12455), .ZN(n12459) );
  OAI22_X1 U14355 ( .A1(n12772), .A2(n14604), .B1(n12634), .B2(n14602), .ZN(
        n12458) );
  AOI21_X1 U14356 ( .B1(n12459), .B2(n16584), .A(n12458), .ZN(n12460) );
  OAI21_X1 U14357 ( .B1(n12639), .B2(n14609), .A(n12460), .ZN(n12640) );
  NAND2_X1 U14358 ( .A1(n12640), .A2(n14610), .ZN(n12461) );
  OAI211_X1 U14359 ( .C1(n12639), .C2(n14613), .A(n12462), .B(n12461), .ZN(
        P2_U3254) );
  XNOR2_X1 U14360 ( .A(n12463), .B(n14244), .ZN(n12464) );
  OR2_X1 U14361 ( .A1(n12634), .A2(n12771), .ZN(n12465) );
  NAND2_X1 U14362 ( .A1(n12464), .A2(n12465), .ZN(n12627) );
  INV_X1 U14363 ( .A(n12464), .ZN(n12467) );
  INV_X1 U14364 ( .A(n12465), .ZN(n12466) );
  NAND2_X1 U14365 ( .A1(n12467), .A2(n12466), .ZN(n12468) );
  AND2_X1 U14366 ( .A1(n12627), .A2(n12468), .ZN(n12472) );
  NAND2_X1 U14367 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  OAI21_X1 U14368 ( .B1(n12472), .B2(n12471), .A(n12628), .ZN(n12473) );
  NAND2_X1 U14369 ( .A1(n12473), .A2(n14352), .ZN(n12479) );
  OAI22_X1 U14370 ( .A1(n14281), .A2(n12475), .B1(n12474), .B2(n14355), .ZN(
        n12476) );
  AOI211_X1 U14371 ( .C1(n14331), .C2(n14378), .A(n12477), .B(n12476), .ZN(
        n12478) );
  OAI211_X1 U14372 ( .C1(n7847), .C2(n14362), .A(n12479), .B(n12478), .ZN(
        P2_U3189) );
  XNOR2_X1 U14373 ( .A(n12480), .B(n13518), .ZN(n12650) );
  OAI211_X1 U14374 ( .C1(n12483), .C2(n12482), .A(n12481), .B(n13979), .ZN(
        n12485) );
  NAND2_X1 U14375 ( .A1(n13713), .A2(n13987), .ZN(n12484) );
  OAI211_X1 U14376 ( .C1(n12850), .C2(n14089), .A(n12485), .B(n12484), .ZN(
        n12486) );
  AOI21_X1 U14377 ( .B1(n12650), .B2(n16428), .A(n12486), .ZN(n12651) );
  OAI22_X1 U14378 ( .A1(n14149), .A2(n13379), .B1(n16615), .B2(n12487), .ZN(
        n12488) );
  AOI21_X1 U14379 ( .B1(n12650), .B2(n16331), .A(n12488), .ZN(n12489) );
  OAI21_X1 U14380 ( .B1(n12651), .B2(n9060), .A(n12489), .ZN(P3_U3463) );
  NAND2_X1 U14381 ( .A1(n12490), .A2(n13512), .ZN(n12491) );
  NAND2_X1 U14382 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  NAND2_X1 U14383 ( .A1(n12493), .A2(n13979), .ZN(n12497) );
  XNOR2_X1 U14384 ( .A(n12494), .B(n13512), .ZN(n12526) );
  NAND2_X1 U14385 ( .A1(n12526), .A2(n16428), .ZN(n12496) );
  AOI22_X1 U14386 ( .A1(n13986), .A2(n13709), .B1(n13712), .B2(n13987), .ZN(
        n12495) );
  NAND3_X1 U14387 ( .A1(n12497), .A2(n12496), .A3(n12495), .ZN(n12667) );
  INV_X1 U14388 ( .A(n12667), .ZN(n12502) );
  INV_X1 U14389 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n12498) );
  OAI22_X1 U14390 ( .A1(n14149), .A2(n12499), .B1(n16615), .B2(n12498), .ZN(
        n12500) );
  AOI21_X1 U14391 ( .B1(n12526), .B2(n16331), .A(n12500), .ZN(n12501) );
  OAI21_X1 U14392 ( .B1(n12502), .B2(n9060), .A(n12501), .ZN(P3_U3464) );
  INV_X1 U14393 ( .A(n12503), .ZN(n12507) );
  AOI21_X1 U14394 ( .B1(n12928), .B2(n16560), .A(n12504), .ZN(n12505) );
  OAI211_X1 U14395 ( .C1(n16628), .C2(n12507), .A(n12506), .B(n12505), .ZN(
        n12510) );
  NAND2_X1 U14396 ( .A1(n12510), .A2(n16635), .ZN(n12508) );
  OAI21_X1 U14397 ( .B1(n16635), .B2(n12509), .A(n12508), .ZN(P1_U3538) );
  NAND2_X1 U14398 ( .A1(n12510), .A2(n16638), .ZN(n12511) );
  OAI21_X1 U14399 ( .B1(n16638), .B2(n9363), .A(n12511), .ZN(P1_U3489) );
  INV_X1 U14400 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U14401 ( .A1(n12512), .A2(P3_U3897), .ZN(n12513) );
  OAI21_X1 U14402 ( .B1(P3_U3897), .B2(n12514), .A(n12513), .ZN(P3_U3520) );
  INV_X1 U14403 ( .A(n14207), .ZN(n14163) );
  AOI22_X1 U14404 ( .A1(n14163), .A2(n12654), .B1(P3_REG0_REG_4__SCAN_IN), 
        .B2(n9044), .ZN(n12517) );
  NAND2_X1 U14405 ( .A1(n12650), .A2(n12515), .ZN(n12516) );
  OAI211_X1 U14406 ( .C1(n12651), .C2(n9044), .A(n12517), .B(n12516), .ZN(
        P3_U3402) );
  INV_X1 U14407 ( .A(n12857), .ZN(n12525) );
  OAI211_X1 U14408 ( .C1(n12520), .C2(n12519), .A(n12518), .B(n13690), .ZN(
        n12524) );
  NAND2_X1 U14409 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n16121) );
  INV_X1 U14410 ( .A(n16121), .ZN(n12522) );
  OAI22_X1 U14411 ( .A1(n12850), .A2(n13681), .B1(n12988), .B2(n13671), .ZN(
        n12521) );
  AOI211_X1 U14412 ( .C1(n13391), .C2(n13673), .A(n12522), .B(n12521), .ZN(
        n12523) );
  OAI211_X1 U14413 ( .C1(n12525), .C2(n13694), .A(n12524), .B(n12523), .ZN(
        P3_U3179) );
  INV_X1 U14414 ( .A(n12526), .ZN(n12673) );
  NAND2_X1 U14415 ( .A1(n12667), .A2(n16618), .ZN(n12528) );
  AOI22_X1 U14416 ( .A1(n14163), .A2(n12670), .B1(P3_REG0_REG_5__SCAN_IN), 
        .B2(n9044), .ZN(n12527) );
  OAI211_X1 U14417 ( .C1(n12673), .C2(n14188), .A(n12528), .B(n12527), .ZN(
        P3_U3405) );
  XOR2_X1 U14418 ( .A(n12530), .B(n12529), .Z(n12536) );
  OAI22_X1 U14419 ( .A1(n13392), .A2(n13671), .B1(n12531), .B2(n13681), .ZN(
        n12532) );
  AOI211_X1 U14420 ( .C1(n12670), .C2(n13673), .A(n12533), .B(n12532), .ZN(
        n12535) );
  NAND2_X1 U14421 ( .A1(n13683), .A2(n12669), .ZN(n12534) );
  OAI211_X1 U14422 ( .C1(n12536), .C2(n13675), .A(n12535), .B(n12534), .ZN(
        P3_U3167) );
  INV_X1 U14423 ( .A(n12537), .ZN(n12539) );
  OAI222_X1 U14424 ( .A1(n15810), .A2(n12538), .B1(n15805), .B2(n12539), .C1(
        n13032), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U14425 ( .A1(n14792), .A2(n12540), .B1(n14775), .B2(n12539), .C1(
        P2_U3088), .C2(n13114), .ZN(P2_U3308) );
  OAI21_X1 U14426 ( .B1(n12542), .B2(n12553), .A(n12541), .ZN(n12818) );
  INV_X1 U14427 ( .A(n12818), .ZN(n12556) );
  AOI22_X1 U14428 ( .A1(n15233), .A2(n14933), .B1(n15234), .B2(n14931), .ZN(
        n13145) );
  INV_X1 U14429 ( .A(n13145), .ZN(n12544) );
  INV_X1 U14430 ( .A(n12543), .ZN(n13147) );
  AOI22_X1 U14431 ( .A1(n7416), .A2(n12544), .B1(n13147), .B2(n16490), .ZN(
        n12545) );
  OAI21_X1 U14432 ( .B1(n12546), .B2(n7416), .A(n12545), .ZN(n12550) );
  NAND2_X1 U14433 ( .A1(n12611), .A2(n12813), .ZN(n12547) );
  NAND3_X1 U14434 ( .A1(n12548), .A2(n16622), .A3(n12547), .ZN(n12814) );
  NOR2_X1 U14435 ( .A1(n12814), .A2(n16644), .ZN(n12549) );
  AOI211_X1 U14436 ( .C1(n16389), .C2(n12813), .A(n12550), .B(n12549), .ZN(
        n12555) );
  NAND2_X1 U14437 ( .A1(n12552), .A2(n12553), .ZN(n12815) );
  NAND3_X1 U14438 ( .A1(n12551), .A2(n12815), .A3(n12966), .ZN(n12554) );
  OAI211_X1 U14439 ( .C1(n12556), .C2(n15247), .A(n12555), .B(n12554), .ZN(
        P1_U3281) );
  INV_X1 U14440 ( .A(n12557), .ZN(n12563) );
  MUX2_X1 U14441 ( .A(n11829), .B(n12558), .S(n16340), .Z(n12562) );
  AOI22_X1 U14442 ( .A1(n14095), .A2(n12560), .B1(n16337), .B2(n12559), .ZN(
        n12561) );
  OAI211_X1 U14443 ( .C1(n12563), .C2(n14080), .A(n12562), .B(n12561), .ZN(
        P3_U3230) );
  OAI21_X1 U14444 ( .B1(n12566), .B2(n12565), .A(n12564), .ZN(n12567) );
  NAND2_X1 U14445 ( .A1(n12567), .A2(n14905), .ZN(n12575) );
  OAI22_X1 U14446 ( .A1(n16558), .A2(n12569), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12568), .ZN(n12572) );
  OAI22_X1 U14447 ( .A1(n12570), .A2(n16543), .B1(n16542), .B2(n12925), .ZN(
        n12571) );
  AOI211_X1 U14448 ( .C1(n12573), .C2(n16554), .A(n12572), .B(n12571), .ZN(
        n12574) );
  NAND2_X1 U14449 ( .A1(n12575), .A2(n12574), .ZN(P1_U3221) );
  INV_X1 U14450 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n16590) );
  OAI21_X1 U14451 ( .B1(n12805), .B2(n12577), .A(n12576), .ZN(n15863) );
  NOR2_X1 U14452 ( .A1(n15859), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12578) );
  AOI21_X1 U14453 ( .B1(n15859), .B2(P2_REG1_REG_14__SCAN_IN), .A(n12578), 
        .ZN(n15862) );
  NAND2_X1 U14454 ( .A1(n15863), .A2(n15862), .ZN(n15861) );
  OAI21_X1 U14455 ( .B1(n16590), .B2(n12579), .A(n15861), .ZN(n12717) );
  XNOR2_X1 U14456 ( .A(n12717), .B(n12725), .ZN(n12580) );
  NAND2_X1 U14457 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n12580), .ZN(n12719) );
  OAI211_X1 U14458 ( .C1(n12580), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15920), 
        .B(n12719), .ZN(n12590) );
  INV_X1 U14459 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U14460 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13061)
         );
  OAI21_X1 U14461 ( .B1(n15928), .B2(n12581), .A(n13061), .ZN(n12588) );
  XNOR2_X1 U14462 ( .A(n15859), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n15858) );
  AOI21_X1 U14463 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n12583), .A(n12582), 
        .ZN(n12584) );
  INV_X1 U14464 ( .A(n12584), .ZN(n15857) );
  OAI22_X1 U14465 ( .A1(n15858), .A2(n15857), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15859), .ZN(n12724) );
  XNOR2_X1 U14466 ( .A(n12724), .B(n12725), .ZN(n12586) );
  INV_X1 U14467 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12585) );
  NOR2_X1 U14468 ( .A1(n12585), .A2(n12586), .ZN(n12726) );
  AOI211_X1 U14469 ( .C1(n12586), .C2(n12585), .A(n12726), .B(n15897), .ZN(
        n12587) );
  AOI211_X1 U14470 ( .C1(n15922), .C2(n12718), .A(n12588), .B(n12587), .ZN(
        n12589) );
  NAND2_X1 U14471 ( .A1(n12590), .A2(n12589), .ZN(P2_U3229) );
  INV_X1 U14472 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U14473 ( .A1(n13829), .A2(P3_U3897), .ZN(n12591) );
  OAI21_X1 U14474 ( .B1(P3_U3897), .B2(n12592), .A(n12591), .ZN(P3_U3519) );
  XNOR2_X1 U14475 ( .A(n12593), .B(n12595), .ZN(n16508) );
  XOR2_X1 U14476 ( .A(n12595), .B(n12594), .Z(n12597) );
  OAI22_X1 U14477 ( .A1(n12784), .A2(n14602), .B1(n12864), .B2(n14604), .ZN(
        n12596) );
  AOI21_X1 U14478 ( .B1(n12597), .B2(n16584), .A(n12596), .ZN(n12598) );
  OAI21_X1 U14479 ( .B1(n16508), .B2(n14609), .A(n12598), .ZN(n16511) );
  NAND2_X1 U14480 ( .A1(n16511), .A2(n14610), .ZN(n12605) );
  OAI22_X1 U14481 ( .A1(n14610), .A2(n12599), .B1(n12783), .B2(n14640), .ZN(
        n12603) );
  INV_X1 U14482 ( .A(n12770), .ZN(n16510) );
  INV_X1 U14483 ( .A(n12600), .ZN(n12711) );
  OAI211_X1 U14484 ( .C1(n12601), .C2(n16510), .A(n12771), .B(n12711), .ZN(
        n16509) );
  NOR2_X1 U14485 ( .A1(n16509), .A2(n16601), .ZN(n12602) );
  AOI211_X1 U14486 ( .C1(n16599), .C2(n12770), .A(n12603), .B(n12602), .ZN(
        n12604) );
  OAI211_X1 U14487 ( .C1(n16508), .C2(n14613), .A(n12605), .B(n12604), .ZN(
        P2_U3253) );
  NAND2_X1 U14488 ( .A1(n12606), .A2(n14212), .ZN(n12607) );
  OAI211_X1 U14489 ( .C1(n12608), .C2(n14223), .A(n12607), .B(n13547), .ZN(
        P3_U3272) );
  INV_X1 U14490 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n12621) );
  OAI21_X1 U14491 ( .B1(n12610), .B2(n10621), .A(n12609), .ZN(n16495) );
  INV_X1 U14492 ( .A(n12611), .ZN(n12612) );
  AOI211_X1 U14493 ( .C1(n12614), .C2(n12613), .A(n16566), .B(n12612), .ZN(
        n16499) );
  AOI21_X1 U14494 ( .B1(n12614), .B2(n16560), .A(n16499), .ZN(n12619) );
  XNOR2_X1 U14495 ( .A(n12615), .B(n12616), .ZN(n12618) );
  AOI22_X1 U14496 ( .A1(n15233), .A2(n14934), .B1(n15234), .B2(n14932), .ZN(
        n13046) );
  INV_X1 U14497 ( .A(n13046), .ZN(n12617) );
  AOI21_X1 U14498 ( .B1(n12618), .B2(n16631), .A(n12617), .ZN(n16501) );
  OAI211_X1 U14499 ( .C1(n16628), .C2(n16495), .A(n12619), .B(n16501), .ZN(
        n15769) );
  NAND2_X1 U14500 ( .A1(n15769), .A2(n16638), .ZN(n12620) );
  OAI21_X1 U14501 ( .B1(n16638), .B2(n12621), .A(n12620), .ZN(P1_U3492) );
  XNOR2_X1 U14502 ( .A(n12644), .B(n14244), .ZN(n12622) );
  NAND2_X1 U14503 ( .A1(n14378), .A2(n11533), .ZN(n12623) );
  NAND2_X1 U14504 ( .A1(n12622), .A2(n12623), .ZN(n12778) );
  INV_X1 U14505 ( .A(n12622), .ZN(n12625) );
  INV_X1 U14506 ( .A(n12623), .ZN(n12624) );
  NAND2_X1 U14507 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  AND2_X1 U14508 ( .A1(n12778), .A2(n12626), .ZN(n12630) );
  OAI21_X1 U14509 ( .B1(n12630), .B2(n12629), .A(n12779), .ZN(n12631) );
  NAND2_X1 U14510 ( .A1(n12631), .A2(n14352), .ZN(n12638) );
  INV_X1 U14511 ( .A(n12632), .ZN(n12636) );
  OAI22_X1 U14512 ( .A1(n14281), .A2(n12634), .B1(n12633), .B2(n14355), .ZN(
        n12635) );
  AOI211_X1 U14513 ( .C1(n14331), .C2(n12702), .A(n12636), .B(n12635), .ZN(
        n12637) );
  OAI211_X1 U14514 ( .C1(n12646), .C2(n14362), .A(n12638), .B(n12637), .ZN(
        P2_U3208) );
  INV_X1 U14515 ( .A(n12639), .ZN(n12642) );
  AOI211_X1 U14516 ( .C1(n16514), .C2(n12642), .A(n12641), .B(n12640), .ZN(
        n12649) );
  AOI22_X1 U14517 ( .A1(n12644), .A2(n12643), .B1(n16589), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n12645) );
  OAI21_X1 U14518 ( .B1(n12649), .B2(n16589), .A(n12645), .ZN(P2_U3510) );
  OAI22_X1 U14519 ( .A1(n12646), .A2(n14764), .B1(n16595), .B2(n10110), .ZN(
        n12647) );
  INV_X1 U14520 ( .A(n12647), .ZN(n12648) );
  OAI21_X1 U14521 ( .B1(n12649), .B2(n16592), .A(n12648), .ZN(P2_U3463) );
  INV_X1 U14522 ( .A(n12650), .ZN(n12657) );
  INV_X1 U14523 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n12652) );
  MUX2_X1 U14524 ( .A(n12652), .B(n12651), .S(n16340), .Z(n12656) );
  AOI22_X1 U14525 ( .A1(n14095), .A2(n12654), .B1(n16337), .B2(n12653), .ZN(
        n12655) );
  OAI211_X1 U14526 ( .C1(n12657), .C2(n14080), .A(n12656), .B(n12655), .ZN(
        P3_U3229) );
  INV_X1 U14527 ( .A(n12658), .ZN(n12743) );
  NAND2_X1 U14528 ( .A1(n12660), .A2(n12659), .ZN(n12790) );
  OAI211_X1 U14529 ( .C1(n12660), .C2(n12659), .A(n12790), .B(n13690), .ZN(
        n12665) );
  OAI22_X1 U14530 ( .A1(n12974), .A2(n13671), .B1(n13392), .B2(n13681), .ZN(
        n12661) );
  AOI211_X1 U14531 ( .C1(n12663), .C2(n13673), .A(n12662), .B(n12661), .ZN(
        n12664) );
  OAI211_X1 U14532 ( .C1(n12743), .C2(n13694), .A(n12665), .B(n12664), .ZN(
        P3_U3153) );
  INV_X1 U14533 ( .A(n12666), .ZN(n12845) );
  OAI222_X1 U14534 ( .A1(n14792), .A2(n8795), .B1(n14775), .B2(n12845), .C1(
        n10329), .C2(P2_U3088), .ZN(P2_U3307) );
  MUX2_X1 U14535 ( .A(n12667), .B(P3_REG2_REG_5__SCAN_IN), .S(n14100), .Z(
        n12668) );
  INV_X1 U14536 ( .A(n12668), .ZN(n12672) );
  AOI22_X1 U14537 ( .A1(n14095), .A2(n12670), .B1(n16337), .B2(n12669), .ZN(
        n12671) );
  OAI211_X1 U14538 ( .C1(n12673), .C2(n14080), .A(n12672), .B(n12671), .ZN(
        P3_U3228) );
  MUX2_X1 U14539 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13791), .Z(n13761) );
  XNOR2_X1 U14540 ( .A(n13761), .B(n13762), .ZN(n13759) );
  NAND2_X1 U14541 ( .A1(n12675), .A2(n12674), .ZN(n12679) );
  INV_X1 U14542 ( .A(n12676), .ZN(n12677) );
  NAND2_X1 U14543 ( .A1(n12677), .A2(n12688), .ZN(n12678) );
  NAND2_X1 U14544 ( .A1(n12679), .A2(n12678), .ZN(n13760) );
  XOR2_X1 U14545 ( .A(n13759), .B(n13760), .Z(n12700) );
  NAND2_X1 U14546 ( .A1(n12681), .A2(n12680), .ZN(n12683) );
  NAND2_X1 U14547 ( .A1(n12683), .A2(n12682), .ZN(n12686) );
  INV_X1 U14548 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12684) );
  MUX2_X1 U14549 ( .A(n12684), .B(P3_REG1_REG_10__SCAN_IN), .S(n13762), .Z(
        n12685) );
  NAND2_X1 U14550 ( .A1(n12686), .A2(n12685), .ZN(n13738) );
  OAI21_X1 U14551 ( .B1(n12686), .B2(n12685), .A(n13738), .ZN(n12698) );
  INV_X1 U14552 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n12687) );
  NOR2_X1 U14553 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12687), .ZN(n12900) );
  NOR2_X1 U14554 ( .A1(n12688), .A2(n7505), .ZN(n12690) );
  INV_X1 U14555 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12691) );
  MUX2_X1 U14556 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n12691), .S(n13762), .Z(
        n12692) );
  NOR2_X1 U14557 ( .A1(n12693), .A2(n12692), .ZN(n13716) );
  AOI21_X1 U14558 ( .B1(n12693), .B2(n12692), .A(n13716), .ZN(n12694) );
  NOR2_X1 U14559 ( .A1(n16250), .A2(n12694), .ZN(n12695) );
  AOI211_X1 U14560 ( .C1(n16252), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n12900), 
        .B(n12695), .ZN(n12696) );
  OAI21_X1 U14561 ( .B1(n13717), .B2(n16244), .A(n12696), .ZN(n12697) );
  AOI21_X1 U14562 ( .B1(n12698), .B2(n16262), .A(n12697), .ZN(n12699) );
  OAI21_X1 U14563 ( .B1(n12700), .B2(n16190), .A(n12699), .ZN(P3_U3192) );
  XNOR2_X1 U14564 ( .A(n12701), .B(n12705), .ZN(n12704) );
  AOI22_X1 U14565 ( .A1(n14376), .A2(n14575), .B1(n12702), .B2(n14578), .ZN(
        n12877) );
  INV_X1 U14566 ( .A(n12877), .ZN(n12703) );
  AOI21_X1 U14567 ( .B1(n12704), .B2(n16584), .A(n12703), .ZN(n12802) );
  NAND2_X1 U14568 ( .A1(n12706), .A2(n12705), .ZN(n12707) );
  NAND2_X1 U14569 ( .A1(n12708), .A2(n12707), .ZN(n12803) );
  NAND2_X1 U14570 ( .A1(n16598), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12709) );
  OAI21_X1 U14571 ( .B1(n14640), .B2(n12875), .A(n12709), .ZN(n12710) );
  AOI21_X1 U14572 ( .B1(n12863), .B2(n16599), .A(n12710), .ZN(n12714) );
  AOI21_X1 U14573 ( .B1(n12863), .B2(n12711), .A(n11533), .ZN(n12712) );
  AND2_X1 U14574 ( .A1(n16575), .A2(n12712), .ZN(n12800) );
  NAND2_X1 U14575 ( .A1(n12800), .A2(n14645), .ZN(n12713) );
  OAI211_X1 U14576 ( .C1(n12803), .C2(n14648), .A(n12714), .B(n12713), .ZN(
        n12715) );
  INV_X1 U14577 ( .A(n12715), .ZN(n12716) );
  OAI21_X1 U14578 ( .B1(n12802), .B2(n16598), .A(n12716), .ZN(P2_U3252) );
  NAND2_X1 U14579 ( .A1(n12718), .A2(n12717), .ZN(n12720) );
  NAND2_X1 U14580 ( .A1(n12720), .A2(n12719), .ZN(n15875) );
  INV_X1 U14581 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12721) );
  XNOR2_X1 U14582 ( .A(n15874), .B(n12721), .ZN(n15876) );
  NAND2_X1 U14583 ( .A1(n15875), .A2(n15876), .ZN(n12723) );
  NAND2_X1 U14584 ( .A1(n15874), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12722) );
  NAND2_X1 U14585 ( .A1(n12723), .A2(n12722), .ZN(n13108) );
  XNOR2_X1 U14586 ( .A(n13105), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13107) );
  XNOR2_X1 U14587 ( .A(n13108), .B(n13107), .ZN(n12737) );
  NOR2_X1 U14588 ( .A1(n12725), .A2(n12724), .ZN(n12727) );
  NAND2_X1 U14589 ( .A1(n15874), .A2(n12729), .ZN(n12728) );
  OAI21_X1 U14590 ( .B1(n15874), .B2(n12729), .A(n12728), .ZN(n15869) );
  NAND2_X1 U14591 ( .A1(n15870), .A2(n15869), .ZN(n15868) );
  OAI21_X1 U14592 ( .B1(n12730), .B2(n12729), .A(n15868), .ZN(n12732) );
  MUX2_X1 U14593 ( .A(n13100), .B(P2_REG2_REG_17__SCAN_IN), .S(n13105), .Z(
        n12731) );
  NAND2_X1 U14594 ( .A1(n12732), .A2(n12731), .ZN(n13099) );
  OAI211_X1 U14595 ( .C1(n12732), .C2(n12731), .A(n13099), .B(n15924), .ZN(
        n12736) );
  INV_X1 U14596 ( .A(n13105), .ZN(n12734) );
  NAND2_X1 U14597 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13189)
         );
  OAI21_X1 U14598 ( .B1(n15928), .B2(n7687), .A(n13189), .ZN(n12733) );
  AOI21_X1 U14599 ( .B1(n12734), .B2(n15922), .A(n12733), .ZN(n12735) );
  OAI211_X1 U14600 ( .C1(n12737), .C2(n15903), .A(n12736), .B(n12735), .ZN(
        P2_U3231) );
  XNOR2_X1 U14601 ( .A(n12738), .B(n13514), .ZN(n16432) );
  OAI211_X1 U14602 ( .C1(n12740), .C2(n13514), .A(n12739), .B(n13979), .ZN(
        n12742) );
  AOI22_X1 U14603 ( .A1(n13986), .A2(n13707), .B1(n13709), .B2(n13987), .ZN(
        n12741) );
  NAND2_X1 U14604 ( .A1(n12742), .A2(n12741), .ZN(n16435) );
  NAND2_X1 U14605 ( .A1(n16435), .A2(n16340), .ZN(n12748) );
  OAI22_X1 U14606 ( .A1(n14046), .A2(n16430), .B1(n12743), .B2(n14073), .ZN(
        n12746) );
  NOR2_X1 U14607 ( .A1(n16340), .A2(n12744), .ZN(n12745) );
  NOR2_X1 U14608 ( .A1(n12746), .A2(n12745), .ZN(n12747) );
  OAI211_X1 U14609 ( .C1(n16432), .C2(n13892), .A(n12748), .B(n12747), .ZN(
        P3_U3226) );
  XNOR2_X1 U14610 ( .A(n15044), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15051) );
  INV_X1 U14611 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12752) );
  AOI21_X1 U14612 ( .B1(n12751), .B2(n12750), .A(n12749), .ZN(n15040) );
  XOR2_X1 U14613 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15037), .Z(n15039) );
  NAND2_X1 U14614 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  OAI21_X1 U14615 ( .B1(n12762), .B2(n12752), .A(n15038), .ZN(n15050) );
  NAND2_X1 U14616 ( .A1(n15051), .A2(n15050), .ZN(n15049) );
  OAI21_X1 U14617 ( .B1(n15044), .B2(n12753), .A(n15049), .ZN(n13014) );
  XOR2_X1 U14618 ( .A(n13019), .B(n13014), .Z(n12754) );
  NAND2_X1 U14619 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n12754), .ZN(n13016) );
  OAI21_X1 U14620 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n12754), .A(n13016), 
        .ZN(n12769) );
  INV_X1 U14621 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n16083) );
  NAND2_X1 U14622 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14887)
         );
  OAI21_X1 U14623 ( .B1(n15046), .B2(n16083), .A(n14887), .ZN(n12767) );
  NOR2_X1 U14624 ( .A1(n15044), .A2(n12755), .ZN(n12756) );
  AOI21_X1 U14625 ( .B1(n12755), .B2(n15044), .A(n12756), .ZN(n15054) );
  INV_X1 U14626 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12761) );
  NOR2_X1 U14627 ( .A1(n12758), .A2(n12757), .ZN(n12760) );
  NOR2_X1 U14628 ( .A1(n12760), .A2(n12759), .ZN(n15033) );
  XOR2_X1 U14629 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n15037), .Z(n15032) );
  NAND2_X1 U14630 ( .A1(n15033), .A2(n15032), .ZN(n15031) );
  OAI21_X1 U14631 ( .B1(n12762), .B2(n12761), .A(n15031), .ZN(n15053) );
  NAND2_X1 U14632 ( .A1(n15054), .A2(n15053), .ZN(n15052) );
  OAI21_X1 U14633 ( .B1(n15044), .B2(n12755), .A(n15052), .ZN(n13018) );
  XNOR2_X1 U14634 ( .A(n12763), .B(n13018), .ZN(n12764) );
  NAND2_X1 U14635 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n12764), .ZN(n13021) );
  OAI21_X1 U14636 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n12764), .A(n13021), 
        .ZN(n12765) );
  NOR2_X1 U14637 ( .A1(n12765), .A2(n13028), .ZN(n12766) );
  AOI211_X1 U14638 ( .C1(n16285), .C2(n13019), .A(n12767), .B(n12766), .ZN(
        n12768) );
  OAI21_X1 U14639 ( .B1(n12769), .B2(n13030), .A(n12768), .ZN(P1_U3261) );
  XNOR2_X1 U14640 ( .A(n12770), .B(n14244), .ZN(n12773) );
  OR2_X1 U14641 ( .A1(n12772), .A2(n12771), .ZN(n12774) );
  NAND2_X1 U14642 ( .A1(n12773), .A2(n12774), .ZN(n12870) );
  INV_X1 U14643 ( .A(n12773), .ZN(n12776) );
  INV_X1 U14644 ( .A(n12774), .ZN(n12775) );
  NAND2_X1 U14645 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  AND2_X1 U14646 ( .A1(n12870), .A2(n12777), .ZN(n12781) );
  OAI21_X1 U14647 ( .B1(n12781), .B2(n12780), .A(n12871), .ZN(n12782) );
  NAND2_X1 U14648 ( .A1(n12782), .A2(n14352), .ZN(n12788) );
  NAND2_X1 U14649 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15909)
         );
  INV_X1 U14650 ( .A(n15909), .ZN(n12786) );
  OAI22_X1 U14651 ( .A1(n14281), .A2(n12784), .B1(n14355), .B2(n12783), .ZN(
        n12785) );
  AOI211_X1 U14652 ( .C1(n14331), .C2(n14377), .A(n12786), .B(n12785), .ZN(
        n12787) );
  OAI211_X1 U14653 ( .C1(n16510), .C2(n14362), .A(n12788), .B(n12787), .ZN(
        P2_U3196) );
  INV_X1 U14654 ( .A(n12990), .ZN(n12799) );
  NAND2_X1 U14655 ( .A1(n12790), .A2(n12789), .ZN(n12794) );
  AND2_X1 U14656 ( .A1(n12821), .A2(n12791), .ZN(n12792) );
  OAI211_X1 U14657 ( .C1(n12794), .C2(n12793), .A(n12792), .B(n13690), .ZN(
        n12798) );
  OAI22_X1 U14658 ( .A1(n13075), .A2(n13671), .B1(n12988), .B2(n13681), .ZN(
        n12795) );
  AOI211_X1 U14659 ( .C1(n12991), .C2(n13673), .A(n12796), .B(n12795), .ZN(
        n12797) );
  OAI211_X1 U14660 ( .C1(n12799), .C2(n13694), .A(n12798), .B(n12797), .ZN(
        P3_U3161) );
  AOI21_X1 U14661 ( .B1(n16418), .B2(n12863), .A(n12800), .ZN(n12801) );
  OAI211_X1 U14662 ( .C1(n14723), .C2(n12803), .A(n12802), .B(n12801), .ZN(
        n12811) );
  NAND2_X1 U14663 ( .A1(n12811), .A2(n16591), .ZN(n12804) );
  OAI21_X1 U14664 ( .B1(n16591), .B2(n12805), .A(n12804), .ZN(P2_U3512) );
  INV_X1 U14665 ( .A(n12806), .ZN(n12809) );
  OAI222_X1 U14666 ( .A1(n14792), .A2(n12807), .B1(n14775), .B2(n12809), .C1(
        P2_U3088), .C2(n10331), .ZN(P2_U3306) );
  OAI222_X1 U14667 ( .A1(n15810), .A2(n12810), .B1(n15805), .B2(n12809), .C1(
        n12808), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U14668 ( .A1(n12811), .A2(n16595), .ZN(n12812) );
  OAI21_X1 U14669 ( .B1(n16595), .B2(n10141), .A(n12812), .ZN(P2_U3469) );
  OAI211_X1 U14670 ( .C1(n7945), .C2(n16624), .A(n12814), .B(n13145), .ZN(
        n12817) );
  AND3_X1 U14671 ( .A1(n12551), .A2(n16631), .A3(n12815), .ZN(n12816) );
  AOI211_X1 U14672 ( .C1(n16568), .C2(n12818), .A(n12817), .B(n12816), .ZN(
        n12860) );
  NAND2_X1 U14673 ( .A1(n16633), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n12819) );
  OAI21_X1 U14674 ( .B1(n12860), .B2(n16633), .A(n12819), .ZN(P1_U3540) );
  NAND2_X1 U14675 ( .A1(n12821), .A2(n12820), .ZN(n12824) );
  INV_X1 U14676 ( .A(n12822), .ZN(n12823) );
  AOI21_X1 U14677 ( .B1(n12825), .B2(n12824), .A(n12823), .ZN(n12831) );
  OAI22_X1 U14678 ( .A1(n12974), .A2(n13681), .B1(n14086), .B2(n13671), .ZN(
        n12826) );
  AOI211_X1 U14679 ( .C1(n12828), .C2(n13673), .A(n12827), .B(n12826), .ZN(
        n12830) );
  NAND2_X1 U14680 ( .A1(n13683), .A2(n12978), .ZN(n12829) );
  OAI211_X1 U14681 ( .C1(n12831), .C2(n13675), .A(n12830), .B(n12829), .ZN(
        P3_U3171) );
  OAI21_X1 U14682 ( .B1(n12833), .B2(n8236), .A(n12832), .ZN(n16528) );
  INV_X1 U14683 ( .A(n16528), .ZN(n12844) );
  OAI21_X1 U14684 ( .B1(n12834), .B2(n12836), .A(n12835), .ZN(n16531) );
  XNOR2_X1 U14685 ( .A(n12837), .B(n13176), .ZN(n12838) );
  NAND2_X1 U14686 ( .A1(n12838), .A2(n16622), .ZN(n16526) );
  AOI22_X1 U14687 ( .A1(n15233), .A2(n14932), .B1(n15234), .B2(n14930), .ZN(
        n16525) );
  OAI22_X1 U14688 ( .A1(n16398), .A2(n16525), .B1(n13171), .B2(n16653), .ZN(
        n12840) );
  NOR2_X1 U14689 ( .A1(n16527), .A2(n16493), .ZN(n12839) );
  AOI211_X1 U14690 ( .C1(n16398), .C2(P1_REG2_REG_13__SCAN_IN), .A(n12840), 
        .B(n12839), .ZN(n12841) );
  OAI21_X1 U14691 ( .B1(n16644), .B2(n16526), .A(n12841), .ZN(n12842) );
  AOI21_X1 U14692 ( .B1(n16531), .B2(n12966), .A(n12842), .ZN(n12843) );
  OAI21_X1 U14693 ( .B1(n12844), .B2(n16646), .A(n12843), .ZN(P1_U3280) );
  OAI222_X1 U14694 ( .A1(n15810), .A2(n8092), .B1(P1_U3086), .B2(n7436), .C1(
        n15805), .C2(n12845), .ZN(P1_U3335) );
  XNOR2_X1 U14695 ( .A(n12847), .B(n13516), .ZN(n12852) );
  INV_X1 U14696 ( .A(n12852), .ZN(n16407) );
  OAI211_X1 U14697 ( .C1(n7578), .C2(n12849), .A(n12848), .B(n13979), .ZN(
        n12855) );
  OAI22_X1 U14698 ( .A1(n12850), .A2(n14087), .B1(n12988), .B2(n14089), .ZN(
        n12851) );
  INV_X1 U14699 ( .A(n12851), .ZN(n12854) );
  NAND2_X1 U14700 ( .A1(n12852), .A2(n16428), .ZN(n12853) );
  NAND3_X1 U14701 ( .A1(n12855), .A2(n12854), .A3(n12853), .ZN(n16409) );
  MUX2_X1 U14702 ( .A(n16409), .B(P3_REG2_REG_6__SCAN_IN), .S(n14100), .Z(
        n12856) );
  INV_X1 U14703 ( .A(n12856), .ZN(n12859) );
  AOI22_X1 U14704 ( .A1(n14095), .A2(n13391), .B1(n16337), .B2(n12857), .ZN(
        n12858) );
  OAI211_X1 U14705 ( .C1(n16407), .C2(n14080), .A(n12859), .B(n12858), .ZN(
        P3_U3227) );
  INV_X1 U14706 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12862) );
  OR2_X1 U14707 ( .A1(n12860), .A2(n16636), .ZN(n12861) );
  OAI21_X1 U14708 ( .B1(n16638), .B2(n12862), .A(n12861), .ZN(P1_U3495) );
  XNOR2_X1 U14709 ( .A(n12863), .B(n14244), .ZN(n12865) );
  OR2_X1 U14710 ( .A1(n12864), .A2(n12771), .ZN(n12866) );
  NAND2_X1 U14711 ( .A1(n12865), .A2(n12866), .ZN(n12937) );
  INV_X1 U14712 ( .A(n12865), .ZN(n12868) );
  INV_X1 U14713 ( .A(n12866), .ZN(n12867) );
  NAND2_X1 U14714 ( .A1(n12868), .A2(n12867), .ZN(n12869) );
  AND2_X1 U14715 ( .A1(n12937), .A2(n12869), .ZN(n12873) );
  NAND2_X1 U14716 ( .A1(n12872), .A2(n12873), .ZN(n12938) );
  OAI21_X1 U14717 ( .B1(n12873), .B2(n12872), .A(n12938), .ZN(n12874) );
  NAND2_X1 U14718 ( .A1(n12874), .A2(n14352), .ZN(n12881) );
  INV_X1 U14719 ( .A(n12875), .ZN(n12879) );
  OAI22_X1 U14720 ( .A1(n14297), .A2(n12877), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12876), .ZN(n12878) );
  AOI21_X1 U14721 ( .B1(n12879), .B2(n14332), .A(n12878), .ZN(n12880) );
  OAI211_X1 U14722 ( .C1(n12882), .C2(n14362), .A(n12881), .B(n12880), .ZN(
        P2_U3206) );
  XOR2_X1 U14723 ( .A(n12883), .B(n12884), .Z(n12893) );
  OAI21_X1 U14724 ( .B1(n16558), .B2(n12886), .A(n12885), .ZN(n12890) );
  OAI22_X1 U14725 ( .A1(n12888), .A2(n16543), .B1(n16542), .B2(n12887), .ZN(
        n12889) );
  AOI211_X1 U14726 ( .C1(n12891), .C2(n16554), .A(n12890), .B(n12889), .ZN(
        n12892) );
  OAI21_X1 U14727 ( .B1(n12893), .B2(n16549), .A(n12892), .ZN(P1_U3231) );
  INV_X1 U14728 ( .A(n12894), .ZN(n13079) );
  AOI21_X1 U14729 ( .B1(n12896), .B2(n12895), .A(n13675), .ZN(n12898) );
  NAND2_X1 U14730 ( .A1(n12898), .A2(n12897), .ZN(n12903) );
  OAI22_X1 U14731 ( .A1(n13075), .A2(n13681), .B1(n8630), .B2(n13671), .ZN(
        n12899) );
  AOI211_X1 U14732 ( .C1(n12901), .C2(n13673), .A(n12900), .B(n12899), .ZN(
        n12902) );
  OAI211_X1 U14733 ( .C1(n13079), .C2(n13694), .A(n12903), .B(n12902), .ZN(
        P3_U3157) );
  INV_X1 U14734 ( .A(n12904), .ZN(n12906) );
  OAI222_X1 U14735 ( .A1(n12907), .A2(P3_U3151), .B1(n14221), .B2(n12906), 
        .C1(n12905), .C2(n14223), .ZN(P3_U3271) );
  XNOR2_X1 U14736 ( .A(n12909), .B(n12908), .ZN(n12910) );
  AOI22_X1 U14737 ( .A1(n14578), .A2(n14376), .B1(n14374), .B2(n14575), .ZN(
        n13062) );
  OAI21_X1 U14738 ( .B1(n12910), .B2(n14510), .A(n13062), .ZN(n13005) );
  INV_X1 U14739 ( .A(n13005), .ZN(n12918) );
  OAI21_X1 U14740 ( .B1(n12913), .B2(n12912), .A(n12911), .ZN(n13007) );
  OAI211_X1 U14741 ( .C1(n13067), .C2(n16578), .A(n12771), .B(n13093), .ZN(
        n13004) );
  AOI22_X1 U14742 ( .A1(n16598), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13064), 
        .B2(n16596), .ZN(n12915) );
  NAND2_X1 U14743 ( .A1(n13050), .A2(n16599), .ZN(n12914) );
  OAI211_X1 U14744 ( .C1(n13004), .C2(n16601), .A(n12915), .B(n12914), .ZN(
        n12916) );
  AOI21_X1 U14745 ( .B1(n13007), .B2(n16604), .A(n12916), .ZN(n12917) );
  OAI21_X1 U14746 ( .B1(n12918), .B2(n16598), .A(n12917), .ZN(P2_U3250) );
  NOR2_X1 U14747 ( .A1(n12920), .A2(n7571), .ZN(n12921) );
  XNOR2_X1 U14748 ( .A(n12919), .B(n12921), .ZN(n12930) );
  OAI21_X1 U14749 ( .B1(n16558), .B2(n12923), .A(n12922), .ZN(n12927) );
  OAI22_X1 U14750 ( .A1(n12925), .A2(n16543), .B1(n16542), .B2(n12924), .ZN(
        n12926) );
  AOI211_X1 U14751 ( .C1(n12928), .C2(n16554), .A(n12927), .B(n12926), .ZN(
        n12929) );
  OAI21_X1 U14752 ( .B1(n12930), .B2(n16549), .A(n12929), .ZN(P1_U3217) );
  XNOR2_X1 U14753 ( .A(n16600), .B(n14244), .ZN(n12932) );
  OR2_X1 U14754 ( .A1(n12931), .A2(n12771), .ZN(n12933) );
  NAND2_X1 U14755 ( .A1(n12932), .A2(n12933), .ZN(n13056) );
  INV_X1 U14756 ( .A(n12932), .ZN(n12935) );
  INV_X1 U14757 ( .A(n12933), .ZN(n12934) );
  NAND2_X1 U14758 ( .A1(n12935), .A2(n12934), .ZN(n12936) );
  AND2_X1 U14759 ( .A1(n13056), .A2(n12936), .ZN(n12940) );
  NAND2_X1 U14760 ( .A1(n12938), .A2(n12937), .ZN(n12939) );
  NAND2_X1 U14761 ( .A1(n12939), .A2(n12940), .ZN(n13057) );
  OAI21_X1 U14762 ( .B1(n12940), .B2(n12939), .A(n13057), .ZN(n12941) );
  NAND2_X1 U14763 ( .A1(n12941), .A2(n14352), .ZN(n12945) );
  AOI22_X1 U14764 ( .A1(n14375), .A2(n14575), .B1(n14377), .B2(n14578), .ZN(
        n16582) );
  OAI22_X1 U14765 ( .A1(n14297), .A2(n16582), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12942), .ZN(n12943) );
  AOI21_X1 U14766 ( .B1(n16597), .B2(n14332), .A(n12943), .ZN(n12944) );
  OAI211_X1 U14767 ( .C1(n7846), .C2(n14362), .A(n12945), .B(n12944), .ZN(
        P2_U3187) );
  NAND2_X1 U14768 ( .A1(n12946), .A2(n12947), .ZN(n13553) );
  OAI211_X1 U14769 ( .C1(n12946), .C2(n12947), .A(n13553), .B(n13690), .ZN(
        n12953) );
  INV_X1 U14770 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12948) );
  NOR2_X1 U14771 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12948), .ZN(n16138) );
  AOI21_X1 U14772 ( .B1(n13697), .B2(n13656), .A(n16138), .ZN(n12950) );
  NAND2_X1 U14773 ( .A1(n14094), .A2(n13673), .ZN(n12949) );
  OAI211_X1 U14774 ( .C1(n14086), .C2(n13681), .A(n12950), .B(n12949), .ZN(
        n12951) );
  AOI21_X1 U14775 ( .B1(n14093), .B2(n13683), .A(n12951), .ZN(n12952) );
  NAND2_X1 U14776 ( .A1(n12953), .A2(n12952), .ZN(P3_U3176) );
  INV_X1 U14777 ( .A(n12954), .ZN(n12955) );
  AOI21_X1 U14778 ( .B1(n12963), .B2(n12956), .A(n12955), .ZN(n16569) );
  AND2_X1 U14779 ( .A1(n16561), .A2(n12957), .ZN(n12958) );
  OR2_X1 U14780 ( .A1(n16623), .A2(n12958), .ZN(n16565) );
  NAND2_X1 U14781 ( .A1(n16498), .A2(n16622), .ZN(n13122) );
  NAND2_X1 U14782 ( .A1(n15234), .A2(n14929), .ZN(n12959) );
  OAI21_X1 U14783 ( .B1(n16544), .B2(n15216), .A(n12959), .ZN(n16559) );
  NAND2_X1 U14784 ( .A1(n7416), .A2(n16559), .ZN(n12961) );
  OR2_X1 U14785 ( .A1(n16653), .A2(n16557), .ZN(n12960) );
  OAI211_X1 U14786 ( .C1(n7416), .C2(n11621), .A(n12961), .B(n12960), .ZN(
        n12962) );
  AOI21_X1 U14787 ( .B1(n16561), .B2(n16389), .A(n12962), .ZN(n12968) );
  OR2_X1 U14788 ( .A1(n12964), .A2(n12963), .ZN(n16562) );
  NAND3_X1 U14789 ( .A1(n16562), .A2(n12966), .A3(n12965), .ZN(n12967) );
  OAI211_X1 U14790 ( .C1(n16565), .C2(n13122), .A(n12968), .B(n12967), .ZN(
        n12969) );
  AOI21_X1 U14791 ( .B1(n16394), .B2(n16569), .A(n12969), .ZN(n12970) );
  INV_X1 U14792 ( .A(n12970), .ZN(P1_U3279) );
  INV_X1 U14793 ( .A(n12971), .ZN(n13410) );
  OR2_X1 U14794 ( .A1(n13410), .A2(n13409), .ZN(n13513) );
  INV_X1 U14795 ( .A(n13513), .ZN(n13407) );
  XNOR2_X1 U14796 ( .A(n12972), .B(n13407), .ZN(n16465) );
  INV_X1 U14797 ( .A(n16465), .ZN(n12983) );
  XNOR2_X1 U14798 ( .A(n12973), .B(n13407), .ZN(n12977) );
  OAI22_X1 U14799 ( .A1(n12974), .A2(n14087), .B1(n14086), .B2(n14089), .ZN(
        n12975) );
  AOI21_X1 U14800 ( .B1(n16465), .B2(n16428), .A(n12975), .ZN(n12976) );
  OAI21_X1 U14801 ( .B1(n12977), .B2(n14084), .A(n12976), .ZN(n16463) );
  NAND2_X1 U14802 ( .A1(n16463), .A2(n16340), .ZN(n12982) );
  INV_X1 U14803 ( .A(n12978), .ZN(n12979) );
  OAI22_X1 U14804 ( .A1(n14046), .A2(n16462), .B1(n12979), .B2(n14073), .ZN(
        n12980) );
  AOI21_X1 U14805 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n14100), .A(n12980), .ZN(
        n12981) );
  OAI211_X1 U14806 ( .C1(n12983), .C2(n14080), .A(n12982), .B(n12981), .ZN(
        P3_U3224) );
  INV_X1 U14807 ( .A(n12984), .ZN(n12985) );
  AOI21_X1 U14808 ( .B1(n13517), .B2(n12986), .A(n12985), .ZN(n12987) );
  OAI222_X1 U14809 ( .A1(n14089), .A2(n13075), .B1(n14087), .B2(n12988), .C1(
        n14084), .C2(n12987), .ZN(n16440) );
  INV_X1 U14810 ( .A(n16440), .ZN(n12996) );
  XNOR2_X1 U14811 ( .A(n12989), .B(n13517), .ZN(n16442) );
  INV_X1 U14812 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U14813 ( .A1(n14095), .A2(n12991), .B1(n16337), .B2(n12990), .ZN(
        n12992) );
  OAI21_X1 U14814 ( .B1(n12993), .B2(n16340), .A(n12992), .ZN(n12994) );
  AOI21_X1 U14815 ( .B1(n16442), .B2(n14098), .A(n12994), .ZN(n12995) );
  OAI21_X1 U14816 ( .B1(n12996), .B2(n14100), .A(n12995), .ZN(P3_U3225) );
  INV_X1 U14817 ( .A(n13000), .ZN(n12999) );
  INV_X1 U14818 ( .A(n15810), .ZN(n15802) );
  NAND2_X1 U14819 ( .A1(n15802), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12997) );
  OAI211_X1 U14820 ( .C1(n12999), .C2(n15805), .A(n12998), .B(n12997), .ZN(
        P1_U3332) );
  NAND2_X1 U14821 ( .A1(n13000), .A2(n14779), .ZN(n13002) );
  OAI211_X1 U14822 ( .C1(n13003), .C2(n14792), .A(n13002), .B(n13001), .ZN(
        P2_U3304) );
  INV_X1 U14823 ( .A(n16418), .ZN(n16579) );
  OAI21_X1 U14824 ( .B1(n13067), .B2(n16579), .A(n13004), .ZN(n13006) );
  AOI211_X1 U14825 ( .C1(n16588), .C2(n13007), .A(n13006), .B(n13005), .ZN(
        n13010) );
  NAND2_X1 U14826 ( .A1(n16592), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n13008) );
  OAI21_X1 U14827 ( .B1(n13010), .B2(n16592), .A(n13008), .ZN(P2_U3475) );
  NAND2_X1 U14828 ( .A1(n16589), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n13009) );
  OAI21_X1 U14829 ( .B1(n13010), .B2(n16589), .A(n13009), .ZN(P2_U3514) );
  INV_X1 U14830 ( .A(n13011), .ZN(n13012) );
  OAI222_X1 U14831 ( .A1(n13013), .A2(P3_U3151), .B1(n14221), .B2(n13012), 
        .C1(n15466), .C2(n14223), .ZN(P3_U3270) );
  NAND2_X1 U14832 ( .A1(n13019), .A2(n13014), .ZN(n13015) );
  NAND2_X1 U14833 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  XNOR2_X1 U14834 ( .A(n13017), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13031) );
  INV_X1 U14835 ( .A(n13031), .ZN(n13027) );
  NAND2_X1 U14836 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  NAND2_X1 U14837 ( .A1(n13021), .A2(n13020), .ZN(n13022) );
  XNOR2_X1 U14838 ( .A(n13022), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n13029) );
  NAND3_X1 U14839 ( .A1(n13029), .A2(n13024), .A3(n13023), .ZN(n13025) );
  OAI211_X1 U14840 ( .C1(n13027), .C2(n13030), .A(n13026), .B(n13025), .ZN(
        n13034) );
  OAI22_X1 U14841 ( .A1(n13031), .A2(n13030), .B1(n13029), .B2(n13028), .ZN(
        n13033) );
  MUX2_X1 U14842 ( .A(n13034), .B(n13033), .S(n13032), .Z(n13035) );
  INV_X1 U14843 ( .A(n13035), .ZN(n13036) );
  NAND2_X1 U14844 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14821)
         );
  OAI211_X1 U14845 ( .C1(n16084), .C2(n15046), .A(n13036), .B(n14821), .ZN(
        P1_U3262) );
  INV_X1 U14846 ( .A(n13037), .ZN(n13038) );
  OAI21_X1 U14847 ( .B1(n13042), .B2(n13040), .A(n13041), .ZN(n13043) );
  NAND2_X1 U14848 ( .A1(n13043), .A2(n14905), .ZN(n13049) );
  INV_X1 U14849 ( .A(n13044), .ZN(n16491) );
  INV_X1 U14850 ( .A(n14899), .ZN(n14912) );
  OAI21_X1 U14851 ( .B1(n14912), .B2(n13046), .A(n13045), .ZN(n13047) );
  AOI21_X1 U14852 ( .B1(n16491), .B2(n14914), .A(n13047), .ZN(n13048) );
  OAI211_X1 U14853 ( .C1(n16494), .C2(n14918), .A(n13049), .B(n13048), .ZN(
        P1_U3236) );
  XNOR2_X1 U14854 ( .A(n13050), .B(n14244), .ZN(n13051) );
  NAND2_X1 U14855 ( .A1(n14375), .A2(n11533), .ZN(n13052) );
  NAND2_X1 U14856 ( .A1(n13051), .A2(n13052), .ZN(n13155) );
  INV_X1 U14857 ( .A(n13051), .ZN(n13054) );
  INV_X1 U14858 ( .A(n13052), .ZN(n13053) );
  NAND2_X1 U14859 ( .A1(n13054), .A2(n13053), .ZN(n13055) );
  AND2_X1 U14860 ( .A1(n13155), .A2(n13055), .ZN(n13059) );
  NAND2_X1 U14861 ( .A1(n13057), .A2(n13056), .ZN(n13058) );
  OAI21_X1 U14862 ( .B1(n13059), .B2(n13058), .A(n13156), .ZN(n13060) );
  NAND2_X1 U14863 ( .A1(n13060), .A2(n14352), .ZN(n13066) );
  OAI21_X1 U14864 ( .B1(n14297), .B2(n13062), .A(n13061), .ZN(n13063) );
  AOI21_X1 U14865 ( .B1(n13064), .B2(n14332), .A(n13063), .ZN(n13065) );
  OAI211_X1 U14866 ( .C1(n13067), .C2(n14362), .A(n13066), .B(n13065), .ZN(
        P2_U3213) );
  OAI222_X1 U14867 ( .A1(P3_U3151), .A2(n13070), .B1(n14223), .B2(n13069), 
        .C1(n14221), .C2(n13068), .ZN(P3_U3269) );
  NAND2_X1 U14868 ( .A1(n13071), .A2(n13403), .ZN(n13072) );
  NAND2_X1 U14869 ( .A1(n13073), .A2(n13072), .ZN(n16472) );
  INV_X1 U14870 ( .A(n16472), .ZN(n13083) );
  XNOR2_X1 U14871 ( .A(n13074), .B(n13403), .ZN(n13078) );
  OAI22_X1 U14872 ( .A1(n13075), .A2(n14087), .B1(n8630), .B2(n14089), .ZN(
        n13076) );
  AOI21_X1 U14873 ( .B1(n16472), .B2(n16428), .A(n13076), .ZN(n13077) );
  OAI21_X1 U14874 ( .B1(n13078), .B2(n14084), .A(n13077), .ZN(n16470) );
  NAND2_X1 U14875 ( .A1(n16470), .A2(n16340), .ZN(n13082) );
  OAI22_X1 U14876 ( .A1(n14046), .A2(n16469), .B1(n13079), .B2(n14073), .ZN(
        n13080) );
  AOI21_X1 U14877 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14100), .A(n13080), 
        .ZN(n13081) );
  OAI211_X1 U14878 ( .C1(n13083), .C2(n14080), .A(n13082), .B(n13081), .ZN(
        P3_U3223) );
  OAI211_X1 U14879 ( .C1(n13086), .C2(n13085), .A(n13084), .B(n16584), .ZN(
        n13087) );
  AOI22_X1 U14880 ( .A1(n14373), .A2(n14575), .B1(n14375), .B2(n14578), .ZN(
        n13161) );
  AND2_X1 U14881 ( .A1(n13087), .A2(n13161), .ZN(n14722) );
  OAI21_X1 U14882 ( .B1(n13090), .B2(n13089), .A(n13088), .ZN(n14724) );
  NAND2_X1 U14883 ( .A1(n16598), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13091) );
  OAI21_X1 U14884 ( .B1(n14640), .B2(n13160), .A(n13091), .ZN(n13092) );
  AOI21_X1 U14885 ( .B1(n14720), .B2(n16599), .A(n13092), .ZN(n13096) );
  AOI21_X1 U14886 ( .B1(n13093), .B2(n14720), .A(n11533), .ZN(n13094) );
  AND2_X1 U14887 ( .A1(n13094), .A2(n14642), .ZN(n14719) );
  NAND2_X1 U14888 ( .A1(n14719), .A2(n14645), .ZN(n13095) );
  OAI211_X1 U14889 ( .C1(n14724), .C2(n14648), .A(n13096), .B(n13095), .ZN(
        n13097) );
  INV_X1 U14890 ( .A(n13097), .ZN(n13098) );
  OAI21_X1 U14891 ( .B1(n16598), .B2(n14722), .A(n13098), .ZN(P2_U3249) );
  OAI21_X1 U14892 ( .B1(n13100), .B2(n13105), .A(n13099), .ZN(n13101) );
  XOR2_X1 U14893 ( .A(n15885), .B(n13101), .Z(n15883) );
  NAND2_X1 U14894 ( .A1(n15883), .A2(n15882), .ZN(n15881) );
  OAI21_X1 U14895 ( .B1(n15885), .B2(n13101), .A(n15881), .ZN(n13103) );
  MUX2_X1 U14896 ( .A(n14596), .B(P2_REG2_REG_19__SCAN_IN), .S(n10696), .Z(
        n13102) );
  XNOR2_X1 U14897 ( .A(n13103), .B(n13102), .ZN(n13118) );
  INV_X1 U14898 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13104) );
  NOR2_X1 U14899 ( .A1(n13105), .A2(n13104), .ZN(n13106) );
  AOI21_X1 U14900 ( .B1(n13108), .B2(n13107), .A(n13106), .ZN(n13109) );
  XNOR2_X1 U14901 ( .A(n13109), .B(n15885), .ZN(n15886) );
  INV_X1 U14902 ( .A(n13109), .ZN(n13110) );
  AOI22_X1 U14903 ( .A1(n15886), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n15885), 
        .B2(n13110), .ZN(n13112) );
  INV_X1 U14904 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14706) );
  XNOR2_X1 U14905 ( .A(n10696), .B(n14706), .ZN(n13111) );
  XNOR2_X1 U14906 ( .A(n13112), .B(n13111), .ZN(n13116) );
  NAND2_X1 U14907 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14280)
         );
  NAND2_X1 U14908 ( .A1(n15880), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n13113) );
  OAI211_X1 U14909 ( .C1(n14418), .C2(n13114), .A(n14280), .B(n13113), .ZN(
        n13115) );
  AOI21_X1 U14910 ( .B1(n13116), .B2(n15920), .A(n13115), .ZN(n13117) );
  OAI21_X1 U14911 ( .B1(n13118), .B2(n15897), .A(n13117), .ZN(P2_U3233) );
  AOI21_X1 U14912 ( .B1(n8228), .B2(n13119), .A(n7564), .ZN(n15768) );
  OAI21_X1 U14913 ( .B1(n13121), .B2(n8228), .A(n13120), .ZN(n15766) );
  XNOR2_X1 U14914 ( .A(n16621), .B(n15762), .ZN(n15764) );
  NOR2_X1 U14915 ( .A1(n15764), .A2(n13122), .ZN(n13128) );
  INV_X1 U14916 ( .A(n15762), .ZN(n13126) );
  OAI22_X1 U14917 ( .A1(n14889), .A2(n15218), .B1(n16541), .B2(n15216), .ZN(
        n15761) );
  INV_X1 U14918 ( .A(n14852), .ZN(n13123) );
  AOI22_X1 U14919 ( .A1(n15761), .A2(n7416), .B1(n13123), .B2(n16490), .ZN(
        n13125) );
  NAND2_X1 U14920 ( .A1(n16398), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13124) );
  OAI211_X1 U14921 ( .C1(n13126), .C2(n16493), .A(n13125), .B(n13124), .ZN(
        n13127) );
  AOI211_X1 U14922 ( .C1(n15766), .C2(n16394), .A(n13128), .B(n13127), .ZN(
        n13129) );
  OAI21_X1 U14923 ( .B1(n15768), .B2(n16647), .A(n13129), .ZN(P1_U3277) );
  OAI222_X1 U14924 ( .A1(n14221), .A2(n13130), .B1(n14223), .B2(n15461), .C1(
        P3_U3151), .C2(n13791), .ZN(P3_U3268) );
  XNOR2_X1 U14925 ( .A(n13132), .B(n13625), .ZN(n13133) );
  XNOR2_X1 U14926 ( .A(n13131), .B(n13133), .ZN(n13139) );
  NOR2_X1 U14927 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15562), .ZN(n16205) );
  AOI21_X1 U14928 ( .B1(n13988), .B2(n13697), .A(n16205), .ZN(n13135) );
  NAND2_X1 U14929 ( .A1(n13683), .A2(n14031), .ZN(n13134) );
  OAI211_X1 U14930 ( .C1(n14055), .C2(n13681), .A(n13135), .B(n13134), .ZN(
        n13136) );
  AOI21_X1 U14931 ( .B1(n13137), .B2(n13673), .A(n13136), .ZN(n13138) );
  OAI21_X1 U14932 ( .B1(n13139), .B2(n13675), .A(n13138), .ZN(P3_U3181) );
  OAI21_X1 U14933 ( .B1(n13142), .B2(n13140), .A(n13141), .ZN(n13143) );
  NAND2_X1 U14934 ( .A1(n13143), .A2(n14905), .ZN(n13149) );
  OAI21_X1 U14935 ( .B1(n14912), .B2(n13145), .A(n13144), .ZN(n13146) );
  AOI21_X1 U14936 ( .B1(n13147), .B2(n14914), .A(n13146), .ZN(n13148) );
  OAI211_X1 U14937 ( .C1(n7945), .C2(n14918), .A(n13149), .B(n13148), .ZN(
        P1_U3224) );
  INV_X1 U14938 ( .A(n14720), .ZN(n13166) );
  XNOR2_X1 U14939 ( .A(n14720), .B(n14244), .ZN(n13150) );
  NAND2_X1 U14940 ( .A1(n14374), .A2(n11533), .ZN(n13151) );
  NAND2_X1 U14941 ( .A1(n13150), .A2(n13151), .ZN(n13184) );
  INV_X1 U14942 ( .A(n13150), .ZN(n13153) );
  INV_X1 U14943 ( .A(n13151), .ZN(n13152) );
  NAND2_X1 U14944 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  AND2_X1 U14945 ( .A1(n13184), .A2(n13154), .ZN(n13158) );
  OAI21_X1 U14946 ( .B1(n13158), .B2(n13157), .A(n13185), .ZN(n13159) );
  NAND2_X1 U14947 ( .A1(n13159), .A2(n14352), .ZN(n13165) );
  INV_X1 U14948 ( .A(n13160), .ZN(n13163) );
  OAI22_X1 U14949 ( .A1(n14297), .A2(n13161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15867), .ZN(n13162) );
  AOI21_X1 U14950 ( .B1(n13163), .B2(n14332), .A(n13162), .ZN(n13164) );
  OAI211_X1 U14951 ( .C1(n13166), .C2(n14362), .A(n13165), .B(n13164), .ZN(
        P2_U3198) );
  NAND2_X1 U14952 ( .A1(n16546), .A2(n13168), .ZN(n13169) );
  XNOR2_X1 U14953 ( .A(n13167), .B(n13169), .ZN(n13178) );
  OAI21_X1 U14954 ( .B1(n16558), .B2(n13171), .A(n13170), .ZN(n13175) );
  OAI22_X1 U14955 ( .A1(n13173), .A2(n16543), .B1(n16542), .B2(n13172), .ZN(
        n13174) );
  AOI211_X1 U14956 ( .C1(n13176), .C2(n16554), .A(n13175), .B(n13174), .ZN(
        n13177) );
  OAI21_X1 U14957 ( .B1(n13178), .B2(n16549), .A(n13177), .ZN(P1_U3234) );
  XNOR2_X1 U14958 ( .A(n14716), .B(n14244), .ZN(n13179) );
  NAND2_X1 U14959 ( .A1(n14373), .A2(n11533), .ZN(n13180) );
  NAND2_X1 U14960 ( .A1(n13179), .A2(n13180), .ZN(n13194) );
  INV_X1 U14961 ( .A(n13179), .ZN(n13182) );
  INV_X1 U14962 ( .A(n13180), .ZN(n13181) );
  NAND2_X1 U14963 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  AND2_X1 U14964 ( .A1(n13194), .A2(n13183), .ZN(n13187) );
  NAND2_X1 U14965 ( .A1(n13186), .A2(n13187), .ZN(n13195) );
  OAI21_X1 U14966 ( .B1(n13187), .B2(n13186), .A(n13195), .ZN(n13188) );
  NAND2_X1 U14967 ( .A1(n13188), .A2(n14352), .ZN(n13193) );
  INV_X1 U14968 ( .A(n14639), .ZN(n13191) );
  AOI22_X1 U14969 ( .A1(n14372), .A2(n14575), .B1(n14578), .B2(n14374), .ZN(
        n14633) );
  OAI21_X1 U14970 ( .B1(n14633), .B2(n14297), .A(n13189), .ZN(n13190) );
  AOI21_X1 U14971 ( .B1(n13191), .B2(n14332), .A(n13190), .ZN(n13192) );
  OAI211_X1 U14972 ( .C1(n8300), .C2(n14362), .A(n13193), .B(n13192), .ZN(
        P2_U3200) );
  NAND2_X1 U14973 ( .A1(n14372), .A2(n11533), .ZN(n14226) );
  XNOR2_X1 U14974 ( .A(n14225), .B(n14226), .ZN(n14230) );
  XNOR2_X1 U14975 ( .A(n14231), .B(n14230), .ZN(n13202) );
  INV_X1 U14976 ( .A(n14619), .ZN(n13199) );
  OAI22_X1 U14977 ( .A1(n13197), .A2(n14604), .B1(n13196), .B2(n14602), .ZN(
        n14615) );
  AOI22_X1 U14978 ( .A1(n14615), .A2(n14358), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13198) );
  OAI21_X1 U14979 ( .B1(n13199), .B2(n14355), .A(n13198), .ZN(n13200) );
  AOI21_X1 U14980 ( .B1(n14710), .B2(n14324), .A(n13200), .ZN(n13201) );
  OAI21_X1 U14981 ( .B1(n13202), .B2(n14326), .A(n13201), .ZN(P2_U3210) );
  INV_X1 U14982 ( .A(n13203), .ZN(n13206) );
  OAI222_X1 U14983 ( .A1(n14792), .A2(n8076), .B1(n14775), .B2(n13206), .C1(
        P2_U3088), .C2(n13204), .ZN(P2_U3303) );
  INV_X1 U14984 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13207) );
  OAI222_X1 U14985 ( .A1(n15810), .A2(n13207), .B1(n15805), .B2(n13206), .C1(
        P1_U3086), .C2(n13205), .ZN(P1_U3331) );
  INV_X1 U14986 ( .A(n13208), .ZN(n14777) );
  OAI222_X1 U14987 ( .A1(n15810), .A2(n13337), .B1(P1_U3086), .B2(n13209), 
        .C1(n15805), .C2(n14777), .ZN(P1_U3326) );
  INV_X1 U14988 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13346) );
  OAI222_X1 U14989 ( .A1(n15805), .A2(n13213), .B1(P1_U3086), .B2(n13210), 
        .C1(n13346), .C2(n15810), .ZN(P1_U3325) );
  OAI222_X1 U14990 ( .A1(n14775), .A2(n13213), .B1(P2_U3088), .B2(n13212), 
        .C1(n13211), .C2(n14792), .ZN(P2_U3297) );
  OAI21_X1 U14991 ( .B1(n7473), .B2(n13215), .A(n13214), .ZN(n13216) );
  NAND2_X1 U14992 ( .A1(n15074), .A2(n13216), .ZN(n13220) );
  NAND2_X1 U14993 ( .A1(n14921), .A2(n15234), .ZN(n13218) );
  INV_X1 U14994 ( .A(n15098), .ZN(n13221) );
  AOI211_X1 U14995 ( .C1(n15691), .C2(n13221), .A(n16566), .B(n15082), .ZN(
        n15690) );
  INV_X1 U14996 ( .A(n14799), .ZN(n13222) );
  AOI22_X1 U14997 ( .A1(n16398), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13222), 
        .B2(n16490), .ZN(n13223) );
  OAI21_X1 U14998 ( .B1(n13224), .B2(n16493), .A(n13223), .ZN(n13230) );
  INV_X1 U14999 ( .A(n13225), .ZN(n13229) );
  INV_X1 U15000 ( .A(n13231), .ZN(n13233) );
  AND2_X1 U15001 ( .A1(n13232), .A2(n13233), .ZN(n13235) );
  XNOR2_X1 U15002 ( .A(n13237), .B(n13236), .ZN(n13238) );
  XNOR2_X1 U15003 ( .A(n13239), .B(n13238), .ZN(n13247) );
  INV_X1 U15004 ( .A(n13821), .ZN(n13241) );
  INV_X1 U15005 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13240) );
  OAI22_X1 U15006 ( .A1(n13241), .A2(n13694), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13240), .ZN(n13244) );
  OAI22_X1 U15007 ( .A1(n13242), .A2(n13671), .B1(n13839), .B2(n13681), .ZN(
        n13243) );
  AOI211_X1 U15008 ( .C1(n13245), .C2(n13673), .A(n13244), .B(n13243), .ZN(
        n13246) );
  OAI21_X1 U15009 ( .B1(n13247), .B2(n13675), .A(n13246), .ZN(P3_U3160) );
  OAI222_X1 U15010 ( .A1(n14221), .A2(n13248), .B1(n14223), .B2(n15459), .C1(
        P3_U3151), .C2(n8956), .ZN(P3_U3267) );
  INV_X1 U15011 ( .A(n13249), .ZN(n13250) );
  NAND2_X1 U15012 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  AOI22_X1 U15013 ( .A1(n15729), .A2(n13313), .B1(n13316), .B2(n15194), .ZN(
        n13254) );
  XNOR2_X1 U15014 ( .A(n13254), .B(n10643), .ZN(n13257) );
  AOI22_X1 U15015 ( .A1(n15729), .A2(n13316), .B1(n13315), .B2(n15194), .ZN(
        n13256) );
  XNOR2_X1 U15016 ( .A(n13257), .B(n13256), .ZN(n14829) );
  INV_X1 U15017 ( .A(n14829), .ZN(n13255) );
  NAND2_X1 U15018 ( .A1(n13257), .A2(n13256), .ZN(n13258) );
  NAND2_X1 U15019 ( .A1(n15726), .A2(n13313), .ZN(n13260) );
  NAND2_X1 U15020 ( .A1(n14925), .A2(n13316), .ZN(n13259) );
  NAND2_X1 U15021 ( .A1(n13260), .A2(n13259), .ZN(n13261) );
  XNOR2_X1 U15022 ( .A(n13261), .B(n13305), .ZN(n13264) );
  NOR2_X1 U15023 ( .A1(n14830), .A2(n10968), .ZN(n13262) );
  AOI21_X1 U15024 ( .B1(n15726), .B2(n13316), .A(n13262), .ZN(n13263) );
  OR2_X1 U15025 ( .A1(n13264), .A2(n13263), .ZN(n14879) );
  NAND2_X1 U15026 ( .A1(n13264), .A2(n13263), .ZN(n14878) );
  NAND2_X1 U15027 ( .A1(n15718), .A2(n13313), .ZN(n13267) );
  NAND2_X1 U15028 ( .A1(n14924), .A2(n13316), .ZN(n13266) );
  NAND2_X1 U15029 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  XNOR2_X1 U15030 ( .A(n13268), .B(n10643), .ZN(n13272) );
  NAND2_X1 U15031 ( .A1(n15718), .A2(n13316), .ZN(n13270) );
  NAND2_X1 U15032 ( .A1(n14924), .A2(n13315), .ZN(n13269) );
  NAND2_X1 U15033 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  NOR2_X1 U15034 ( .A1(n13272), .A2(n13271), .ZN(n14867) );
  AOI21_X1 U15035 ( .B1(n13272), .B2(n13271), .A(n14867), .ZN(n14807) );
  NAND2_X1 U15036 ( .A1(n15711), .A2(n13313), .ZN(n13274) );
  NAND2_X1 U15037 ( .A1(n15114), .A2(n13316), .ZN(n13273) );
  NAND2_X1 U15038 ( .A1(n13274), .A2(n13273), .ZN(n13275) );
  XNOR2_X1 U15039 ( .A(n13275), .B(n13305), .ZN(n13277) );
  AND2_X1 U15040 ( .A1(n15114), .A2(n13315), .ZN(n13276) );
  AOI21_X1 U15041 ( .B1(n15711), .B2(n13316), .A(n13276), .ZN(n13278) );
  NAND2_X1 U15042 ( .A1(n13277), .A2(n13278), .ZN(n14837) );
  INV_X1 U15043 ( .A(n13277), .ZN(n13280) );
  INV_X1 U15044 ( .A(n13278), .ZN(n13279) );
  NAND2_X1 U15045 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U15046 ( .A1(n15123), .A2(n13313), .ZN(n13283) );
  NAND2_X1 U15047 ( .A1(n13316), .A2(n14923), .ZN(n13282) );
  NAND2_X1 U15048 ( .A1(n13283), .A2(n13282), .ZN(n13284) );
  XNOR2_X1 U15049 ( .A(n13284), .B(n13305), .ZN(n13286) );
  NOR2_X1 U15050 ( .A1(n10968), .A2(n14898), .ZN(n13285) );
  AOI21_X1 U15051 ( .B1(n15123), .B2(n13316), .A(n13285), .ZN(n13287) );
  NAND2_X1 U15052 ( .A1(n13286), .A2(n13287), .ZN(n13292) );
  INV_X1 U15053 ( .A(n13286), .ZN(n13289) );
  INV_X1 U15054 ( .A(n13287), .ZN(n13288) );
  NAND2_X1 U15055 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  NAND2_X1 U15056 ( .A1(n15696), .A2(n13313), .ZN(n13294) );
  NAND2_X1 U15057 ( .A1(n13316), .A2(n14922), .ZN(n13293) );
  NAND2_X1 U15058 ( .A1(n13294), .A2(n13293), .ZN(n13295) );
  XNOR2_X1 U15059 ( .A(n13295), .B(n13305), .ZN(n13298) );
  INV_X1 U15060 ( .A(n13298), .ZN(n13300) );
  NOR2_X1 U15061 ( .A1(n10968), .A2(n15112), .ZN(n13296) );
  AOI21_X1 U15062 ( .B1(n15696), .B2(n13316), .A(n13296), .ZN(n13297) );
  INV_X1 U15063 ( .A(n13297), .ZN(n13299) );
  AND2_X1 U15064 ( .A1(n13298), .A2(n13297), .ZN(n13301) );
  AOI21_X1 U15065 ( .B1(n13300), .B2(n13299), .A(n13301), .ZN(n14896) );
  NAND2_X1 U15066 ( .A1(n15691), .A2(n13302), .ZN(n13304) );
  NAND2_X1 U15067 ( .A1(n13316), .A2(n15076), .ZN(n13303) );
  NAND2_X1 U15068 ( .A1(n13304), .A2(n13303), .ZN(n13306) );
  XNOR2_X1 U15069 ( .A(n13306), .B(n13305), .ZN(n13309) );
  INV_X1 U15070 ( .A(n13309), .ZN(n13311) );
  NOR2_X1 U15071 ( .A1(n10968), .A2(n14897), .ZN(n13307) );
  AOI21_X1 U15072 ( .B1(n15691), .B2(n13316), .A(n13307), .ZN(n13308) );
  INV_X1 U15073 ( .A(n13308), .ZN(n13310) );
  AND2_X1 U15074 ( .A1(n13309), .A2(n13308), .ZN(n13312) );
  AOI21_X1 U15075 ( .B1(n13311), .B2(n13310), .A(n13312), .ZN(n14796) );
  AOI22_X1 U15076 ( .A1(n15686), .A2(n13313), .B1(n13316), .B2(n14921), .ZN(
        n13314) );
  XNOR2_X1 U15077 ( .A(n13314), .B(n10643), .ZN(n13318) );
  AOI22_X1 U15078 ( .A1(n15686), .A2(n13316), .B1(n13315), .B2(n14921), .ZN(
        n13317) );
  XNOR2_X1 U15079 ( .A(n13318), .B(n13317), .ZN(n13319) );
  XNOR2_X1 U15080 ( .A(n13320), .B(n13319), .ZN(n13326) );
  OAI22_X1 U15081 ( .A1(n16558), .A2(n15086), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13321), .ZN(n13324) );
  OAI22_X1 U15082 ( .A1(n14897), .A2(n16543), .B1(n16542), .B2(n13322), .ZN(
        n13323) );
  AOI211_X1 U15083 ( .C1(n15686), .C2(n16554), .A(n13324), .B(n13323), .ZN(
        n13325) );
  OAI21_X1 U15084 ( .B1(n13326), .B2(n16549), .A(n13325), .ZN(P1_U3220) );
  NAND2_X1 U15085 ( .A1(n13328), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13331) );
  NAND2_X1 U15086 ( .A1(n7437), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U15087 ( .A1(n8498), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13329) );
  AND3_X1 U15088 ( .A1(n13331), .A2(n13330), .A3(n13329), .ZN(n13332) );
  NAND2_X1 U15089 ( .A1(n13333), .A2(n13332), .ZN(n13806) );
  INV_X1 U15090 ( .A(n13806), .ZN(n13501) );
  INV_X1 U15091 ( .A(n13334), .ZN(n13335) );
  NAND2_X1 U15092 ( .A1(n13336), .A2(n13335), .ZN(n13339) );
  NAND2_X1 U15093 ( .A1(n13337), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13338) );
  NAND2_X1 U15094 ( .A1(n13339), .A2(n13338), .ZN(n13345) );
  XNOR2_X1 U15095 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n13344) );
  INV_X1 U15096 ( .A(n13344), .ZN(n13340) );
  XNOR2_X1 U15097 ( .A(n13345), .B(n13340), .ZN(n13548) );
  NAND2_X1 U15098 ( .A1(n13548), .A2(n13353), .ZN(n13342) );
  INV_X1 U15099 ( .A(SI_30_), .ZN(n13550) );
  OR2_X1 U15100 ( .A1(n13351), .A2(n13550), .ZN(n13341) );
  NAND2_X1 U15101 ( .A1(n13342), .A2(n13341), .ZN(n13810) );
  INV_X1 U15102 ( .A(n13701), .ZN(n13354) );
  NAND2_X1 U15103 ( .A1(n13810), .A2(n13354), .ZN(n13534) );
  NAND2_X1 U15104 ( .A1(n13534), .A2(n13343), .ZN(n13500) );
  NAND2_X1 U15105 ( .A1(n13345), .A2(n13344), .ZN(n13348) );
  NAND2_X1 U15106 ( .A1(n13346), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U15107 ( .A1(n13348), .A2(n13347), .ZN(n13350) );
  XNOR2_X1 U15108 ( .A(n14771), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n13349) );
  XNOR2_X1 U15109 ( .A(n13350), .B(n13349), .ZN(n14213) );
  INV_X1 U15110 ( .A(SI_31_), .ZN(n14218) );
  NOR2_X1 U15111 ( .A1(n13351), .A2(n14218), .ZN(n13352) );
  AND2_X1 U15112 ( .A1(n14152), .A2(n13806), .ZN(n13538) );
  AOI211_X1 U15113 ( .C1(n13501), .C2(n13810), .A(n13500), .B(n13538), .ZN(
        n13356) );
  OR2_X1 U15114 ( .A1(n13810), .A2(n13354), .ZN(n13503) );
  AOI21_X1 U15115 ( .B1(n13806), .B2(n13503), .A(n14152), .ZN(n13355) );
  NOR2_X1 U15116 ( .A1(n13841), .A2(n13855), .ZN(n13359) );
  NAND2_X1 U15117 ( .A1(n13361), .A2(n13487), .ZN(n13362) );
  OAI211_X1 U15118 ( .C1(n13364), .C2(n13363), .A(n8970), .B(n13362), .ZN(
        n13373) );
  NAND2_X1 U15119 ( .A1(n13366), .A2(n13365), .ZN(n13369) );
  NAND3_X1 U15120 ( .A1(n13369), .A2(n13466), .A3(n13367), .ZN(n13368) );
  OAI21_X1 U15121 ( .B1(n13369), .B2(n13544), .A(n13368), .ZN(n13372) );
  AND2_X1 U15122 ( .A1(n13378), .A2(n13370), .ZN(n13371) );
  OAI22_X1 U15123 ( .A1(n13373), .A2(n13372), .B1(n13371), .B2(n13487), .ZN(
        n13377) );
  AOI21_X1 U15124 ( .B1(n13376), .B2(n13374), .A(n13466), .ZN(n13375) );
  AOI21_X1 U15125 ( .B1(n13377), .B2(n13376), .A(n13375), .ZN(n13384) );
  OAI21_X1 U15126 ( .B1(n13466), .B2(n13378), .A(n13518), .ZN(n13383) );
  NAND2_X1 U15127 ( .A1(n13712), .A2(n13379), .ZN(n13380) );
  MUX2_X1 U15128 ( .A(n13381), .B(n13380), .S(n13466), .Z(n13382) );
  OAI21_X1 U15129 ( .B1(n13384), .B2(n13383), .A(n13382), .ZN(n13385) );
  NAND2_X1 U15130 ( .A1(n13385), .A2(n13512), .ZN(n13386) );
  NAND2_X1 U15131 ( .A1(n13386), .A2(n13516), .ZN(n13394) );
  INV_X1 U15132 ( .A(n13387), .ZN(n13389) );
  OAI21_X1 U15133 ( .B1(n13394), .B2(n13389), .A(n13388), .ZN(n13396) );
  INV_X1 U15134 ( .A(n13390), .ZN(n13393) );
  OAI22_X1 U15135 ( .A1(n13394), .A2(n13393), .B1(n13392), .B2(n13391), .ZN(
        n13395) );
  MUX2_X1 U15136 ( .A(n13396), .B(n13395), .S(n13487), .Z(n13398) );
  NAND2_X1 U15137 ( .A1(n13398), .A2(n13397), .ZN(n13402) );
  MUX2_X1 U15138 ( .A(n13400), .B(n13399), .S(n13466), .Z(n13401) );
  NAND3_X1 U15139 ( .A1(n13402), .A2(n13517), .A3(n13401), .ZN(n13408) );
  INV_X1 U15140 ( .A(n13403), .ZN(n13521) );
  NAND2_X1 U15141 ( .A1(n13707), .A2(n16439), .ZN(n13404) );
  MUX2_X1 U15142 ( .A(n13405), .B(n13404), .S(n13466), .Z(n13406) );
  NAND4_X1 U15143 ( .A1(n13408), .A2(n13407), .A3(n13521), .A4(n13406), .ZN(
        n13417) );
  MUX2_X1 U15144 ( .A(n13410), .B(n13409), .S(n13466), .Z(n13411) );
  NAND2_X1 U15145 ( .A1(n13411), .A2(n13521), .ZN(n13415) );
  MUX2_X1 U15146 ( .A(n13413), .B(n13412), .S(n13466), .Z(n13414) );
  AND3_X1 U15147 ( .A1(n13415), .A2(n14091), .A3(n13414), .ZN(n13416) );
  NAND2_X1 U15148 ( .A1(n13417), .A2(n13416), .ZN(n13425) );
  NAND3_X1 U15149 ( .A1(n13425), .A2(n13426), .A3(n13418), .ZN(n13419) );
  NAND3_X1 U15150 ( .A1(n13419), .A2(n13423), .A3(n13487), .ZN(n13420) );
  NAND2_X1 U15151 ( .A1(n13420), .A2(n14051), .ZN(n13422) );
  NAND3_X1 U15152 ( .A1(n16517), .A2(n14036), .A3(n13487), .ZN(n13421) );
  NAND2_X1 U15153 ( .A1(n13422), .A2(n13421), .ZN(n13429) );
  NAND3_X1 U15154 ( .A1(n13425), .A2(n13424), .A3(n13423), .ZN(n13427) );
  NAND3_X1 U15155 ( .A1(n13427), .A2(n13466), .A3(n13426), .ZN(n13428) );
  NAND4_X1 U15156 ( .A1(n13429), .A2(n8691), .A3(n13527), .A4(n13428), .ZN(
        n13437) );
  MUX2_X1 U15157 ( .A(n13430), .B(n13947), .S(n13466), .Z(n13436) );
  AOI21_X1 U15158 ( .B1(n13431), .B2(n14040), .A(n13487), .ZN(n13433) );
  NAND2_X1 U15159 ( .A1(n16534), .A2(n13655), .ZN(n13432) );
  MUX2_X1 U15160 ( .A(n13487), .B(n13433), .S(n13432), .Z(n13434) );
  NAND2_X1 U15161 ( .A1(n8691), .A2(n13434), .ZN(n13435) );
  NAND3_X1 U15162 ( .A1(n13437), .A2(n13436), .A3(n13435), .ZN(n13444) );
  MUX2_X1 U15163 ( .A(n14208), .B(n14028), .S(n13466), .Z(n13440) );
  INV_X1 U15164 ( .A(n13440), .ZN(n13439) );
  NAND2_X1 U15165 ( .A1(n13439), .A2(n13438), .ZN(n13443) );
  NAND2_X1 U15166 ( .A1(n13440), .A2(n13984), .ZN(n13441) );
  NAND4_X1 U15167 ( .A1(n13994), .A2(n13452), .A3(n13450), .A4(n13441), .ZN(
        n13442) );
  AOI21_X1 U15168 ( .B1(n13444), .B2(n13443), .A(n13442), .ZN(n13457) );
  NAND2_X1 U15169 ( .A1(n13450), .A2(n13445), .ZN(n13446) );
  AND2_X1 U15170 ( .A1(n13446), .A2(n13452), .ZN(n13448) );
  OR2_X1 U15171 ( .A1(n13448), .A2(n13447), .ZN(n13454) );
  NAND3_X1 U15172 ( .A1(n13450), .A2(n14203), .A3(n13705), .ZN(n13451) );
  NAND3_X1 U15173 ( .A1(n13510), .A2(n13452), .A3(n13451), .ZN(n13453) );
  MUX2_X1 U15174 ( .A(n13454), .B(n13453), .S(n13466), .Z(n13456) );
  MUX2_X1 U15175 ( .A(n13510), .B(n13511), .S(n13466), .Z(n13455) );
  OAI211_X1 U15176 ( .C1(n13457), .C2(n13456), .A(n13931), .B(n13455), .ZN(
        n13460) );
  INV_X1 U15177 ( .A(n13907), .ZN(n13911) );
  MUX2_X1 U15178 ( .A(n13906), .B(n13458), .S(n13466), .Z(n13459) );
  NAND3_X1 U15179 ( .A1(n13460), .A2(n13911), .A3(n13459), .ZN(n13465) );
  INV_X1 U15180 ( .A(n13461), .ZN(n13468) );
  MUX2_X1 U15181 ( .A(n13463), .B(n13462), .S(n13466), .Z(n13464) );
  NAND4_X1 U15182 ( .A1(n13465), .A2(n13895), .A3(n13881), .A4(n13464), .ZN(
        n13476) );
  MUX2_X1 U15183 ( .A(n13468), .B(n13467), .S(n13466), .Z(n13469) );
  INV_X1 U15184 ( .A(n13469), .ZN(n13470) );
  NAND2_X1 U15185 ( .A1(n13881), .A2(n13470), .ZN(n13474) );
  MUX2_X1 U15186 ( .A(n13472), .B(n13471), .S(n13487), .Z(n13473) );
  NAND2_X1 U15187 ( .A1(n13474), .A2(n13473), .ZN(n13475) );
  NAND2_X1 U15188 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  NAND2_X1 U15189 ( .A1(n13478), .A2(n13840), .ZN(n13479) );
  NAND3_X1 U15190 ( .A1(n13481), .A2(n13480), .A3(n13479), .ZN(n13483) );
  NAND2_X1 U15191 ( .A1(n13483), .A2(n13482), .ZN(n13489) );
  INV_X1 U15192 ( .A(n13489), .ZN(n13484) );
  NAND2_X1 U15193 ( .A1(n13488), .A2(n13466), .ZN(n13495) );
  AOI21_X1 U15194 ( .B1(n13533), .B2(n13490), .A(n13489), .ZN(n13491) );
  NAND2_X1 U15195 ( .A1(n13495), .A2(n13494), .ZN(n13499) );
  OAI211_X1 U15196 ( .C1(n13499), .C2(n8054), .A(n13498), .B(n13497), .ZN(
        n13506) );
  INV_X1 U15197 ( .A(n13500), .ZN(n13505) );
  INV_X1 U15198 ( .A(n14152), .ZN(n13502) );
  NAND2_X1 U15199 ( .A1(n13502), .A2(n13501), .ZN(n13504) );
  NAND2_X1 U15200 ( .A1(n13504), .A2(n13503), .ZN(n13536) );
  AOI21_X1 U15201 ( .B1(n13506), .B2(n13505), .A(n13536), .ZN(n13507) );
  NOR4_X1 U15202 ( .A1(n13515), .A2(n8515), .A3(n13514), .A4(n13513), .ZN(
        n13519) );
  NAND4_X1 U15203 ( .A1(n13519), .A2(n13518), .A3(n13517), .A4(n13516), .ZN(
        n13525) );
  INV_X1 U15204 ( .A(n14091), .ZN(n14083) );
  INV_X1 U15205 ( .A(n14068), .ZN(n13524) );
  NAND4_X1 U15206 ( .A1(n13522), .A2(n13521), .A3(n8970), .A4(n13520), .ZN(
        n13523) );
  NOR4_X1 U15207 ( .A1(n13525), .A2(n14083), .A3(n13524), .A4(n13523), .ZN(
        n13526) );
  NAND4_X1 U15208 ( .A1(n8691), .A2(n13527), .A3(n14051), .A4(n13526), .ZN(
        n13528) );
  NOR4_X1 U15209 ( .A1(n13961), .A2(n13528), .A3(n8711), .A4(n13983), .ZN(
        n13529) );
  NAND4_X1 U15210 ( .A1(n13911), .A2(n13931), .A3(n13950), .A4(n13529), .ZN(
        n13530) );
  NOR4_X1 U15211 ( .A1(n13873), .A2(n7935), .A3(n13531), .A4(n13530), .ZN(
        n13532) );
  NAND4_X1 U15212 ( .A1(n8994), .A2(n9063), .A3(n13533), .A4(n13532), .ZN(
        n13537) );
  INV_X1 U15213 ( .A(n13534), .ZN(n13535) );
  XNOR2_X1 U15214 ( .A(n13539), .B(n13799), .ZN(n13540) );
  NOR3_X1 U15215 ( .A1(n13543), .A2(n13542), .A3(n8956), .ZN(n13546) );
  OAI21_X1 U15216 ( .B1(n13547), .B2(n13544), .A(P3_B_REG_SCAN_IN), .ZN(n13545) );
  INV_X1 U15217 ( .A(n13548), .ZN(n13549) );
  OAI222_X1 U15218 ( .A1(n8418), .A2(P3_U3151), .B1(n14223), .B2(n13550), .C1(
        n14221), .C2(n13549), .ZN(P3_U3265) );
  INV_X1 U15219 ( .A(n13551), .ZN(n13663) );
  NAND2_X1 U15220 ( .A1(n13553), .A2(n13552), .ZN(n13605) );
  INV_X1 U15221 ( .A(n13554), .ZN(n13603) );
  NOR2_X1 U15222 ( .A1(n13605), .A2(n13603), .ZN(n13660) );
  NOR3_X1 U15223 ( .A1(n13660), .A2(n13659), .A3(n13663), .ZN(n13661) );
  AOI21_X1 U15224 ( .B1(n14036), .B2(n13663), .A(n13661), .ZN(n13557) );
  OAI21_X1 U15225 ( .B1(n13557), .B2(n13556), .A(n13555), .ZN(n13558) );
  NAND2_X1 U15226 ( .A1(n13558), .A2(n13690), .ZN(n13562) );
  NAND2_X1 U15227 ( .A1(n13692), .A2(n14036), .ZN(n13559) );
  NAND2_X1 U15228 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n16182)
         );
  OAI211_X1 U15229 ( .C1(n14039), .C2(n13671), .A(n13559), .B(n16182), .ZN(
        n13560) );
  AOI21_X1 U15230 ( .B1(n14044), .B2(n13683), .A(n13560), .ZN(n13561) );
  OAI211_X1 U15231 ( .C1(n13700), .C2(n16534), .A(n13562), .B(n13561), .ZN(
        P3_U3155) );
  OAI21_X1 U15232 ( .B1(n13897), .B2(n13564), .A(n13640), .ZN(n13565) );
  NAND2_X1 U15233 ( .A1(n13565), .A2(n13690), .ZN(n13569) );
  AOI22_X1 U15234 ( .A1(n13914), .A2(n13692), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13566) );
  OAI21_X1 U15235 ( .B1(n13859), .B2(n13671), .A(n13566), .ZN(n13567) );
  AOI21_X1 U15236 ( .B1(n13887), .B2(n13683), .A(n13567), .ZN(n13568) );
  OAI211_X1 U15237 ( .C1(n14175), .C2(n13700), .A(n13569), .B(n13568), .ZN(
        P3_U3156) );
  OAI211_X1 U15238 ( .C1(n13571), .C2(n13573), .A(n13572), .B(n13690), .ZN(
        n13577) );
  NAND2_X1 U15239 ( .A1(n13692), .A2(n13985), .ZN(n13574) );
  NAND2_X1 U15240 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13798)
         );
  OAI211_X1 U15241 ( .C1(n13945), .C2(n13671), .A(n13574), .B(n13798), .ZN(
        n13575) );
  AOI21_X1 U15242 ( .B1(n13952), .B2(n13683), .A(n13575), .ZN(n13576) );
  OAI211_X1 U15243 ( .C1(n14195), .C2(n13700), .A(n13577), .B(n13576), .ZN(
        P3_U3159) );
  OAI21_X1 U15244 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n13581) );
  NAND2_X1 U15245 ( .A1(n13581), .A2(n13690), .ZN(n13589) );
  OAI22_X1 U15246 ( .A1(n13582), .A2(n13671), .B1(n8448), .B2(n13700), .ZN(
        n13583) );
  INV_X1 U15247 ( .A(n13583), .ZN(n13588) );
  NAND2_X1 U15248 ( .A1(n13584), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n13587) );
  NAND2_X1 U15249 ( .A1(n13692), .A2(n13585), .ZN(n13586) );
  NAND4_X1 U15250 ( .A1(n13589), .A2(n13588), .A3(n13587), .A4(n13586), .ZN(
        P3_U3162) );
  NAND2_X1 U15251 ( .A1(n13591), .A2(n13590), .ZN(n13593) );
  XOR2_X1 U15252 ( .A(n13593), .B(n13592), .Z(n13599) );
  AOI22_X1 U15253 ( .A1(n13915), .A2(n13692), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13595) );
  NAND2_X1 U15254 ( .A1(n13683), .A2(n13920), .ZN(n13594) );
  OAI211_X1 U15255 ( .C1(n13596), .C2(n13671), .A(n13595), .B(n13594), .ZN(
        n13597) );
  AOI21_X1 U15256 ( .B1(n13921), .B2(n13673), .A(n13597), .ZN(n13598) );
  OAI21_X1 U15257 ( .B1(n13599), .B2(n13675), .A(n13598), .ZN(P3_U3163) );
  INV_X1 U15258 ( .A(n13600), .ZN(n14074) );
  NOR2_X1 U15259 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15335), .ZN(n16156) );
  AOI21_X1 U15260 ( .B1(n13697), .B2(n14036), .A(n16156), .ZN(n13602) );
  NAND2_X1 U15261 ( .A1(n13692), .A2(n13706), .ZN(n13601) );
  OAI211_X1 U15262 ( .C1(n14074), .C2(n13694), .A(n13602), .B(n13601), .ZN(
        n13608) );
  NOR2_X1 U15263 ( .A1(n13659), .A2(n13603), .ZN(n13604) );
  XNOR2_X1 U15264 ( .A(n13605), .B(n13604), .ZN(n13606) );
  NOR2_X1 U15265 ( .A1(n13606), .A2(n13675), .ZN(n13607) );
  AOI211_X1 U15266 ( .C1(n14077), .C2(n13673), .A(n13608), .B(n13607), .ZN(
        n13609) );
  INV_X1 U15267 ( .A(n13609), .ZN(P3_U3164) );
  INV_X1 U15268 ( .A(n14164), .ZN(n13620) );
  INV_X1 U15269 ( .A(n13610), .ZN(n13614) );
  NOR3_X1 U15270 ( .A1(n13642), .A2(n13612), .A3(n13611), .ZN(n13613) );
  OAI21_X1 U15271 ( .B1(n13614), .B2(n13613), .A(n13690), .ZN(n13619) );
  AOI22_X1 U15272 ( .A1(n13884), .A2(n13692), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13615) );
  OAI21_X1 U15273 ( .B1(n13616), .B2(n13671), .A(n13615), .ZN(n13617) );
  AOI21_X1 U15274 ( .B1(n13865), .B2(n13683), .A(n13617), .ZN(n13618) );
  OAI211_X1 U15275 ( .C1(n13620), .C2(n13700), .A(n13619), .B(n13618), .ZN(
        P3_U3165) );
  OAI211_X1 U15276 ( .C1(n13623), .C2(n13622), .A(n13621), .B(n13690), .ZN(
        n13629) );
  INV_X1 U15277 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13624) );
  NOR2_X1 U15278 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13624), .ZN(n16222) );
  AOI21_X1 U15279 ( .B1(n13692), .B2(n13625), .A(n16222), .ZN(n13626) );
  OAI21_X1 U15280 ( .B1(n14012), .B2(n13671), .A(n13626), .ZN(n13627) );
  AOI21_X1 U15281 ( .B1(n14016), .B2(n13683), .A(n13627), .ZN(n13628) );
  OAI211_X1 U15282 ( .C1(n14208), .C2(n13700), .A(n13629), .B(n13628), .ZN(
        P3_U3166) );
  OAI211_X1 U15283 ( .C1(n13632), .C2(n13631), .A(n13630), .B(n13690), .ZN(
        n13636) );
  AND2_X1 U15284 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n16248) );
  AOI21_X1 U15285 ( .B1(n13697), .B2(n13985), .A(n16248), .ZN(n13633) );
  OAI21_X1 U15286 ( .B1(n14028), .B2(n13681), .A(n13633), .ZN(n13634) );
  AOI21_X1 U15287 ( .B1(n13996), .B2(n13683), .A(n13634), .ZN(n13635) );
  OAI211_X1 U15288 ( .C1(n14203), .C2(n13700), .A(n13636), .B(n13635), .ZN(
        P3_U3168) );
  AND3_X1 U15289 ( .A1(n13640), .A2(n13639), .A3(n13638), .ZN(n13641) );
  OAI21_X1 U15290 ( .B1(n13642), .B2(n13641), .A(n13690), .ZN(n13646) );
  AOI22_X1 U15291 ( .A1(n13871), .A2(n13692), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13643) );
  OAI21_X1 U15292 ( .B1(n13838), .B2(n13671), .A(n13643), .ZN(n13644) );
  AOI21_X1 U15293 ( .B1(n13876), .B2(n13683), .A(n13644), .ZN(n13645) );
  OAI211_X1 U15294 ( .C1(n14171), .C2(n13700), .A(n13646), .B(n13645), .ZN(
        P3_U3169) );
  INV_X1 U15295 ( .A(n13940), .ZN(n14187) );
  OAI211_X1 U15296 ( .C1(n13649), .C2(n13648), .A(n13647), .B(n13690), .ZN(
        n13653) );
  AOI22_X1 U15297 ( .A1(n13703), .A2(n13697), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13650) );
  OAI21_X1 U15298 ( .B1(n13965), .B2(n13681), .A(n13650), .ZN(n13651) );
  AOI21_X1 U15299 ( .B1(n13939), .B2(n13683), .A(n13651), .ZN(n13652) );
  OAI211_X1 U15300 ( .C1(n14187), .C2(n13700), .A(n13653), .B(n13652), .ZN(
        P3_U3173) );
  INV_X1 U15301 ( .A(n13654), .ZN(n14059) );
  NOR2_X1 U15302 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15554), .ZN(n16168) );
  AOI21_X1 U15303 ( .B1(n13697), .B2(n13655), .A(n16168), .ZN(n13658) );
  NAND2_X1 U15304 ( .A1(n13692), .A2(n13656), .ZN(n13657) );
  OAI211_X1 U15305 ( .C1(n14059), .C2(n13694), .A(n13658), .B(n13657), .ZN(
        n13665) );
  OR2_X1 U15306 ( .A1(n13660), .A2(n13659), .ZN(n13662) );
  AOI211_X1 U15307 ( .C1(n13663), .C2(n13662), .A(n13675), .B(n13661), .ZN(
        n13664) );
  AOI211_X1 U15308 ( .C1(n14061), .C2(n13673), .A(n13665), .B(n13664), .ZN(
        n13666) );
  INV_X1 U15309 ( .A(n13666), .ZN(P3_U3174) );
  AOI21_X1 U15310 ( .B1(n13914), .B2(n13668), .A(n13667), .ZN(n13676) );
  AOI22_X1 U15311 ( .A1(n13703), .A2(n13692), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13670) );
  NAND2_X1 U15312 ( .A1(n13683), .A2(n13902), .ZN(n13669) );
  OAI211_X1 U15313 ( .C1(n13897), .C2(n13671), .A(n13670), .B(n13669), .ZN(
        n13672) );
  AOI21_X1 U15314 ( .B1(n13903), .B2(n13673), .A(n13672), .ZN(n13674) );
  OAI21_X1 U15315 ( .B1(n13676), .B2(n13675), .A(n13674), .ZN(P3_U3175) );
  OAI211_X1 U15316 ( .C1(n13679), .C2(n13678), .A(n13677), .B(n13690), .ZN(
        n13685) );
  AND2_X1 U15317 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n16264) );
  AOI21_X1 U15318 ( .B1(n13697), .B2(n13704), .A(n16264), .ZN(n13680) );
  OAI21_X1 U15319 ( .B1(n14012), .B2(n13681), .A(n13680), .ZN(n13682) );
  AOI21_X1 U15320 ( .B1(n13974), .B2(n13683), .A(n13682), .ZN(n13684) );
  OAI211_X1 U15321 ( .C1(n14199), .C2(n13700), .A(n13685), .B(n13684), .ZN(
        P3_U3178) );
  OAI21_X1 U15322 ( .B1(n13689), .B2(n13688), .A(n13687), .ZN(n13691) );
  NAND2_X1 U15323 ( .A1(n13691), .A2(n13690), .ZN(n13699) );
  INV_X1 U15324 ( .A(n13845), .ZN(n13695) );
  AOI22_X1 U15325 ( .A1(n13870), .A2(n13692), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13693) );
  OAI21_X1 U15326 ( .B1(n13695), .B2(n13694), .A(n13693), .ZN(n13696) );
  AOI21_X1 U15327 ( .B1(n13697), .B2(n13702), .A(n13696), .ZN(n13698) );
  OAI211_X1 U15328 ( .C1(n14160), .C2(n13700), .A(n13699), .B(n13698), .ZN(
        P3_U3180) );
  MUX2_X1 U15329 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13806), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15330 ( .A(n13701), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13711), .Z(
        P3_U3521) );
  MUX2_X1 U15331 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13702), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15332 ( .A(n13857), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13711), .Z(
        P3_U3517) );
  MUX2_X1 U15333 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13870), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15334 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13884), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15335 ( .A(n13871), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13711), .Z(
        P3_U3514) );
  MUX2_X1 U15336 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13914), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15337 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13703), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15338 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13915), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15339 ( .A(n13704), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13711), .Z(
        P3_U3510) );
  MUX2_X1 U15340 ( .A(n13985), .B(P3_DATAO_REG_18__SCAN_IN), .S(n13711), .Z(
        P3_U3509) );
  MUX2_X1 U15341 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13705), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15342 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13988), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15343 ( .A(n14036), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13711), .Z(
        P3_U3504) );
  MUX2_X1 U15344 ( .A(n13706), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13711), .Z(
        P3_U3502) );
  MUX2_X1 U15345 ( .A(n13707), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13711), .Z(
        P3_U3499) );
  MUX2_X1 U15346 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13708), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15347 ( .A(n13709), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13711), .Z(
        P3_U3497) );
  MUX2_X1 U15348 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13710), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15349 ( .A(n13712), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13711), .Z(
        P3_U3495) );
  MUX2_X1 U15350 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13713), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15351 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13714), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15352 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13715), .S(P3_U3897), .Z(
        P3_U3492) );
  INV_X1 U15353 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n16233) );
  INV_X1 U15354 ( .A(n13776), .ZN(n16159) );
  INV_X1 U15355 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14075) );
  OR2_X1 U15356 ( .A1(n13741), .A2(n14075), .ZN(n13774) );
  INV_X1 U15357 ( .A(n13774), .ZN(n13721) );
  AOI21_X1 U15358 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13717), .A(n13716), 
        .ZN(n13718) );
  NOR2_X1 U15359 ( .A1(n13768), .A2(n13718), .ZN(n13719) );
  INV_X1 U15360 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U15361 ( .A1(n13741), .A2(n14075), .ZN(n13720) );
  NAND2_X1 U15362 ( .A1(n13774), .A2(n13720), .ZN(n16142) );
  INV_X1 U15363 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n16170) );
  INV_X1 U15364 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13723) );
  OR2_X1 U15365 ( .A1(n16185), .A2(n13723), .ZN(n13725) );
  NAND2_X1 U15366 ( .A1(n16185), .A2(n13723), .ZN(n13724) );
  AND2_X1 U15367 ( .A1(n13725), .A2(n13724), .ZN(n16177) );
  NOR2_X1 U15368 ( .A1(n16178), .A2(n16177), .ZN(n16176) );
  INV_X1 U15369 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n16207) );
  NAND2_X1 U15370 ( .A1(n13758), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n13728) );
  INV_X1 U15371 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U15372 ( .A1(n16213), .A2(n13757), .ZN(n13727) );
  NAND2_X1 U15373 ( .A1(n13728), .A2(n13727), .ZN(n16224) );
  NOR2_X1 U15374 ( .A1(n13756), .A2(n13730), .ZN(n13731) );
  OR2_X1 U15375 ( .A1(n16253), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U15376 ( .A1(n16253), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13732) );
  AND2_X1 U15377 ( .A1(n13733), .A2(n13732), .ZN(n16266) );
  AOI21_X1 U15378 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13793), .A(n16267), 
        .ZN(n13735) );
  INV_X1 U15379 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13734) );
  MUX2_X1 U15380 ( .A(n13734), .B(P3_REG2_REG_19__SCAN_IN), .S(n13736), .Z(
        n13755) );
  XNOR2_X1 U15381 ( .A(n13735), .B(n13755), .ZN(n13804) );
  XNOR2_X1 U15382 ( .A(n13736), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13754) );
  NAND2_X1 U15383 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13758), .ZN(n13750) );
  XNOR2_X1 U15384 ( .A(n16213), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n16218) );
  INV_X1 U15385 ( .A(n16185), .ZN(n13747) );
  INV_X1 U15386 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n16538) );
  INV_X1 U15387 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13737) );
  OR2_X1 U15388 ( .A1(n13741), .A2(n13737), .ZN(n13773) );
  NAND2_X1 U15389 ( .A1(n16134), .A2(n13739), .ZN(n13740) );
  NAND2_X1 U15390 ( .A1(n13741), .A2(n13737), .ZN(n13742) );
  NAND2_X1 U15391 ( .A1(n13773), .A2(n13742), .ZN(n13772) );
  INV_X1 U15392 ( .A(n13772), .ZN(n16145) );
  NAND2_X1 U15393 ( .A1(n16144), .A2(n16145), .ZN(n16143) );
  NAND2_X1 U15394 ( .A1(n13773), .A2(n16143), .ZN(n13743) );
  NAND2_X1 U15395 ( .A1(n13776), .A2(n13743), .ZN(n13744) );
  XNOR2_X1 U15396 ( .A(n16159), .B(n13743), .ZN(n16161) );
  NAND2_X1 U15397 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n16161), .ZN(n16160) );
  OR2_X1 U15398 ( .A1(n16185), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13746) );
  NAND2_X1 U15399 ( .A1(n16185), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13745) );
  AND2_X1 U15400 ( .A1(n13746), .A2(n13745), .ZN(n16181) );
  NAND2_X1 U15401 ( .A1(n13785), .A2(n13748), .ZN(n13749) );
  NAND2_X1 U15402 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n16199), .ZN(n16198) );
  NAND2_X1 U15403 ( .A1(n13749), .A2(n16198), .ZN(n16219) );
  NAND2_X1 U15404 ( .A1(n16218), .A2(n16219), .ZN(n16217) );
  NAND2_X1 U15405 ( .A1(n16243), .A2(n13751), .ZN(n13752) );
  XNOR2_X1 U15406 ( .A(n16253), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n16255) );
  AOI22_X1 U15407 ( .A1(n16256), .A2(n16255), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n13793), .ZN(n13753) );
  XOR2_X1 U15408 ( .A(n13754), .B(n13753), .Z(n13802) );
  MUX2_X1 U15409 ( .A(n13755), .B(n13754), .S(n13791), .Z(n13795) );
  MUX2_X1 U15410 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13791), .Z(n13789) );
  XNOR2_X1 U15411 ( .A(n13789), .B(n13756), .ZN(n16239) );
  INV_X1 U15412 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n14147) );
  MUX2_X1 U15413 ( .A(n13757), .B(n14147), .S(n13791), .Z(n13788) );
  XNOR2_X1 U15414 ( .A(n13788), .B(n13758), .ZN(n16215) );
  MUX2_X1 U15415 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13791), .Z(n13781) );
  AND2_X1 U15416 ( .A1(n13781), .A2(n16185), .ZN(n13782) );
  NAND2_X1 U15417 ( .A1(n13760), .A2(n13759), .ZN(n13765) );
  INV_X1 U15418 ( .A(n13761), .ZN(n13763) );
  NAND2_X1 U15419 ( .A1(n13763), .A2(n13762), .ZN(n13764) );
  NAND2_X1 U15420 ( .A1(n13765), .A2(n13764), .ZN(n16130) );
  MUX2_X1 U15421 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n7414), .Z(n13767) );
  XNOR2_X1 U15422 ( .A(n13767), .B(n13768), .ZN(n16131) );
  NAND2_X1 U15423 ( .A1(n16130), .A2(n16131), .ZN(n13771) );
  INV_X1 U15424 ( .A(n13767), .ZN(n13769) );
  NAND2_X1 U15425 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  NAND2_X1 U15426 ( .A1(n13771), .A2(n13770), .ZN(n16149) );
  MUX2_X1 U15427 ( .A(n16142), .B(n13772), .S(n13791), .Z(n16150) );
  OR2_X1 U15428 ( .A1(n16149), .A2(n16150), .ZN(n16147) );
  MUX2_X1 U15429 ( .A(n13774), .B(n13773), .S(n13791), .Z(n13775) );
  NAND2_X1 U15430 ( .A1(n16147), .A2(n13775), .ZN(n16163) );
  MUX2_X1 U15431 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13791), .Z(n13777) );
  XNOR2_X1 U15432 ( .A(n13777), .B(n13776), .ZN(n16162) );
  INV_X1 U15433 ( .A(n13777), .ZN(n13778) );
  NAND2_X1 U15434 ( .A1(n13778), .A2(n16159), .ZN(n13779) );
  INV_X1 U15435 ( .A(n13782), .ZN(n13780) );
  OAI21_X1 U15436 ( .B1(n13781), .B2(n16185), .A(n13780), .ZN(n16188) );
  NOR2_X1 U15437 ( .A1(n16189), .A2(n16188), .ZN(n16192) );
  NAND2_X1 U15438 ( .A1(n16197), .A2(n13784), .ZN(n13786) );
  INV_X1 U15439 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13783) );
  MUX2_X1 U15440 ( .A(n16207), .B(n13783), .S(n13791), .Z(n16201) );
  XNOR2_X1 U15441 ( .A(n13785), .B(n13784), .ZN(n16202) );
  NAND2_X1 U15442 ( .A1(n16201), .A2(n16202), .ZN(n16200) );
  NAND2_X1 U15443 ( .A1(n13786), .A2(n16200), .ZN(n16216) );
  NAND2_X1 U15444 ( .A1(n16215), .A2(n16216), .ZN(n16214) );
  INV_X1 U15445 ( .A(n16214), .ZN(n13787) );
  NAND2_X1 U15446 ( .A1(n16239), .A2(n16238), .ZN(n16237) );
  NAND2_X1 U15447 ( .A1(n13789), .A2(n16243), .ZN(n13790) );
  NAND2_X1 U15448 ( .A1(n16237), .A2(n13790), .ZN(n13794) );
  XNOR2_X1 U15449 ( .A(n13794), .B(n16253), .ZN(n16259) );
  INV_X1 U15450 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13792) );
  INV_X1 U15451 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14139) );
  MUX2_X1 U15452 ( .A(n13792), .B(n14139), .S(n13791), .Z(n16258) );
  NAND2_X1 U15453 ( .A1(n16259), .A2(n16258), .ZN(n16257) );
  NOR2_X1 U15454 ( .A1(n13796), .A2(n16190), .ZN(n13801) );
  NAND2_X1 U15455 ( .A1(n16252), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13797) );
  OAI211_X1 U15456 ( .C1(n16244), .C2(n13799), .A(n13798), .B(n13797), .ZN(
        n13800) );
  OAI21_X1 U15457 ( .B1(n13804), .B2(n16250), .A(n13803), .ZN(P3_U3201) );
  NAND2_X1 U15458 ( .A1(n13806), .A2(n13805), .ZN(n14150) );
  INV_X1 U15459 ( .A(n14150), .ZN(n13808) );
  NOR2_X1 U15460 ( .A1(n13807), .A2(n14073), .ZN(n13817) );
  NOR3_X1 U15461 ( .A1(n13808), .A2(n14100), .A3(n13817), .ZN(n13812) );
  NOR2_X1 U15462 ( .A1(n16340), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13809) );
  OAI22_X1 U15463 ( .A1(n14152), .A2(n14046), .B1(n13812), .B2(n13809), .ZN(
        P3_U3202) );
  INV_X1 U15464 ( .A(n13810), .ZN(n14155) );
  NOR2_X1 U15465 ( .A1(n16340), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13811) );
  OAI22_X1 U15466 ( .A1(n14155), .A2(n14046), .B1(n13812), .B2(n13811), .ZN(
        P3_U3203) );
  INV_X1 U15467 ( .A(n13813), .ZN(n13820) );
  NAND2_X1 U15468 ( .A1(n13814), .A2(n16340), .ZN(n13819) );
  NOR2_X1 U15469 ( .A1(n13815), .A2(n14046), .ZN(n13816) );
  AOI211_X1 U15470 ( .C1(n14100), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13817), 
        .B(n13816), .ZN(n13818) );
  OAI211_X1 U15471 ( .C1(n13820), .C2(n13892), .A(n13819), .B(n13818), .ZN(
        P3_U3204) );
  AOI22_X1 U15472 ( .A1(n13821), .A2(n16337), .B1(n14100), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13822) );
  OAI21_X1 U15473 ( .B1(n13823), .B2(n14046), .A(n13822), .ZN(n13824) );
  AOI21_X1 U15474 ( .B1(n13825), .B2(n14098), .A(n13824), .ZN(n13826) );
  OAI21_X1 U15475 ( .B1(n13827), .B2(n14100), .A(n13826), .ZN(P3_U3205) );
  XNOR2_X1 U15476 ( .A(n13830), .B(n8914), .ZN(n14106) );
  AOI22_X1 U15477 ( .A1(n13831), .A2(n16337), .B1(n14100), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13832) );
  OAI21_X1 U15478 ( .B1(n13833), .B2(n14046), .A(n13832), .ZN(n13834) );
  AOI21_X1 U15479 ( .B1(n14106), .B2(n14098), .A(n13834), .ZN(n13835) );
  OAI21_X1 U15480 ( .B1(n14108), .B2(n14100), .A(n13835), .ZN(P3_U3206) );
  XNOR2_X1 U15481 ( .A(n13836), .B(n13841), .ZN(n13837) );
  OAI222_X1 U15482 ( .A1(n14089), .A2(n13839), .B1(n14087), .B2(n13838), .C1(
        n13837), .C2(n14084), .ZN(n14109) );
  NAND2_X1 U15483 ( .A1(n13853), .A2(n13840), .ZN(n13842) );
  NAND2_X1 U15484 ( .A1(n13842), .A2(n13841), .ZN(n13843) );
  NAND2_X1 U15485 ( .A1(n14110), .A2(n14098), .ZN(n13847) );
  AOI22_X1 U15486 ( .A1(n13845), .A2(n16337), .B1(n14100), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13846) );
  OAI211_X1 U15487 ( .C1(n14160), .C2(n14046), .A(n13847), .B(n13846), .ZN(
        n13848) );
  AOI21_X1 U15488 ( .B1(n14109), .B2(n16340), .A(n13848), .ZN(n13849) );
  INV_X1 U15489 ( .A(n13849), .ZN(P3_U3207) );
  OR2_X1 U15490 ( .A1(n13851), .A2(n13850), .ZN(n13852) );
  NAND2_X1 U15491 ( .A1(n13853), .A2(n13852), .ZN(n13861) );
  OAI211_X1 U15492 ( .C1(n13856), .C2(n13855), .A(n13854), .B(n13979), .ZN(
        n13863) );
  NAND2_X1 U15493 ( .A1(n13857), .A2(n13986), .ZN(n13858) );
  OAI21_X1 U15494 ( .B1(n13859), .B2(n14087), .A(n13858), .ZN(n13860) );
  AOI21_X1 U15495 ( .B1(n13861), .B2(n16428), .A(n13860), .ZN(n13862) );
  NAND2_X1 U15496 ( .A1(n13863), .A2(n13862), .ZN(n14113) );
  MUX2_X1 U15497 ( .A(n14113), .B(P3_REG2_REG_25__SCAN_IN), .S(n14100), .Z(
        n13864) );
  INV_X1 U15498 ( .A(n13864), .ZN(n13867) );
  AOI22_X1 U15499 ( .A1(n14164), .A2(n14095), .B1(n16337), .B2(n13865), .ZN(
        n13866) );
  OAI211_X1 U15500 ( .C1(n14167), .C2(n14080), .A(n13867), .B(n13866), .ZN(
        P3_U3208) );
  OAI21_X1 U15501 ( .B1(n13869), .B2(n13873), .A(n13868), .ZN(n13872) );
  AOI222_X1 U15502 ( .A1(n13979), .A2(n13872), .B1(n13871), .B2(n13987), .C1(
        n13870), .C2(n13986), .ZN(n14117) );
  OAI21_X1 U15503 ( .B1(n13875), .B2(n8991), .A(n13874), .ZN(n14119) );
  AOI22_X1 U15504 ( .A1(n13876), .A2(n16337), .B1(n14100), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13877) );
  OAI21_X1 U15505 ( .B1(n14171), .B2(n14046), .A(n13877), .ZN(n13878) );
  AOI21_X1 U15506 ( .B1(n14119), .B2(n14098), .A(n13878), .ZN(n13879) );
  OAI21_X1 U15507 ( .B1(n14117), .B2(n14100), .A(n13879), .ZN(P3_U3209) );
  XNOR2_X1 U15508 ( .A(n13880), .B(n13881), .ZN(n14123) );
  INV_X1 U15509 ( .A(n14123), .ZN(n13891) );
  OAI211_X1 U15510 ( .C1(n7934), .C2(n7935), .A(n13979), .B(n7938), .ZN(n13886) );
  AOI22_X1 U15511 ( .A1(n13884), .A2(n13986), .B1(n13987), .B2(n13914), .ZN(
        n13885) );
  NAND2_X1 U15512 ( .A1(n13886), .A2(n13885), .ZN(n14122) );
  AOI22_X1 U15513 ( .A1(n14100), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n16337), 
        .B2(n13887), .ZN(n13888) );
  OAI21_X1 U15514 ( .B1(n14175), .B2(n14046), .A(n13888), .ZN(n13889) );
  AOI21_X1 U15515 ( .B1(n14122), .B2(n16340), .A(n13889), .ZN(n13890) );
  OAI21_X1 U15516 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(P3_U3210) );
  XNOR2_X1 U15517 ( .A(n13893), .B(n13895), .ZN(n14178) );
  INV_X1 U15518 ( .A(n16428), .ZN(n13918) );
  XNOR2_X1 U15519 ( .A(n13894), .B(n13895), .ZN(n13896) );
  NAND2_X1 U15520 ( .A1(n13896), .A2(n13979), .ZN(n13900) );
  OAI22_X1 U15521 ( .A1(n13897), .A2(n14089), .B1(n13933), .B2(n14087), .ZN(
        n13898) );
  INV_X1 U15522 ( .A(n13898), .ZN(n13899) );
  OAI211_X1 U15523 ( .C1(n14178), .C2(n13918), .A(n13900), .B(n13899), .ZN(
        n14176) );
  MUX2_X1 U15524 ( .A(P3_REG2_REG_22__SCAN_IN), .B(n14176), .S(n16340), .Z(
        n13901) );
  INV_X1 U15525 ( .A(n13901), .ZN(n13905) );
  AOI22_X1 U15526 ( .A1(n13903), .A2(n14095), .B1(n16337), .B2(n13902), .ZN(
        n13904) );
  OAI211_X1 U15527 ( .C1(n14178), .C2(n14080), .A(n13905), .B(n13904), .ZN(
        P3_U3211) );
  NAND2_X1 U15528 ( .A1(n13927), .A2(n13906), .ZN(n13908) );
  NAND2_X1 U15529 ( .A1(n13908), .A2(n13907), .ZN(n13910) );
  NAND2_X1 U15530 ( .A1(n13910), .A2(n13909), .ZN(n14183) );
  XNOR2_X1 U15531 ( .A(n13912), .B(n13911), .ZN(n13913) );
  NAND2_X1 U15532 ( .A1(n13913), .A2(n13979), .ZN(n13917) );
  AOI22_X1 U15533 ( .A1(n13915), .A2(n13987), .B1(n13914), .B2(n13986), .ZN(
        n13916) );
  OAI211_X1 U15534 ( .C1(n13918), .C2(n14183), .A(n13917), .B(n13916), .ZN(
        n14181) );
  MUX2_X1 U15535 ( .A(P3_REG2_REG_21__SCAN_IN), .B(n14181), .S(n16340), .Z(
        n13919) );
  INV_X1 U15536 ( .A(n13919), .ZN(n13923) );
  AOI22_X1 U15537 ( .A1(n13921), .A2(n14095), .B1(n16337), .B2(n13920), .ZN(
        n13922) );
  OAI211_X1 U15538 ( .C1(n14183), .C2(n14080), .A(n13923), .B(n13922), .ZN(
        P3_U3212) );
  NAND2_X1 U15539 ( .A1(n13925), .A2(n13924), .ZN(n13926) );
  NAND2_X1 U15540 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  NAND2_X1 U15541 ( .A1(n13928), .A2(n16428), .ZN(n13937) );
  NAND2_X1 U15542 ( .A1(n13930), .A2(n13931), .ZN(n13932) );
  NAND3_X1 U15543 ( .A1(n13929), .A2(n13979), .A3(n13932), .ZN(n13936) );
  OAI22_X1 U15544 ( .A1(n13933), .A2(n14089), .B1(n13965), .B2(n14087), .ZN(
        n13934) );
  INV_X1 U15545 ( .A(n13934), .ZN(n13935) );
  NAND3_X1 U15546 ( .A1(n13937), .A2(n13936), .A3(n13935), .ZN(n14186) );
  MUX2_X1 U15547 ( .A(P3_REG2_REG_20__SCAN_IN), .B(n14186), .S(n16340), .Z(
        n13938) );
  INV_X1 U15548 ( .A(n13938), .ZN(n13942) );
  AOI22_X1 U15549 ( .A1(n13940), .A2(n14095), .B1(n16337), .B2(n13939), .ZN(
        n13941) );
  OAI211_X1 U15550 ( .C1(n14189), .C2(n14080), .A(n13942), .B(n13941), .ZN(
        P3_U3213) );
  XNOR2_X1 U15551 ( .A(n13943), .B(n13950), .ZN(n13944) );
  OAI222_X1 U15552 ( .A1(n14087), .A2(n13946), .B1(n14089), .B2(n13945), .C1(
        n14084), .C2(n13944), .ZN(n14133) );
  INV_X1 U15553 ( .A(n14133), .ZN(n13956) );
  NAND2_X1 U15554 ( .A1(n14029), .A2(n13947), .ZN(n14015) );
  NAND2_X1 U15555 ( .A1(n14015), .A2(n13948), .ZN(n13970) );
  NAND2_X1 U15556 ( .A1(n13970), .A2(n13949), .ZN(n13951) );
  XNOR2_X1 U15557 ( .A(n13951), .B(n13950), .ZN(n14134) );
  AOI22_X1 U15558 ( .A1(n14100), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n16337), 
        .B2(n13952), .ZN(n13953) );
  OAI21_X1 U15559 ( .B1(n14195), .B2(n14046), .A(n13953), .ZN(n13954) );
  AOI21_X1 U15560 ( .B1(n14134), .B2(n14098), .A(n13954), .ZN(n13955) );
  OAI21_X1 U15561 ( .B1(n13956), .B2(n14100), .A(n13955), .ZN(P3_U3214) );
  NAND2_X1 U15562 ( .A1(n14002), .A2(n13959), .ZN(n13982) );
  NAND2_X1 U15563 ( .A1(n13982), .A2(n13960), .ZN(n13980) );
  AOI21_X1 U15564 ( .B1(n13980), .B2(n13962), .A(n13961), .ZN(n13963) );
  NOR2_X1 U15565 ( .A1(n7561), .A2(n13963), .ZN(n13964) );
  OAI222_X1 U15566 ( .A1(n14089), .A2(n13965), .B1(n14087), .B2(n14012), .C1(
        n14084), .C2(n13964), .ZN(n14137) );
  INV_X1 U15567 ( .A(n14137), .ZN(n13978) );
  NAND2_X1 U15568 ( .A1(n14015), .A2(n13966), .ZN(n13968) );
  NAND2_X1 U15569 ( .A1(n13968), .A2(n13967), .ZN(n13973) );
  AND2_X1 U15570 ( .A1(n13970), .A2(n13969), .ZN(n13971) );
  OAI21_X1 U15571 ( .B1(n13973), .B2(n13972), .A(n13971), .ZN(n14138) );
  AOI22_X1 U15572 ( .A1(n14100), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n16337), 
        .B2(n13974), .ZN(n13975) );
  OAI21_X1 U15573 ( .B1(n14199), .B2(n14046), .A(n13975), .ZN(n13976) );
  AOI21_X1 U15574 ( .B1(n14138), .B2(n14098), .A(n13976), .ZN(n13977) );
  OAI21_X1 U15575 ( .B1(n13978), .B2(n14100), .A(n13977), .ZN(P3_U3215) );
  NAND2_X1 U15576 ( .A1(n13980), .A2(n13979), .ZN(n13991) );
  AND2_X1 U15577 ( .A1(n13982), .A2(n13981), .ZN(n14008) );
  AOI21_X1 U15578 ( .B1(n14008), .B2(n13984), .A(n13983), .ZN(n13990) );
  AOI22_X1 U15579 ( .A1(n13988), .A2(n13987), .B1(n13986), .B2(n13985), .ZN(
        n13989) );
  OAI21_X1 U15580 ( .B1(n13991), .B2(n13990), .A(n13989), .ZN(n14141) );
  INV_X1 U15581 ( .A(n14141), .ZN(n14000) );
  NAND2_X1 U15582 ( .A1(n14015), .A2(n14014), .ZN(n14013) );
  NAND2_X1 U15583 ( .A1(n14013), .A2(n13992), .ZN(n13995) );
  NAND2_X1 U15584 ( .A1(n13995), .A2(n13994), .ZN(n13993) );
  OAI21_X1 U15585 ( .B1(n13995), .B2(n13994), .A(n13993), .ZN(n14142) );
  AOI22_X1 U15586 ( .A1(n14100), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n16337), 
        .B2(n13996), .ZN(n13997) );
  OAI21_X1 U15587 ( .B1(n14203), .B2(n14046), .A(n13997), .ZN(n13998) );
  AOI21_X1 U15588 ( .B1(n14142), .B2(n14098), .A(n13998), .ZN(n13999) );
  OAI21_X1 U15589 ( .B1(n14000), .B2(n14100), .A(n13999), .ZN(P3_U3216) );
  NAND2_X1 U15590 ( .A1(n14002), .A2(n14001), .ZN(n14054) );
  NAND2_X1 U15591 ( .A1(n14054), .A2(n14003), .ZN(n14005) );
  AND2_X1 U15592 ( .A1(n14005), .A2(n14004), .ZN(n14007) );
  NAND2_X1 U15593 ( .A1(n14007), .A2(n14006), .ZN(n14010) );
  INV_X1 U15594 ( .A(n14008), .ZN(n14009) );
  AOI21_X1 U15595 ( .B1(n14014), .B2(n14010), .A(n14009), .ZN(n14011) );
  OAI222_X1 U15596 ( .A1(n14087), .A2(n14039), .B1(n14089), .B2(n14012), .C1(
        n14084), .C2(n14011), .ZN(n14145) );
  INV_X1 U15597 ( .A(n14145), .ZN(n14020) );
  OAI21_X1 U15598 ( .B1(n14015), .B2(n14014), .A(n14013), .ZN(n14146) );
  AOI22_X1 U15599 ( .A1(n14100), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n16337), 
        .B2(n14016), .ZN(n14017) );
  OAI21_X1 U15600 ( .B1(n14208), .B2(n14046), .A(n14017), .ZN(n14018) );
  AOI21_X1 U15601 ( .B1(n14146), .B2(n14098), .A(n14018), .ZN(n14019) );
  OAI21_X1 U15602 ( .B1(n14020), .B2(n14100), .A(n14019), .ZN(P3_U3217) );
  NAND2_X1 U15603 ( .A1(n14054), .A2(n14053), .ZN(n14022) );
  NAND2_X1 U15604 ( .A1(n14022), .A2(n14021), .ZN(n14037) );
  NAND2_X1 U15605 ( .A1(n14037), .A2(n14041), .ZN(n14024) );
  NAND2_X1 U15606 ( .A1(n14024), .A2(n14023), .ZN(n14026) );
  XNOR2_X1 U15607 ( .A(n14026), .B(n14025), .ZN(n14027) );
  OAI222_X1 U15608 ( .A1(n14089), .A2(n14028), .B1(n14087), .B2(n14055), .C1(
        n14027), .C2(n14084), .ZN(n16611) );
  INV_X1 U15609 ( .A(n16611), .ZN(n14035) );
  OAI21_X1 U15610 ( .B1(n14030), .B2(n8691), .A(n14029), .ZN(n16613) );
  AOI22_X1 U15611 ( .A1(n14100), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n16337), 
        .B2(n14031), .ZN(n14032) );
  OAI21_X1 U15612 ( .B1(n16610), .B2(n14046), .A(n14032), .ZN(n14033) );
  AOI21_X1 U15613 ( .B1(n16613), .B2(n14098), .A(n14033), .ZN(n14034) );
  OAI21_X1 U15614 ( .B1(n14035), .B2(n14100), .A(n14034), .ZN(P3_U3218) );
  INV_X1 U15615 ( .A(n14036), .ZN(n14069) );
  XNOR2_X1 U15616 ( .A(n14037), .B(n14041), .ZN(n14038) );
  OAI222_X1 U15617 ( .A1(n14089), .A2(n14039), .B1(n14087), .B2(n14069), .C1(
        n14038), .C2(n14084), .ZN(n16535) );
  INV_X1 U15618 ( .A(n16535), .ZN(n14049) );
  NAND3_X1 U15619 ( .A1(n14050), .A2(n14041), .A3(n14040), .ZN(n14042) );
  NAND2_X1 U15620 ( .A1(n14043), .A2(n14042), .ZN(n16537) );
  AOI22_X1 U15621 ( .A1(n14100), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n16337), 
        .B2(n14044), .ZN(n14045) );
  OAI21_X1 U15622 ( .B1(n16534), .B2(n14046), .A(n14045), .ZN(n14047) );
  AOI21_X1 U15623 ( .B1(n16537), .B2(n14098), .A(n14047), .ZN(n14048) );
  OAI21_X1 U15624 ( .B1(n14049), .B2(n14100), .A(n14048), .ZN(P3_U3219) );
  OAI21_X1 U15625 ( .B1(n14052), .B2(n14051), .A(n14050), .ZN(n16520) );
  INV_X1 U15626 ( .A(n16520), .ZN(n14064) );
  XNOR2_X1 U15627 ( .A(n14054), .B(n14053), .ZN(n14058) );
  OAI22_X1 U15628 ( .A1(n14088), .A2(n14087), .B1(n14055), .B2(n14089), .ZN(
        n14056) );
  AOI21_X1 U15629 ( .B1(n16520), .B2(n16428), .A(n14056), .ZN(n14057) );
  OAI21_X1 U15630 ( .B1(n14058), .B2(n14084), .A(n14057), .ZN(n16518) );
  NAND2_X1 U15631 ( .A1(n16518), .A2(n16340), .ZN(n14063) );
  OAI22_X1 U15632 ( .A1(n16340), .A2(n16170), .B1(n14059), .B2(n14073), .ZN(
        n14060) );
  AOI21_X1 U15633 ( .B1(n14061), .B2(n14095), .A(n14060), .ZN(n14062) );
  OAI211_X1 U15634 ( .C1(n14064), .C2(n14080), .A(n14063), .B(n14062), .ZN(
        P3_U3220) );
  OAI21_X1 U15635 ( .B1(n14066), .B2(n14068), .A(n14065), .ZN(n16505) );
  INV_X1 U15636 ( .A(n16505), .ZN(n14081) );
  XNOR2_X1 U15637 ( .A(n14067), .B(n14068), .ZN(n14072) );
  OAI22_X1 U15638 ( .A1(n8630), .A2(n14087), .B1(n14069), .B2(n14089), .ZN(
        n14070) );
  AOI21_X1 U15639 ( .B1(n16505), .B2(n16428), .A(n14070), .ZN(n14071) );
  OAI21_X1 U15640 ( .B1(n14072), .B2(n14084), .A(n14071), .ZN(n16503) );
  NAND2_X1 U15641 ( .A1(n16503), .A2(n16340), .ZN(n14079) );
  OAI22_X1 U15642 ( .A1(n16340), .A2(n14075), .B1(n14074), .B2(n14073), .ZN(
        n14076) );
  AOI21_X1 U15643 ( .B1(n14077), .B2(n14095), .A(n14076), .ZN(n14078) );
  OAI211_X1 U15644 ( .C1(n14081), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        P3_U3221) );
  XNOR2_X1 U15645 ( .A(n14082), .B(n14083), .ZN(n14085) );
  OAI222_X1 U15646 ( .A1(n14089), .A2(n14088), .B1(n14087), .B2(n14086), .C1(
        n14085), .C2(n14084), .ZN(n16484) );
  INV_X1 U15647 ( .A(n16484), .ZN(n14101) );
  OAI21_X1 U15648 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n16486) );
  AOI22_X1 U15649 ( .A1(n14095), .A2(n14094), .B1(n16337), .B2(n14093), .ZN(
        n14096) );
  OAI21_X1 U15650 ( .B1(n16126), .B2(n16340), .A(n14096), .ZN(n14097) );
  AOI21_X1 U15651 ( .B1(n16486), .B2(n14098), .A(n14097), .ZN(n14099) );
  OAI21_X1 U15652 ( .B1(n14101), .B2(n14100), .A(n14099), .ZN(P3_U3222) );
  NOR2_X1 U15653 ( .A1(n14150), .A2(n9060), .ZN(n14103) );
  AOI21_X1 U15654 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n9060), .A(n14103), .ZN(
        n14102) );
  OAI21_X1 U15655 ( .B1(n14152), .B2(n14149), .A(n14102), .ZN(P3_U3490) );
  AOI21_X1 U15656 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n9060), .A(n14103), .ZN(
        n14104) );
  OAI21_X1 U15657 ( .B1(n14155), .B2(n14149), .A(n14104), .ZN(P3_U3489) );
  AOI22_X1 U15658 ( .A1(n14106), .A2(n16614), .B1(n14105), .B2(n8915), .ZN(
        n14107) );
  NAND2_X1 U15659 ( .A1(n14108), .A2(n14107), .ZN(n14156) );
  MUX2_X1 U15660 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n14156), .S(n16615), .Z(
        P3_U3486) );
  AOI21_X1 U15661 ( .B1(n14110), .B2(n16614), .A(n14109), .ZN(n14157) );
  MUX2_X1 U15662 ( .A(n14111), .B(n14157), .S(n16615), .Z(n14112) );
  OAI21_X1 U15663 ( .B1(n14160), .B2(n14149), .A(n14112), .ZN(P3_U3485) );
  INV_X1 U15664 ( .A(n14113), .ZN(n14162) );
  MUX2_X1 U15665 ( .A(n14162), .B(n14114), .S(n9060), .Z(n14116) );
  NAND2_X1 U15666 ( .A1(n14164), .A2(n9056), .ZN(n14115) );
  OAI211_X1 U15667 ( .C1(n14167), .C2(n14130), .A(n14116), .B(n14115), .ZN(
        P3_U3484) );
  INV_X1 U15668 ( .A(n14117), .ZN(n14118) );
  AOI21_X1 U15669 ( .B1(n16614), .B2(n14119), .A(n14118), .ZN(n14168) );
  MUX2_X1 U15670 ( .A(n14120), .B(n14168), .S(n16615), .Z(n14121) );
  OAI21_X1 U15671 ( .B1(n14171), .B2(n14149), .A(n14121), .ZN(P3_U3483) );
  INV_X1 U15672 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14124) );
  AOI21_X1 U15673 ( .B1(n14123), .B2(n16614), .A(n14122), .ZN(n14172) );
  MUX2_X1 U15674 ( .A(n14124), .B(n14172), .S(n16615), .Z(n14125) );
  OAI21_X1 U15675 ( .B1(n14175), .B2(n14149), .A(n14125), .ZN(P3_U3482) );
  MUX2_X1 U15676 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n14176), .S(n16615), .Z(
        n14127) );
  OAI22_X1 U15677 ( .A1(n14178), .A2(n14130), .B1(n14177), .B2(n14149), .ZN(
        n14126) );
  OR2_X1 U15678 ( .A1(n14127), .A2(n14126), .ZN(P3_U3481) );
  MUX2_X1 U15679 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n14181), .S(n16615), .Z(
        n14129) );
  OAI22_X1 U15680 ( .A1(n14183), .A2(n14130), .B1(n14182), .B2(n14149), .ZN(
        n14128) );
  OR2_X1 U15681 ( .A1(n14129), .A2(n14128), .ZN(P3_U3480) );
  MUX2_X1 U15682 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n14186), .S(n16615), .Z(
        n14132) );
  OAI22_X1 U15683 ( .A1(n14189), .A2(n14130), .B1(n14187), .B2(n14149), .ZN(
        n14131) );
  OR2_X1 U15684 ( .A1(n14132), .A2(n14131), .ZN(P3_U3479) );
  INV_X1 U15685 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14135) );
  AOI21_X1 U15686 ( .B1(n14134), .B2(n16614), .A(n14133), .ZN(n14192) );
  MUX2_X1 U15687 ( .A(n14135), .B(n14192), .S(n16615), .Z(n14136) );
  OAI21_X1 U15688 ( .B1(n14195), .B2(n14149), .A(n14136), .ZN(P3_U3478) );
  AOI21_X1 U15689 ( .B1(n16614), .B2(n14138), .A(n14137), .ZN(n14196) );
  MUX2_X1 U15690 ( .A(n14139), .B(n14196), .S(n16615), .Z(n14140) );
  OAI21_X1 U15691 ( .B1(n14199), .B2(n14149), .A(n14140), .ZN(P3_U3477) );
  INV_X1 U15692 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14143) );
  AOI21_X1 U15693 ( .B1(n16614), .B2(n14142), .A(n14141), .ZN(n14200) );
  MUX2_X1 U15694 ( .A(n14143), .B(n14200), .S(n16615), .Z(n14144) );
  OAI21_X1 U15695 ( .B1(n14203), .B2(n14149), .A(n14144), .ZN(P3_U3476) );
  AOI21_X1 U15696 ( .B1(n16614), .B2(n14146), .A(n14145), .ZN(n14204) );
  MUX2_X1 U15697 ( .A(n14147), .B(n14204), .S(n16615), .Z(n14148) );
  OAI21_X1 U15698 ( .B1(n14208), .B2(n14149), .A(n14148), .ZN(P3_U3475) );
  NOR2_X1 U15699 ( .A1(n14150), .A2(n9044), .ZN(n14153) );
  AOI21_X1 U15700 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n9044), .A(n14153), .ZN(
        n14151) );
  OAI21_X1 U15701 ( .B1(n14152), .B2(n14207), .A(n14151), .ZN(P3_U3458) );
  AOI21_X1 U15702 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(n9044), .A(n14153), .ZN(
        n14154) );
  OAI21_X1 U15703 ( .B1(n14155), .B2(n14207), .A(n14154), .ZN(P3_U3457) );
  MUX2_X1 U15704 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n14156), .S(n16618), .Z(
        P3_U3454) );
  INV_X1 U15705 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14158) );
  MUX2_X1 U15706 ( .A(n14158), .B(n14157), .S(n16618), .Z(n14159) );
  OAI21_X1 U15707 ( .B1(n14160), .B2(n14207), .A(n14159), .ZN(P3_U3453) );
  INV_X1 U15708 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14161) );
  MUX2_X1 U15709 ( .A(n14162), .B(n14161), .S(n9044), .Z(n14166) );
  NAND2_X1 U15710 ( .A1(n14164), .A2(n14163), .ZN(n14165) );
  OAI211_X1 U15711 ( .C1(n14167), .C2(n14188), .A(n14166), .B(n14165), .ZN(
        P3_U3452) );
  INV_X1 U15712 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14169) );
  MUX2_X1 U15713 ( .A(n14169), .B(n14168), .S(n16618), .Z(n14170) );
  OAI21_X1 U15714 ( .B1(n14171), .B2(n14207), .A(n14170), .ZN(P3_U3451) );
  INV_X1 U15715 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14173) );
  MUX2_X1 U15716 ( .A(n14173), .B(n14172), .S(n16618), .Z(n14174) );
  OAI21_X1 U15717 ( .B1(n14175), .B2(n14207), .A(n14174), .ZN(P3_U3450) );
  MUX2_X1 U15718 ( .A(n14176), .B(P3_REG0_REG_22__SCAN_IN), .S(n9044), .Z(
        n14180) );
  OAI22_X1 U15719 ( .A1(n14178), .A2(n14188), .B1(n14177), .B2(n14207), .ZN(
        n14179) );
  OR2_X1 U15720 ( .A1(n14180), .A2(n14179), .ZN(P3_U3449) );
  MUX2_X1 U15721 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n14181), .S(n16618), .Z(
        n14185) );
  OAI22_X1 U15722 ( .A1(n14183), .A2(n14188), .B1(n14182), .B2(n14207), .ZN(
        n14184) );
  OR2_X1 U15723 ( .A1(n14185), .A2(n14184), .ZN(P3_U3448) );
  MUX2_X1 U15724 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n14186), .S(n16618), .Z(
        n14191) );
  OAI22_X1 U15725 ( .A1(n14189), .A2(n14188), .B1(n14187), .B2(n14207), .ZN(
        n14190) );
  OR2_X1 U15726 ( .A1(n14191), .A2(n14190), .ZN(P3_U3447) );
  INV_X1 U15727 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14193) );
  MUX2_X1 U15728 ( .A(n14193), .B(n14192), .S(n16618), .Z(n14194) );
  OAI21_X1 U15729 ( .B1(n14195), .B2(n14207), .A(n14194), .ZN(P3_U3446) );
  INV_X1 U15730 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n14197) );
  MUX2_X1 U15731 ( .A(n14197), .B(n14196), .S(n16618), .Z(n14198) );
  OAI21_X1 U15732 ( .B1(n14199), .B2(n14207), .A(n14198), .ZN(P3_U3444) );
  INV_X1 U15733 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14201) );
  MUX2_X1 U15734 ( .A(n14201), .B(n14200), .S(n16618), .Z(n14202) );
  OAI21_X1 U15735 ( .B1(n14203), .B2(n14207), .A(n14202), .ZN(P3_U3441) );
  INV_X1 U15736 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14205) );
  MUX2_X1 U15737 ( .A(n14205), .B(n14204), .S(n16618), .Z(n14206) );
  OAI21_X1 U15738 ( .B1(n14208), .B2(n14207), .A(n14206), .ZN(P3_U3438) );
  MUX2_X1 U15739 ( .A(P3_D_REG_1__SCAN_IN), .B(n14209), .S(n14210), .Z(
        P3_U3377) );
  MUX2_X1 U15740 ( .A(P3_D_REG_0__SCAN_IN), .B(n14211), .S(n14210), .Z(
        P3_U3376) );
  NAND2_X1 U15741 ( .A1(n14213), .A2(n14212), .ZN(n14217) );
  NAND4_X1 U15742 ( .A1(n8414), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n14215), .ZN(n14216) );
  OAI211_X1 U15743 ( .C1(n14218), .C2(n14223), .A(n14217), .B(n14216), .ZN(
        P3_U3264) );
  INV_X1 U15744 ( .A(n14219), .ZN(n14220) );
  OAI222_X1 U15745 ( .A1(n14223), .A2(n15460), .B1(P3_U3151), .B2(n14222), 
        .C1(n14221), .C2(n14220), .ZN(P3_U3266) );
  MUX2_X1 U15746 ( .A(n14224), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  NOR2_X1 U15747 ( .A1(n14512), .A2(n12771), .ZN(n14272) );
  XOR2_X1 U15748 ( .A(n11490), .B(n14551), .Z(n14250) );
  INV_X1 U15749 ( .A(n14225), .ZN(n14228) );
  INV_X1 U15750 ( .A(n14226), .ZN(n14227) );
  NAND2_X1 U15751 ( .A1(n14228), .A2(n14227), .ZN(n14229) );
  XNOR2_X1 U15752 ( .A(n14594), .B(n14244), .ZN(n14232) );
  NAND2_X1 U15753 ( .A1(n14579), .A2(n11533), .ZN(n14233) );
  NAND2_X1 U15754 ( .A1(n14232), .A2(n14233), .ZN(n14237) );
  INV_X1 U15755 ( .A(n14232), .ZN(n14235) );
  INV_X1 U15756 ( .A(n14233), .ZN(n14234) );
  NAND2_X1 U15757 ( .A1(n14235), .A2(n14234), .ZN(n14236) );
  NAND2_X1 U15758 ( .A1(n14237), .A2(n14236), .ZN(n14278) );
  XNOR2_X1 U15759 ( .A(n14698), .B(n14244), .ZN(n14238) );
  NAND2_X1 U15760 ( .A1(n14371), .A2(n11533), .ZN(n14239) );
  NAND2_X1 U15761 ( .A1(n14238), .A2(n14239), .ZN(n14243) );
  INV_X1 U15762 ( .A(n14238), .ZN(n14241) );
  INV_X1 U15763 ( .A(n14239), .ZN(n14240) );
  NAND2_X1 U15764 ( .A1(n14241), .A2(n14240), .ZN(n14242) );
  AND2_X1 U15765 ( .A1(n14243), .A2(n14242), .ZN(n14330) );
  NAND2_X1 U15766 ( .A1(n14328), .A2(n14243), .ZN(n14302) );
  XNOR2_X1 U15767 ( .A(n14566), .B(n14244), .ZN(n14245) );
  NAND2_X1 U15768 ( .A1(n14576), .A2(n11533), .ZN(n14246) );
  XNOR2_X1 U15769 ( .A(n14245), .B(n14246), .ZN(n14303) );
  INV_X1 U15770 ( .A(n14245), .ZN(n14248) );
  INV_X1 U15771 ( .A(n14246), .ZN(n14247) );
  NAND2_X1 U15772 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  NAND2_X1 U15773 ( .A1(n14370), .A2(n11533), .ZN(n14340) );
  INV_X1 U15774 ( .A(n14250), .ZN(n14251) );
  OR2_X1 U15775 ( .A1(n14252), .A2(n14251), .ZN(n14253) );
  NAND2_X1 U15776 ( .A1(n14339), .A2(n14253), .ZN(n14254) );
  XNOR2_X1 U15777 ( .A(n14527), .B(n11490), .ZN(n14255) );
  XNOR2_X1 U15778 ( .A(n14254), .B(n14255), .ZN(n14271) );
  INV_X1 U15779 ( .A(n14254), .ZN(n14256) );
  NAND2_X1 U15780 ( .A1(n14492), .A2(n11533), .ZN(n14258) );
  XNOR2_X1 U15781 ( .A(n14676), .B(n11490), .ZN(n14257) );
  XOR2_X1 U15782 ( .A(n14258), .B(n14257), .Z(n14319) );
  XNOR2_X1 U15783 ( .A(n14498), .B(n11490), .ZN(n14260) );
  NAND2_X1 U15784 ( .A1(n14368), .A2(n11533), .ZN(n14259) );
  XNOR2_X1 U15785 ( .A(n14260), .B(n14259), .ZN(n14311) );
  INV_X1 U15786 ( .A(n14259), .ZN(n14261) );
  AND2_X1 U15787 ( .A1(n14493), .A2(n11533), .ZN(n14263) );
  XNOR2_X1 U15788 ( .A(n14480), .B(n11490), .ZN(n14262) );
  NOR2_X1 U15789 ( .A1(n14262), .A2(n14263), .ZN(n14264) );
  AOI21_X1 U15790 ( .B1(n14263), .B2(n14262), .A(n14264), .ZN(n14351) );
  INV_X1 U15791 ( .A(n14264), .ZN(n14265) );
  XNOR2_X1 U15792 ( .A(n14467), .B(n11490), .ZN(n14286) );
  NOR2_X1 U15793 ( .A1(n14266), .A2(n12771), .ZN(n14287) );
  XNOR2_X1 U15794 ( .A(n14286), .B(n14287), .ZN(n14290) );
  XNOR2_X1 U15795 ( .A(n14291), .B(n14290), .ZN(n14270) );
  AOI22_X1 U15796 ( .A1(n14366), .A2(n14575), .B1(n14578), .B2(n14493), .ZN(
        n14461) );
  AOI22_X1 U15797 ( .A1(n14468), .A2(n14332), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14267) );
  OAI21_X1 U15798 ( .B1(n14461), .B2(n14297), .A(n14267), .ZN(n14268) );
  AOI21_X1 U15799 ( .B1(n14467), .B2(n14324), .A(n14268), .ZN(n14269) );
  OAI21_X1 U15800 ( .B1(n14270), .B2(n14326), .A(n14269), .ZN(P2_U3186) );
  XNOR2_X1 U15801 ( .A(n14271), .B(n14272), .ZN(n14277) );
  OAI22_X1 U15802 ( .A1(n14535), .A2(n14320), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14273), .ZN(n14275) );
  OAI22_X1 U15803 ( .A1(n14534), .A2(n14281), .B1(n14355), .B2(n14529), .ZN(
        n14274) );
  AOI211_X1 U15804 ( .C1(n14527), .C2(n14324), .A(n14275), .B(n14274), .ZN(
        n14276) );
  OAI21_X1 U15805 ( .B1(n14277), .B2(n14326), .A(n14276), .ZN(P2_U3188) );
  AOI21_X1 U15806 ( .B1(n14279), .B2(n14278), .A(n7563), .ZN(n14285) );
  OAI21_X1 U15807 ( .B1(n14320), .B2(n14605), .A(n14280), .ZN(n14283) );
  OAI22_X1 U15808 ( .A1(n14281), .A2(n14603), .B1(n14595), .B2(n14355), .ZN(
        n14282) );
  AOI211_X1 U15809 ( .C1(n14594), .C2(n14324), .A(n14283), .B(n14282), .ZN(
        n14284) );
  OAI21_X1 U15810 ( .B1(n14285), .B2(n14326), .A(n14284), .ZN(P2_U3191) );
  INV_X1 U15811 ( .A(n14286), .ZN(n14289) );
  INV_X1 U15812 ( .A(n14287), .ZN(n14288) );
  NAND2_X1 U15813 ( .A1(n14366), .A2(n11533), .ZN(n14292) );
  XNOR2_X1 U15814 ( .A(n14292), .B(n11490), .ZN(n14293) );
  XNOR2_X1 U15815 ( .A(n14453), .B(n14293), .ZN(n14294) );
  INV_X1 U15816 ( .A(n14451), .ZN(n14295) );
  AOI22_X1 U15817 ( .A1(n14295), .A2(n14332), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14296) );
  OAI21_X1 U15818 ( .B1(n14298), .B2(n14297), .A(n14296), .ZN(n14299) );
  AOI21_X1 U15819 ( .B1(n14453), .B2(n14324), .A(n14299), .ZN(n14300) );
  OAI21_X1 U15820 ( .B1(n14301), .B2(n14326), .A(n14300), .ZN(P2_U3192) );
  XNOR2_X1 U15821 ( .A(n14302), .B(n14303), .ZN(n14309) );
  NOR2_X1 U15822 ( .A1(n14605), .A2(n14602), .ZN(n14304) );
  AOI21_X1 U15823 ( .B1(n14370), .B2(n14575), .A(n14304), .ZN(n14560) );
  INV_X1 U15824 ( .A(n14560), .ZN(n14305) );
  AOI22_X1 U15825 ( .A1(n14305), .A2(n14358), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14306) );
  OAI21_X1 U15826 ( .B1(n14564), .B2(n14355), .A(n14306), .ZN(n14307) );
  AOI21_X1 U15827 ( .B1(n14566), .B2(n14324), .A(n14307), .ZN(n14308) );
  OAI21_X1 U15828 ( .B1(n14309), .B2(n14326), .A(n14308), .ZN(P2_U3195) );
  XNOR2_X1 U15829 ( .A(n14310), .B(n14311), .ZN(n14317) );
  NOR2_X1 U15830 ( .A1(n14312), .A2(n14320), .ZN(n14315) );
  AOI22_X1 U15831 ( .A1(n14492), .A2(n14333), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14313) );
  OAI21_X1 U15832 ( .B1(n14500), .B2(n14355), .A(n14313), .ZN(n14314) );
  AOI211_X1 U15833 ( .C1(n14498), .C2(n14324), .A(n14315), .B(n14314), .ZN(
        n14316) );
  OAI21_X1 U15834 ( .B1(n14317), .B2(n14326), .A(n14316), .ZN(P2_U3197) );
  XNOR2_X1 U15835 ( .A(n14318), .B(n14319), .ZN(n14327) );
  NOR2_X1 U15836 ( .A1(n14513), .A2(n14320), .ZN(n14323) );
  AOI22_X1 U15837 ( .A1(n14369), .A2(n14333), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14321) );
  OAI21_X1 U15838 ( .B1(n14517), .B2(n14355), .A(n14321), .ZN(n14322) );
  OAI21_X1 U15839 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(P2_U3201) );
  OAI21_X1 U15840 ( .B1(n14330), .B2(n14329), .A(n14328), .ZN(n14337) );
  AOI22_X1 U15841 ( .A1(n14331), .A2(n14576), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14335) );
  AOI22_X1 U15842 ( .A1(n14333), .A2(n14579), .B1(n14584), .B2(n14332), .ZN(
        n14334) );
  OAI211_X1 U15843 ( .C1(n14587), .C2(n14362), .A(n14335), .B(n14334), .ZN(
        n14336) );
  AOI21_X1 U15844 ( .B1(n14337), .B2(n14352), .A(n14336), .ZN(n14338) );
  INV_X1 U15845 ( .A(n14338), .ZN(P2_U3205) );
  OAI21_X1 U15846 ( .B1(n14341), .B2(n14340), .A(n14339), .ZN(n14342) );
  NAND2_X1 U15847 ( .A1(n14342), .A2(n14352), .ZN(n14348) );
  OAI22_X1 U15848 ( .A1(n14512), .A2(n14604), .B1(n14343), .B2(n14602), .ZN(
        n14544) );
  INV_X1 U15849 ( .A(n14552), .ZN(n14345) );
  OAI22_X1 U15850 ( .A1(n14345), .A2(n14355), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14344), .ZN(n14346) );
  AOI21_X1 U15851 ( .B1(n14544), .B2(n14358), .A(n14346), .ZN(n14347) );
  OAI211_X1 U15852 ( .C1(n7856), .C2(n14362), .A(n14348), .B(n14347), .ZN(
        P2_U3207) );
  OAI21_X1 U15853 ( .B1(n14351), .B2(n14350), .A(n14349), .ZN(n14353) );
  NAND2_X1 U15854 ( .A1(n14353), .A2(n14352), .ZN(n14361) );
  AOI22_X1 U15855 ( .A1(n14367), .A2(n14575), .B1(n14578), .B2(n14368), .ZN(
        n14475) );
  INV_X1 U15856 ( .A(n14475), .ZN(n14359) );
  INV_X1 U15857 ( .A(n14481), .ZN(n14356) );
  OAI22_X1 U15858 ( .A1(n14356), .A2(n14355), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14354), .ZN(n14357) );
  AOI21_X1 U15859 ( .B1(n14359), .B2(n14358), .A(n14357), .ZN(n14360) );
  OAI211_X1 U15860 ( .C1(n14744), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        P2_U3212) );
  MUX2_X1 U15861 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14363), .S(P2_U3947), .Z(
        P2_U3562) );
  MUX2_X1 U15862 ( .A(n14364), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14385), .Z(
        P2_U3561) );
  MUX2_X1 U15863 ( .A(n14365), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14385), .Z(
        P2_U3560) );
  MUX2_X1 U15864 ( .A(n14366), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14385), .Z(
        P2_U3559) );
  MUX2_X1 U15865 ( .A(n14367), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14385), .Z(
        P2_U3558) );
  MUX2_X1 U15866 ( .A(n14493), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14385), .Z(
        P2_U3557) );
  MUX2_X1 U15867 ( .A(n14368), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14385), .Z(
        P2_U3556) );
  MUX2_X1 U15868 ( .A(n14492), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14385), .Z(
        P2_U3555) );
  MUX2_X1 U15869 ( .A(n14369), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14385), .Z(
        P2_U3554) );
  MUX2_X1 U15870 ( .A(n14370), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14385), .Z(
        P2_U3553) );
  MUX2_X1 U15871 ( .A(n14576), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14385), .Z(
        P2_U3552) );
  MUX2_X1 U15872 ( .A(n14371), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14385), .Z(
        P2_U3551) );
  MUX2_X1 U15873 ( .A(n14579), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14385), .Z(
        P2_U3550) );
  MUX2_X1 U15874 ( .A(n14372), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14385), .Z(
        P2_U3549) );
  MUX2_X1 U15875 ( .A(n14373), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14385), .Z(
        P2_U3548) );
  MUX2_X1 U15876 ( .A(n14374), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14385), .Z(
        P2_U3547) );
  MUX2_X1 U15877 ( .A(n14375), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14385), .Z(
        P2_U3546) );
  MUX2_X1 U15878 ( .A(n14376), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14385), .Z(
        P2_U3545) );
  MUX2_X1 U15879 ( .A(n14377), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14385), .Z(
        P2_U3544) );
  MUX2_X1 U15880 ( .A(n14378), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14385), .Z(
        P2_U3542) );
  MUX2_X1 U15881 ( .A(n14379), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14385), .Z(
        P2_U3540) );
  MUX2_X1 U15882 ( .A(n14380), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14385), .Z(
        P2_U3539) );
  MUX2_X1 U15883 ( .A(n14381), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14385), .Z(
        P2_U3537) );
  MUX2_X1 U15884 ( .A(n14382), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14385), .Z(
        P2_U3536) );
  MUX2_X1 U15885 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n14383), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15886 ( .A(n14384), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14385), .Z(
        P2_U3534) );
  MUX2_X1 U15887 ( .A(n14386), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14385), .Z(
        P2_U3533) );
  MUX2_X1 U15888 ( .A(n7435), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14385), .Z(
        P2_U3532) );
  MUX2_X1 U15889 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n14387), .S(P2_U3947), .Z(
        P2_U3531) );
  INV_X1 U15890 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14389) );
  INV_X1 U15891 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14388) );
  OAI22_X1 U15892 ( .A1(n15928), .A2(n14389), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14388), .ZN(n14390) );
  AOI21_X1 U15893 ( .B1(n14391), .B2(n15922), .A(n14390), .ZN(n14400) );
  OAI211_X1 U15894 ( .C1(n14394), .C2(n14393), .A(n15924), .B(n14392), .ZN(
        n14399) );
  OR3_X1 U15895 ( .A1(n15850), .A2(n14396), .A3(n14395), .ZN(n14397) );
  NAND3_X1 U15896 ( .A1(n15920), .A2(n14410), .A3(n14397), .ZN(n14398) );
  NAND3_X1 U15897 ( .A1(n14400), .A2(n14399), .A3(n14398), .ZN(P2_U3217) );
  INV_X1 U15898 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14402) );
  OAI21_X1 U15899 ( .B1(n15928), .B2(n14402), .A(n14401), .ZN(n14403) );
  AOI21_X1 U15900 ( .B1(n14404), .B2(n15922), .A(n14403), .ZN(n14415) );
  OAI211_X1 U15901 ( .C1(n14407), .C2(n14406), .A(n15924), .B(n14405), .ZN(
        n14414) );
  INV_X1 U15902 ( .A(n14430), .ZN(n14412) );
  NAND3_X1 U15903 ( .A1(n14410), .A2(n14409), .A3(n14408), .ZN(n14411) );
  NAND3_X1 U15904 ( .A1(n14412), .A2(n15920), .A3(n14411), .ZN(n14413) );
  NAND3_X1 U15905 ( .A1(n14415), .A2(n14414), .A3(n14413), .ZN(P2_U3218) );
  INV_X1 U15906 ( .A(n14416), .ZN(n14420) );
  NOR2_X1 U15907 ( .A1(n14418), .A2(n14417), .ZN(n14419) );
  AOI211_X1 U15908 ( .C1(n15880), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n14420), .B(
        n14419), .ZN(n14433) );
  OAI211_X1 U15909 ( .C1(n14423), .C2(n14422), .A(n15924), .B(n14421), .ZN(
        n14432) );
  MUX2_X1 U15910 ( .A(n11295), .B(P2_REG1_REG_5__SCAN_IN), .S(n14424), .Z(
        n14427) );
  INV_X1 U15911 ( .A(n14425), .ZN(n14426) );
  NAND2_X1 U15912 ( .A1(n14427), .A2(n14426), .ZN(n14429) );
  OAI211_X1 U15913 ( .C1(n14430), .C2(n14429), .A(n14428), .B(n15920), .ZN(
        n14431) );
  NAND3_X1 U15914 ( .A1(n14433), .A2(n14432), .A3(n14431), .ZN(P2_U3219) );
  NAND2_X1 U15915 ( .A1(n14443), .A2(n14732), .ZN(n14442) );
  XNOR2_X1 U15916 ( .A(n14442), .B(n14728), .ZN(n14435) );
  NAND2_X1 U15917 ( .A1(n14435), .A2(n12771), .ZN(n14651) );
  NOR2_X1 U15918 ( .A1(n14610), .A2(n14436), .ZN(n14440) );
  INV_X1 U15919 ( .A(n14437), .ZN(n14439) );
  OR2_X1 U15920 ( .A1(n14439), .A2(n14438), .ZN(n14654) );
  NOR2_X1 U15921 ( .A1(n16598), .A2(n14654), .ZN(n14445) );
  AOI211_X1 U15922 ( .C1(n14434), .C2(n16599), .A(n14440), .B(n14445), .ZN(
        n14441) );
  OAI21_X1 U15923 ( .B1(n14651), .B2(n16601), .A(n14441), .ZN(P2_U3234) );
  OAI211_X1 U15924 ( .C1(n14443), .C2(n14732), .A(n12771), .B(n14442), .ZN(
        n14655) );
  NOR2_X1 U15925 ( .A1(n14610), .A2(n14444), .ZN(n14446) );
  AOI211_X1 U15926 ( .C1(n14447), .C2(n16599), .A(n14446), .B(n14445), .ZN(
        n14448) );
  OAI21_X1 U15927 ( .B1(n14655), .B2(n16601), .A(n14448), .ZN(P2_U3235) );
  NAND2_X1 U15928 ( .A1(n14449), .A2(n14610), .ZN(n14459) );
  OAI22_X1 U15929 ( .A1(n14451), .A2(n14640), .B1(n14450), .B2(n14610), .ZN(
        n14452) );
  AOI21_X1 U15930 ( .B1(n14453), .B2(n16599), .A(n14452), .ZN(n14458) );
  NAND2_X1 U15931 ( .A1(n14454), .A2(n16604), .ZN(n14457) );
  NAND2_X1 U15932 ( .A1(n14455), .A2(n14645), .ZN(n14456) );
  NAND4_X1 U15933 ( .A1(n14459), .A2(n14458), .A3(n14457), .A4(n14456), .ZN(
        P2_U3237) );
  OAI21_X1 U15934 ( .B1(n14462), .B2(n14510), .A(n14461), .ZN(n14660) );
  INV_X1 U15935 ( .A(n14660), .ZN(n14473) );
  XNOR2_X1 U15936 ( .A(n14464), .B(n14463), .ZN(n14662) );
  INV_X1 U15937 ( .A(n14465), .ZN(n14466) );
  AOI211_X1 U15938 ( .C1(n14467), .C2(n7861), .A(n11533), .B(n14466), .ZN(
        n14661) );
  NAND2_X1 U15939 ( .A1(n14661), .A2(n14645), .ZN(n14470) );
  AOI22_X1 U15940 ( .A1(n14468), .A2(n16596), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n16598), .ZN(n14469) );
  OAI211_X1 U15941 ( .C1(n14740), .C2(n14621), .A(n14470), .B(n14469), .ZN(
        n14471) );
  AOI21_X1 U15942 ( .B1(n14662), .B2(n16604), .A(n14471), .ZN(n14472) );
  OAI21_X1 U15943 ( .B1(n14473), .B2(n16598), .A(n14472), .ZN(P2_U3238) );
  XNOR2_X1 U15944 ( .A(n14474), .B(n14477), .ZN(n14476) );
  OAI21_X1 U15945 ( .B1(n14476), .B2(n14510), .A(n14475), .ZN(n14664) );
  INV_X1 U15946 ( .A(n14664), .ZN(n14486) );
  XOR2_X1 U15947 ( .A(n14478), .B(n14477), .Z(n14666) );
  AOI211_X1 U15948 ( .C1(n14480), .C2(n14496), .A(n11533), .B(n14479), .ZN(
        n14665) );
  NAND2_X1 U15949 ( .A1(n14665), .A2(n14645), .ZN(n14483) );
  AOI22_X1 U15950 ( .A1(n14481), .A2(n16596), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n16598), .ZN(n14482) );
  OAI211_X1 U15951 ( .C1(n14744), .C2(n14621), .A(n14483), .B(n14482), .ZN(
        n14484) );
  AOI21_X1 U15952 ( .B1(n14666), .B2(n16604), .A(n14484), .ZN(n14485) );
  OAI21_X1 U15953 ( .B1(n14486), .B2(n16598), .A(n14485), .ZN(P2_U3239) );
  AOI21_X1 U15954 ( .B1(n14490), .B2(n14488), .A(n14487), .ZN(n14671) );
  INV_X1 U15955 ( .A(n14671), .ZN(n14505) );
  OAI211_X1 U15956 ( .C1(n14491), .C2(n14490), .A(n14489), .B(n16584), .ZN(
        n14495) );
  AOI22_X1 U15957 ( .A1(n14493), .A2(n14575), .B1(n14578), .B2(n14492), .ZN(
        n14494) );
  NAND2_X1 U15958 ( .A1(n14495), .A2(n14494), .ZN(n14669) );
  NAND2_X1 U15959 ( .A1(n14669), .A2(n14610), .ZN(n14504) );
  INV_X1 U15960 ( .A(n14496), .ZN(n14497) );
  AOI211_X1 U15961 ( .C1(n14498), .C2(n14514), .A(n11533), .B(n14497), .ZN(
        n14670) );
  NOR2_X1 U15962 ( .A1(n10368), .A2(n14621), .ZN(n14502) );
  OAI22_X1 U15963 ( .A1(n14500), .A2(n14640), .B1(n14499), .B2(n14610), .ZN(
        n14501) );
  AOI211_X1 U15964 ( .C1(n14670), .C2(n14645), .A(n14502), .B(n14501), .ZN(
        n14503) );
  OAI211_X1 U15965 ( .C1(n14648), .C2(n14505), .A(n14504), .B(n14503), .ZN(
        P2_U3240) );
  XNOR2_X1 U15966 ( .A(n14509), .B(n14506), .ZN(n14678) );
  AOI21_X1 U15967 ( .B1(n14509), .B2(n14508), .A(n14507), .ZN(n14511) );
  OAI222_X1 U15968 ( .A1(n14604), .A2(n14513), .B1(n14602), .B2(n14512), .C1(
        n14511), .C2(n14510), .ZN(n14674) );
  AOI21_X1 U15969 ( .B1(n14676), .B2(n14524), .A(n11533), .ZN(n14515) );
  AND2_X1 U15970 ( .A1(n14515), .A2(n14514), .ZN(n14675) );
  NAND2_X1 U15971 ( .A1(n14675), .A2(n14645), .ZN(n14520) );
  OAI22_X1 U15972 ( .A1(n14517), .A2(n14640), .B1(n14516), .B2(n14610), .ZN(
        n14518) );
  AOI21_X1 U15973 ( .B1(n14676), .B2(n16599), .A(n14518), .ZN(n14519) );
  NAND2_X1 U15974 ( .A1(n14520), .A2(n14519), .ZN(n14521) );
  AOI21_X1 U15975 ( .B1(n14674), .B2(n14610), .A(n14521), .ZN(n14522) );
  OAI21_X1 U15976 ( .B1(n14648), .B2(n14678), .A(n14522), .ZN(P2_U3241) );
  XNOR2_X1 U15977 ( .A(n14523), .B(n14532), .ZN(n14679) );
  INV_X1 U15978 ( .A(n14550), .ZN(n14526) );
  INV_X1 U15979 ( .A(n14524), .ZN(n14525) );
  AOI211_X1 U15980 ( .C1(n14527), .C2(n14526), .A(n11533), .B(n14525), .ZN(
        n14680) );
  NOR2_X1 U15981 ( .A1(n14752), .A2(n14621), .ZN(n14531) );
  OAI22_X1 U15982 ( .A1(n14529), .A2(n14640), .B1(n14528), .B2(n14610), .ZN(
        n14530) );
  AOI211_X1 U15983 ( .C1(n14680), .C2(n14645), .A(n14531), .B(n14530), .ZN(
        n14540) );
  XNOR2_X1 U15984 ( .A(n14533), .B(n14532), .ZN(n14537) );
  OAI22_X1 U15985 ( .A1(n14535), .A2(n14604), .B1(n14534), .B2(n14602), .ZN(
        n14536) );
  AOI21_X1 U15986 ( .B1(n14537), .B2(n16584), .A(n14536), .ZN(n14538) );
  OAI21_X1 U15987 ( .B1(n14679), .B2(n14609), .A(n14538), .ZN(n14681) );
  NAND2_X1 U15988 ( .A1(n14681), .A2(n14610), .ZN(n14539) );
  OAI211_X1 U15989 ( .C1(n14679), .C2(n14613), .A(n14540), .B(n14539), .ZN(
        P2_U3242) );
  OAI211_X1 U15990 ( .C1(n14549), .C2(n14542), .A(n14541), .B(n16584), .ZN(
        n14543) );
  INV_X1 U15991 ( .A(n14543), .ZN(n14545) );
  INV_X1 U15992 ( .A(n14686), .ZN(n14557) );
  INV_X1 U15993 ( .A(n14546), .ZN(n14547) );
  AOI21_X1 U15994 ( .B1(n14549), .B2(n14548), .A(n14547), .ZN(n14687) );
  AOI211_X1 U15995 ( .C1(n14551), .C2(n14562), .A(n11533), .B(n14550), .ZN(
        n14685) );
  NAND2_X1 U15996 ( .A1(n14685), .A2(n14645), .ZN(n14554) );
  AOI22_X1 U15997 ( .A1(n14552), .A2(n16596), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n16598), .ZN(n14553) );
  OAI211_X1 U15998 ( .C1(n7856), .C2(n14621), .A(n14554), .B(n14553), .ZN(
        n14555) );
  AOI21_X1 U15999 ( .B1(n14687), .B2(n16604), .A(n14555), .ZN(n14556) );
  OAI21_X1 U16000 ( .B1(n16598), .B2(n14557), .A(n14556), .ZN(P2_U3243) );
  OAI211_X1 U16001 ( .C1(n14570), .C2(n14559), .A(n14558), .B(n16584), .ZN(
        n14561) );
  NAND2_X1 U16002 ( .A1(n14561), .A2(n14560), .ZN(n14691) );
  INV_X1 U16003 ( .A(n14691), .ZN(n14573) );
  AOI21_X1 U16004 ( .B1(n14583), .B2(n14566), .A(n11533), .ZN(n14563) );
  AND2_X1 U16005 ( .A1(n14563), .A2(n14562), .ZN(n14690) );
  OAI22_X1 U16006 ( .A1(n14610), .A2(n14565), .B1(n14564), .B2(n14640), .ZN(
        n14568) );
  INV_X1 U16007 ( .A(n14566), .ZN(n14759) );
  NOR2_X1 U16008 ( .A1(n14759), .A2(n14621), .ZN(n14567) );
  AOI211_X1 U16009 ( .C1(n14690), .C2(n14645), .A(n14568), .B(n14567), .ZN(
        n14572) );
  XNOR2_X1 U16010 ( .A(n14569), .B(n14570), .ZN(n14692) );
  NAND2_X1 U16011 ( .A1(n14692), .A2(n16604), .ZN(n14571) );
  OAI211_X1 U16012 ( .C1(n14573), .C2(n16598), .A(n14572), .B(n14571), .ZN(
        P2_U3244) );
  XOR2_X1 U16013 ( .A(n14574), .B(n14580), .Z(n14577) );
  AOI222_X1 U16014 ( .A1(n14579), .A2(n14578), .B1(n16584), .B2(n14577), .C1(
        n14576), .C2(n14575), .ZN(n14700) );
  XNOR2_X1 U16015 ( .A(n14581), .B(n14580), .ZN(n14701) );
  INV_X1 U16016 ( .A(n14701), .ZN(n14589) );
  OR2_X1 U16017 ( .A1(n14587), .A2(n14593), .ZN(n14582) );
  AND3_X1 U16018 ( .A1(n14583), .A2(n12771), .A3(n14582), .ZN(n14697) );
  NAND2_X1 U16019 ( .A1(n14697), .A2(n14645), .ZN(n14586) );
  AOI22_X1 U16020 ( .A1(n16598), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14584), 
        .B2(n16596), .ZN(n14585) );
  OAI211_X1 U16021 ( .C1(n14587), .C2(n14621), .A(n14586), .B(n14585), .ZN(
        n14588) );
  AOI21_X1 U16022 ( .B1(n14589), .B2(n16604), .A(n14588), .ZN(n14590) );
  OAI21_X1 U16023 ( .B1(n14700), .B2(n16598), .A(n14590), .ZN(P2_U3245) );
  OAI21_X1 U16024 ( .B1(n7548), .B2(n14592), .A(n14591), .ZN(n14702) );
  AOI211_X1 U16025 ( .C1(n14594), .C2(n14617), .A(n11533), .B(n14593), .ZN(
        n14704) );
  INV_X1 U16026 ( .A(n14594), .ZN(n14765) );
  NOR2_X1 U16027 ( .A1(n14765), .A2(n14621), .ZN(n14598) );
  OAI22_X1 U16028 ( .A1(n14610), .A2(n14596), .B1(n14595), .B2(n14640), .ZN(
        n14597) );
  AOI211_X1 U16029 ( .C1(n14704), .C2(n14645), .A(n14598), .B(n14597), .ZN(
        n14612) );
  OAI21_X1 U16030 ( .B1(n14601), .B2(n14600), .A(n14599), .ZN(n14607) );
  OAI22_X1 U16031 ( .A1(n14605), .A2(n14604), .B1(n14603), .B2(n14602), .ZN(
        n14606) );
  AOI21_X1 U16032 ( .B1(n14607), .B2(n16584), .A(n14606), .ZN(n14608) );
  OAI21_X1 U16033 ( .B1(n14702), .B2(n14609), .A(n14608), .ZN(n14703) );
  NAND2_X1 U16034 ( .A1(n14703), .A2(n14610), .ZN(n14611) );
  OAI211_X1 U16035 ( .C1(n14702), .C2(n14613), .A(n14612), .B(n14611), .ZN(
        P2_U3246) );
  XOR2_X1 U16036 ( .A(n14614), .B(n14626), .Z(n14616) );
  AOI21_X1 U16037 ( .B1(n14616), .B2(n16584), .A(n14615), .ZN(n14711) );
  INV_X1 U16038 ( .A(n14617), .ZN(n14618) );
  AOI211_X1 U16039 ( .C1(n14710), .C2(n14643), .A(n11533), .B(n14618), .ZN(
        n14709) );
  INV_X1 U16040 ( .A(n14710), .ZN(n14622) );
  AOI22_X1 U16041 ( .A1(n16598), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14619), 
        .B2(n16596), .ZN(n14620) );
  OAI21_X1 U16042 ( .B1(n14622), .B2(n14621), .A(n14620), .ZN(n14628) );
  INV_X1 U16043 ( .A(n14623), .ZN(n14624) );
  AOI21_X1 U16044 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14713) );
  NOR2_X1 U16045 ( .A1(n14713), .A2(n14648), .ZN(n14627) );
  AOI211_X1 U16046 ( .C1(n14709), .C2(n14645), .A(n14628), .B(n14627), .ZN(
        n14629) );
  OAI21_X1 U16047 ( .B1(n16598), .B2(n14711), .A(n14629), .ZN(P2_U3247) );
  OAI211_X1 U16048 ( .C1(n14630), .C2(n14632), .A(n14631), .B(n16584), .ZN(
        n14634) );
  NAND2_X1 U16049 ( .A1(n14634), .A2(n14633), .ZN(n14714) );
  OAI21_X1 U16050 ( .B1(n14637), .B2(n14636), .A(n14635), .ZN(n14718) );
  NAND2_X1 U16051 ( .A1(n16598), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14638) );
  OAI21_X1 U16052 ( .B1(n14640), .B2(n14639), .A(n14638), .ZN(n14641) );
  AOI21_X1 U16053 ( .B1(n14716), .B2(n16599), .A(n14641), .ZN(n14647) );
  AOI21_X1 U16054 ( .B1(n14716), .B2(n14642), .A(n11533), .ZN(n14644) );
  AND2_X1 U16055 ( .A1(n14644), .A2(n14643), .ZN(n14715) );
  NAND2_X1 U16056 ( .A1(n14715), .A2(n14645), .ZN(n14646) );
  OAI211_X1 U16057 ( .C1(n14718), .C2(n14648), .A(n14647), .B(n14646), .ZN(
        n14649) );
  AOI21_X1 U16058 ( .B1(n14610), .B2(n14714), .A(n14649), .ZN(n14650) );
  INV_X1 U16059 ( .A(n14650), .ZN(P2_U3248) );
  OAI21_X1 U16060 ( .B1(n14728), .B2(n14708), .A(n14653), .ZN(P2_U3530) );
  INV_X1 U16061 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14656) );
  AND2_X1 U16062 ( .A1(n14655), .A2(n14654), .ZN(n14729) );
  MUX2_X1 U16063 ( .A(n14656), .B(n14729), .S(n16591), .Z(n14657) );
  OAI21_X1 U16064 ( .B1(n14732), .B2(n14708), .A(n14657), .ZN(P2_U3529) );
  INV_X1 U16065 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14663) );
  INV_X1 U16066 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14667) );
  AOI211_X1 U16067 ( .C1(n16588), .C2(n14666), .A(n14665), .B(n14664), .ZN(
        n14741) );
  MUX2_X1 U16068 ( .A(n14667), .B(n14741), .S(n16591), .Z(n14668) );
  OAI21_X1 U16069 ( .B1(n14744), .B2(n14708), .A(n14668), .ZN(P2_U3525) );
  INV_X1 U16070 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14672) );
  AOI211_X1 U16071 ( .C1(n14671), .C2(n16588), .A(n14670), .B(n14669), .ZN(
        n14745) );
  MUX2_X1 U16072 ( .A(n14672), .B(n14745), .S(n16591), .Z(n14673) );
  OAI21_X1 U16073 ( .B1(n10368), .B2(n14708), .A(n14673), .ZN(P2_U3524) );
  AOI211_X1 U16074 ( .C1(n16418), .C2(n14676), .A(n14675), .B(n14674), .ZN(
        n14677) );
  OAI21_X1 U16075 ( .B1(n14723), .B2(n14678), .A(n14677), .ZN(n14748) );
  MUX2_X1 U16076 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14748), .S(n16591), .Z(
        P2_U3523) );
  INV_X1 U16077 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14683) );
  INV_X1 U16078 ( .A(n14679), .ZN(n14682) );
  AOI211_X1 U16079 ( .C1(n16514), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        n14749) );
  MUX2_X1 U16080 ( .A(n14683), .B(n14749), .S(n16591), .Z(n14684) );
  OAI21_X1 U16081 ( .B1(n14752), .B2(n14708), .A(n14684), .ZN(P2_U3522) );
  INV_X1 U16082 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14688) );
  AOI211_X1 U16083 ( .C1(n14687), .C2(n16588), .A(n14686), .B(n14685), .ZN(
        n14753) );
  MUX2_X1 U16084 ( .A(n14688), .B(n14753), .S(n16591), .Z(n14689) );
  OAI21_X1 U16085 ( .B1(n7856), .B2(n14708), .A(n14689), .ZN(P2_U3521) );
  INV_X1 U16086 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14695) );
  NOR2_X1 U16087 ( .A1(n14691), .A2(n14690), .ZN(n14694) );
  NAND2_X1 U16088 ( .A1(n14692), .A2(n16588), .ZN(n14693) );
  AND2_X1 U16089 ( .A1(n14694), .A2(n14693), .ZN(n14756) );
  MUX2_X1 U16090 ( .A(n14695), .B(n14756), .S(n16591), .Z(n14696) );
  OAI21_X1 U16091 ( .B1(n14759), .B2(n14708), .A(n14696), .ZN(P2_U3520) );
  AOI21_X1 U16092 ( .B1(n16418), .B2(n14698), .A(n14697), .ZN(n14699) );
  OAI211_X1 U16093 ( .C1(n14723), .C2(n14701), .A(n14700), .B(n14699), .ZN(
        n14760) );
  MUX2_X1 U16094 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14760), .S(n16591), .Z(
        P2_U3519) );
  INV_X1 U16095 ( .A(n14702), .ZN(n14705) );
  AOI211_X1 U16096 ( .C1(n14705), .C2(n16514), .A(n14704), .B(n14703), .ZN(
        n14761) );
  MUX2_X1 U16097 ( .A(n14706), .B(n14761), .S(n16591), .Z(n14707) );
  OAI21_X1 U16098 ( .B1(n14765), .B2(n14708), .A(n14707), .ZN(P2_U3518) );
  AOI21_X1 U16099 ( .B1(n16418), .B2(n14710), .A(n14709), .ZN(n14712) );
  OAI211_X1 U16100 ( .C1(n14713), .C2(n14723), .A(n14712), .B(n14711), .ZN(
        n14766) );
  MUX2_X1 U16101 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14766), .S(n16591), .Z(
        P2_U3517) );
  AOI211_X1 U16102 ( .C1(n16418), .C2(n14716), .A(n14715), .B(n14714), .ZN(
        n14717) );
  OAI21_X1 U16103 ( .B1(n14723), .B2(n14718), .A(n14717), .ZN(n14767) );
  MUX2_X1 U16104 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14767), .S(n16591), .Z(
        P2_U3516) );
  AOI21_X1 U16105 ( .B1(n16418), .B2(n14720), .A(n14719), .ZN(n14721) );
  OAI211_X1 U16106 ( .C1(n14724), .C2(n14723), .A(n14722), .B(n14721), .ZN(
        n14768) );
  MUX2_X1 U16107 ( .A(n14768), .B(P2_REG1_REG_16__SCAN_IN), .S(n16589), .Z(
        P2_U3515) );
  MUX2_X1 U16108 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14725), .S(n16591), .Z(
        P2_U3499) );
  OAI21_X1 U16109 ( .B1(n14728), .B2(n14764), .A(n14727), .ZN(P2_U3498) );
  INV_X1 U16110 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14730) );
  MUX2_X1 U16111 ( .A(n14730), .B(n14729), .S(n16595), .Z(n14731) );
  OAI21_X1 U16112 ( .B1(n14732), .B2(n14764), .A(n14731), .ZN(P2_U3497) );
  INV_X1 U16113 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14734) );
  MUX2_X1 U16114 ( .A(n14734), .B(n14733), .S(n16595), .Z(n14735) );
  OAI21_X1 U16115 ( .B1(n14736), .B2(n14764), .A(n14735), .ZN(P2_U3495) );
  INV_X1 U16116 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14738) );
  MUX2_X1 U16117 ( .A(n14738), .B(n14737), .S(n16595), .Z(n14739) );
  OAI21_X1 U16118 ( .B1(n14740), .B2(n14764), .A(n14739), .ZN(P2_U3494) );
  INV_X1 U16119 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14742) );
  MUX2_X1 U16120 ( .A(n14742), .B(n14741), .S(n16595), .Z(n14743) );
  OAI21_X1 U16121 ( .B1(n14744), .B2(n14764), .A(n14743), .ZN(P2_U3493) );
  INV_X1 U16122 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14746) );
  MUX2_X1 U16123 ( .A(n14746), .B(n14745), .S(n16595), .Z(n14747) );
  OAI21_X1 U16124 ( .B1(n10368), .B2(n14764), .A(n14747), .ZN(P2_U3492) );
  MUX2_X1 U16125 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14748), .S(n16595), .Z(
        P2_U3491) );
  INV_X1 U16126 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14750) );
  MUX2_X1 U16127 ( .A(n14750), .B(n14749), .S(n16595), .Z(n14751) );
  OAI21_X1 U16128 ( .B1(n14752), .B2(n14764), .A(n14751), .ZN(P2_U3490) );
  INV_X1 U16129 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14754) );
  MUX2_X1 U16130 ( .A(n14754), .B(n14753), .S(n16595), .Z(n14755) );
  OAI21_X1 U16131 ( .B1(n7856), .B2(n14764), .A(n14755), .ZN(P2_U3489) );
  INV_X1 U16132 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14757) );
  MUX2_X1 U16133 ( .A(n14757), .B(n14756), .S(n16595), .Z(n14758) );
  OAI21_X1 U16134 ( .B1(n14759), .B2(n14764), .A(n14758), .ZN(P2_U3488) );
  MUX2_X1 U16135 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14760), .S(n16595), .Z(
        P2_U3487) );
  INV_X1 U16136 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14762) );
  MUX2_X1 U16137 ( .A(n14762), .B(n14761), .S(n16595), .Z(n14763) );
  OAI21_X1 U16138 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(P2_U3486) );
  MUX2_X1 U16139 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14766), .S(n16595), .Z(
        P2_U3484) );
  MUX2_X1 U16140 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14767), .S(n16595), .Z(
        P2_U3481) );
  MUX2_X1 U16141 ( .A(n14768), .B(P2_REG0_REG_16__SCAN_IN), .S(n16592), .Z(
        P2_U3478) );
  INV_X1 U16142 ( .A(n10872), .ZN(n15795) );
  NAND3_X1 U16143 ( .A1(n14770), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14772) );
  OAI22_X1 U16144 ( .A1(n14769), .A2(n14772), .B1(n14771), .B2(n14792), .ZN(
        n14773) );
  INV_X1 U16145 ( .A(n14773), .ZN(n14774) );
  OAI21_X1 U16146 ( .B1(n15795), .B2(n14775), .A(n14774), .ZN(P2_U3296) );
  OAI222_X1 U16147 ( .A1(n14792), .A2(n14778), .B1(n14775), .B2(n14777), .C1(
        n14776), .C2(P2_U3088), .ZN(P2_U3298) );
  NAND2_X1 U16148 ( .A1(n15796), .A2(n14779), .ZN(n14781) );
  OAI211_X1 U16149 ( .C1(n14792), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        P2_U3299) );
  INV_X1 U16150 ( .A(n14783), .ZN(n15801) );
  OAI222_X1 U16151 ( .A1(n14792), .A2(n14785), .B1(n14775), .B2(n15801), .C1(
        P2_U3088), .C2(n14784), .ZN(P2_U3300) );
  INV_X1 U16152 ( .A(n14786), .ZN(n15806) );
  OAI222_X1 U16153 ( .A1(P2_U3088), .A2(n14788), .B1(n14775), .B2(n15806), 
        .C1(n14787), .C2(n14792), .ZN(P2_U3301) );
  INV_X1 U16154 ( .A(n14789), .ZN(n15808) );
  OAI222_X1 U16155 ( .A1(n14792), .A2(n14791), .B1(n14775), .B2(n15808), .C1(
        P2_U3088), .C2(n14790), .ZN(P2_U3302) );
  INV_X1 U16156 ( .A(n14793), .ZN(n14794) );
  MUX2_X1 U16157 ( .A(n14794), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16158 ( .A1(n14797), .A2(n14905), .ZN(n14804) );
  OAI22_X1 U16159 ( .A1(n16558), .A2(n14799), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14798), .ZN(n14802) );
  OAI22_X1 U16160 ( .A1(n15112), .A2(n16543), .B1(n16542), .B2(n14800), .ZN(
        n14801) );
  AOI211_X1 U16161 ( .C1(n15691), .C2(n16554), .A(n14802), .B(n14801), .ZN(
        n14803) );
  NAND2_X1 U16162 ( .A1(n14804), .A2(n14803), .ZN(P1_U3214) );
  INV_X1 U16163 ( .A(n15718), .ZN(n14815) );
  OAI21_X1 U16164 ( .B1(n14807), .B2(n14805), .A(n14806), .ZN(n14808) );
  NAND2_X1 U16165 ( .A1(n14808), .A2(n14905), .ZN(n14814) );
  NAND2_X1 U16166 ( .A1(n15114), .A2(n15234), .ZN(n14810) );
  NAND2_X1 U16167 ( .A1(n14925), .A2(n15233), .ZN(n14809) );
  NAND2_X1 U16168 ( .A1(n14810), .A2(n14809), .ZN(n15717) );
  INV_X1 U16169 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14811) );
  OAI22_X1 U16170 ( .A1(n15145), .A2(n16558), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14811), .ZN(n14812) );
  AOI21_X1 U16171 ( .B1(n15717), .B2(n14899), .A(n14812), .ZN(n14813) );
  OAI211_X1 U16172 ( .C1(n14815), .C2(n14918), .A(n14814), .B(n14813), .ZN(
        P1_U3216) );
  NAND2_X1 U16173 ( .A1(n14816), .A2(n14886), .ZN(n14818) );
  NAND2_X1 U16174 ( .A1(n14818), .A2(n14817), .ZN(n14819) );
  XOR2_X1 U16175 ( .A(n14820), .B(n14819), .Z(n14825) );
  OAI21_X1 U16176 ( .B1(n16558), .B2(n15219), .A(n14821), .ZN(n14823) );
  OAI22_X1 U16177 ( .A1(n15217), .A2(n16542), .B1(n16543), .B2(n15215), .ZN(
        n14822) );
  AOI211_X1 U16178 ( .C1(n15748), .C2(n16554), .A(n14823), .B(n14822), .ZN(
        n14824) );
  OAI21_X1 U16179 ( .B1(n14825), .B2(n16549), .A(n14824), .ZN(P1_U3219) );
  INV_X1 U16180 ( .A(n14826), .ZN(n14827) );
  AOI21_X1 U16181 ( .B1(n14829), .B2(n14828), .A(n14827), .ZN(n14835) );
  INV_X1 U16182 ( .A(n15186), .ZN(n14832) );
  OAI22_X1 U16183 ( .A1(n14830), .A2(n15218), .B1(n15217), .B2(n15216), .ZN(
        n15178) );
  AOI22_X1 U16184 ( .A1(n15178), .A2(n14899), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14831) );
  OAI21_X1 U16185 ( .B1(n14832), .B2(n16558), .A(n14831), .ZN(n14833) );
  AOI21_X1 U16186 ( .B1(n15729), .B2(n16554), .A(n14833), .ZN(n14834) );
  OAI21_X1 U16187 ( .B1(n14835), .B2(n16549), .A(n14834), .ZN(P1_U3223) );
  INV_X1 U16188 ( .A(n15123), .ZN(n15704) );
  INV_X1 U16189 ( .A(n14836), .ZN(n14869) );
  INV_X1 U16190 ( .A(n14837), .ZN(n14839) );
  NOR3_X1 U16191 ( .A1(n14869), .A2(n14839), .A3(n14838), .ZN(n14842) );
  INV_X1 U16192 ( .A(n14840), .ZN(n14841) );
  OAI21_X1 U16193 ( .B1(n14842), .B2(n14841), .A(n14905), .ZN(n14847) );
  NOR2_X1 U16194 ( .A1(n16558), .A2(n15120), .ZN(n14845) );
  OAI22_X1 U16195 ( .A1(n14843), .A2(n16543), .B1(n15112), .B2(n16542), .ZN(
        n14844) );
  AOI211_X1 U16196 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n14845), 
        .B(n14844), .ZN(n14846) );
  OAI211_X1 U16197 ( .C1(n15704), .C2(n14918), .A(n14847), .B(n14846), .ZN(
        P1_U3225) );
  INV_X1 U16198 ( .A(n14849), .ZN(n14850) );
  AOI21_X1 U16199 ( .B1(n14851), .B2(n14848), .A(n14850), .ZN(n14856) );
  NAND2_X1 U16200 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15034)
         );
  OAI21_X1 U16201 ( .B1(n16558), .B2(n14852), .A(n15034), .ZN(n14854) );
  OAI22_X1 U16202 ( .A1(n16541), .A2(n16543), .B1(n16542), .B2(n14889), .ZN(
        n14853) );
  AOI211_X1 U16203 ( .C1(n15762), .C2(n16554), .A(n14854), .B(n14853), .ZN(
        n14855) );
  OAI21_X1 U16204 ( .B1(n14856), .B2(n16549), .A(n14855), .ZN(P1_U3226) );
  OAI21_X1 U16205 ( .B1(n14859), .B2(n14857), .A(n14858), .ZN(n14860) );
  NAND2_X1 U16206 ( .A1(n14860), .A2(n14905), .ZN(n14865) );
  INV_X1 U16207 ( .A(n14861), .ZN(n15254) );
  AND2_X1 U16208 ( .A1(n14928), .A2(n15233), .ZN(n14862) );
  AOI21_X1 U16209 ( .B1(n14927), .B2(n15234), .A(n14862), .ZN(n15250) );
  NAND2_X1 U16210 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15045)
         );
  OAI21_X1 U16211 ( .B1(n14912), .B2(n15250), .A(n15045), .ZN(n14863) );
  AOI21_X1 U16212 ( .B1(n15254), .B2(n14914), .A(n14863), .ZN(n14864) );
  OAI211_X1 U16213 ( .C1(n7950), .C2(n14918), .A(n14865), .B(n14864), .ZN(
        P1_U3228) );
  INV_X1 U16214 ( .A(n15711), .ZN(n15138) );
  INV_X1 U16215 ( .A(n14806), .ZN(n14868) );
  NOR3_X1 U16216 ( .A1(n14868), .A2(n14867), .A3(n14866), .ZN(n14870) );
  OAI21_X1 U16217 ( .B1(n14870), .B2(n14869), .A(n14905), .ZN(n14876) );
  NAND2_X1 U16218 ( .A1(n14924), .A2(n15233), .ZN(n14872) );
  NAND2_X1 U16219 ( .A1(n15234), .A2(n14923), .ZN(n14871) );
  NAND2_X1 U16220 ( .A1(n14872), .A2(n14871), .ZN(n15710) );
  INV_X1 U16221 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14873) );
  OAI22_X1 U16222 ( .A1(n15134), .A2(n16558), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14873), .ZN(n14874) );
  AOI21_X1 U16223 ( .B1(n15710), .B2(n14899), .A(n14874), .ZN(n14875) );
  OAI211_X1 U16224 ( .C1(n15138), .C2(n14918), .A(n14876), .B(n14875), .ZN(
        P1_U3229) );
  NAND2_X1 U16225 ( .A1(n14879), .A2(n14878), .ZN(n14880) );
  XNOR2_X1 U16226 ( .A(n14877), .B(n14880), .ZN(n14885) );
  OAI22_X1 U16227 ( .A1(n15167), .A2(n16558), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14881), .ZN(n14883) );
  OAI22_X1 U16228 ( .A1(n15162), .A2(n16542), .B1(n15161), .B2(n16543), .ZN(
        n14882) );
  AOI211_X1 U16229 ( .C1(n15726), .C2(n16554), .A(n14883), .B(n14882), .ZN(
        n14884) );
  OAI21_X1 U16230 ( .B1(n14885), .B2(n16549), .A(n14884), .ZN(P1_U3235) );
  XOR2_X1 U16231 ( .A(n14816), .B(n14886), .Z(n14893) );
  OAI21_X1 U16232 ( .B1(n16558), .B2(n15240), .A(n14887), .ZN(n14891) );
  OAI22_X1 U16233 ( .A1(n14889), .A2(n16543), .B1(n16542), .B2(n14888), .ZN(
        n14890) );
  AOI211_X1 U16234 ( .C1(n15753), .C2(n16554), .A(n14891), .B(n14890), .ZN(
        n14892) );
  OAI21_X1 U16235 ( .B1(n14893), .B2(n16549), .A(n14892), .ZN(P1_U3238) );
  OAI21_X1 U16236 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14903) );
  NAND2_X1 U16237 ( .A1(n15696), .A2(n16554), .ZN(n14901) );
  OAI22_X1 U16238 ( .A1(n14898), .A2(n15216), .B1(n15218), .B2(n14897), .ZN(
        n15096) );
  AOI22_X1 U16239 ( .A1(n14899), .A2(n15096), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14900) );
  OAI211_X1 U16240 ( .C1(n16558), .C2(n15099), .A(n14901), .B(n14900), .ZN(
        n14902) );
  AOI21_X1 U16241 ( .B1(n14903), .B2(n14905), .A(n14902), .ZN(n14904) );
  INV_X1 U16242 ( .A(n14904), .ZN(P1_U3240) );
  OAI211_X1 U16243 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n14917) );
  INV_X1 U16244 ( .A(n16652), .ZN(n14915) );
  NAND2_X1 U16245 ( .A1(n14928), .A2(n15234), .ZN(n14910) );
  NAND2_X1 U16246 ( .A1(n15233), .A2(n14930), .ZN(n14909) );
  AND2_X1 U16247 ( .A1(n14910), .A2(n14909), .ZN(n16639) );
  OAI22_X1 U16248 ( .A1(n14912), .A2(n16639), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14911), .ZN(n14913) );
  AOI21_X1 U16249 ( .B1(n14915), .B2(n14914), .A(n14913), .ZN(n14916) );
  OAI211_X1 U16250 ( .C1(n16641), .C2(n14918), .A(n14917), .B(n14916), .ZN(
        P1_U3241) );
  MUX2_X1 U16251 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14919), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16252 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14920), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16253 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15077), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16254 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14921), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16255 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15076), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16256 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14922), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16257 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14923), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16258 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15114), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16259 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14924), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16260 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14925), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16261 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15194), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16262 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14926), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16263 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15235), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16264 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14927), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16265 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15232), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16266 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14928), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16267 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14929), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16268 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14930), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16269 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14931), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16270 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14932), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16271 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14933), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16272 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14934), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16273 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14935), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16274 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14936), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16275 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14937), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16276 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14938), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16277 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14939), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16278 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14940), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16279 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14941), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16280 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14942), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16281 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10603), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16282 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14943), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16283 ( .C1(n14956), .C2(n14945), .A(n16277), .B(n14944), .ZN(
        n14953) );
  OAI211_X1 U16284 ( .C1(n14948), .C2(n14947), .A(n16283), .B(n14946), .ZN(
        n14952) );
  AOI22_X1 U16285 ( .A1(n16287), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14951) );
  NAND2_X1 U16286 ( .A1(n16285), .A2(n14949), .ZN(n14950) );
  NAND4_X1 U16287 ( .A1(n14953), .A2(n14952), .A3(n14951), .A4(n14950), .ZN(
        P1_U3244) );
  MUX2_X1 U16288 ( .A(n14956), .B(n14955), .S(n14954), .Z(n14958) );
  NAND2_X1 U16289 ( .A1(n14958), .A2(n14957), .ZN(n14960) );
  OAI211_X1 U16290 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14961), .A(n14960), .B(
        P1_U4016), .ZN(n16292) );
  INV_X1 U16291 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14963) );
  OAI22_X1 U16292 ( .A1(n15046), .A2(n14963), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14962), .ZN(n14964) );
  AOI21_X1 U16293 ( .B1(n16285), .B2(n14965), .A(n14964), .ZN(n14972) );
  OAI211_X1 U16294 ( .C1(n14967), .C2(n14966), .A(n16277), .B(n14977), .ZN(
        n14971) );
  OAI211_X1 U16295 ( .C1(n14969), .C2(n14968), .A(n16283), .B(n14982), .ZN(
        n14970) );
  NAND4_X1 U16296 ( .A1(n16292), .A2(n14972), .A3(n14971), .A4(n14970), .ZN(
        P1_U3245) );
  OAI22_X1 U16297 ( .A1(n15046), .A2(n15947), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14973), .ZN(n14974) );
  AOI21_X1 U16298 ( .B1(n16285), .B2(n14979), .A(n14974), .ZN(n14986) );
  MUX2_X1 U16299 ( .A(n11153), .B(P1_REG2_REG_3__SCAN_IN), .S(n14979), .Z(
        n14975) );
  NAND3_X1 U16300 ( .A1(n14977), .A2(n14976), .A3(n14975), .ZN(n14978) );
  NAND3_X1 U16301 ( .A1(n16277), .A2(n16274), .A3(n14978), .ZN(n14985) );
  MUX2_X1 U16302 ( .A(n11129), .B(P1_REG1_REG_3__SCAN_IN), .S(n14979), .Z(
        n14980) );
  NAND3_X1 U16303 ( .A1(n14982), .A2(n14981), .A3(n14980), .ZN(n14983) );
  NAND3_X1 U16304 ( .A1(n16283), .A2(n16280), .A3(n14983), .ZN(n14984) );
  NAND3_X1 U16305 ( .A1(n14986), .A2(n14985), .A3(n14984), .ZN(P1_U3246) );
  INV_X1 U16306 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14988) );
  OAI21_X1 U16307 ( .B1(n15046), .B2(n14988), .A(n14987), .ZN(n14989) );
  AOI21_X1 U16308 ( .B1(n16285), .B2(n14994), .A(n14989), .ZN(n15001) );
  OAI21_X1 U16309 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n14993) );
  NAND2_X1 U16310 ( .A1(n16283), .A2(n14993), .ZN(n15000) );
  MUX2_X1 U16311 ( .A(n14995), .B(P1_REG2_REG_5__SCAN_IN), .S(n14994), .Z(
        n14996) );
  NAND3_X1 U16312 ( .A1(n16276), .A2(n14997), .A3(n14996), .ZN(n14998) );
  NAND3_X1 U16313 ( .A1(n16277), .A2(n15009), .A3(n14998), .ZN(n14999) );
  NAND3_X1 U16314 ( .A1(n15001), .A2(n15000), .A3(n14999), .ZN(P1_U3248) );
  OAI21_X1 U16315 ( .B1(n15046), .B2(n15973), .A(n15002), .ZN(n15003) );
  AOI21_X1 U16316 ( .B1(n16285), .B2(n15006), .A(n15003), .ZN(n15013) );
  OAI211_X1 U16317 ( .C1(n15005), .C2(n15004), .A(n16283), .B(n15025), .ZN(
        n15012) );
  MUX2_X1 U16318 ( .A(n11161), .B(P1_REG2_REG_6__SCAN_IN), .S(n15006), .Z(
        n15007) );
  NAND3_X1 U16319 ( .A1(n15009), .A2(n15008), .A3(n15007), .ZN(n15010) );
  NAND3_X1 U16320 ( .A1(n16277), .A2(n15018), .A3(n15010), .ZN(n15011) );
  NAND3_X1 U16321 ( .A1(n15013), .A2(n15012), .A3(n15011), .ZN(P1_U3249) );
  INV_X1 U16322 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15978) );
  OAI21_X1 U16323 ( .B1(n15046), .B2(n15978), .A(n15014), .ZN(n15015) );
  AOI21_X1 U16324 ( .B1(n16285), .B2(n15021), .A(n15015), .ZN(n15030) );
  MUX2_X1 U16325 ( .A(n11164), .B(P1_REG2_REG_7__SCAN_IN), .S(n15021), .Z(
        n15016) );
  NAND3_X1 U16326 ( .A1(n15018), .A2(n15017), .A3(n15016), .ZN(n15019) );
  NAND3_X1 U16327 ( .A1(n16277), .A2(n15020), .A3(n15019), .ZN(n15029) );
  MUX2_X1 U16328 ( .A(n15022), .B(P1_REG1_REG_7__SCAN_IN), .S(n15021), .Z(
        n15023) );
  NAND3_X1 U16329 ( .A1(n15025), .A2(n15024), .A3(n15023), .ZN(n15026) );
  NAND3_X1 U16330 ( .A1(n16283), .A2(n15027), .A3(n15026), .ZN(n15028) );
  NAND3_X1 U16331 ( .A1(n15030), .A2(n15029), .A3(n15028), .ZN(P1_U3250) );
  OAI211_X1 U16332 ( .C1(n15033), .C2(n15032), .A(n16277), .B(n15031), .ZN(
        n15043) );
  INV_X1 U16333 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15035) );
  OAI21_X1 U16334 ( .B1(n15046), .B2(n15035), .A(n15034), .ZN(n15036) );
  AOI21_X1 U16335 ( .B1(n16285), .B2(n15037), .A(n15036), .ZN(n15042) );
  OAI211_X1 U16336 ( .C1(n15040), .C2(n15039), .A(n16283), .B(n15038), .ZN(
        n15041) );
  NAND3_X1 U16337 ( .A1(n15043), .A2(n15042), .A3(n15041), .ZN(P1_U3259) );
  INV_X1 U16338 ( .A(n15044), .ZN(n15048) );
  OAI21_X1 U16339 ( .B1(n15046), .B2(n7688), .A(n15045), .ZN(n15047) );
  AOI21_X1 U16340 ( .B1(n16285), .B2(n15048), .A(n15047), .ZN(n15057) );
  OAI211_X1 U16341 ( .C1(n15051), .C2(n15050), .A(n16283), .B(n15049), .ZN(
        n15056) );
  OAI211_X1 U16342 ( .C1(n15054), .C2(n15053), .A(n16277), .B(n15052), .ZN(
        n15055) );
  NAND3_X1 U16343 ( .A1(n15057), .A2(n15056), .A3(n15055), .ZN(P1_U3260) );
  INV_X1 U16344 ( .A(n15262), .ZN(n15063) );
  XOR2_X1 U16345 ( .A(n15262), .B(n15066), .Z(n15058) );
  NOR2_X1 U16346 ( .A1(n15058), .A2(n16566), .ZN(n15265) );
  NAND2_X1 U16347 ( .A1(n15265), .A2(n16498), .ZN(n15062) );
  NOR2_X1 U16348 ( .A1(n16398), .A2(n8390), .ZN(n15070) );
  AOI21_X1 U16349 ( .B1(n16398), .B2(P1_REG2_REG_31__SCAN_IN), .A(n15070), 
        .ZN(n15061) );
  OAI211_X1 U16350 ( .C1(n15063), .C2(n16493), .A(n15062), .B(n15061), .ZN(
        P1_U3263) );
  INV_X1 U16351 ( .A(n15064), .ZN(n15068) );
  INV_X1 U16352 ( .A(n15066), .ZN(n15067) );
  OAI211_X1 U16353 ( .C1(n15068), .C2(n15674), .A(n15067), .B(n16622), .ZN(
        n15673) );
  NOR2_X1 U16354 ( .A1(n15674), .A2(n16493), .ZN(n15069) );
  AOI211_X1 U16355 ( .C1(n16398), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15070), 
        .B(n15069), .ZN(n15071) );
  OAI21_X1 U16356 ( .B1(n15673), .B2(n16644), .A(n15071), .ZN(P1_U3264) );
  NAND3_X1 U16357 ( .A1(n15074), .A2(n15090), .A3(n15073), .ZN(n15075) );
  NAND2_X1 U16358 ( .A1(n15072), .A2(n15075), .ZN(n15081) );
  NAND2_X1 U16359 ( .A1(n15076), .A2(n15233), .ZN(n15079) );
  NAND2_X1 U16360 ( .A1(n15077), .A2(n15234), .ZN(n15078) );
  OAI21_X1 U16361 ( .B1(n15082), .B2(n15085), .A(n16622), .ZN(n15084) );
  NOR2_X1 U16362 ( .A1(n15084), .A2(n15083), .ZN(n15685) );
  NOR2_X1 U16363 ( .A1(n15085), .A2(n16493), .ZN(n15089) );
  OAI22_X1 U16364 ( .A1(n7416), .A2(n15087), .B1(n15086), .B2(n16653), .ZN(
        n15088) );
  AOI211_X1 U16365 ( .C1(n15685), .C2(n16498), .A(n15089), .B(n15088), .ZN(
        n15094) );
  OR2_X2 U16366 ( .A1(n15091), .A2(n15090), .ZN(n15684) );
  NAND3_X1 U16367 ( .A1(n15684), .A2(n16394), .A3(n15092), .ZN(n15093) );
  OAI211_X1 U16368 ( .C1(n15688), .C2(n16398), .A(n15094), .B(n15093), .ZN(
        P1_U3265) );
  AOI211_X1 U16369 ( .C1(n15103), .C2(n15095), .A(n16351), .B(n7473), .ZN(
        n15097) );
  NOR2_X1 U16370 ( .A1(n15097), .A2(n15096), .ZN(n15698) );
  AOI211_X1 U16371 ( .C1(n15696), .C2(n7494), .A(n16566), .B(n15098), .ZN(
        n15695) );
  INV_X1 U16372 ( .A(n15696), .ZN(n15102) );
  INV_X1 U16373 ( .A(n15099), .ZN(n15100) );
  AOI22_X1 U16374 ( .A1(n16398), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15100), 
        .B2(n16490), .ZN(n15101) );
  OAI21_X1 U16375 ( .B1(n15102), .B2(n16493), .A(n15101), .ZN(n15108) );
  OR2_X1 U16376 ( .A1(n15104), .A2(n15103), .ZN(n15105) );
  NAND2_X1 U16377 ( .A1(n15106), .A2(n15105), .ZN(n15699) );
  NOR2_X1 U16378 ( .A1(n15699), .A2(n16646), .ZN(n15107) );
  AOI211_X1 U16379 ( .C1(n15695), .C2(n16498), .A(n15108), .B(n15107), .ZN(
        n15109) );
  OAI21_X1 U16380 ( .B1(n15698), .B2(n16398), .A(n15109), .ZN(P1_U3267) );
  XNOR2_X1 U16381 ( .A(n15110), .B(n15118), .ZN(n15111) );
  NAND2_X1 U16382 ( .A1(n15111), .A2(n16631), .ZN(n15116) );
  NOR2_X1 U16383 ( .A1(n15218), .A2(n15112), .ZN(n15113) );
  AOI21_X1 U16384 ( .B1(n15114), .B2(n15233), .A(n15113), .ZN(n15115) );
  NAND2_X1 U16385 ( .A1(n15116), .A2(n15115), .ZN(n15706) );
  AOI21_X1 U16386 ( .B1(n15123), .B2(n15131), .A(n16566), .ZN(n15117) );
  NAND2_X1 U16387 ( .A1(n15117), .A2(n7494), .ZN(n15702) );
  NAND2_X1 U16388 ( .A1(n15119), .A2(n15118), .ZN(n15700) );
  NAND3_X1 U16389 ( .A1(n15701), .A2(n15700), .A3(n16394), .ZN(n15125) );
  INV_X1 U16390 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15121) );
  OAI22_X1 U16391 ( .A1(n7416), .A2(n15121), .B1(n15120), .B2(n16653), .ZN(
        n15122) );
  AOI21_X1 U16392 ( .B1(n15123), .B2(n16389), .A(n15122), .ZN(n15124) );
  OAI211_X1 U16393 ( .C1(n15702), .C2(n16644), .A(n15125), .B(n15124), .ZN(
        n15126) );
  AOI21_X1 U16394 ( .B1(n15706), .B2(n7416), .A(n15126), .ZN(n15127) );
  INV_X1 U16395 ( .A(n15127), .ZN(P1_U3268) );
  XOR2_X1 U16396 ( .A(n7536), .B(n15130), .Z(n15715) );
  OAI21_X1 U16397 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(n15712) );
  AOI21_X1 U16398 ( .B1(n15711), .B2(n15142), .A(n16566), .ZN(n15132) );
  AND2_X1 U16399 ( .A1(n15132), .A2(n15131), .ZN(n15709) );
  NAND2_X1 U16400 ( .A1(n15709), .A2(n16498), .ZN(n15137) );
  INV_X1 U16401 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15133) );
  OAI22_X1 U16402 ( .A1(n15134), .A2(n16653), .B1(n15133), .B2(n7416), .ZN(
        n15135) );
  AOI21_X1 U16403 ( .B1(n15710), .B2(n7416), .A(n15135), .ZN(n15136) );
  OAI211_X1 U16404 ( .C1(n15138), .C2(n16493), .A(n15137), .B(n15136), .ZN(
        n15139) );
  AOI21_X1 U16405 ( .B1(n16394), .B2(n15712), .A(n15139), .ZN(n15140) );
  OAI21_X1 U16406 ( .B1(n15715), .B2(n16647), .A(n15140), .ZN(P1_U3269) );
  XNOR2_X1 U16407 ( .A(n15141), .B(n15151), .ZN(n15716) );
  INV_X1 U16408 ( .A(n15716), .ZN(n15154) );
  AOI21_X1 U16409 ( .B1(n15165), .B2(n15718), .A(n16566), .ZN(n15143) );
  NAND2_X1 U16410 ( .A1(n15143), .A2(n15142), .ZN(n15720) );
  INV_X1 U16411 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15144) );
  OAI22_X1 U16412 ( .A1(n15145), .A2(n16653), .B1(n15144), .B2(n7416), .ZN(
        n15146) );
  AOI21_X1 U16413 ( .B1(n15717), .B2(n7416), .A(n15146), .ZN(n15148) );
  NAND2_X1 U16414 ( .A1(n15718), .A2(n16389), .ZN(n15147) );
  OAI211_X1 U16415 ( .C1(n15720), .C2(n16644), .A(n15148), .B(n15147), .ZN(
        n15149) );
  INV_X1 U16416 ( .A(n15149), .ZN(n15153) );
  NAND2_X1 U16417 ( .A1(n15150), .A2(n15151), .ZN(n15719) );
  NAND3_X1 U16418 ( .A1(n8166), .A2(n15719), .A3(n16394), .ZN(n15152) );
  OAI211_X1 U16419 ( .C1(n15154), .C2(n16647), .A(n15153), .B(n15152), .ZN(
        P1_U3270) );
  XNOR2_X1 U16420 ( .A(n15155), .B(n10570), .ZN(n15728) );
  INV_X1 U16421 ( .A(n15156), .ZN(n15157) );
  AOI21_X1 U16422 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15160) );
  OAI222_X1 U16423 ( .A1(n15218), .A2(n15162), .B1(n15216), .B2(n15161), .C1(
        n16351), .C2(n15160), .ZN(n15724) );
  AOI21_X1 U16424 ( .B1(n15726), .B2(n15185), .A(n16566), .ZN(n15164) );
  AND2_X1 U16425 ( .A1(n15165), .A2(n15164), .ZN(n15725) );
  NAND2_X1 U16426 ( .A1(n15725), .A2(n16498), .ZN(n15170) );
  INV_X1 U16427 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15166) );
  OAI22_X1 U16428 ( .A1(n15167), .A2(n16653), .B1(n15166), .B2(n7416), .ZN(
        n15168) );
  AOI21_X1 U16429 ( .B1(n15726), .B2(n16389), .A(n15168), .ZN(n15169) );
  NAND2_X1 U16430 ( .A1(n15170), .A2(n15169), .ZN(n15171) );
  AOI21_X1 U16431 ( .B1(n15724), .B2(n7416), .A(n15171), .ZN(n15172) );
  OAI21_X1 U16432 ( .B1(n15728), .B2(n16646), .A(n15172), .ZN(P1_U3271) );
  NAND3_X1 U16433 ( .A1(n15173), .A2(n15175), .A3(n15174), .ZN(n15176) );
  NAND3_X1 U16434 ( .A1(n15177), .A2(n16631), .A3(n15176), .ZN(n15180) );
  INV_X1 U16435 ( .A(n15178), .ZN(n15179) );
  NAND2_X1 U16436 ( .A1(n15180), .A2(n15179), .ZN(n15735) );
  INV_X1 U16437 ( .A(n15735), .ZN(n15191) );
  NAND2_X1 U16438 ( .A1(n15181), .A2(n9854), .ZN(n15182) );
  NAND2_X1 U16439 ( .A1(n15183), .A2(n15182), .ZN(n15730) );
  NAND2_X1 U16440 ( .A1(n15198), .A2(n15729), .ZN(n15184) );
  NAND3_X1 U16441 ( .A1(n15185), .A2(n16622), .A3(n15184), .ZN(n15731) );
  AOI22_X1 U16442 ( .A1(n15186), .A2(n16490), .B1(n16398), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U16443 ( .A1(n15729), .A2(n16389), .ZN(n15187) );
  OAI211_X1 U16444 ( .C1(n15731), .C2(n16644), .A(n15188), .B(n15187), .ZN(
        n15189) );
  AOI21_X1 U16445 ( .B1(n15730), .B2(n16394), .A(n15189), .ZN(n15190) );
  OAI21_X1 U16446 ( .B1(n15191), .B2(n16398), .A(n15190), .ZN(P1_U3272) );
  OAI211_X1 U16447 ( .C1(n15193), .C2(n15192), .A(n16631), .B(n15173), .ZN(
        n15745) );
  NAND2_X1 U16448 ( .A1(n15194), .A2(n15234), .ZN(n15196) );
  NAND2_X1 U16449 ( .A1(n15235), .A2(n15233), .ZN(n15195) );
  NAND2_X1 U16450 ( .A1(n15196), .A2(n15195), .ZN(n15738) );
  INV_X1 U16451 ( .A(n15738), .ZN(n15197) );
  AOI21_X1 U16452 ( .B1(n15745), .B2(n15197), .A(n16398), .ZN(n15208) );
  OAI211_X1 U16453 ( .C1(n15199), .C2(n15221), .A(n16622), .B(n15198), .ZN(
        n15742) );
  OR2_X1 U16454 ( .A1(n15201), .A2(n15200), .ZN(n15740) );
  NAND3_X1 U16455 ( .A1(n15740), .A2(n15741), .A3(n16394), .ZN(n15206) );
  INV_X1 U16456 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15203) );
  OAI22_X1 U16457 ( .A1(n7416), .A2(n15203), .B1(n15202), .B2(n16653), .ZN(
        n15204) );
  AOI21_X1 U16458 ( .B1(n15739), .B2(n16389), .A(n15204), .ZN(n15205) );
  OAI211_X1 U16459 ( .C1(n15742), .C2(n16644), .A(n15206), .B(n15205), .ZN(
        n15207) );
  OR2_X1 U16460 ( .A1(n15208), .A2(n15207), .ZN(P1_U3273) );
  XOR2_X1 U16461 ( .A(n15209), .B(n15213), .Z(n15750) );
  INV_X1 U16462 ( .A(n15210), .ZN(n15211) );
  AOI21_X1 U16463 ( .B1(n15213), .B2(n15212), .A(n15211), .ZN(n15214) );
  OAI222_X1 U16464 ( .A1(n15218), .A2(n15217), .B1(n15216), .B2(n15215), .C1(
        n16351), .C2(n15214), .ZN(n15746) );
  NOR2_X1 U16465 ( .A1(n15219), .A2(n16653), .ZN(n15220) );
  OAI21_X1 U16466 ( .B1(n15746), .B2(n15220), .A(n7416), .ZN(n15226) );
  AOI211_X1 U16467 ( .C1(n15748), .C2(n15238), .A(n16566), .B(n15221), .ZN(
        n15747) );
  INV_X1 U16468 ( .A(n15748), .ZN(n15223) );
  INV_X1 U16469 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15222) );
  OAI22_X1 U16470 ( .A1(n15223), .A2(n16493), .B1(n15222), .B2(n7416), .ZN(
        n15224) );
  AOI21_X1 U16471 ( .B1(n15747), .B2(n16498), .A(n15224), .ZN(n15225) );
  OAI211_X1 U16472 ( .C1(n15750), .C2(n16646), .A(n15226), .B(n15225), .ZN(
        P1_U3274) );
  XNOR2_X1 U16473 ( .A(n15228), .B(n15227), .ZN(n15755) );
  OAI211_X1 U16474 ( .C1(n15231), .C2(n15230), .A(n15229), .B(n16631), .ZN(
        n15237) );
  AOI22_X1 U16475 ( .A1(n15235), .A2(n15234), .B1(n15233), .B2(n15232), .ZN(
        n15236) );
  NAND2_X1 U16476 ( .A1(n15237), .A2(n15236), .ZN(n15751) );
  AOI21_X1 U16477 ( .B1(n15753), .B2(n15252), .A(n16566), .ZN(n15239) );
  AND2_X1 U16478 ( .A1(n15239), .A2(n15238), .ZN(n15752) );
  NAND2_X1 U16479 ( .A1(n15752), .A2(n16498), .ZN(n15244) );
  OAI22_X1 U16480 ( .A1(n7416), .A2(n15241), .B1(n15240), .B2(n16653), .ZN(
        n15242) );
  AOI21_X1 U16481 ( .B1(n15753), .B2(n16389), .A(n15242), .ZN(n15243) );
  NAND2_X1 U16482 ( .A1(n15244), .A2(n15243), .ZN(n15245) );
  AOI21_X1 U16483 ( .B1(n15751), .B2(n7416), .A(n15245), .ZN(n15246) );
  OAI21_X1 U16484 ( .B1(n15247), .B2(n15755), .A(n15246), .ZN(P1_U3275) );
  OAI211_X1 U16485 ( .C1(n15249), .C2(n15256), .A(n15248), .B(n16631), .ZN(
        n15251) );
  AOI211_X1 U16486 ( .C1(n15757), .C2(n15253), .A(n16566), .B(n7949), .ZN(
        n15756) );
  AOI22_X1 U16487 ( .A1(n16398), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15254), 
        .B2(n16490), .ZN(n15255) );
  OAI21_X1 U16488 ( .B1(n7950), .B2(n16493), .A(n15255), .ZN(n15260) );
  OAI21_X1 U16489 ( .B1(n15258), .B2(n7696), .A(n15257), .ZN(n15760) );
  NOR2_X1 U16490 ( .A1(n15760), .A2(n16646), .ZN(n15259) );
  AOI211_X1 U16491 ( .C1(n15756), .C2(n16498), .A(n15260), .B(n15259), .ZN(
        n15261) );
  OAI21_X1 U16492 ( .B1(n16398), .B2(n15759), .A(n15261), .ZN(P1_U3276) );
  NOR2_X2 U16493 ( .A1(n15265), .A2(n15264), .ZN(n15771) );
  NAND2_X1 U16494 ( .A1(n16633), .A2(n15266), .ZN(n15267) );
  XNOR2_X1 U16495 ( .A(n15663), .B(keyinput_254), .ZN(n15670) );
  XOR2_X1 U16496 ( .A(SI_31_), .B(keyinput_129), .Z(n15271) );
  XOR2_X1 U16497 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n15270) );
  XOR2_X1 U16498 ( .A(SI_30_), .B(keyinput_130), .Z(n15269) );
  AOI21_X1 U16499 ( .B1(n15271), .B2(n15270), .A(n15269), .ZN(n15275) );
  XNOR2_X1 U16500 ( .A(n15461), .B(keyinput_133), .ZN(n15274) );
  XNOR2_X1 U16501 ( .A(n15459), .B(keyinput_132), .ZN(n15273) );
  XNOR2_X1 U16502 ( .A(SI_29_), .B(keyinput_131), .ZN(n15272) );
  NOR4_X1 U16503 ( .A1(n15275), .A2(n15274), .A3(n15273), .A4(n15272), .ZN(
        n15279) );
  XOR2_X1 U16504 ( .A(SI_26_), .B(keyinput_134), .Z(n15278) );
  XNOR2_X1 U16505 ( .A(n15466), .B(keyinput_135), .ZN(n15277) );
  XOR2_X1 U16506 ( .A(SI_24_), .B(keyinput_136), .Z(n15276) );
  OAI211_X1 U16507 ( .C1(n15279), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15282) );
  XOR2_X1 U16508 ( .A(SI_23_), .B(keyinput_137), .Z(n15281) );
  XOR2_X1 U16509 ( .A(SI_22_), .B(keyinput_138), .Z(n15280) );
  NAND3_X1 U16510 ( .A1(n15282), .A2(n15281), .A3(n15280), .ZN(n15286) );
  XOR2_X1 U16511 ( .A(SI_20_), .B(keyinput_140), .Z(n15285) );
  XNOR2_X1 U16512 ( .A(SI_21_), .B(keyinput_139), .ZN(n15284) );
  XNOR2_X1 U16513 ( .A(SI_19_), .B(keyinput_141), .ZN(n15283) );
  NAND4_X1 U16514 ( .A1(n15286), .A2(n15285), .A3(n15284), .A4(n15283), .ZN(
        n15292) );
  XNOR2_X1 U16515 ( .A(SI_18_), .B(keyinput_142), .ZN(n15291) );
  XNOR2_X1 U16516 ( .A(n15480), .B(keyinput_143), .ZN(n15289) );
  XNOR2_X1 U16517 ( .A(SI_16_), .B(keyinput_144), .ZN(n15288) );
  XNOR2_X1 U16518 ( .A(SI_15_), .B(keyinput_145), .ZN(n15287) );
  NAND3_X1 U16519 ( .A1(n15289), .A2(n15288), .A3(n15287), .ZN(n15290) );
  AOI21_X1 U16520 ( .B1(n15292), .B2(n15291), .A(n15290), .ZN(n15296) );
  XNOR2_X1 U16521 ( .A(SI_12_), .B(keyinput_148), .ZN(n15295) );
  XNOR2_X1 U16522 ( .A(SI_13_), .B(keyinput_147), .ZN(n15294) );
  XNOR2_X1 U16523 ( .A(SI_14_), .B(keyinput_146), .ZN(n15293) );
  NOR4_X1 U16524 ( .A1(n15296), .A2(n15295), .A3(n15294), .A4(n15293), .ZN(
        n15300) );
  XOR2_X1 U16525 ( .A(SI_10_), .B(keyinput_150), .Z(n15299) );
  XNOR2_X1 U16526 ( .A(n15493), .B(keyinput_149), .ZN(n15298) );
  XNOR2_X1 U16527 ( .A(SI_9_), .B(keyinput_151), .ZN(n15297) );
  NOR4_X1 U16528 ( .A1(n15300), .A2(n15299), .A3(n15298), .A4(n15297), .ZN(
        n15317) );
  XNOR2_X1 U16529 ( .A(SI_8_), .B(keyinput_152), .ZN(n15316) );
  INV_X1 U16530 ( .A(keyinput_153), .ZN(n15305) );
  AOI22_X1 U16531 ( .A1(SI_6_), .A2(keyinput_154), .B1(n15309), .B2(
        keyinput_157), .ZN(n15303) );
  AOI22_X1 U16532 ( .A1(SI_0_), .A2(keyinput_160), .B1(SI_7_), .B2(
        keyinput_153), .ZN(n15302) );
  AOI22_X1 U16533 ( .A1(SI_4_), .A2(keyinput_156), .B1(SI_5_), .B2(
        keyinput_155), .ZN(n15301) );
  NAND3_X1 U16534 ( .A1(n15303), .A2(n15302), .A3(n15301), .ZN(n15304) );
  AOI21_X1 U16535 ( .B1(n15306), .B2(n15305), .A(n15304), .ZN(n15307) );
  OAI21_X1 U16536 ( .B1(SI_6_), .B2(keyinput_154), .A(n15307), .ZN(n15313) );
  XNOR2_X1 U16537 ( .A(n15308), .B(keyinput_158), .ZN(n15312) );
  OAI22_X1 U16538 ( .A1(n15309), .A2(keyinput_157), .B1(SI_4_), .B2(
        keyinput_156), .ZN(n15311) );
  OAI22_X1 U16539 ( .A1(SI_5_), .A2(keyinput_155), .B1(SI_0_), .B2(
        keyinput_160), .ZN(n15310) );
  NOR4_X1 U16540 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15315) );
  XNOR2_X1 U16541 ( .A(SI_1_), .B(keyinput_159), .ZN(n15314) );
  OAI211_X1 U16542 ( .C1(n15317), .C2(n15316), .A(n15315), .B(n15314), .ZN(
        n15321) );
  XOR2_X1 U16543 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_161), .Z(n15320) );
  XNOR2_X1 U16544 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n15319)
         );
  XNOR2_X1 U16545 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n15318) );
  AOI211_X1 U16546 ( .C1(n15321), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        n15330) );
  XOR2_X1 U16547 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n15327)
         );
  XNOR2_X1 U16548 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n15326)
         );
  XNOR2_X1 U16549 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n15325)
         );
  XNOR2_X1 U16550 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n15323)
         );
  XNOR2_X1 U16551 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n15322)
         );
  NAND2_X1 U16552 ( .A1(n15323), .A2(n15322), .ZN(n15324) );
  OR4_X1 U16553 ( .A1(n15327), .A2(n15326), .A3(n15325), .A4(n15324), .ZN(
        n15329) );
  XNOR2_X1 U16554 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n15328)
         );
  OAI21_X1 U16555 ( .B1(n15330), .B2(n15329), .A(n15328), .ZN(n15334) );
  XOR2_X1 U16556 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .Z(n15333)
         );
  XOR2_X1 U16557 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_171), .Z(n15332) );
  XOR2_X1 U16558 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n15331) );
  AOI211_X1 U16559 ( .C1(n15334), .C2(n15333), .A(n15332), .B(n15331), .ZN(
        n15339) );
  XNOR2_X1 U16560 ( .A(n15532), .B(keyinput_173), .ZN(n15338) );
  XNOR2_X1 U16561 ( .A(n15335), .B(keyinput_174), .ZN(n15337) );
  XNOR2_X1 U16562 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n15336)
         );
  OAI211_X1 U16563 ( .C1(n15339), .C2(n15338), .A(n15337), .B(n15336), .ZN(
        n15342) );
  XNOR2_X1 U16564 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n15341)
         );
  XNOR2_X1 U16565 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n15340)
         );
  NAND3_X1 U16566 ( .A1(n15342), .A2(n15341), .A3(n15340), .ZN(n15348) );
  XNOR2_X1 U16567 ( .A(n15541), .B(keyinput_178), .ZN(n15347) );
  XNOR2_X1 U16568 ( .A(n15543), .B(keyinput_181), .ZN(n15345) );
  XNOR2_X1 U16569 ( .A(n15544), .B(keyinput_179), .ZN(n15344) );
  XNOR2_X1 U16570 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n15343)
         );
  NAND3_X1 U16571 ( .A1(n15345), .A2(n15344), .A3(n15343), .ZN(n15346) );
  AOI21_X1 U16572 ( .B1(n15348), .B2(n15347), .A(n15346), .ZN(n15351) );
  XNOR2_X1 U16573 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n15350)
         );
  XOR2_X1 U16574 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_183), .Z(n15349)
         );
  OAI21_X1 U16575 ( .B1(n15351), .B2(n15350), .A(n15349), .ZN(n15355) );
  XNOR2_X1 U16576 ( .A(P3_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n15354)
         );
  XOR2_X1 U16577 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_185), .Z(n15353)
         );
  XNOR2_X1 U16578 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n15352)
         );
  AOI211_X1 U16579 ( .C1(n15355), .C2(n15354), .A(n15353), .B(n15352), .ZN(
        n15358) );
  XNOR2_X1 U16580 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n15357)
         );
  XNOR2_X1 U16581 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n15356)
         );
  OAI21_X1 U16582 ( .B1(n15358), .B2(n15357), .A(n15356), .ZN(n15366) );
  XOR2_X1 U16583 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .Z(n15365) );
  XOR2_X1 U16584 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_190), .Z(n15364)
         );
  XNOR2_X1 U16585 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n15362) );
  XNOR2_X1 U16586 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n15361) );
  XNOR2_X1 U16587 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n15360)
         );
  XNOR2_X1 U16588 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n15359) );
  NOR4_X1 U16589 ( .A1(n15362), .A2(n15361), .A3(n15360), .A4(n15359), .ZN(
        n15363) );
  NAND4_X1 U16590 ( .A1(n15366), .A2(n15365), .A3(n15364), .A4(n15363), .ZN(
        n15369) );
  XOR2_X1 U16591 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .Z(n15368)
         );
  XOR2_X1 U16592 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n15367)
         );
  NAND3_X1 U16593 ( .A1(n15369), .A2(n15368), .A3(n15367), .ZN(n15372) );
  XOR2_X1 U16594 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n15371)
         );
  XOR2_X1 U16595 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .Z(n15370)
         );
  AOI21_X1 U16596 ( .B1(n15372), .B2(n15371), .A(n15370), .ZN(n15375) );
  XNOR2_X1 U16597 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n15374) );
  XNOR2_X1 U16598 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n15373) );
  OAI21_X1 U16599 ( .B1(n15375), .B2(n15374), .A(n15373), .ZN(n15378) );
  XNOR2_X1 U16600 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .ZN(n15377) );
  XOR2_X1 U16601 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .Z(n15376)
         );
  AOI21_X1 U16602 ( .B1(n15378), .B2(n15377), .A(n15376), .ZN(n15381) );
  XOR2_X1 U16603 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .Z(n15380)
         );
  XNOR2_X1 U16604 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .ZN(n15379) );
  NOR3_X1 U16605 ( .A1(n15381), .A2(n15380), .A3(n15379), .ZN(n15384) );
  XOR2_X1 U16606 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .Z(n15383)
         );
  XNOR2_X1 U16607 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n15382) );
  OAI21_X1 U16608 ( .B1(n15384), .B2(n15383), .A(n15382), .ZN(n15387) );
  XNOR2_X1 U16609 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n15386) );
  XNOR2_X1 U16610 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n15385) );
  NAND3_X1 U16611 ( .A1(n15387), .A2(n15386), .A3(n15385), .ZN(n15400) );
  AOI22_X1 U16612 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput_215), .B1(
        n15389), .B2(keyinput_214), .ZN(n15388) );
  OAI221_X1 U16613 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_215), .C1(
        n15389), .C2(keyinput_214), .A(n15388), .ZN(n15397) );
  INV_X1 U16614 ( .A(keyinput_209), .ZN(n15393) );
  XNOR2_X1 U16615 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n15392) );
  OAI22_X1 U16616 ( .A1(P3_DATAO_REG_14__SCAN_IN), .A2(keyinput_210), .B1(
        P3_DATAO_REG_15__SCAN_IN), .B2(keyinput_209), .ZN(n15390) );
  AOI21_X1 U16617 ( .B1(keyinput_210), .B2(P3_DATAO_REG_14__SCAN_IN), .A(
        n15390), .ZN(n15391) );
  OAI211_X1 U16618 ( .C1(n15393), .C2(n15596), .A(n15392), .B(n15391), .ZN(
        n15396) );
  XNOR2_X1 U16619 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n15395) );
  XNOR2_X1 U16620 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n15394) );
  NOR4_X1 U16621 ( .A1(n15397), .A2(n15396), .A3(n15395), .A4(n15394), .ZN(
        n15399) );
  XOR2_X1 U16622 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .Z(n15398)
         );
  AOI21_X1 U16623 ( .B1(n15400), .B2(n15399), .A(n15398), .ZN(n15404) );
  XOR2_X1 U16624 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .Z(n15403)
         );
  XNOR2_X1 U16625 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_219), .ZN(n15402)
         );
  XNOR2_X1 U16626 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n15401)
         );
  OAI211_X1 U16627 ( .C1(n15404), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        n15407) );
  XNOR2_X1 U16628 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_220), .ZN(n15406)
         );
  XNOR2_X1 U16629 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n15405)
         );
  NAND3_X1 U16630 ( .A1(n15407), .A2(n15406), .A3(n15405), .ZN(n15411) );
  XNOR2_X1 U16631 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_222), .ZN(n15410)
         );
  XOR2_X1 U16632 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_223), .Z(n15409)
         );
  XNOR2_X1 U16633 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_224), .ZN(n15408)
         );
  AOI211_X1 U16634 ( .C1(n15411), .C2(n15410), .A(n15409), .B(n15408), .ZN(
        n15415) );
  XNOR2_X1 U16635 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_227), .ZN(n15414)
         );
  XNOR2_X1 U16636 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_225), .ZN(n15413)
         );
  XNOR2_X1 U16637 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_226), .ZN(n15412)
         );
  NOR4_X1 U16638 ( .A1(n15415), .A2(n15414), .A3(n15413), .A4(n15412), .ZN(
        n15418) );
  XOR2_X1 U16639 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_228), .Z(n15417) );
  XOR2_X1 U16640 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_229), .Z(n15416) );
  OAI21_X1 U16641 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15421) );
  XOR2_X1 U16642 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_230), .Z(n15420) );
  XNOR2_X1 U16643 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_231), .ZN(n15419)
         );
  NAND3_X1 U16644 ( .A1(n15421), .A2(n15420), .A3(n15419), .ZN(n15425) );
  XOR2_X1 U16645 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_232), .Z(n15424) );
  XNOR2_X1 U16646 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n15423)
         );
  XNOR2_X1 U16647 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_233), .ZN(n15422)
         );
  AOI211_X1 U16648 ( .C1(n15425), .C2(n15424), .A(n15423), .B(n15422), .ZN(
        n15436) );
  XOR2_X1 U16649 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .Z(n15429) );
  XOR2_X1 U16650 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .Z(n15428) );
  XNOR2_X1 U16651 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_237), .ZN(n15427) );
  XNOR2_X1 U16652 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_235), .ZN(n15426) );
  NAND4_X1 U16653 ( .A1(n15429), .A2(n15428), .A3(n15427), .A4(n15426), .ZN(
        n15435) );
  XOR2_X1 U16654 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_242), .Z(n15433) );
  XNOR2_X1 U16655 ( .A(n15637), .B(keyinput_240), .ZN(n15432) );
  XNOR2_X1 U16656 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n15431) );
  XNOR2_X1 U16657 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n15430) );
  NOR4_X1 U16658 ( .A1(n15433), .A2(n15432), .A3(n15431), .A4(n15430), .ZN(
        n15434) );
  OAI21_X1 U16659 ( .B1(n15436), .B2(n15435), .A(n15434), .ZN(n15444) );
  XNOR2_X1 U16660 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_243), .ZN(n15443) );
  XNOR2_X1 U16661 ( .A(n15437), .B(keyinput_246), .ZN(n15441) );
  XNOR2_X1 U16662 ( .A(n15438), .B(keyinput_245), .ZN(n15440) );
  XNOR2_X1 U16663 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n15439) );
  NAND3_X1 U16664 ( .A1(n15441), .A2(n15440), .A3(n15439), .ZN(n15442) );
  AOI21_X1 U16665 ( .B1(n15444), .B2(n15443), .A(n15442), .ZN(n15448) );
  XNOR2_X1 U16666 ( .A(n15651), .B(keyinput_247), .ZN(n15447) );
  XNOR2_X1 U16667 ( .A(n15652), .B(keyinput_248), .ZN(n15446) );
  XNOR2_X1 U16668 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_249), .ZN(n15445)
         );
  NOR4_X1 U16669 ( .A1(n15448), .A2(n15447), .A3(n15446), .A4(n15445), .ZN(
        n15455) );
  XNOR2_X1 U16670 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_250), .ZN(n15454)
         );
  XOR2_X1 U16671 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .Z(n15452) );
  XNOR2_X1 U16672 ( .A(n15449), .B(keyinput_251), .ZN(n15451) );
  XNOR2_X1 U16673 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_252), .ZN(n15450)
         );
  NOR3_X1 U16674 ( .A1(n15452), .A2(n15451), .A3(n15450), .ZN(n15453) );
  OAI21_X1 U16675 ( .B1(n15455), .B2(n15454), .A(n15453), .ZN(n15669) );
  XNOR2_X1 U16676 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n15668)
         );
  XOR2_X1 U16677 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n15458) );
  XOR2_X1 U16678 ( .A(SI_31_), .B(keyinput_1), .Z(n15457) );
  XOR2_X1 U16679 ( .A(SI_30_), .B(keyinput_2), .Z(n15456) );
  AOI21_X1 U16680 ( .B1(n15458), .B2(n15457), .A(n15456), .ZN(n15465) );
  XNOR2_X1 U16681 ( .A(n15459), .B(keyinput_4), .ZN(n15464) );
  XNOR2_X1 U16682 ( .A(n15460), .B(keyinput_3), .ZN(n15463) );
  XNOR2_X1 U16683 ( .A(n15461), .B(keyinput_5), .ZN(n15462) );
  NOR4_X1 U16684 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        n15470) );
  XNOR2_X1 U16685 ( .A(SI_26_), .B(keyinput_6), .ZN(n15469) );
  XOR2_X1 U16686 ( .A(SI_24_), .B(keyinput_8), .Z(n15468) );
  XNOR2_X1 U16687 ( .A(n15466), .B(keyinput_7), .ZN(n15467) );
  OAI211_X1 U16688 ( .C1(n15470), .C2(n15469), .A(n15468), .B(n15467), .ZN(
        n15473) );
  XNOR2_X1 U16689 ( .A(SI_23_), .B(keyinput_9), .ZN(n15472) );
  XNOR2_X1 U16690 ( .A(SI_22_), .B(keyinput_10), .ZN(n15471) );
  NAND3_X1 U16691 ( .A1(n15473), .A2(n15472), .A3(n15471), .ZN(n15478) );
  XNOR2_X1 U16692 ( .A(n15474), .B(keyinput_13), .ZN(n15477) );
  XOR2_X1 U16693 ( .A(SI_21_), .B(keyinput_11), .Z(n15476) );
  XNOR2_X1 U16694 ( .A(SI_20_), .B(keyinput_12), .ZN(n15475) );
  NAND4_X1 U16695 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        n15486) );
  XNOR2_X1 U16696 ( .A(SI_18_), .B(keyinput_14), .ZN(n15485) );
  XNOR2_X1 U16697 ( .A(n15479), .B(keyinput_16), .ZN(n15483) );
  XNOR2_X1 U16698 ( .A(n15480), .B(keyinput_15), .ZN(n15482) );
  XNOR2_X1 U16699 ( .A(SI_15_), .B(keyinput_17), .ZN(n15481) );
  NAND3_X1 U16700 ( .A1(n15483), .A2(n15482), .A3(n15481), .ZN(n15484) );
  AOI21_X1 U16701 ( .B1(n15486), .B2(n15485), .A(n15484), .ZN(n15492) );
  XNOR2_X1 U16702 ( .A(n15487), .B(keyinput_20), .ZN(n15491) );
  XNOR2_X1 U16703 ( .A(n15488), .B(keyinput_19), .ZN(n15490) );
  XNOR2_X1 U16704 ( .A(SI_14_), .B(keyinput_18), .ZN(n15489) );
  NOR4_X1 U16705 ( .A1(n15492), .A2(n15491), .A3(n15490), .A4(n15489), .ZN(
        n15497) );
  XOR2_X1 U16706 ( .A(SI_9_), .B(keyinput_23), .Z(n15496) );
  XOR2_X1 U16707 ( .A(SI_10_), .B(keyinput_22), .Z(n15495) );
  XNOR2_X1 U16708 ( .A(n15493), .B(keyinput_21), .ZN(n15494) );
  NOR4_X1 U16709 ( .A1(n15497), .A2(n15496), .A3(n15495), .A4(n15494), .ZN(
        n15511) );
  XOR2_X1 U16710 ( .A(SI_8_), .B(keyinput_24), .Z(n15510) );
  XOR2_X1 U16711 ( .A(SI_6_), .B(keyinput_26), .Z(n15501) );
  XOR2_X1 U16712 ( .A(SI_0_), .B(keyinput_32), .Z(n15500) );
  XOR2_X1 U16713 ( .A(SI_3_), .B(keyinput_29), .Z(n15499) );
  XOR2_X1 U16714 ( .A(SI_5_), .B(keyinput_27), .Z(n15498) );
  NAND4_X1 U16715 ( .A1(n15501), .A2(n15500), .A3(n15499), .A4(n15498), .ZN(
        n15508) );
  XNOR2_X1 U16716 ( .A(n15502), .B(keyinput_31), .ZN(n15507) );
  XNOR2_X1 U16717 ( .A(SI_4_), .B(keyinput_28), .ZN(n15504) );
  XNOR2_X1 U16718 ( .A(SI_2_), .B(keyinput_30), .ZN(n15503) );
  NAND2_X1 U16719 ( .A1(n15504), .A2(n15503), .ZN(n15506) );
  XNOR2_X1 U16720 ( .A(SI_7_), .B(keyinput_25), .ZN(n15505) );
  NOR4_X1 U16721 ( .A1(n15508), .A2(n15507), .A3(n15506), .A4(n15505), .ZN(
        n15509) );
  OAI21_X1 U16722 ( .B1(n15511), .B2(n15510), .A(n15509), .ZN(n15516) );
  XOR2_X1 U16723 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .Z(n15515) );
  XNOR2_X1 U16724 ( .A(n15512), .B(keyinput_35), .ZN(n15514) );
  XNOR2_X1 U16725 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n15513) );
  AOI211_X1 U16726 ( .C1(n15516), .C2(n15515), .A(n15514), .B(n15513), .ZN(
        n15527) );
  XNOR2_X1 U16727 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n15518)
         );
  XNOR2_X1 U16728 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n15517)
         );
  NOR2_X1 U16729 ( .A1(n15518), .A2(n15517), .ZN(n15523) );
  INV_X1 U16730 ( .A(keyinput_39), .ZN(n15519) );
  XNOR2_X1 U16731 ( .A(n15519), .B(P3_REG3_REG_10__SCAN_IN), .ZN(n15522) );
  XNOR2_X1 U16732 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n15521)
         );
  XNOR2_X1 U16733 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n15520)
         );
  NAND4_X1 U16734 ( .A1(n15523), .A2(n15522), .A3(n15521), .A4(n15520), .ZN(
        n15526) );
  XNOR2_X1 U16735 ( .A(n15524), .B(keyinput_41), .ZN(n15525) );
  OAI21_X1 U16736 ( .B1(n15527), .B2(n15526), .A(n15525), .ZN(n15531) );
  XOR2_X1 U16737 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .Z(n15530) );
  XOR2_X1 U16738 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_43), .Z(n15529) );
  XNOR2_X1 U16739 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n15528)
         );
  AOI211_X1 U16740 ( .C1(n15531), .C2(n15530), .A(n15529), .B(n15528), .ZN(
        n15537) );
  XNOR2_X1 U16741 ( .A(n15532), .B(keyinput_45), .ZN(n15536) );
  XNOR2_X1 U16742 ( .A(n15533), .B(keyinput_47), .ZN(n15535) );
  XNOR2_X1 U16743 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n15534)
         );
  OAI211_X1 U16744 ( .C1(n15537), .C2(n15536), .A(n15535), .B(n15534), .ZN(
        n15540) );
  XNOR2_X1 U16745 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n15539)
         );
  XNOR2_X1 U16746 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n15538)
         );
  NAND3_X1 U16747 ( .A1(n15540), .A2(n15539), .A3(n15538), .ZN(n15550) );
  XNOR2_X1 U16748 ( .A(n15541), .B(keyinput_50), .ZN(n15549) );
  XNOR2_X1 U16749 ( .A(n15542), .B(keyinput_52), .ZN(n15547) );
  XNOR2_X1 U16750 ( .A(n15543), .B(keyinput_53), .ZN(n15546) );
  XNOR2_X1 U16751 ( .A(n15544), .B(keyinput_51), .ZN(n15545) );
  NAND3_X1 U16752 ( .A1(n15547), .A2(n15546), .A3(n15545), .ZN(n15548) );
  AOI21_X1 U16753 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15553) );
  XOR2_X1 U16754 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n15552) );
  XNOR2_X1 U16755 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n15551)
         );
  OAI21_X1 U16756 ( .B1(n15553), .B2(n15552), .A(n15551), .ZN(n15558) );
  XNOR2_X1 U16757 ( .A(n15554), .B(keyinput_56), .ZN(n15557) );
  XOR2_X1 U16758 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n15556) );
  XNOR2_X1 U16759 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n15555)
         );
  AOI211_X1 U16760 ( .C1(n15558), .C2(n15557), .A(n15556), .B(n15555), .ZN(
        n15561) );
  XOR2_X1 U16761 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n15560) );
  XNOR2_X1 U16762 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n15559)
         );
  OAI21_X1 U16763 ( .B1(n15561), .B2(n15560), .A(n15559), .ZN(n15570) );
  XOR2_X1 U16764 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_62), .Z(n15569) );
  XOR2_X1 U16765 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_61), .Z(n15568) );
  XOR2_X1 U16766 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n15566)
         );
  XOR2_X1 U16767 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_64), .Z(n15565) );
  XOR2_X1 U16768 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n15564)
         );
  XNOR2_X1 U16769 ( .A(n15562), .B(keyinput_63), .ZN(n15563) );
  NOR4_X1 U16770 ( .A1(n15566), .A2(n15565), .A3(n15564), .A4(n15563), .ZN(
        n15567) );
  NAND4_X1 U16771 ( .A1(n15570), .A2(n15569), .A3(n15568), .A4(n15567), .ZN(
        n15573) );
  XOR2_X1 U16772 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n15572)
         );
  XOR2_X1 U16773 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n15571)
         );
  NAND3_X1 U16774 ( .A1(n15573), .A2(n15572), .A3(n15571), .ZN(n15576) );
  XNOR2_X1 U16775 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n15575)
         );
  XOR2_X1 U16776 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n15574)
         );
  AOI21_X1 U16777 ( .B1(n15576), .B2(n15575), .A(n15574), .ZN(n15579) );
  XNOR2_X1 U16778 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n15578)
         );
  XOR2_X1 U16779 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n15577)
         );
  OAI21_X1 U16780 ( .B1(n15579), .B2(n15578), .A(n15577), .ZN(n15582) );
  XOR2_X1 U16781 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .Z(n15581)
         );
  XOR2_X1 U16782 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n15580)
         );
  AOI21_X1 U16783 ( .B1(n15582), .B2(n15581), .A(n15580), .ZN(n15585) );
  XOR2_X1 U16784 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n15584)
         );
  XOR2_X1 U16785 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .Z(n15583)
         );
  NOR3_X1 U16786 ( .A1(n15585), .A2(n15584), .A3(n15583), .ZN(n15588) );
  XOR2_X1 U16787 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n15587)
         );
  XNOR2_X1 U16788 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n15586)
         );
  OAI21_X1 U16789 ( .B1(n15588), .B2(n15587), .A(n15586), .ZN(n15591) );
  XNOR2_X1 U16790 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n15590)
         );
  XNOR2_X1 U16791 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n15589)
         );
  NAND3_X1 U16792 ( .A1(n15591), .A2(n15590), .A3(n15589), .ZN(n15603) );
  OAI22_X1 U16793 ( .A1(n15594), .A2(keyinput_82), .B1(n15593), .B2(
        keyinput_84), .ZN(n15592) );
  AOI221_X1 U16794 ( .B1(n15594), .B2(keyinput_82), .C1(keyinput_84), .C2(
        n15593), .A(n15592), .ZN(n15602) );
  OAI22_X1 U16795 ( .A1(n15596), .A2(keyinput_81), .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_87), .ZN(n15595) );
  AOI221_X1 U16796 ( .B1(n15596), .B2(keyinput_81), .C1(keyinput_87), .C2(
        P3_DATAO_REG_9__SCAN_IN), .A(n15595), .ZN(n15601) );
  XNOR2_X1 U16797 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n15599)
         );
  XNOR2_X1 U16798 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n15598)
         );
  XNOR2_X1 U16799 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n15597)
         );
  NOR3_X1 U16800 ( .A1(n15599), .A2(n15598), .A3(n15597), .ZN(n15600) );
  NAND4_X1 U16801 ( .A1(n15603), .A2(n15602), .A3(n15601), .A4(n15600), .ZN(
        n15606) );
  XOR2_X1 U16802 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n15605) );
  XOR2_X1 U16803 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n15604) );
  AOI21_X1 U16804 ( .B1(n15606), .B2(n15605), .A(n15604), .ZN(n15612) );
  XNOR2_X1 U16805 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_91), .ZN(n15608)
         );
  XNOR2_X1 U16806 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n15607)
         );
  NAND2_X1 U16807 ( .A1(n15608), .A2(n15607), .ZN(n15611) );
  XOR2_X1 U16808 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .Z(n15610) );
  XNOR2_X1 U16809 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_92), .ZN(n15609)
         );
  OAI211_X1 U16810 ( .C1(n15612), .C2(n15611), .A(n15610), .B(n15609), .ZN(
        n15616) );
  XNOR2_X1 U16811 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_94), .ZN(n15615)
         );
  XNOR2_X1 U16812 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .ZN(n15614)
         );
  XNOR2_X1 U16813 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .ZN(n15613)
         );
  AOI211_X1 U16814 ( .C1(n15616), .C2(n15615), .A(n15614), .B(n15613), .ZN(
        n15620) );
  XOR2_X1 U16815 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .Z(n15619) );
  XNOR2_X1 U16816 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .ZN(n15618)
         );
  XNOR2_X1 U16817 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .ZN(n15617)
         );
  NOR4_X1 U16818 ( .A1(n15620), .A2(n15619), .A3(n15618), .A4(n15617), .ZN(
        n15623) );
  XNOR2_X1 U16819 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_100), .ZN(n15622)
         );
  XNOR2_X1 U16820 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .ZN(n15621)
         );
  OAI21_X1 U16821 ( .B1(n15623), .B2(n15622), .A(n15621), .ZN(n15626) );
  XNOR2_X1 U16822 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .ZN(n15625)
         );
  XNOR2_X1 U16823 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_102), .ZN(n15624)
         );
  NAND3_X1 U16824 ( .A1(n15626), .A2(n15625), .A3(n15624), .ZN(n15630) );
  XNOR2_X1 U16825 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .ZN(n15629)
         );
  XNOR2_X1 U16826 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n15628)
         );
  XNOR2_X1 U16827 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .ZN(n15627)
         );
  AOI211_X1 U16828 ( .C1(n15630), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        n15644) );
  XOR2_X1 U16829 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .Z(n15635) );
  XNOR2_X1 U16830 ( .A(n15631), .B(keyinput_109), .ZN(n15634) );
  XNOR2_X1 U16831 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n15633) );
  XNOR2_X1 U16832 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_107), .ZN(n15632) );
  NAND4_X1 U16833 ( .A1(n15635), .A2(n15634), .A3(n15633), .A4(n15632), .ZN(
        n15643) );
  XNOR2_X1 U16834 ( .A(n15636), .B(keyinput_113), .ZN(n15641) );
  XNOR2_X1 U16835 ( .A(n15637), .B(keyinput_112), .ZN(n15640) );
  XNOR2_X1 U16836 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n15639) );
  XNOR2_X1 U16837 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .ZN(n15638) );
  NOR4_X1 U16838 ( .A1(n15641), .A2(n15640), .A3(n15639), .A4(n15638), .ZN(
        n15642) );
  OAI21_X1 U16839 ( .B1(n15644), .B2(n15643), .A(n15642), .ZN(n15650) );
  XNOR2_X1 U16840 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .ZN(n15649) );
  XNOR2_X1 U16841 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_118), .ZN(n15647)
         );
  XNOR2_X1 U16842 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_116), .ZN(n15646) );
  XNOR2_X1 U16843 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_117), .ZN(n15645)
         );
  NAND3_X1 U16844 ( .A1(n15647), .A2(n15646), .A3(n15645), .ZN(n15648) );
  AOI21_X1 U16845 ( .B1(n15650), .B2(n15649), .A(n15648), .ZN(n15656) );
  XNOR2_X1 U16846 ( .A(n15651), .B(keyinput_119), .ZN(n15655) );
  XNOR2_X1 U16847 ( .A(n15652), .B(keyinput_120), .ZN(n15654) );
  XNOR2_X1 U16848 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_121), .ZN(n15653)
         );
  NOR4_X1 U16849 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        n15662) );
  XNOR2_X1 U16850 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_122), .ZN(n15661)
         );
  XNOR2_X1 U16851 ( .A(n9081), .B(keyinput_124), .ZN(n15659) );
  XNOR2_X1 U16852 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .ZN(n15658)
         );
  XNOR2_X1 U16853 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n15657)
         );
  NOR3_X1 U16854 ( .A1(n15659), .A2(n15658), .A3(n15657), .ZN(n15660) );
  OAI21_X1 U16855 ( .B1(n15662), .B2(n15661), .A(n15660), .ZN(n15666) );
  XNOR2_X1 U16856 ( .A(n15663), .B(keyinput_126), .ZN(n15665) );
  XNOR2_X1 U16857 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_127), .ZN(n15664)
         );
  AOI21_X1 U16858 ( .B1(n15666), .B2(n15665), .A(n15664), .ZN(n15667) );
  AOI211_X1 U16859 ( .C1(n15670), .C2(n15669), .A(n15668), .B(n15667), .ZN(
        n15671) );
  XNOR2_X1 U16860 ( .A(n15672), .B(n15671), .ZN(P1_U3559) );
  OAI211_X1 U16861 ( .C1(n16624), .C2(n15674), .A(n15673), .B(n8390), .ZN(
        n15772) );
  MUX2_X1 U16862 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15772), .S(n16635), .Z(
        P1_U3558) );
  NAND2_X1 U16863 ( .A1(n15675), .A2(n16568), .ZN(n15683) );
  NAND2_X1 U16864 ( .A1(n15677), .A2(n15676), .ZN(n15678) );
  AOI21_X1 U16865 ( .B1(n15679), .B2(n16560), .A(n15678), .ZN(n15680) );
  MUX2_X1 U16866 ( .A(n15773), .B(P1_REG1_REG_29__SCAN_IN), .S(n16633), .Z(
        P1_U3557) );
  NAND3_X1 U16867 ( .A1(n15684), .A2(n16568), .A3(n15092), .ZN(n15689) );
  AOI21_X1 U16868 ( .B1(n15686), .B2(n16560), .A(n15685), .ZN(n15687) );
  NAND3_X1 U16869 ( .A1(n15689), .A2(n15688), .A3(n15687), .ZN(n15774) );
  MUX2_X1 U16870 ( .A(n15774), .B(P1_REG1_REG_28__SCAN_IN), .S(n16633), .Z(
        P1_U3556) );
  AOI21_X1 U16871 ( .B1(n15691), .B2(n16560), .A(n15690), .ZN(n15692) );
  OAI211_X1 U16872 ( .C1(n16628), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        n15775) );
  MUX2_X1 U16873 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15775), .S(n16635), .Z(
        P1_U3555) );
  AOI21_X1 U16874 ( .B1(n15696), .B2(n16560), .A(n15695), .ZN(n15697) );
  OAI211_X1 U16875 ( .C1(n16628), .C2(n15699), .A(n15698), .B(n15697), .ZN(
        n15776) );
  MUX2_X1 U16876 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15776), .S(n16635), .Z(
        P1_U3554) );
  NAND3_X1 U16877 ( .A1(n15701), .A2(n15700), .A3(n16568), .ZN(n15703) );
  OAI211_X1 U16878 ( .C1(n15704), .C2(n16624), .A(n15703), .B(n15702), .ZN(
        n15705) );
  NOR2_X1 U16879 ( .A1(n15706), .A2(n15705), .ZN(n15777) );
  MUX2_X1 U16880 ( .A(n15707), .B(n15777), .S(n16635), .Z(n15708) );
  INV_X1 U16881 ( .A(n15708), .ZN(P1_U3553) );
  AOI211_X1 U16882 ( .C1(n15711), .C2(n16560), .A(n15710), .B(n15709), .ZN(
        n15714) );
  NAND2_X1 U16883 ( .A1(n15712), .A2(n16568), .ZN(n15713) );
  OAI211_X1 U16884 ( .C1(n15715), .C2(n16351), .A(n15714), .B(n15713), .ZN(
        n15780) );
  MUX2_X1 U16885 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15780), .S(n16635), .Z(
        P1_U3552) );
  NAND2_X1 U16886 ( .A1(n15716), .A2(n16631), .ZN(n15723) );
  AOI21_X1 U16887 ( .B1(n15718), .B2(n16560), .A(n15717), .ZN(n15722) );
  NAND3_X1 U16888 ( .A1(n8166), .A2(n15719), .A3(n16568), .ZN(n15721) );
  NAND4_X1 U16889 ( .A1(n15723), .A2(n15722), .A3(n15721), .A4(n15720), .ZN(
        n15781) );
  MUX2_X1 U16890 ( .A(n15781), .B(P1_REG1_REG_23__SCAN_IN), .S(n16633), .Z(
        P1_U3551) );
  AOI211_X1 U16891 ( .C1(n15726), .C2(n16560), .A(n15725), .B(n15724), .ZN(
        n15727) );
  OAI21_X1 U16892 ( .B1(n16628), .B2(n15728), .A(n15727), .ZN(n15782) );
  MUX2_X1 U16893 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15782), .S(n16635), .Z(
        P1_U3550) );
  INV_X1 U16894 ( .A(n15729), .ZN(n15733) );
  NAND2_X1 U16895 ( .A1(n15730), .A2(n16568), .ZN(n15732) );
  OAI211_X1 U16896 ( .C1(n15733), .C2(n16624), .A(n15732), .B(n15731), .ZN(
        n15734) );
  NOR2_X1 U16897 ( .A1(n15735), .A2(n15734), .ZN(n15783) );
  MUX2_X1 U16898 ( .A(n15736), .B(n15783), .S(n16635), .Z(n15737) );
  INV_X1 U16899 ( .A(n15737), .ZN(P1_U3549) );
  AOI21_X1 U16900 ( .B1(n15739), .B2(n16560), .A(n15738), .ZN(n15744) );
  NAND3_X1 U16901 ( .A1(n15741), .A2(n15740), .A3(n16568), .ZN(n15743) );
  NAND4_X1 U16902 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        n15786) );
  MUX2_X1 U16903 ( .A(n15786), .B(P1_REG1_REG_20__SCAN_IN), .S(n16633), .Z(
        P1_U3548) );
  AOI211_X1 U16904 ( .C1(n15748), .C2(n16560), .A(n15747), .B(n15746), .ZN(
        n15749) );
  OAI21_X1 U16905 ( .B1(n16628), .B2(n15750), .A(n15749), .ZN(n15787) );
  MUX2_X1 U16906 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15787), .S(n16635), .Z(
        P1_U3547) );
  AOI211_X1 U16907 ( .C1(n15753), .C2(n16560), .A(n15752), .B(n15751), .ZN(
        n15754) );
  OAI21_X1 U16908 ( .B1(n16628), .B2(n15755), .A(n15754), .ZN(n15788) );
  MUX2_X1 U16909 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15788), .S(n16635), .Z(
        P1_U3546) );
  AOI21_X1 U16910 ( .B1(n15757), .B2(n16560), .A(n15756), .ZN(n15758) );
  OAI211_X1 U16911 ( .C1(n16628), .C2(n15760), .A(n15759), .B(n15758), .ZN(
        n15789) );
  MUX2_X1 U16912 ( .A(n15789), .B(P1_REG1_REG_17__SCAN_IN), .S(n16633), .Z(
        P1_U3545) );
  AOI21_X1 U16913 ( .B1(n15762), .B2(n16560), .A(n15761), .ZN(n15763) );
  OAI21_X1 U16914 ( .B1(n15764), .B2(n16566), .A(n15763), .ZN(n15765) );
  AOI21_X1 U16915 ( .B1(n15766), .B2(n16568), .A(n15765), .ZN(n15767) );
  OAI21_X1 U16916 ( .B1(n15768), .B2(n16351), .A(n15767), .ZN(n15790) );
  MUX2_X1 U16917 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15790), .S(n16635), .Z(
        P1_U3544) );
  MUX2_X1 U16918 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15769), .S(n16635), .Z(
        P1_U3539) );
  NAND2_X1 U16919 ( .A1(n16636), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n15770) );
  OAI21_X1 U16920 ( .B1(n15771), .B2(n16636), .A(n15770), .ZN(P1_U3527) );
  MUX2_X1 U16921 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15772), .S(n16638), .Z(
        P1_U3526) );
  MUX2_X1 U16922 ( .A(n15774), .B(P1_REG0_REG_28__SCAN_IN), .S(n16636), .Z(
        P1_U3524) );
  MUX2_X1 U16923 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15775), .S(n16638), .Z(
        P1_U3523) );
  MUX2_X1 U16924 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15776), .S(n16638), .Z(
        P1_U3522) );
  MUX2_X1 U16925 ( .A(n15778), .B(n15777), .S(n16638), .Z(n15779) );
  INV_X1 U16926 ( .A(n15779), .ZN(P1_U3521) );
  MUX2_X1 U16927 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15780), .S(n16638), .Z(
        P1_U3520) );
  MUX2_X1 U16928 ( .A(n15781), .B(P1_REG0_REG_23__SCAN_IN), .S(n16636), .Z(
        P1_U3519) );
  MUX2_X1 U16929 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15782), .S(n16638), .Z(
        P1_U3518) );
  INV_X1 U16930 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15784) );
  MUX2_X1 U16931 ( .A(n15784), .B(n15783), .S(n16638), .Z(n15785) );
  INV_X1 U16932 ( .A(n15785), .ZN(P1_U3517) );
  MUX2_X1 U16933 ( .A(n15786), .B(P1_REG0_REG_20__SCAN_IN), .S(n16636), .Z(
        P1_U3516) );
  MUX2_X1 U16934 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15787), .S(n16638), .Z(
        P1_U3515) );
  MUX2_X1 U16935 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15788), .S(n16638), .Z(
        P1_U3513) );
  MUX2_X1 U16936 ( .A(n15789), .B(P1_REG0_REG_17__SCAN_IN), .S(n16636), .Z(
        P1_U3510) );
  MUX2_X1 U16937 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15790), .S(n16638), .Z(
        P1_U3507) );
  NOR4_X1 U16938 ( .A1(n15792), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7761), .A4(
        P1_U3086), .ZN(n15793) );
  AOI21_X1 U16939 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15802), .A(n15793), 
        .ZN(n15794) );
  OAI21_X1 U16940 ( .B1(n15795), .B2(n15805), .A(n15794), .ZN(P1_U3324) );
  INV_X1 U16941 ( .A(n15796), .ZN(n15797) );
  OAI222_X1 U16942 ( .A1(n15810), .A2(n15798), .B1(n15805), .B2(n15797), .C1(
        n9908), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U16943 ( .A1(n15802), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n15800) );
  OAI211_X1 U16944 ( .C1(n15801), .C2(n15805), .A(n15800), .B(n15799), .ZN(
        P1_U3328) );
  AOI22_X1 U16945 ( .A1(n15803), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n15802), .ZN(n15804) );
  OAI21_X1 U16946 ( .B1(n15806), .B2(n15805), .A(n15804), .ZN(P1_U3329) );
  OAI222_X1 U16947 ( .A1(n15810), .A2(n15809), .B1(n15805), .B2(n15808), .C1(
        P1_U3086), .C2(n15807), .ZN(P1_U3330) );
  MUX2_X1 U16948 ( .A(n15811), .B(n9824), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16949 ( .A(n15812), .ZN(n15813) );
  MUX2_X1 U16950 ( .A(n15813), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16951 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15814), .ZN(P1_U3323) );
  AND2_X1 U16952 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15814), .ZN(P1_U3322) );
  AND2_X1 U16953 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15814), .ZN(P1_U3321) );
  AND2_X1 U16954 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15814), .ZN(P1_U3320) );
  AND2_X1 U16955 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15814), .ZN(P1_U3319) );
  AND2_X1 U16956 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15814), .ZN(P1_U3318) );
  AND2_X1 U16957 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15814), .ZN(P1_U3317) );
  AND2_X1 U16958 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15814), .ZN(P1_U3316) );
  AND2_X1 U16959 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15814), .ZN(P1_U3315) );
  AND2_X1 U16960 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15814), .ZN(P1_U3314) );
  AND2_X1 U16961 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15814), .ZN(P1_U3313) );
  AND2_X1 U16962 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15814), .ZN(P1_U3312) );
  AND2_X1 U16963 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15814), .ZN(P1_U3311) );
  AND2_X1 U16964 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15814), .ZN(P1_U3310) );
  AND2_X1 U16965 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15814), .ZN(P1_U3309) );
  AND2_X1 U16966 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15814), .ZN(P1_U3308) );
  AND2_X1 U16967 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15814), .ZN(P1_U3307) );
  AND2_X1 U16968 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15814), .ZN(P1_U3306) );
  AND2_X1 U16969 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15814), .ZN(P1_U3305) );
  AND2_X1 U16970 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15814), .ZN(P1_U3304) );
  AND2_X1 U16971 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15814), .ZN(P1_U3303) );
  AND2_X1 U16972 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15814), .ZN(P1_U3302) );
  AND2_X1 U16973 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15814), .ZN(P1_U3301) );
  AND2_X1 U16974 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15814), .ZN(P1_U3300) );
  AND2_X1 U16975 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15814), .ZN(P1_U3299) );
  AND2_X1 U16976 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15814), .ZN(P1_U3298) );
  AND2_X1 U16977 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15814), .ZN(P1_U3297) );
  AND2_X1 U16978 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15814), .ZN(P1_U3296) );
  AND2_X1 U16979 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15814), .ZN(P1_U3295) );
  AND2_X1 U16980 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15814), .ZN(P1_U3294) );
  INV_X1 U16981 ( .A(n15815), .ZN(n15816) );
  AOI21_X1 U16982 ( .B1(n15817), .B2(n15820), .A(n15816), .ZN(P2_U3417) );
  AND2_X1 U16983 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15819), .ZN(P2_U3295) );
  AND2_X1 U16984 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15819), .ZN(P2_U3294) );
  AND2_X1 U16985 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15819), .ZN(P2_U3293) );
  AND2_X1 U16986 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15819), .ZN(P2_U3292) );
  AND2_X1 U16987 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15819), .ZN(P2_U3291) );
  AND2_X1 U16988 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15819), .ZN(P2_U3290) );
  AND2_X1 U16989 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15819), .ZN(P2_U3289) );
  AND2_X1 U16990 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15819), .ZN(P2_U3288) );
  AND2_X1 U16991 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15819), .ZN(P2_U3287) );
  AND2_X1 U16992 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15819), .ZN(P2_U3286) );
  AND2_X1 U16993 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15819), .ZN(P2_U3285) );
  AND2_X1 U16994 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15819), .ZN(P2_U3284) );
  AND2_X1 U16995 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15819), .ZN(P2_U3283) );
  AND2_X1 U16996 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15819), .ZN(P2_U3282) );
  AND2_X1 U16997 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15819), .ZN(P2_U3281) );
  AND2_X1 U16998 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15819), .ZN(P2_U3280) );
  AND2_X1 U16999 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15819), .ZN(P2_U3279) );
  AND2_X1 U17000 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15819), .ZN(P2_U3278) );
  AND2_X1 U17001 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15819), .ZN(P2_U3277) );
  AND2_X1 U17002 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15819), .ZN(P2_U3276) );
  AND2_X1 U17003 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15819), .ZN(P2_U3275) );
  AND2_X1 U17004 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15819), .ZN(P2_U3274) );
  AND2_X1 U17005 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15819), .ZN(P2_U3273) );
  AND2_X1 U17006 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15819), .ZN(P2_U3272) );
  AND2_X1 U17007 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15819), .ZN(P2_U3271) );
  AND2_X1 U17008 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15819), .ZN(P2_U3270) );
  AND2_X1 U17009 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15819), .ZN(P2_U3269) );
  AND2_X1 U17010 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15819), .ZN(P2_U3268) );
  AND2_X1 U17011 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15819), .ZN(P2_U3267) );
  AND2_X1 U17012 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15819), .ZN(P2_U3266) );
  NOR2_X1 U17013 ( .A1(n15880), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17014 ( .A1(P3_U3897), .A2(n16252), .ZN(P3_U3150) );
  INV_X1 U17015 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15821) );
  AOI22_X1 U17016 ( .A1(n15823), .A2(n15822), .B1(n15821), .B2(n15820), .ZN(
        P2_U3416) );
  AOI22_X1 U17017 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15920), .B1(n15924), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n15827) );
  AOI22_X1 U17018 ( .A1(n15880), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15826) );
  OAI22_X1 U17019 ( .A1(n15903), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15897), .ZN(n15824) );
  OAI21_X1 U17020 ( .B1(n15922), .B2(n15824), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15825) );
  OAI211_X1 U17021 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15827), .A(n15826), .B(
        n15825), .ZN(P2_U3214) );
  OAI21_X1 U17022 ( .B1(n15830), .B2(n15829), .A(n15828), .ZN(n15835) );
  NOR2_X1 U17023 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12053), .ZN(n15831) );
  AOI21_X1 U17024 ( .B1(n15922), .B2(n15832), .A(n15831), .ZN(n15834) );
  NAND2_X1 U17025 ( .A1(n15880), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n15833) );
  OAI211_X1 U17026 ( .C1(n15897), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        n15836) );
  INV_X1 U17027 ( .A(n15836), .ZN(n15842) );
  AOI211_X1 U17028 ( .C1(n15839), .C2(n15838), .A(n15837), .B(n15903), .ZN(
        n15840) );
  INV_X1 U17029 ( .A(n15840), .ZN(n15841) );
  NAND2_X1 U17030 ( .A1(n15842), .A2(n15841), .ZN(P2_U3215) );
  AOI22_X1 U17031 ( .A1(n15880), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15856) );
  OAI21_X1 U17032 ( .B1(n15845), .B2(n15844), .A(n15843), .ZN(n15848) );
  NAND2_X1 U17033 ( .A1(n15922), .A2(n15846), .ZN(n15847) );
  OAI21_X1 U17034 ( .B1(n15897), .B2(n15848), .A(n15847), .ZN(n15849) );
  INV_X1 U17035 ( .A(n15849), .ZN(n15855) );
  AOI211_X1 U17036 ( .C1(n15852), .C2(n15851), .A(n15850), .B(n15903), .ZN(
        n15853) );
  INV_X1 U17037 ( .A(n15853), .ZN(n15854) );
  NAND3_X1 U17038 ( .A1(n15856), .A2(n15855), .A3(n15854), .ZN(P2_U3216) );
  AOI22_X1 U17039 ( .A1(n15880), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n15866) );
  XNOR2_X1 U17040 ( .A(n15858), .B(n15857), .ZN(n15860) );
  AOI22_X1 U17041 ( .A1(n15924), .A2(n15860), .B1(n15859), .B2(n15922), .ZN(
        n15865) );
  OAI211_X1 U17042 ( .C1(n15863), .C2(n15862), .A(n15861), .B(n15920), .ZN(
        n15864) );
  NAND3_X1 U17043 ( .A1(n15866), .A2(n15865), .A3(n15864), .ZN(P2_U3228) );
  INV_X1 U17044 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n16066) );
  NOR2_X1 U17045 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15867), .ZN(n15873) );
  OAI211_X1 U17046 ( .C1(n15870), .C2(n15869), .A(n15868), .B(n15924), .ZN(
        n15871) );
  INV_X1 U17047 ( .A(n15871), .ZN(n15872) );
  AOI211_X1 U17048 ( .C1(n15922), .C2(n15874), .A(n15873), .B(n15872), .ZN(
        n15879) );
  XOR2_X1 U17049 ( .A(n15876), .B(n15875), .Z(n15877) );
  NAND2_X1 U17050 ( .A1(n15877), .A2(n15920), .ZN(n15878) );
  OAI211_X1 U17051 ( .C1(n15928), .C2(n16066), .A(n15879), .B(n15878), .ZN(
        P2_U3230) );
  AOI22_X1 U17052 ( .A1(n15880), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(P2_U3088), .ZN(n15891) );
  OAI21_X1 U17053 ( .B1(n15883), .B2(n15882), .A(n15881), .ZN(n15884) );
  NAND2_X1 U17054 ( .A1(n15884), .A2(n15924), .ZN(n15890) );
  NAND2_X1 U17055 ( .A1(n15922), .A2(n15885), .ZN(n15889) );
  XOR2_X1 U17056 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n15886), .Z(n15887) );
  NAND2_X1 U17057 ( .A1(n15887), .A2(n15920), .ZN(n15888) );
  NAND4_X1 U17058 ( .A1(n15891), .A2(n15890), .A3(n15889), .A4(n15888), .ZN(
        P2_U3232) );
  INV_X1 U17059 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n16028) );
  INV_X1 U17060 ( .A(n15892), .ZN(n15895) );
  AOI21_X1 U17061 ( .B1(n15896), .B2(P2_REG2_REG_12__SCAN_IN), .A(n15893), 
        .ZN(n15894) );
  OAI211_X1 U17062 ( .C1(P2_REG2_REG_12__SCAN_IN), .C2(n15896), .A(n15895), 
        .B(n15894), .ZN(n15898) );
  AOI21_X1 U17063 ( .B1(n15899), .B2(n15898), .A(n15897), .ZN(n15907) );
  INV_X1 U17064 ( .A(n15900), .ZN(n15905) );
  NAND2_X1 U17065 ( .A1(n15908), .A2(n16515), .ZN(n15901) );
  OAI211_X1 U17066 ( .C1(n15908), .C2(n16515), .A(n15902), .B(n15901), .ZN(
        n15904) );
  AOI21_X1 U17067 ( .B1(n15905), .B2(n15904), .A(n15903), .ZN(n15906) );
  AOI211_X1 U17068 ( .C1(n15922), .C2(n15908), .A(n15907), .B(n15906), .ZN(
        n15910) );
  OAI211_X1 U17069 ( .C1(n16028), .C2(n15928), .A(n15910), .B(n15909), .ZN(
        P2_U3226) );
  INV_X1 U17070 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n16001) );
  INV_X1 U17071 ( .A(n15911), .ZN(n15916) );
  OAI21_X1 U17072 ( .B1(n15914), .B2(n15913), .A(n15912), .ZN(n15915) );
  NAND2_X1 U17073 ( .A1(n15916), .A2(n15915), .ZN(n15925) );
  OAI21_X1 U17074 ( .B1(n15919), .B2(n15918), .A(n15917), .ZN(n15921) );
  AOI222_X1 U17075 ( .A1(n15925), .A2(n15924), .B1(n15923), .B2(n15922), .C1(
        n15921), .C2(n15920), .ZN(n15927) );
  OAI211_X1 U17076 ( .C1(n16001), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P2_U3223) );
  AOI21_X1 U17077 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n16105), .A(n15934), .ZN(
        n15930) );
  INV_X1 U17078 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15929) );
  AOI21_X1 U17079 ( .B1(n15930), .B2(n15929), .A(n16096), .ZN(SUB_1596_U53) );
  XNOR2_X1 U17080 ( .A(n15935), .B(n15934), .ZN(n16097) );
  NOR2_X1 U17081 ( .A1(n16096), .A2(n16097), .ZN(n15932) );
  INV_X1 U17082 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15931) );
  NAND2_X1 U17083 ( .A1(n16096), .A2(n16097), .ZN(n16095) );
  OAI21_X1 U17084 ( .B1(n15932), .B2(n15931), .A(n16095), .ZN(n15933) );
  INV_X1 U17085 ( .A(n15933), .ZN(n15938) );
  XOR2_X1 U17086 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15944), .Z(n15937) );
  AND2_X1 U17087 ( .A1(n15938), .A2(n15937), .ZN(n15942) );
  NOR2_X1 U17088 ( .A1(n15942), .A2(n15940), .ZN(n15939) );
  XOR2_X1 U17089 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n15939), .Z(SUB_1596_U61) );
  NOR2_X1 U17090 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n15940), .ZN(n15941) );
  NOR2_X1 U17091 ( .A1(n15942), .A2(n15941), .ZN(n15952) );
  NAND2_X1 U17092 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n15943), .ZN(n15945) );
  XNOR2_X1 U17093 ( .A(n15947), .B(n15948), .ZN(n15951) );
  XNOR2_X1 U17094 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15953), .ZN(SUB_1596_U60)
         );
  NAND2_X1 U17095 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15946), .ZN(n15949) );
  NOR2_X1 U17096 ( .A1(n15952), .A2(n15951), .ZN(n15955) );
  NOR2_X1 U17097 ( .A1(n15955), .A2(n15954), .ZN(n15957) );
  XOR2_X1 U17098 ( .A(n15958), .B(n15957), .Z(SUB_1596_U59) );
  NAND2_X1 U17099 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15956), .ZN(n15959) );
  NAND2_X1 U17100 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15960), .ZN(n15963) );
  NAND2_X1 U17101 ( .A1(n15961), .A2(n15950), .ZN(n15962) );
  NAND2_X1 U17102 ( .A1(n15963), .A2(n15962), .ZN(n15968) );
  NOR2_X1 U17103 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15971), .ZN(n15964) );
  AOI21_X1 U17104 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(n15971), .A(n15964), .ZN(
        n15969) );
  XNOR2_X1 U17105 ( .A(n15968), .B(n15969), .ZN(n15965) );
  XNOR2_X1 U17106 ( .A(n15966), .B(n15965), .ZN(n15967) );
  XNOR2_X1 U17107 ( .A(n15967), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  INV_X1 U17108 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n16093) );
  NAND2_X1 U17109 ( .A1(n15969), .A2(n15968), .ZN(n15970) );
  XNOR2_X1 U17110 ( .A(n16123), .B(n15972), .ZN(n15974) );
  XNOR2_X1 U17111 ( .A(n15973), .B(n15974), .ZN(n16091) );
  XNOR2_X1 U17112 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n15981), .ZN(n15983) );
  NAND2_X1 U17113 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n15972), .ZN(n15976) );
  NAND2_X1 U17114 ( .A1(n15974), .A2(n15973), .ZN(n15975) );
  XNOR2_X1 U17115 ( .A(n15978), .B(n15979), .ZN(n15982) );
  XNOR2_X1 U17116 ( .A(n15983), .B(n15982), .ZN(SUB_1596_U56) );
  NAND2_X1 U17117 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15977), .ZN(n15980) );
  XNOR2_X1 U17118 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n15993), .ZN(n15987) );
  NOR2_X1 U17119 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15981), .ZN(n15985) );
  NOR2_X1 U17120 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  XNOR2_X1 U17121 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n15988), .ZN(SUB_1596_U55)
         );
  NOR2_X1 U17122 ( .A1(n15987), .A2(n15986), .ZN(n15990) );
  NOR2_X1 U17123 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n15991), .ZN(n15995) );
  NOR2_X1 U17124 ( .A1(n15993), .A2(n15992), .ZN(n15994) );
  NAND2_X1 U17125 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16005), .ZN(n15996) );
  OAI21_X1 U17126 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16005), .A(n15996), .ZN(
        n16002) );
  XOR2_X1 U17127 ( .A(n16003), .B(n16002), .Z(n15999) );
  AOI21_X1 U17128 ( .B1(n15998), .B2(n15999), .A(n16000), .ZN(n15997) );
  XNOR2_X1 U17129 ( .A(n15997), .B(n16001), .ZN(SUB_1596_U54) );
  NOR2_X1 U17130 ( .A1(n16003), .A2(n16002), .ZN(n16004) );
  XNOR2_X1 U17131 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n16009) );
  XOR2_X1 U17132 ( .A(n16010), .B(n16009), .Z(n16007) );
  NOR2_X1 U17133 ( .A1(n16015), .A2(n16014), .ZN(n16008) );
  XOR2_X1 U17134 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n16008), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U17135 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n16013) );
  INV_X1 U17136 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n16012) );
  XNOR2_X1 U17137 ( .A(n16013), .B(n16018), .ZN(n16020) );
  AOI21_X1 U17138 ( .B1(n16020), .B2(n16021), .A(n16022), .ZN(n16016) );
  INV_X1 U17139 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n16023) );
  XNOR2_X1 U17140 ( .A(n16016), .B(n16023), .ZN(SUB_1596_U69) );
  XOR2_X1 U17141 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n16031) );
  INV_X1 U17142 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n16133) );
  NOR2_X1 U17143 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n16133), .ZN(n16019) );
  XNOR2_X1 U17144 ( .A(n16031), .B(n16030), .ZN(n16025) );
  NAND2_X1 U17145 ( .A1(n16026), .A2(n16025), .ZN(n16027) );
  OAI21_X1 U17146 ( .B1(n16025), .B2(n16026), .A(n16027), .ZN(n16024) );
  XNOR2_X1 U17147 ( .A(n16024), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U17148 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n16037) );
  XOR2_X1 U17149 ( .A(n16036), .B(n16037), .Z(n16034) );
  XNOR2_X1 U17150 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n16035), .ZN(SUB_1596_U67)
         );
  XNOR2_X1 U17151 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n16046) );
  XOR2_X1 U17152 ( .A(n16045), .B(n16046), .Z(n16041) );
  AOI21_X1 U17153 ( .B1(n16040), .B2(n16041), .A(n16042), .ZN(n16039) );
  INV_X1 U17154 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n16044) );
  XNOR2_X1 U17155 ( .A(n16039), .B(n16044), .ZN(SUB_1596_U66) );
  NAND2_X1 U17156 ( .A1(n16041), .A2(n16040), .ZN(n16043) );
  AOI21_X2 U17157 ( .B1(n16044), .B2(n16043), .A(n16042), .ZN(n16053) );
  INV_X1 U17158 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n16051) );
  XNOR2_X1 U17159 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(n16051), .ZN(n16050) );
  XNOR2_X1 U17160 ( .A(n16050), .B(n16049), .ZN(n16052) );
  AOI21_X1 U17161 ( .B1(n16053), .B2(n16052), .A(n16054), .ZN(n16048) );
  XNOR2_X1 U17162 ( .A(n16048), .B(n12581), .ZN(SUB_1596_U65) );
  XOR2_X1 U17163 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n16057), .Z(n16059) );
  XNOR2_X1 U17164 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n16059), .ZN(n16062) );
  NAND2_X1 U17165 ( .A1(n16053), .A2(n16052), .ZN(n16055) );
  NOR2_X1 U17166 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  AOI21_X1 U17167 ( .B1(n16062), .B2(n16063), .A(n16064), .ZN(n16056) );
  XNOR2_X1 U17168 ( .A(n16056), .B(n16066), .ZN(SUB_1596_U64) );
  NAND2_X1 U17169 ( .A1(n16057), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n16061) );
  INV_X1 U17170 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n16058) );
  NAND2_X1 U17171 ( .A1(n16059), .A2(n16058), .ZN(n16060) );
  NAND2_X1 U17172 ( .A1(n16063), .A2(n16062), .ZN(n16065) );
  XOR2_X1 U17173 ( .A(n16069), .B(n16068), .Z(SUB_1596_U63) );
  NAND2_X1 U17174 ( .A1(n16067), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n16070) );
  NAND2_X1 U17175 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n16071), .ZN(n16074) );
  INV_X1 U17176 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n16242) );
  NAND2_X1 U17177 ( .A1(n16072), .A2(n16242), .ZN(n16073) );
  NAND2_X1 U17178 ( .A1(n16074), .A2(n16073), .ZN(n16080) );
  XNOR2_X1 U17179 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n16081) );
  XOR2_X1 U17180 ( .A(n16080), .B(n16081), .Z(n16077) );
  XOR2_X1 U17181 ( .A(n16075), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  NAND2_X1 U17182 ( .A1(n16075), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U17183 ( .A1(n16077), .A2(n16076), .ZN(n16078) );
  NAND2_X1 U17184 ( .A1(n16079), .A2(n16078), .ZN(n16089) );
  NAND2_X1 U17185 ( .A1(n16081), .A2(n16080), .ZN(n16082) );
  OAI21_X1 U17186 ( .B1(n16083), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n16082), 
        .ZN(n16087) );
  XNOR2_X1 U17187 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n16085) );
  XNOR2_X1 U17188 ( .A(n16085), .B(n16084), .ZN(n16086) );
  XNOR2_X1 U17189 ( .A(n16087), .B(n16086), .ZN(n16088) );
  XNOR2_X1 U17190 ( .A(n16089), .B(n16088), .ZN(SUB_1596_U4) );
  AOI21_X1 U17191 ( .B1(n16092), .B2(n16091), .A(n16090), .ZN(n16094) );
  XNOR2_X1 U17192 ( .A(n16094), .B(n16093), .ZN(SUB_1596_U57) );
  OAI21_X1 U17193 ( .B1(n16097), .B2(n16096), .A(n16095), .ZN(n16098) );
  XNOR2_X1 U17194 ( .A(n16098), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(SUB_1596_U5)
         );
  AOI22_X1 U17195 ( .A1(n16254), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n16104) );
  NAND3_X1 U17196 ( .A1(n16250), .A2(n16116), .A3(n16190), .ZN(n16102) );
  OAI21_X1 U17197 ( .B1(n16100), .B2(P3_IR_REG_0__SCAN_IN), .A(n16099), .ZN(
        n16101) );
  NAND2_X1 U17198 ( .A1(n16102), .A2(n16101), .ZN(n16103) );
  OAI211_X1 U17199 ( .C1(n16241), .C2(n16105), .A(n16104), .B(n16103), .ZN(
        P3_U3182) );
  XNOR2_X1 U17200 ( .A(n16107), .B(n16106), .ZN(n16120) );
  INV_X1 U17201 ( .A(n16190), .ZN(n16261) );
  NOR2_X1 U17202 ( .A1(n16244), .A2(n16108), .ZN(n16119) );
  INV_X1 U17203 ( .A(n16109), .ZN(n16110) );
  AOI21_X1 U17204 ( .B1(n16112), .B2(n16111), .A(n16110), .ZN(n16117) );
  XOR2_X1 U17205 ( .A(n16114), .B(n16113), .Z(n16115) );
  OAI22_X1 U17206 ( .A1(n16117), .A2(n16250), .B1(n16116), .B2(n16115), .ZN(
        n16118) );
  AOI211_X1 U17207 ( .C1(n16120), .C2(n16261), .A(n16119), .B(n16118), .ZN(
        n16122) );
  OAI211_X1 U17208 ( .C1(n16241), .C2(n16123), .A(n16122), .B(n16121), .ZN(
        P3_U3188) );
  AOI21_X1 U17209 ( .B1(n16126), .B2(n16125), .A(n16124), .ZN(n16140) );
  OAI21_X1 U17210 ( .B1(n16128), .B2(P3_REG1_REG_11__SCAN_IN), .A(n16127), 
        .ZN(n16129) );
  AND2_X1 U17211 ( .A1(n16129), .A2(n16262), .ZN(n16137) );
  XOR2_X1 U17212 ( .A(n16130), .B(n16131), .Z(n16132) );
  NOR2_X1 U17213 ( .A1(n16132), .A2(n16190), .ZN(n16136) );
  OAI22_X1 U17214 ( .A1(n16244), .A2(n16134), .B1(n16133), .B2(n16241), .ZN(
        n16135) );
  NOR4_X1 U17215 ( .A1(n16138), .A2(n16137), .A3(n16136), .A4(n16135), .ZN(
        n16139) );
  OAI21_X1 U17216 ( .B1(n16140), .B2(n16250), .A(n16139), .ZN(P3_U3193) );
  AOI21_X1 U17217 ( .B1(n7574), .B2(n16142), .A(n16141), .ZN(n16158) );
  OAI21_X1 U17218 ( .B1(n16145), .B2(n16144), .A(n16143), .ZN(n16146) );
  AND2_X1 U17219 ( .A1(n16146), .A2(n16262), .ZN(n16155) );
  INV_X1 U17220 ( .A(n16147), .ZN(n16148) );
  AOI211_X1 U17221 ( .C1(n16150), .C2(n16149), .A(n16190), .B(n16148), .ZN(
        n16154) );
  INV_X1 U17222 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n16151) );
  OAI22_X1 U17223 ( .A1(n16244), .A2(n16152), .B1(n16151), .B2(n16241), .ZN(
        n16153) );
  NOR4_X1 U17224 ( .A1(n16156), .A2(n16155), .A3(n16154), .A4(n16153), .ZN(
        n16157) );
  OAI21_X1 U17225 ( .B1(n16158), .B2(n16250), .A(n16157), .ZN(P3_U3194) );
  AOI22_X1 U17226 ( .A1(n16254), .A2(n16159), .B1(n16252), .B2(
        P3_ADDR_REG_13__SCAN_IN), .ZN(n16175) );
  OAI21_X1 U17227 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n16161), .A(n16160), 
        .ZN(n16167) );
  NAND2_X1 U17228 ( .A1(n16163), .A2(n16162), .ZN(n16164) );
  AOI21_X1 U17229 ( .B1(n16165), .B2(n16164), .A(n16190), .ZN(n16166) );
  AOI21_X1 U17230 ( .B1(n16167), .B2(n16262), .A(n16166), .ZN(n16174) );
  INV_X1 U17231 ( .A(n16168), .ZN(n16173) );
  OAI221_X1 U17232 ( .B1(n16171), .B2(n16170), .C1(n16171), .C2(n16169), .A(
        n16265), .ZN(n16172) );
  NAND4_X1 U17233 ( .A1(n16175), .A2(n16174), .A3(n16173), .A4(n16172), .ZN(
        P3_U3195) );
  AOI21_X1 U17234 ( .B1(n16178), .B2(n16177), .A(n16176), .ZN(n16196) );
  OAI21_X1 U17235 ( .B1(n16181), .B2(n16180), .A(n16179), .ZN(n16187) );
  INV_X1 U17236 ( .A(n16182), .ZN(n16183) );
  AOI21_X1 U17237 ( .B1(n16252), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n16183), 
        .ZN(n16184) );
  OAI21_X1 U17238 ( .B1(n16244), .B2(n16185), .A(n16184), .ZN(n16186) );
  AOI21_X1 U17239 ( .B1(n16187), .B2(n16262), .A(n16186), .ZN(n16194) );
  AND2_X1 U17240 ( .A1(n16189), .A2(n16188), .ZN(n16191) );
  OR3_X1 U17241 ( .A1(n16192), .A2(n16191), .A3(n16190), .ZN(n16193) );
  AND2_X1 U17242 ( .A1(n16194), .A2(n16193), .ZN(n16195) );
  OAI21_X1 U17243 ( .B1(n16196), .B2(n16250), .A(n16195), .ZN(P3_U3196) );
  AOI22_X1 U17244 ( .A1(n16254), .A2(n16197), .B1(n16252), .B2(
        P3_ADDR_REG_15__SCAN_IN), .ZN(n16212) );
  OAI21_X1 U17245 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n16199), .A(n16198), 
        .ZN(n16204) );
  OAI21_X1 U17246 ( .B1(n16202), .B2(n16201), .A(n16200), .ZN(n16203) );
  AOI22_X1 U17247 ( .A1(n16204), .A2(n16262), .B1(n16261), .B2(n16203), .ZN(
        n16211) );
  INV_X1 U17248 ( .A(n16205), .ZN(n16210) );
  OAI221_X1 U17249 ( .B1(n16208), .B2(n16207), .C1(n16208), .C2(n16206), .A(
        n16265), .ZN(n16209) );
  NAND4_X1 U17250 ( .A1(n16212), .A2(n16211), .A3(n16210), .A4(n16209), .ZN(
        P3_U3197) );
  AOI22_X1 U17251 ( .A1(n16254), .A2(n16213), .B1(n16252), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n16230) );
  OAI21_X1 U17252 ( .B1(n16216), .B2(n16215), .A(n16214), .ZN(n16221) );
  OAI21_X1 U17253 ( .B1(n16219), .B2(n16218), .A(n16217), .ZN(n16220) );
  AOI22_X1 U17254 ( .A1(n16221), .A2(n16261), .B1(n16262), .B2(n16220), .ZN(
        n16229) );
  INV_X1 U17255 ( .A(n16222), .ZN(n16228) );
  INV_X1 U17256 ( .A(n16223), .ZN(n16226) );
  OAI221_X1 U17257 ( .B1(n16226), .B2(n16225), .C1(n16226), .C2(n16224), .A(
        n16265), .ZN(n16227) );
  NAND4_X1 U17258 ( .A1(n16230), .A2(n16229), .A3(n16228), .A4(n16227), .ZN(
        P3_U3198) );
  AOI21_X1 U17259 ( .B1(n16233), .B2(n16232), .A(n16231), .ZN(n16251) );
  OAI21_X1 U17260 ( .B1(n16235), .B2(P3_REG1_REG_17__SCAN_IN), .A(n16234), 
        .ZN(n16236) );
  AND2_X1 U17261 ( .A1(n16262), .A2(n16236), .ZN(n16247) );
  OAI211_X1 U17262 ( .C1(n16239), .C2(n16238), .A(n16261), .B(n16237), .ZN(
        n16240) );
  INV_X1 U17263 ( .A(n16240), .ZN(n16246) );
  OAI22_X1 U17264 ( .A1(n16244), .A2(n16243), .B1(n16242), .B2(n16241), .ZN(
        n16245) );
  NOR4_X1 U17265 ( .A1(n16248), .A2(n16247), .A3(n16246), .A4(n16245), .ZN(
        n16249) );
  OAI21_X1 U17266 ( .B1(n16251), .B2(n16250), .A(n16249), .ZN(P3_U3199) );
  AOI22_X1 U17267 ( .A1(n16254), .A2(n16253), .B1(n16252), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n16271) );
  XNOR2_X1 U17268 ( .A(n16256), .B(n16255), .ZN(n16263) );
  OAI21_X1 U17269 ( .B1(n16259), .B2(n16258), .A(n16257), .ZN(n16260) );
  AOI22_X1 U17270 ( .A1(n16263), .A2(n16262), .B1(n16261), .B2(n16260), .ZN(
        n16270) );
  INV_X1 U17271 ( .A(n16264), .ZN(n16269) );
  OAI221_X1 U17272 ( .B1(n16267), .B2(n7509), .C1(n16267), .C2(n16266), .A(
        n16265), .ZN(n16268) );
  NAND4_X1 U17273 ( .A1(n16271), .A2(n16270), .A3(n16269), .A4(n16268), .ZN(
        P3_U3200) );
  MUX2_X1 U17274 ( .A(n11156), .B(P1_REG2_REG_4__SCAN_IN), .S(n16284), .Z(
        n16272) );
  NAND3_X1 U17275 ( .A1(n16274), .A2(n16273), .A3(n16272), .ZN(n16275) );
  NAND3_X1 U17276 ( .A1(n16277), .A2(n16276), .A3(n16275), .ZN(n16291) );
  MUX2_X1 U17277 ( .A(n11132), .B(P1_REG1_REG_4__SCAN_IN), .S(n16284), .Z(
        n16278) );
  NAND3_X1 U17278 ( .A1(n16280), .A2(n16279), .A3(n16278), .ZN(n16281) );
  NAND3_X1 U17279 ( .A1(n16283), .A2(n16282), .A3(n16281), .ZN(n16290) );
  NAND2_X1 U17280 ( .A1(n16285), .A2(n16284), .ZN(n16289) );
  AND2_X1 U17281 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n16286) );
  AOI21_X1 U17282 ( .B1(n16287), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n16286), .ZN(
        n16288) );
  AND4_X1 U17283 ( .A1(n16291), .A2(n16290), .A3(n16289), .A4(n16288), .ZN(
        n16293) );
  NAND2_X1 U17284 ( .A1(n16293), .A2(n16292), .ZN(P1_U3247) );
  AOI22_X1 U17285 ( .A1(n16638), .A2(n16294), .B1(n9098), .B2(n16636), .ZN(
        P1_U3459) );
  INV_X1 U17286 ( .A(n16295), .ZN(n16298) );
  AOI22_X1 U17287 ( .A1(n16299), .A2(n16298), .B1(n16297), .B2(n16296), .ZN(
        n16301) );
  AOI22_X1 U17288 ( .A1(n16490), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n16398), .ZN(n16300) );
  OAI221_X1 U17289 ( .B1(n16398), .B2(n16302), .C1(n16398), .C2(n16301), .A(
        n16300), .ZN(P1_U3293) );
  AOI211_X1 U17290 ( .C1(n16305), .C2(n16614), .A(n16304), .B(n16303), .ZN(
        n16308) );
  INV_X1 U17291 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n16306) );
  AOI22_X1 U17292 ( .A1(n16615), .A2(n16308), .B1(n16306), .B2(n9060), .ZN(
        P3_U3460) );
  INV_X1 U17293 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16307) );
  AOI22_X1 U17294 ( .A1(n16618), .A2(n16308), .B1(n16307), .B2(n9044), .ZN(
        P3_U3393) );
  XNOR2_X1 U17295 ( .A(n10602), .B(n16309), .ZN(n16321) );
  NOR2_X1 U17296 ( .A1(n16314), .A2(n16310), .ZN(n16311) );
  OR2_X1 U17297 ( .A1(n16343), .A2(n16311), .ZN(n16312) );
  NOR2_X1 U17298 ( .A1(n16566), .A2(n16312), .ZN(n16328) );
  INV_X1 U17299 ( .A(n16328), .ZN(n16313) );
  OAI21_X1 U17300 ( .B1(n16314), .B2(n16624), .A(n16313), .ZN(n16319) );
  XNOR2_X1 U17301 ( .A(n16315), .B(n10602), .ZN(n16318) );
  INV_X1 U17302 ( .A(n16316), .ZN(n16317) );
  OAI21_X1 U17303 ( .B1(n16351), .B2(n16318), .A(n16317), .ZN(n16326) );
  AOI211_X1 U17304 ( .C1(n16568), .C2(n16321), .A(n16319), .B(n16326), .ZN(
        n16320) );
  AOI22_X1 U17305 ( .A1(n16635), .A2(n16320), .B1(n11126), .B2(n16633), .ZN(
        P1_U3529) );
  AOI22_X1 U17306 ( .A1(n16638), .A2(n16320), .B1(n9130), .B2(n16636), .ZN(
        P1_U3462) );
  INV_X1 U17307 ( .A(n16321), .ZN(n16322) );
  AOI21_X1 U17308 ( .B1(n16324), .B2(n16323), .A(n16322), .ZN(n16325) );
  AOI211_X1 U17309 ( .C1(n16327), .C2(n9154), .A(n16326), .B(n16325), .ZN(
        n16330) );
  AOI22_X1 U17310 ( .A1(n16498), .A2(n16328), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n16490), .ZN(n16329) );
  OAI221_X1 U17311 ( .B1(n16398), .B2(n16330), .C1(n7416), .C2(n11150), .A(
        n16329), .ZN(P1_U3292) );
  AOI22_X1 U17312 ( .A1(n16338), .A2(n16615), .B1(n16331), .B2(n16336), .ZN(
        n16332) );
  OAI21_X1 U17313 ( .B1(n16615), .B2(n11766), .A(n16332), .ZN(P3_U3461) );
  NAND2_X1 U17314 ( .A1(n16334), .A2(n16333), .ZN(n16339) );
  AOI222_X1 U17315 ( .A1(n16339), .A2(n16338), .B1(n16337), .B2(
        P3_REG3_REG_2__SCAN_IN), .C1(n16336), .C2(n16335), .ZN(n16341) );
  AOI22_X1 U17316 ( .A1(n14100), .A2(n11775), .B1(n16341), .B2(n16340), .ZN(
        P3_U3231) );
  XNOR2_X1 U17317 ( .A(n16342), .B(n16349), .ZN(n16360) );
  INV_X1 U17318 ( .A(n16343), .ZN(n16346) );
  INV_X1 U17319 ( .A(n16344), .ZN(n16345) );
  INV_X1 U17320 ( .A(n16359), .ZN(n16347) );
  OAI21_X1 U17321 ( .B1(n16348), .B2(n16624), .A(n16347), .ZN(n16356) );
  XNOR2_X1 U17322 ( .A(n16350), .B(n16349), .ZN(n16352) );
  NOR2_X1 U17323 ( .A1(n16352), .A2(n16351), .ZN(n16353) );
  AOI211_X1 U17324 ( .C1(n16370), .C2(n16360), .A(n16354), .B(n16353), .ZN(
        n16364) );
  INV_X1 U17325 ( .A(n16364), .ZN(n16355) );
  AOI211_X1 U17326 ( .C1(n16452), .C2(n16360), .A(n16356), .B(n16355), .ZN(
        n16357) );
  AOI22_X1 U17327 ( .A1(n16635), .A2(n16357), .B1(n11128), .B2(n16633), .ZN(
        P1_U3530) );
  AOI22_X1 U17328 ( .A1(n16638), .A2(n16357), .B1(n9175), .B2(n16636), .ZN(
        P1_U3465) );
  AOI222_X1 U17329 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n16398), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n16490), .C1(n16358), .C2(n16389), .ZN(
        n16363) );
  AOI22_X1 U17330 ( .A1(n16361), .A2(n16360), .B1(n16498), .B2(n16359), .ZN(
        n16362) );
  OAI211_X1 U17331 ( .C1(n16398), .C2(n16364), .A(n16363), .B(n16362), .ZN(
        P1_U3291) );
  AND2_X1 U17332 ( .A1(n16560), .A2(n16365), .ZN(n16366) );
  NOR2_X1 U17333 ( .A1(n16367), .A2(n16366), .ZN(n16372) );
  INV_X1 U17334 ( .A(n16368), .ZN(n16369) );
  OAI21_X1 U17335 ( .B1(n16452), .B2(n16370), .A(n16369), .ZN(n16371) );
  AND3_X1 U17336 ( .A1(n16373), .A2(n16372), .A3(n16371), .ZN(n16375) );
  AOI22_X1 U17337 ( .A1(n16635), .A2(n16375), .B1(n11129), .B2(n16633), .ZN(
        P1_U3531) );
  INV_X1 U17338 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n16374) );
  AOI22_X1 U17339 ( .A1(n16638), .A2(n16375), .B1(n16374), .B2(n16636), .ZN(
        P1_U3468) );
  XNOR2_X1 U17340 ( .A(n16376), .B(n16377), .ZN(n16393) );
  OAI211_X1 U17341 ( .C1(n9860), .C2(n16379), .A(n16378), .B(n16622), .ZN(
        n16391) );
  OAI21_X1 U17342 ( .B1(n9860), .B2(n16624), .A(n16391), .ZN(n16385) );
  XNOR2_X1 U17343 ( .A(n16380), .B(n16381), .ZN(n16383) );
  AOI21_X1 U17344 ( .B1(n16383), .B2(n16631), .A(n16382), .ZN(n16397) );
  INV_X1 U17345 ( .A(n16397), .ZN(n16384) );
  AOI211_X1 U17346 ( .C1(n16393), .C2(n16568), .A(n16385), .B(n16384), .ZN(
        n16387) );
  AOI22_X1 U17347 ( .A1(n16635), .A2(n16387), .B1(n11132), .B2(n16633), .ZN(
        P1_U3532) );
  INV_X1 U17348 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16386) );
  AOI22_X1 U17349 ( .A1(n16638), .A2(n16387), .B1(n16386), .B2(n16636), .ZN(
        P1_U3471) );
  AOI222_X1 U17350 ( .A1(n16390), .A2(n16389), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n16398), .C1(n16490), .C2(n16388), .ZN(n16396) );
  INV_X1 U17351 ( .A(n16391), .ZN(n16392) );
  AOI22_X1 U17352 ( .A1(n16394), .A2(n16393), .B1(n16498), .B2(n16392), .ZN(
        n16395) );
  OAI211_X1 U17353 ( .C1(n16398), .C2(n16397), .A(n16396), .B(n16395), .ZN(
        P1_U3289) );
  INV_X1 U17354 ( .A(n16399), .ZN(n16400) );
  OAI21_X1 U17355 ( .B1(n16401), .B2(n16624), .A(n16400), .ZN(n16403) );
  AOI211_X1 U17356 ( .C1(n16452), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        n16405) );
  AOI22_X1 U17357 ( .A1(n16635), .A2(n16405), .B1(n9250), .B2(n16633), .ZN(
        P1_U3533) );
  AOI22_X1 U17358 ( .A1(n16638), .A2(n16405), .B1(n9255), .B2(n16636), .ZN(
        P1_U3474) );
  INV_X1 U17359 ( .A(n16521), .ZN(n16431) );
  OAI22_X1 U17360 ( .A1(n16407), .A2(n16431), .B1(n16406), .B2(n16609), .ZN(
        n16408) );
  NOR2_X1 U17361 ( .A1(n16409), .A2(n16408), .ZN(n16411) );
  AOI22_X1 U17362 ( .A1(n16615), .A2(n16411), .B1(n11940), .B2(n9060), .ZN(
        P3_U3465) );
  INV_X1 U17363 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n16410) );
  AOI22_X1 U17364 ( .A1(n16618), .A2(n16411), .B1(n16410), .B2(n9044), .ZN(
        P3_U3408) );
  INV_X1 U17365 ( .A(n16412), .ZN(n16416) );
  OAI21_X1 U17366 ( .B1(n7943), .B2(n16624), .A(n16413), .ZN(n16415) );
  AOI211_X1 U17367 ( .C1(n16452), .C2(n16416), .A(n16415), .B(n16414), .ZN(
        n16417) );
  AOI22_X1 U17368 ( .A1(n16635), .A2(n16417), .B1(n11137), .B2(n16633), .ZN(
        P1_U3534) );
  AOI22_X1 U17369 ( .A1(n16638), .A2(n16417), .B1(n9282), .B2(n16636), .ZN(
        P1_U3477) );
  NAND2_X1 U17370 ( .A1(n16419), .A2(n16418), .ZN(n16420) );
  NAND2_X1 U17371 ( .A1(n16421), .A2(n16420), .ZN(n16422) );
  AOI21_X1 U17372 ( .B1(n16423), .B2(n16514), .A(n16422), .ZN(n16424) );
  AND2_X1 U17373 ( .A1(n16425), .A2(n16424), .ZN(n16427) );
  AOI22_X1 U17374 ( .A1(n16591), .A2(n16427), .B1(n16426), .B2(n16589), .ZN(
        P2_U3505) );
  AOI22_X1 U17375 ( .A1(n16595), .A2(n16427), .B1(n10036), .B2(n16592), .ZN(
        P2_U3448) );
  INV_X1 U17376 ( .A(n16432), .ZN(n16429) );
  AND2_X1 U17377 ( .A1(n16429), .A2(n16428), .ZN(n16434) );
  OAI22_X1 U17378 ( .A1(n16432), .A2(n16431), .B1(n16609), .B2(n16430), .ZN(
        n16433) );
  NOR3_X1 U17379 ( .A1(n16435), .A2(n16434), .A3(n16433), .ZN(n16438) );
  INV_X1 U17380 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U17381 ( .A1(n16615), .A2(n16438), .B1(n16436), .B2(n9060), .ZN(
        P3_U3466) );
  INV_X1 U17382 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16437) );
  AOI22_X1 U17383 ( .A1(n16618), .A2(n16438), .B1(n16437), .B2(n9044), .ZN(
        P3_U3411) );
  NOR2_X1 U17384 ( .A1(n16439), .A2(n16609), .ZN(n16441) );
  AOI211_X1 U17385 ( .C1(n16614), .C2(n16442), .A(n16441), .B(n16440), .ZN(
        n16444) );
  AOI22_X1 U17386 ( .A1(n16615), .A2(n16444), .B1(n12104), .B2(n9060), .ZN(
        P3_U3467) );
  INV_X1 U17387 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16443) );
  AOI22_X1 U17388 ( .A1(n16618), .A2(n16444), .B1(n16443), .B2(n9044), .ZN(
        P3_U3414) );
  INV_X1 U17389 ( .A(n16445), .ZN(n16451) );
  INV_X1 U17390 ( .A(n16446), .ZN(n16447) );
  OAI21_X1 U17391 ( .B1(n16448), .B2(n16624), .A(n16447), .ZN(n16450) );
  AOI211_X1 U17392 ( .C1(n16452), .C2(n16451), .A(n16450), .B(n16449), .ZN(
        n16454) );
  AOI22_X1 U17393 ( .A1(n16635), .A2(n16454), .B1(n11141), .B2(n16633), .ZN(
        P1_U3536) );
  INV_X1 U17394 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n16453) );
  AOI22_X1 U17395 ( .A1(n16638), .A2(n16454), .B1(n16453), .B2(n16636), .ZN(
        P1_U3483) );
  INV_X1 U17396 ( .A(n16455), .ZN(n16459) );
  OAI21_X1 U17397 ( .B1(n8299), .B2(n16579), .A(n16456), .ZN(n16458) );
  AOI211_X1 U17398 ( .C1(n16514), .C2(n16459), .A(n16458), .B(n16457), .ZN(
        n16461) );
  AOI22_X1 U17399 ( .A1(n16591), .A2(n16461), .B1(n10068), .B2(n16589), .ZN(
        P2_U3507) );
  INV_X1 U17400 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n16460) );
  AOI22_X1 U17401 ( .A1(n16595), .A2(n16461), .B1(n16460), .B2(n16592), .ZN(
        P2_U3454) );
  NOR2_X1 U17402 ( .A1(n16462), .A2(n16609), .ZN(n16464) );
  AOI211_X1 U17403 ( .C1(n16465), .C2(n16521), .A(n16464), .B(n16463), .ZN(
        n16468) );
  INV_X1 U17404 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16466) );
  AOI22_X1 U17405 ( .A1(n16615), .A2(n16468), .B1(n16466), .B2(n9060), .ZN(
        P3_U3468) );
  INV_X1 U17406 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U17407 ( .A1(n16618), .A2(n16468), .B1(n16467), .B2(n9044), .ZN(
        P3_U3417) );
  NOR2_X1 U17408 ( .A1(n16469), .A2(n16609), .ZN(n16471) );
  AOI211_X1 U17409 ( .C1(n16521), .C2(n16472), .A(n16471), .B(n16470), .ZN(
        n16474) );
  AOI22_X1 U17410 ( .A1(n16615), .A2(n16474), .B1(n12684), .B2(n9060), .ZN(
        P3_U3469) );
  INV_X1 U17411 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16473) );
  AOI22_X1 U17412 ( .A1(n16618), .A2(n16474), .B1(n16473), .B2(n9044), .ZN(
        P3_U3420) );
  INV_X1 U17413 ( .A(n16475), .ZN(n16479) );
  OAI21_X1 U17414 ( .B1(n7847), .B2(n16579), .A(n16476), .ZN(n16478) );
  AOI211_X1 U17415 ( .C1(n16514), .C2(n16479), .A(n16478), .B(n16477), .ZN(
        n16482) );
  AOI22_X1 U17416 ( .A1(n16591), .A2(n16482), .B1(n16480), .B2(n16589), .ZN(
        P2_U3509) );
  INV_X1 U17417 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n16481) );
  AOI22_X1 U17418 ( .A1(n16595), .A2(n16482), .B1(n16481), .B2(n16592), .ZN(
        P2_U3460) );
  NOR2_X1 U17419 ( .A1(n16483), .A2(n16609), .ZN(n16485) );
  AOI211_X1 U17420 ( .C1(n16614), .C2(n16486), .A(n16485), .B(n16484), .ZN(
        n16489) );
  INV_X1 U17421 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16487) );
  AOI22_X1 U17422 ( .A1(n16615), .A2(n16489), .B1(n16487), .B2(n9060), .ZN(
        P3_U3470) );
  INV_X1 U17423 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16488) );
  AOI22_X1 U17424 ( .A1(n16618), .A2(n16489), .B1(n16488), .B2(n9044), .ZN(
        P3_U3423) );
  AOI22_X1 U17425 ( .A1(n16398), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n16491), 
        .B2(n16490), .ZN(n16492) );
  OAI21_X1 U17426 ( .B1(n16494), .B2(n16493), .A(n16492), .ZN(n16497) );
  NOR2_X1 U17427 ( .A1(n16495), .A2(n16646), .ZN(n16496) );
  AOI211_X1 U17428 ( .C1(n16499), .C2(n16498), .A(n16497), .B(n16496), .ZN(
        n16500) );
  OAI21_X1 U17429 ( .B1(n16398), .B2(n16501), .A(n16500), .ZN(P1_U3282) );
  NOR2_X1 U17430 ( .A1(n16502), .A2(n16609), .ZN(n16504) );
  AOI211_X1 U17431 ( .C1(n16521), .C2(n16505), .A(n16504), .B(n16503), .ZN(
        n16507) );
  AOI22_X1 U17432 ( .A1(n16615), .A2(n16507), .B1(n13737), .B2(n9060), .ZN(
        P3_U3471) );
  INV_X1 U17433 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16506) );
  AOI22_X1 U17434 ( .A1(n16618), .A2(n16507), .B1(n16506), .B2(n9044), .ZN(
        P3_U3426) );
  INV_X1 U17435 ( .A(n16508), .ZN(n16513) );
  OAI21_X1 U17436 ( .B1(n16510), .B2(n16579), .A(n16509), .ZN(n16512) );
  AOI211_X1 U17437 ( .C1(n16514), .C2(n16513), .A(n16512), .B(n16511), .ZN(
        n16516) );
  AOI22_X1 U17438 ( .A1(n16591), .A2(n16516), .B1(n16515), .B2(n16589), .ZN(
        P2_U3511) );
  AOI22_X1 U17439 ( .A1(n16595), .A2(n16516), .B1(n10126), .B2(n16592), .ZN(
        P2_U3466) );
  NOR2_X1 U17440 ( .A1(n16517), .A2(n16609), .ZN(n16519) );
  AOI211_X1 U17441 ( .C1(n16521), .C2(n16520), .A(n16519), .B(n16518), .ZN(
        n16524) );
  INV_X1 U17442 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n16522) );
  AOI22_X1 U17443 ( .A1(n16615), .A2(n16524), .B1(n16522), .B2(n9060), .ZN(
        P3_U3472) );
  INV_X1 U17444 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16523) );
  AOI22_X1 U17445 ( .A1(n16618), .A2(n16524), .B1(n16523), .B2(n9044), .ZN(
        P3_U3429) );
  OAI211_X1 U17446 ( .C1(n16527), .C2(n16624), .A(n16526), .B(n16525), .ZN(
        n16530) );
  AND2_X1 U17447 ( .A1(n16528), .A2(n16568), .ZN(n16529) );
  AOI211_X1 U17448 ( .C1(n16631), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16533) );
  AOI22_X1 U17449 ( .A1(n16635), .A2(n16533), .B1(n11561), .B2(n16633), .ZN(
        P1_U3541) );
  INV_X1 U17450 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n16532) );
  AOI22_X1 U17451 ( .A1(n16638), .A2(n16533), .B1(n16532), .B2(n16636), .ZN(
        P1_U3498) );
  NOR2_X1 U17452 ( .A1(n16534), .A2(n16609), .ZN(n16536) );
  AOI211_X1 U17453 ( .C1(n16614), .C2(n16537), .A(n16536), .B(n16535), .ZN(
        n16540) );
  AOI22_X1 U17454 ( .A1(n16615), .A2(n16540), .B1(n16538), .B2(n9060), .ZN(
        P3_U3473) );
  INV_X1 U17455 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n16539) );
  AOI22_X1 U17456 ( .A1(n16618), .A2(n16540), .B1(n16539), .B2(n9044), .ZN(
        P3_U3432) );
  OAI22_X1 U17457 ( .A1(n16544), .A2(n16543), .B1(n16542), .B2(n16541), .ZN(
        n16553) );
  AOI21_X1 U17458 ( .B1(n16547), .B2(n16546), .A(n16545), .ZN(n16548) );
  INV_X1 U17459 ( .A(n16548), .ZN(n16551) );
  AOI21_X1 U17460 ( .B1(n16551), .B2(n16550), .A(n16549), .ZN(n16552) );
  AOI211_X1 U17461 ( .C1(n16561), .C2(n16554), .A(n16553), .B(n16552), .ZN(
        n16556) );
  OAI211_X1 U17462 ( .C1(n16558), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        P1_U3215) );
  AOI21_X1 U17463 ( .B1(n16561), .B2(n16560), .A(n16559), .ZN(n16564) );
  NAND3_X1 U17464 ( .A1(n16562), .A2(n16631), .A3(n12965), .ZN(n16563) );
  OAI211_X1 U17465 ( .C1(n16566), .C2(n16565), .A(n16564), .B(n16563), .ZN(
        n16567) );
  AOI21_X1 U17466 ( .B1(n16569), .B2(n16568), .A(n16567), .ZN(n16571) );
  AOI22_X1 U17467 ( .A1(n16635), .A2(n16571), .B1(n16570), .B2(n16633), .ZN(
        P1_U3542) );
  AOI22_X1 U17468 ( .A1(n16638), .A2(n16571), .B1(n9460), .B2(n16636), .ZN(
        P1_U3501) );
  OR2_X1 U17469 ( .A1(n16572), .A2(n16581), .ZN(n16573) );
  AND2_X1 U17470 ( .A1(n16574), .A2(n16573), .ZN(n16605) );
  NAND2_X1 U17471 ( .A1(n16600), .A2(n16575), .ZN(n16576) );
  NAND2_X1 U17472 ( .A1(n16576), .A2(n12771), .ZN(n16577) );
  OR2_X1 U17473 ( .A1(n16578), .A2(n16577), .ZN(n16602) );
  OAI21_X1 U17474 ( .B1(n7846), .B2(n16579), .A(n16602), .ZN(n16587) );
  XOR2_X1 U17475 ( .A(n16580), .B(n16581), .Z(n16585) );
  INV_X1 U17476 ( .A(n16582), .ZN(n16583) );
  AOI21_X1 U17477 ( .B1(n16585), .B2(n16584), .A(n16583), .ZN(n16608) );
  INV_X1 U17478 ( .A(n16608), .ZN(n16586) );
  AOI211_X1 U17479 ( .C1(n16605), .C2(n16588), .A(n16587), .B(n16586), .ZN(
        n16594) );
  AOI22_X1 U17480 ( .A1(n16591), .A2(n16594), .B1(n16590), .B2(n16589), .ZN(
        P2_U3513) );
  INV_X1 U17481 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U17482 ( .A1(n16595), .A2(n16594), .B1(n16593), .B2(n16592), .ZN(
        P2_U3472) );
  AOI222_X1 U17483 ( .A1(n16600), .A2(n16599), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n16598), .C1(n16597), .C2(n16596), .ZN(n16607) );
  NOR2_X1 U17484 ( .A1(n16602), .A2(n16601), .ZN(n16603) );
  AOI21_X1 U17485 ( .B1(n16605), .B2(n16604), .A(n16603), .ZN(n16606) );
  OAI211_X1 U17486 ( .C1(n16598), .C2(n16608), .A(n16607), .B(n16606), .ZN(
        P2_U3251) );
  NOR2_X1 U17487 ( .A1(n16610), .A2(n16609), .ZN(n16612) );
  AOI211_X1 U17488 ( .C1(n16614), .C2(n16613), .A(n16612), .B(n16611), .ZN(
        n16617) );
  AOI22_X1 U17489 ( .A1(n16615), .A2(n16617), .B1(n13783), .B2(n9060), .ZN(
        P3_U3474) );
  INV_X1 U17490 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U17491 ( .A1(n16618), .A2(n16617), .B1(n16616), .B2(n9044), .ZN(
        P3_U3435) );
  OAI21_X1 U17492 ( .B1(n16620), .B2(n16625), .A(n16619), .ZN(n16648) );
  INV_X1 U17493 ( .A(n16648), .ZN(n16632) );
  OAI211_X1 U17494 ( .C1(n16641), .C2(n16623), .A(n16622), .B(n16621), .ZN(
        n16643) );
  OAI211_X1 U17495 ( .C1(n16641), .C2(n16624), .A(n16643), .B(n16639), .ZN(
        n16630) );
  INV_X1 U17496 ( .A(n16625), .ZN(n16626) );
  XNOR2_X1 U17497 ( .A(n16627), .B(n16626), .ZN(n16645) );
  NOR2_X1 U17498 ( .A1(n16645), .A2(n16628), .ZN(n16629) );
  AOI211_X1 U17499 ( .C1(n16632), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        n16637) );
  INV_X1 U17500 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n16634) );
  AOI22_X1 U17501 ( .A1(n16635), .A2(n16637), .B1(n16634), .B2(n16633), .ZN(
        P1_U3543) );
  AOI22_X1 U17502 ( .A1(n16638), .A2(n16637), .B1(n9480), .B2(n16636), .ZN(
        P1_U3504) );
  OAI211_X1 U17503 ( .C1(n16641), .C2(n16640), .A(n16639), .B(n7416), .ZN(
        n16642) );
  OAI21_X1 U17504 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n7416), .A(n16642), .ZN(
        n16651) );
  OAI222_X1 U17505 ( .A1(n16648), .A2(n16647), .B1(n16646), .B2(n16645), .C1(
        n16644), .C2(n16643), .ZN(n16649) );
  INV_X1 U17506 ( .A(n16649), .ZN(n16650) );
  OAI211_X1 U17507 ( .C1(n16653), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        P1_U3278) );
  AOI21_X1 U17508 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16654) );
  OAI21_X1 U17509 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16654), 
        .ZN(U28) );
  CLKBUF_X2 U7520 ( .A(n11144), .Z(n7443) );
  CLKBUF_X1 U7538 ( .A(n7437), .Z(n8958) );
  CLKBUF_X1 U9158 ( .A(n7433), .Z(n9689) );
endmodule

