

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9690, n9691, n9692, n9693, n9696, n9697, n9698, n9699, n9701, n9703,
         n9704, n9705, n9706, n9707, n9709, n9710, n9711, n9712, n9713, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9766,
         n9767, n9768, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020;

  NOR2_X1 U11134 ( .A1(n15190), .A2(n20823), .ZN(n15443) );
  NAND2_X2 U11135 ( .A1(n10872), .A2(n10116), .ZN(n15190) );
  INV_X1 U11136 ( .A(n19991), .ZN(n20013) );
  INV_X1 U11137 ( .A(n15212), .ZN(n10872) );
  NOR2_X1 U11138 ( .A1(n16603), .A2(n16604), .ZN(n16602) );
  XNOR2_X1 U11139 ( .A(n14438), .B(n10121), .ZN(n15015) );
  NAND2_X1 U11140 ( .A1(n15022), .A2(n14424), .ZN(n14438) );
  AOI211_X1 U11141 ( .C1(n13207), .C2(n13464), .A(n13463), .B(n13462), .ZN(
        n15640) );
  NOR2_X1 U11142 ( .A1(n16624), .A2(n17537), .ZN(n16623) );
  NAND2_X1 U11143 ( .A1(n10564), .A2(n9782), .ZN(n15314) );
  INV_X2 U11144 ( .A(n9749), .ZN(n16056) );
  BUF_X1 U11145 ( .A(n11299), .Z(n9749) );
  NAND2_X1 U11146 ( .A1(n13942), .A2(n19016), .ZN(n13869) );
  INV_X2 U11147 ( .A(n10032), .ZN(n10012) );
  NOR2_X1 U11148 ( .A1(n10316), .A2(n10317), .ZN(n10492) );
  NOR2_X1 U11149 ( .A1(n10319), .A2(n10315), .ZN(n10483) );
  AND2_X2 U11151 ( .A1(n10333), .A2(n10334), .ZN(n10354) );
  CLKBUF_X2 U11152 ( .A(n12484), .Z(n17160) );
  INV_X1 U11153 ( .A(n12410), .ZN(n17140) );
  NAND3_X1 U11154 ( .A1(n10265), .A2(n10264), .A3(n10263), .ZN(n10299) );
  CLKBUF_X2 U11155 ( .A(n11087), .Z(n11052) );
  AND2_X1 U11156 ( .A1(n10328), .A2(n10334), .ZN(n10379) );
  AND2_X1 U11157 ( .A1(n10327), .A2(n10334), .ZN(n12265) );
  AND2_X1 U11158 ( .A1(n14400), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10405) );
  AND2_X1 U11159 ( .A1(n9698), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10454) );
  INV_X1 U11160 ( .A(n9793), .ZN(n17184) );
  INV_X1 U11161 ( .A(n16878), .ZN(n15740) );
  AND2_X1 U11162 ( .A1(n9743), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10254) );
  AND2_X1 U11164 ( .A1(n13429), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10333) );
  NAND2_X1 U11166 ( .A1(n18821), .A2(n12634), .ZN(n16910) );
  CLKBUF_X2 U11167 ( .A(n9974), .Z(n9761) );
  CLKBUF_X2 U11168 ( .A(n11132), .Z(n11180) );
  CLKBUF_X2 U11169 ( .A(n11081), .Z(n11044) );
  CLKBUF_X2 U11170 ( .A(n11086), .Z(n12082) );
  AND4_X1 U11171 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10913) );
  AND2_X1 U11172 ( .A1(n10887), .A2(n13502), .ZN(n11081) );
  AND2_X2 U11173 ( .A1(n11112), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10886) );
  AOI22_X2 U11174 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13700), .B1(DATAI_28_), 
        .B2(n13699), .ZN(n20466) );
  NOR2_X4 U11175 ( .A1(n20076), .A2(n13564), .ZN(n13700) );
  NOR2_X4 U11176 ( .A1(n13565), .A2(n20076), .ZN(n13699) );
  AND2_X1 U11178 ( .A1(n10889), .A2(n13502), .ZN(n11087) );
  AOI22_X1 U11179 ( .A1(n20908), .A2(keyinput66), .B1(n20907), .B2(keyinput56), 
        .ZN(n20906) );
  INV_X2 U11180 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10129) );
  INV_X2 U11182 ( .A(n14514), .ZN(n11548) );
  AND2_X1 U11183 ( .A1(n14389), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10360) );
  AND2_X1 U11184 ( .A1(n9693), .A2(n10334), .ZN(n10359) );
  AND2_X2 U11185 ( .A1(n13429), .A2(n10129), .ZN(n14467) );
  NOR2_X1 U11186 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15766), .ZN(
        n12572) );
  NAND2_X1 U11187 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12634), .ZN(
        n12419) );
  AND2_X2 U11188 ( .A1(n10888), .A2(n10889), .ZN(n10970) );
  INV_X1 U11189 ( .A(n20677), .ZN(n11502) );
  NOR2_X1 U11190 ( .A1(n11588), .A2(n10014), .ZN(n10835) );
  INV_X2 U11191 ( .A(n10286), .ZN(n10813) );
  NOR2_X1 U11192 ( .A1(n17545), .A2(n17546), .ZN(n17525) );
  OR2_X1 U11193 ( .A1(n17356), .A2(n12520), .ZN(n12523) );
  CLKBUF_X2 U11194 ( .A(n12463), .Z(n9697) );
  NAND2_X1 U11195 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12415) );
  NAND2_X1 U11196 ( .A1(n11145), .A2(n11022), .ZN(n11400) );
  NAND2_X1 U11197 ( .A1(n11016), .A2(n11008), .ZN(n11010) );
  NOR2_X1 U11199 ( .A1(n16169), .A2(n16168), .ZN(n20101) );
  AOI21_X1 U11201 ( .B1(n10001), .B2(n9774), .A(n14456), .ZN(n14459) );
  NOR2_X1 U11202 ( .A1(n13869), .A2(n9836), .ZN(n15041) );
  OR2_X1 U11203 ( .A1(n9862), .A2(n9860), .ZN(n9859) );
  NAND2_X1 U11204 ( .A1(n13107), .A2(n13106), .ZN(n13772) );
  NAND2_X2 U11205 ( .A1(n10193), .A2(n10192), .ZN(n10243) );
  NAND2_X1 U11206 ( .A1(n12143), .A2(n12142), .ZN(n13773) );
  NOR2_X1 U11207 ( .A1(n16582), .A2(n16583), .ZN(n16581) );
  NOR2_X1 U11208 ( .A1(n16647), .A2(n17568), .ZN(n16646) );
  INV_X1 U11210 ( .A(n18227), .ZN(n17235) );
  NOR2_X1 U11211 ( .A1(n17612), .A2(n17611), .ZN(n17589) );
  AOI221_X1 U11212 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17624), 
        .C1(n17626), .C2(n17635), .A(n17563), .ZN(n17616) );
  NOR2_X1 U11213 ( .A1(n17780), .A2(n18103), .ZN(n17779) );
  AND2_X1 U11214 ( .A1(n14995), .A2(n14996), .ZN(n15054) );
  NAND2_X1 U11215 ( .A1(n15029), .A2(n15028), .ZN(n14420) );
  AND2_X1 U11216 ( .A1(n14132), .A2(n14133), .ZN(n14135) );
  OR2_X1 U11217 ( .A1(n14278), .A2(n14277), .ZN(n15137) );
  AND2_X1 U11218 ( .A1(n14240), .A2(n14244), .ZN(n15626) );
  NOR2_X1 U11219 ( .A1(n12631), .A2(n12630), .ZN(n18203) );
  NAND2_X1 U11220 ( .A1(n16416), .A2(n16417), .ZN(n17770) );
  AOI221_X1 U11221 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n15888), .C1(n15887), 
        .C2(n15888), .A(n15886), .ZN(n15889) );
  INV_X1 U11222 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19668) );
  AOI211_X1 U11223 ( .C1(n16577), .C2(n16905), .A(n16576), .B(n16575), .ZN(
        n16580) );
  INV_X1 U11224 ( .A(n17844), .ZN(n17867) );
  AND2_X1 U11225 ( .A1(n14190), .A2(n15955), .ZN(n14566) );
  XNOR2_X2 U11226 ( .A(n11160), .B(n11161), .ZN(n13281) );
  NOR2_X4 U11227 ( .A1(n14080), .A2(n10102), .ZN(n14182) );
  NAND2_X2 U11228 ( .A1(n16384), .A2(n18022), .ZN(n17694) );
  NOR2_X2 U11229 ( .A1(n17652), .A2(n17651), .ZN(n16700) );
  NOR2_X2 U11230 ( .A1(n11025), .A2(n11145), .ZN(n11014) );
  AND2_X4 U11231 ( .A1(n10158), .A2(n10157), .ZN(n15658) );
  NAND2_X1 U11232 ( .A1(n10448), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13799) );
  OR2_X2 U11233 ( .A1(n12634), .A2(n12415), .ZN(n15766) );
  NOR2_X2 U11234 ( .A1(n17739), .A2(n17998), .ZN(n17697) );
  AND2_X1 U11235 ( .A1(n13530), .A2(n13513), .ZN(n9690) );
  AND2_X1 U11236 ( .A1(n13530), .A2(n13513), .ZN(n9691) );
  AND2_X1 U11237 ( .A1(n13530), .A2(n13513), .ZN(n11086) );
  OAI222_X1 U11238 ( .A1(n14635), .A2(n15885), .B1(n20023), .B2(n14600), .C1(
        n15884), .C2(n14629), .ZN(P1_U2846) );
  BUF_X1 U11239 ( .A(n15851), .Z(n9692) );
  AND2_X2 U11240 ( .A1(n15445), .A2(n9731), .ZN(n9940) );
  NAND2_X2 U11241 ( .A1(n13255), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11160) );
  NOR2_X2 U11242 ( .A1(n12756), .A2(n16342), .ZN(n12757) );
  XNOR2_X2 U11243 ( .A(n11164), .B(n20107), .ZN(n13422) );
  AND2_X2 U11244 ( .A1(n13440), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9693) );
  NAND2_X2 U11245 ( .A1(n13282), .A2(n11163), .ZN(n11164) );
  INV_X2 U11246 ( .A(n21020), .ZN(n9696) );
  NOR2_X2 U11248 ( .A1(n17649), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17648) );
  NOR2_X1 U11249 ( .A1(n12420), .A2(n12419), .ZN(n12463) );
  AND2_X2 U11250 ( .A1(n13429), .A2(n10129), .ZN(n9698) );
  NAND2_X2 U11251 ( .A1(n11072), .A2(n11071), .ZN(n11150) );
  CLKBUF_X1 U11252 ( .A(n14769), .Z(n15845) );
  AOI21_X1 U11253 ( .B1(n15294), .B2(n10084), .A(n10639), .ZN(n10085) );
  OR3_X1 U11254 ( .A1(n14949), .A2(n9967), .A3(n12907), .ZN(n9966) );
  XNOR2_X1 U11255 ( .A(n14378), .B(n14379), .ZN(n15035) );
  XNOR2_X1 U11256 ( .A(n10562), .B(n14033), .ZN(n14038) );
  NAND2_X1 U11257 ( .A1(n11277), .A2(n11289), .ZN(n11299) );
  AND2_X1 U11258 ( .A1(n10560), .A2(n10861), .ZN(n10071) );
  XNOR2_X1 U11259 ( .A(n10526), .B(n10530), .ZN(n10851) );
  INV_X1 U11260 ( .A(n13797), .ZN(n9716) );
  NOR2_X2 U11261 ( .A1(n9794), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10667) );
  INV_X2 U11262 ( .A(n17687), .ZN(n17722) );
  NAND2_X1 U11263 ( .A1(n17773), .A2(n17871), .ZN(n17798) );
  BUF_X1 U11264 ( .A(n10490), .Z(n19302) );
  INV_X2 U11265 ( .A(n19451), .ZN(n9699) );
  NOR2_X1 U11266 ( .A1(n9742), .A2(n16550), .ZN(n16677) );
  NAND2_X1 U11267 ( .A1(n12377), .A2(n12164), .ZN(n15629) );
  OR2_X1 U11268 ( .A1(n9953), .A2(n9951), .ZN(n10574) );
  NOR2_X1 U11269 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  NAND4_X2 U11270 ( .A1(n10266), .A2(n9795), .A3(n12145), .A4(n10247), .ZN(
        n10248) );
  CLKBUF_X2 U11271 ( .A(n10273), .Z(n10785) );
  NAND4_X1 U11272 ( .A1(n12707), .A2(n18218), .A3(n12656), .A4(n12662), .ZN(
        n18650) );
  CLKBUF_X1 U11273 ( .A(n11006), .Z(n12385) );
  OR2_X1 U11274 ( .A1(n12558), .A2(n12559), .ZN(n18835) );
  CLKBUF_X2 U11275 ( .A(n11050), .Z(n12081) );
  AND4_X1 U11276 ( .A1(n10954), .A2(n10953), .A3(n10952), .A4(n10951), .ZN(
        n9723) );
  AND4_X1 U11277 ( .A1(n10893), .A2(n10892), .A3(n10891), .A4(n10890), .ZN(
        n10894) );
  CLKBUF_X2 U11278 ( .A(n12549), .Z(n15745) );
  CLKBUF_X2 U11279 ( .A(n11079), .Z(n11051) );
  CLKBUF_X2 U11280 ( .A(n10970), .Z(n12080) );
  BUF_X2 U11281 ( .A(n11887), .Z(n12087) );
  CLKBUF_X2 U11282 ( .A(n11131), .Z(n12079) );
  BUF_X2 U11283 ( .A(n12059), .Z(n11928) );
  CLKBUF_X2 U11284 ( .A(n10152), .Z(n9763) );
  BUF_X2 U11285 ( .A(n11133), .Z(n9703) );
  OR2_X1 U11287 ( .A1(n12416), .A2(n16910), .ZN(n9791) );
  CLKBUF_X1 U11288 ( .A(n10147), .Z(n9757) );
  AND2_X2 U11289 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13429) );
  AND2_X1 U11290 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12761) );
  NOR2_X4 U11291 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13432) );
  OR2_X1 U11292 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U11293 ( .A1(n10040), .A2(n14708), .ZN(n11605) );
  AND2_X1 U11294 ( .A1(n14280), .A2(n14279), .ZN(n14287) );
  AND2_X1 U11295 ( .A1(n14589), .A2(n14545), .ZN(n16010) );
  NAND2_X1 U11296 ( .A1(n10039), .A2(n9926), .ZN(n10041) );
  NAND2_X1 U11297 ( .A1(n11580), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9926) );
  NOR2_X1 U11298 ( .A1(n15054), .A2(n14487), .ZN(n14503) );
  OAI21_X1 U11299 ( .B1(n12194), .B2(n9784), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U11300 ( .A1(n12200), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12382) );
  OR2_X1 U11301 ( .A1(n15392), .A2(n19179), .ZN(n11598) );
  OR2_X1 U11302 ( .A1(n14768), .A2(n10046), .ZN(n11309) );
  NAND2_X1 U11303 ( .A1(n9892), .A2(n15568), .ZN(n9878) );
  NAND2_X1 U11304 ( .A1(n9927), .A2(n11305), .ZN(n14768) );
  OR2_X1 U11305 ( .A1(n15312), .A2(n9877), .ZN(n9780) );
  AOI211_X1 U11306 ( .C1(n16343), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        n14285) );
  OAI21_X1 U11307 ( .B1(n15294), .B2(n10083), .A(n10080), .ZN(n10086) );
  AOI21_X1 U11308 ( .B1(n10867), .B2(n15618), .A(n9886), .ZN(n9885) );
  OR2_X1 U11309 ( .A1(n14950), .A2(n12792), .ZN(n15374) );
  NAND2_X1 U11310 ( .A1(n14423), .A2(n14422), .ZN(n14424) );
  CLKBUF_X1 U11311 ( .A(n15338), .Z(n9717) );
  OAI21_X1 U11312 ( .B1(n12792), .B2(n12793), .A(n12908), .ZN(n15001) );
  OR2_X1 U11313 ( .A1(n14949), .A2(n9967), .ZN(n12908) );
  CLKBUF_X1 U11314 ( .A(n15303), .Z(n9732) );
  NAND2_X1 U11315 ( .A1(n11591), .A2(n10804), .ZN(n14949) );
  NAND2_X1 U11316 ( .A1(n14021), .A2(n10859), .ZN(n10866) );
  AOI211_X1 U11317 ( .C1(n14271), .C2(n20703), .A(n14270), .B(n14269), .ZN(
        n14272) );
  OR2_X1 U11318 ( .A1(n12911), .A2(n12818), .ZN(n15059) );
  NOR2_X1 U11319 ( .A1(n15016), .A2(n15018), .ZN(n11591) );
  AND2_X1 U11320 ( .A1(n10043), .A2(n11273), .ZN(n10042) );
  AND3_X1 U11321 ( .A1(n14779), .A2(n16053), .A3(n9930), .ZN(n9739) );
  AND2_X1 U11322 ( .A1(n16426), .A2(n10052), .ZN(n15775) );
  AND2_X1 U11323 ( .A1(n10681), .A2(n15165), .ZN(n11596) );
  NAND2_X1 U11324 ( .A1(n15041), .A2(n14349), .ZN(n14378) );
  NAND2_X1 U11325 ( .A1(n20057), .A2(n11223), .ZN(n13765) );
  OR2_X1 U11326 ( .A1(n15353), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10117) );
  AND2_X1 U11327 ( .A1(n11299), .A2(n11292), .ZN(n14114) );
  XNOR2_X1 U11328 ( .A(n9750), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16053) );
  XNOR2_X1 U11329 ( .A(n10868), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16338) );
  OAI22_X1 U11330 ( .A1(n13883), .A2(n13884), .B1(n14006), .B2(n13688), .ZN(
        n14000) );
  NOR2_X1 U11331 ( .A1(n15050), .A2(n15051), .ZN(n15049) );
  AND2_X1 U11332 ( .A1(n11270), .A2(n11269), .ZN(n16095) );
  NAND2_X1 U11333 ( .A1(n10561), .A2(n18971), .ZN(n10562) );
  NAND2_X1 U11334 ( .A1(n9810), .A2(n11659), .ZN(n13729) );
  NAND2_X1 U11335 ( .A1(n10860), .A2(n10687), .ZN(n10868) );
  NAND2_X1 U11336 ( .A1(n10862), .A2(n10071), .ZN(n10561) );
  NAND2_X1 U11337 ( .A1(n9963), .A2(n9962), .ZN(n15050) );
  XNOR2_X1 U11338 ( .A(n11277), .B(n11276), .ZN(n11674) );
  NAND2_X1 U11339 ( .A1(n11666), .A2(n11665), .ZN(n13845) );
  NAND2_X1 U11340 ( .A1(n10558), .A2(n10557), .ZN(n10862) );
  OR2_X1 U11341 ( .A1(n10851), .A2(n9891), .ZN(n13995) );
  AND2_X1 U11342 ( .A1(n10851), .A2(n9891), .ZN(n13996) );
  OR2_X1 U11343 ( .A1(n13823), .A2(n13939), .ZN(n14137) );
  AND2_X1 U11344 ( .A1(n10854), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9889) );
  AOI21_X1 U11345 ( .B1(n16201), .B2(n11563), .A(n14856), .ZN(n11577) );
  NAND2_X1 U11346 ( .A1(n10532), .A2(n10531), .ZN(n10559) );
  OR2_X1 U11347 ( .A1(n9792), .A2(n14616), .ZN(n14618) );
  NOR2_X1 U11348 ( .A1(n17604), .A2(n12729), .ZN(n17562) );
  INV_X1 U11349 ( .A(n10531), .ZN(n10526) );
  AND3_X1 U11350 ( .A1(n10478), .A2(n10477), .A3(n12248), .ZN(n10531) );
  CLKBUF_X1 U11351 ( .A(n11609), .Z(n20115) );
  OR2_X1 U11352 ( .A1(n10543), .A2(n10542), .ZN(n10556) );
  OR2_X1 U11353 ( .A1(n14194), .A2(n14195), .ZN(n15959) );
  NAND2_X1 U11354 ( .A1(n11617), .A2(n11616), .ZN(n14902) );
  AND2_X1 U11355 ( .A1(n10024), .A2(n10022), .ZN(n16258) );
  AND2_X1 U11356 ( .A1(n13217), .A2(n13243), .ZN(n13222) );
  AND2_X1 U11357 ( .A1(n13296), .A2(n10744), .ZN(n13656) );
  OR2_X1 U11358 ( .A1(n16270), .A2(n10032), .ZN(n10024) );
  NOR2_X1 U11360 ( .A1(n14641), .A2(n11462), .ZN(n14186) );
  AND2_X1 U11361 ( .A1(n13190), .A2(n13220), .ZN(n13219) );
  NOR2_X2 U11362 ( .A1(n18835), .A2(n16522), .ZN(n17839) );
  NOR2_X1 U11363 ( .A1(n16667), .A2(n17601), .ZN(n16666) );
  NAND2_X1 U11364 ( .A1(n10611), .A2(n10669), .ZN(n10615) );
  NAND2_X1 U11365 ( .A1(n14209), .A2(n9822), .ZN(n14641) );
  AOI21_X1 U11366 ( .B1(n16168), .B2(n13284), .A(n14895), .ZN(n20100) );
  INV_X2 U11367 ( .A(n19513), .ZN(n9701) );
  NAND2_X1 U11368 ( .A1(n11189), .A2(n11188), .ZN(n13587) );
  AND2_X1 U11369 ( .A1(n13621), .A2(n9826), .ZN(n15587) );
  AND2_X1 U11370 ( .A1(n10030), .A2(n10029), .ZN(n15785) );
  AND2_X1 U11371 ( .A1(n14109), .A2(n11445), .ZN(n14209) );
  NAND2_X2 U11372 ( .A1(n14695), .A2(n13546), .ZN(n16009) );
  NAND2_X1 U11373 ( .A1(n20125), .A2(n16236), .ZN(n11189) );
  OAI21_X1 U11374 ( .B1(n11622), .B2(n11239), .A(n11154), .ZN(n13255) );
  XNOR2_X1 U11375 ( .A(n11169), .B(n13604), .ZN(n20125) );
  NOR2_X1 U11376 ( .A1(n14108), .A2(n14107), .ZN(n14109) );
  OR2_X1 U11377 ( .A1(n14983), .A2(n10032), .ZN(n10030) );
  AND2_X1 U11378 ( .A1(n11393), .A2(n13171), .ZN(n11521) );
  OAI21_X1 U11379 ( .B1(n13948), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11108), 
        .ZN(n11614) );
  AOI21_X1 U11380 ( .B1(n13195), .B2(n13194), .A(n13193), .ZN(n13218) );
  NAND2_X1 U11381 ( .A1(n9899), .A2(n9898), .ZN(n14108) );
  INV_X1 U11382 ( .A(n13180), .ZN(n13197) );
  XNOR2_X1 U11383 ( .A(n13772), .B(n13191), .ZN(n13194) );
  INV_X1 U11384 ( .A(n13895), .ZN(n9899) );
  NAND2_X1 U11385 ( .A1(n10295), .A2(n10294), .ZN(n10285) );
  NAND2_X1 U11386 ( .A1(n10302), .A2(n19008), .ZN(n10315) );
  NAND2_X1 U11387 ( .A1(n11106), .A2(n11105), .ZN(n13562) );
  NAND2_X2 U11388 ( .A1(n18076), .A2(n18082), .ZN(n18100) );
  NOR2_X1 U11389 ( .A1(n9985), .A2(n12252), .ZN(n9984) );
  NAND2_X1 U11390 ( .A1(n10298), .A2(n10272), .ZN(n10295) );
  NAND2_X1 U11391 ( .A1(n16220), .A2(n13783), .ZN(n13895) );
  INV_X2 U11392 ( .A(n19048), .ZN(n19052) );
  INV_X1 U11393 ( .A(n13311), .ZN(n9986) );
  NAND2_X1 U11394 ( .A1(n9983), .A2(n13648), .ZN(n9985) );
  NAND2_X2 U11395 ( .A1(n11367), .A2(n11366), .ZN(n13537) );
  NAND2_X1 U11396 ( .A1(n11174), .A2(n11173), .ZN(n13604) );
  NOR2_X1 U11397 ( .A1(n19977), .A2(n13731), .ZN(n16218) );
  OR2_X1 U11398 ( .A1(n13027), .A2(n19793), .ZN(n12147) );
  CLKBUF_X1 U11399 ( .A(n15335), .Z(n16346) );
  NAND2_X1 U11400 ( .A1(n11034), .A2(n11033), .ZN(n11103) );
  INV_X1 U11401 ( .A(n12242), .ZN(n9983) );
  OR2_X1 U11402 ( .A1(n10281), .A2(n10282), .ZN(n10284) );
  OAI21_X1 U11403 ( .B1(n9754), .B2(n10256), .A(n10255), .ZN(n10257) );
  NAND2_X1 U11404 ( .A1(n19869), .A2(n19621), .ZN(n15652) );
  INV_X1 U11405 ( .A(n13894), .ZN(n9898) );
  NOR2_X1 U11406 ( .A1(n10443), .A2(n9937), .ZN(n10439) );
  AND2_X1 U11407 ( .A1(n12718), .A2(n9895), .ZN(n18649) );
  AND4_X1 U11408 ( .A1(n10262), .A2(n10261), .A3(n10267), .A4(n10260), .ZN(
        n10264) );
  AND2_X1 U11409 ( .A1(n13158), .A2(n13159), .ZN(n12232) );
  NOR2_X1 U11410 ( .A1(n12782), .A2(n15168), .ZN(n12784) );
  AND2_X1 U11411 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12518), .ZN(
        n12519) );
  NAND2_X1 U11412 ( .A1(n12222), .A2(n12221), .ZN(n13158) );
  NAND2_X1 U11413 ( .A1(n11076), .A2(n11075), .ZN(n11151) );
  AND3_X1 U11414 ( .A1(n11506), .A2(n13498), .A3(n13908), .ZN(n11029) );
  INV_X1 U11415 ( .A(n10273), .ZN(n10815) );
  NAND3_X1 U11416 ( .A1(n10233), .A2(n13475), .A3(n10234), .ZN(n12145) );
  NOR2_X1 U11417 ( .A1(n18854), .A2(n15764), .ZN(n18661) );
  NAND3_X1 U11418 ( .A1(n16700), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17612) );
  AND2_X1 U11419 ( .A1(n10246), .A2(n10223), .ZN(n10234) );
  AND2_X1 U11420 ( .A1(n17362), .A2(n12515), .ZN(n12517) );
  NAND2_X1 U11421 ( .A1(n10225), .A2(n10224), .ZN(n10717) );
  INV_X1 U11422 ( .A(n9734), .ZN(n13494) );
  OR2_X1 U11423 ( .A1(n10469), .A2(n10468), .ZN(n12248) );
  AND2_X1 U11424 ( .A1(n10944), .A2(n11040), .ZN(n10959) );
  NAND2_X1 U11425 ( .A1(n11007), .A2(n11374), .ZN(n11009) );
  NOR2_X1 U11426 ( .A1(n17367), .A2(n12496), .ZN(n12515) );
  NOR2_X2 U11427 ( .A1(n11175), .A2(n16236), .ZN(n11359) );
  NAND2_X1 U11428 ( .A1(n11175), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11338) );
  OR2_X1 U11429 ( .A1(n11369), .A2(n11027), .ZN(n14257) );
  AND2_X1 U11430 ( .A1(n11371), .A2(n12385), .ZN(n11035) );
  CLKBUF_X1 U11431 ( .A(n13114), .Z(n13904) );
  NAND2_X1 U11432 ( .A1(n13335), .A2(n11328), .ZN(n20677) );
  XNOR2_X1 U11433 ( .A(n12496), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17860) );
  INV_X1 U11434 ( .A(n12512), .ZN(n17367) );
  INV_X2 U11435 ( .A(n18236), .ZN(n17280) );
  INV_X1 U11436 ( .A(n10218), .ZN(n9747) );
  AND2_X1 U11437 ( .A1(n19215), .A2(n19668), .ZN(n12229) );
  INV_X2 U11438 ( .A(U212), .ZN(n16472) );
  INV_X1 U11439 ( .A(n11020), .ZN(n13911) );
  INV_X2 U11440 ( .A(n10218), .ZN(n12214) );
  CLKBUF_X1 U11441 ( .A(n11005), .Z(n9725) );
  NAND2_X2 U11442 ( .A1(n9720), .A2(n9721), .ZN(n11145) );
  NAND2_X2 U11443 ( .A1(n10170), .A2(n10169), .ZN(n19215) );
  MUX2_X1 U11444 ( .A(n10180), .B(n10179), .S(n10334), .Z(n15654) );
  NAND2_X2 U11445 ( .A1(n10955), .A2(n9723), .ZN(n11025) );
  NAND4_X2 U11446 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n11020) );
  NAND2_X1 U11447 ( .A1(n16747), .A2(n12870), .ZN(n17691) );
  OR3_X2 U11448 ( .A1(n12472), .A2(n12471), .A3(n12470), .ZN(n12511) );
  OR2_X1 U11449 ( .A1(n11069), .A2(n11068), .ZN(n11156) );
  NAND2_X2 U11450 ( .A1(n10914), .A2(n10913), .ZN(n11016) );
  AND4_X1 U11451 ( .A1(n10968), .A2(n10967), .A3(n10966), .A4(n10965), .ZN(
        n10981) );
  NAND2_X1 U11452 ( .A1(n10128), .A2(n10894), .ZN(n10945) );
  NAND4_X2 U11453 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(
        n11144) );
  AND4_X1 U11454 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10980) );
  NAND2_X1 U11455 ( .A1(n10124), .A2(n9797), .ZN(n9870) );
  NAND3_X2 U11456 ( .A1(n10904), .A2(n10903), .A3(n10902), .ZN(n11008) );
  NOR2_X1 U11457 ( .A1(n17734), .A2(n17737), .ZN(n16747) );
  AND4_X1 U11458 ( .A1(n10931), .A2(n10930), .A3(n10929), .A4(n10928), .ZN(
        n10942) );
  AND4_X1 U11459 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10940) );
  AND4_X1 U11460 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        n10979) );
  AND4_X1 U11461 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n11004) );
  AND4_X1 U11462 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11001) );
  AND4_X1 U11463 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10215) );
  AND4_X1 U11464 ( .A1(n10964), .A2(n10963), .A3(n10962), .A4(n10961), .ZN(
        n10982) );
  INV_X2 U11465 ( .A(n17093), .ZN(n17161) );
  AND4_X1 U11466 ( .A1(n10923), .A2(n10922), .A3(n10921), .A4(n10920), .ZN(
        n9721) );
  AND4_X1 U11467 ( .A1(n10908), .A2(n10907), .A3(n10906), .A4(n10905), .ZN(
        n10914) );
  AND3_X1 U11468 ( .A1(n10140), .A2(n10334), .A3(n10142), .ZN(n9872) );
  AND3_X1 U11469 ( .A1(n10901), .A2(n10900), .A3(n10899), .ZN(n10902) );
  INV_X1 U11470 ( .A(n18933), .ZN(n18985) );
  AND4_X1 U11471 ( .A1(n10927), .A2(n10926), .A3(n10925), .A4(n10924), .ZN(
        n10943) );
  INV_X2 U11473 ( .A(n16509), .ZN(U215) );
  CLKBUF_X1 U11474 ( .A(n10988), .Z(n11771) );
  NAND2_X2 U11475 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19901), .ZN(n19840) );
  NAND2_X2 U11476 ( .A1(n19901), .A2(n19802), .ZN(n19842) );
  AOI22_X1 U11477 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10920) );
  AND3_X1 U11478 ( .A1(n10131), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10130), .ZN(n10124) );
  NAND2_X2 U11479 ( .A1(n18848), .A2(n18721), .ZN(n18772) );
  NAND2_X2 U11480 ( .A1(n18848), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18776) );
  CLKBUF_X1 U11481 ( .A(n10988), .Z(n9770) );
  CLKBUF_X2 U11482 ( .A(n10969), .Z(n9773) );
  OAI221_X1 U11483 ( .B1(n20908), .B2(keyinput66), .C1(n20907), .C2(keyinput56), .A(n20906), .ZN(n20913) );
  INV_X1 U11484 ( .A(n12428), .ZN(n16878) );
  BUF_X2 U11485 ( .A(n10152), .Z(n9762) );
  INV_X2 U11486 ( .A(n16511), .ZN(n16513) );
  BUF_X2 U11487 ( .A(n10152), .Z(n9764) );
  BUF_X4 U11488 ( .A(n12503), .Z(n9704) );
  CLKBUF_X1 U11489 ( .A(n12635), .Z(n18807) );
  NAND2_X1 U11490 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12635), .ZN(
        n12418) );
  NAND2_X1 U11491 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18821), .ZN(
        n12417) );
  NAND2_X1 U11492 ( .A1(n20947), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12420) );
  NAND2_X2 U11493 ( .A1(n20592), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20689) );
  NOR2_X1 U11494 ( .A1(n17828), .A2(n17830), .ZN(n17809) );
  AND2_X2 U11495 ( .A1(n13429), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9753) );
  AND2_X2 U11496 ( .A1(n13440), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14389) );
  AND2_X1 U11497 ( .A1(n13429), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9752) );
  NAND2_X2 U11498 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18657) );
  INV_X1 U11499 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20947) );
  CLKBUF_X1 U11500 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n14352) );
  AND2_X1 U11501 ( .A1(n10250), .A2(n10251), .ZN(n9743) );
  NAND2_X1 U11502 ( .A1(n9734), .A2(n10251), .ZN(n10273) );
  NAND2_X1 U11504 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17828) );
  NOR2_X1 U11505 ( .A1(n16677), .A2(n17615), .ZN(n16676) );
  OR2_X1 U11506 ( .A1(n10267), .A2(n19890), .ZN(n9705) );
  NAND2_X1 U11507 ( .A1(n9705), .A2(n10726), .ZN(n10268) );
  INV_X1 U11508 ( .A(n10216), .ZN(n9706) );
  AND2_X1 U11509 ( .A1(n11293), .A2(n16090), .ZN(n9707) );
  OAI21_X1 U11512 ( .B1(n13113), .B2(n11377), .A(n11394), .ZN(n11012) );
  NOR2_X2 U11513 ( .A1(n11009), .A2(n13911), .ZN(n13131) );
  NAND2_X1 U11514 ( .A1(n10959), .A2(n10958), .ZN(n11013) );
  NAND2_X2 U11515 ( .A1(n11421), .A2(n11400), .ZN(n11401) );
  NAND2_X1 U11516 ( .A1(n10296), .A2(n10300), .ZN(n9709) );
  INV_X1 U11517 ( .A(n13460), .ZN(n9710) );
  NAND2_X1 U11518 ( .A1(n10296), .A2(n10300), .ZN(n10298) );
  AND2_X1 U11519 ( .A1(n11328), .A2(n11022), .ZN(n13909) );
  NAND2_X1 U11520 ( .A1(n15314), .A2(n10586), .ZN(n9711) );
  CLKBUF_X1 U11521 ( .A(n10296), .Z(n10297) );
  NOR2_X2 U11522 ( .A1(n17940), .A2(n12723), .ZN(n17920) );
  NOR2_X2 U11523 ( .A1(n12416), .A2(n18657), .ZN(n12503) );
  NOR2_X2 U11524 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U11525 ( .A1(n10044), .A2(n10042), .ZN(n16088) );
  NAND2_X1 U11526 ( .A1(n14036), .A2(n14038), .ZN(n9712) );
  NAND2_X1 U11527 ( .A1(n14036), .A2(n14038), .ZN(n10564) );
  CLKBUF_X1 U11528 ( .A(n13880), .Z(n9713) );
  XNOR2_X1 U11529 ( .A(n9862), .B(n9861), .ZN(n13880) );
  INV_X1 U11530 ( .A(n12217), .ZN(n9974) );
  NAND2_X1 U11532 ( .A1(n10304), .A2(n10303), .ZN(n19480) );
  NAND2_X1 U11533 ( .A1(n9713), .A2(n14006), .ZN(n9715) );
  NAND2_X1 U11534 ( .A1(n12913), .A2(n12912), .ZN(n15356) );
  XNOR2_X1 U11536 ( .A(n10866), .B(n10864), .ZN(n15338) );
  NAND2_X1 U11537 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  NAND2_X2 U11538 ( .A1(n14190), .A2(n9718), .ZN(n14567) );
  AND2_X1 U11539 ( .A1(n15955), .A2(n14568), .ZN(n9718) );
  CLKBUF_X1 U11540 ( .A(n13883), .Z(n9719) );
  NAND2_X1 U11541 ( .A1(n10451), .A2(n13800), .ZN(n13883) );
  OR2_X1 U11542 ( .A1(n13449), .A2(n13104), .ZN(n13107) );
  INV_X1 U11543 ( .A(n13449), .ZN(n19008) );
  AND4_X2 U11544 ( .A1(n10919), .A2(n10918), .A3(n10917), .A4(n10916), .ZN(
        n9720) );
  AOI21_X2 U11545 ( .B1(n10970), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n10915), .ZN(n10919) );
  CLKBUF_X1 U11546 ( .A(n14036), .Z(n9722) );
  NAND2_X1 U11547 ( .A1(n12890), .A2(n13114), .ZN(n12384) );
  NAND2_X1 U11548 ( .A1(n15445), .A2(n15446), .ZN(n15175) );
  BUF_X2 U11549 ( .A(n13180), .Z(n13181) );
  AND2_X2 U11550 ( .A1(n10284), .A2(n10283), .ZN(n10294) );
  NOR2_X2 U11551 ( .A1(n13941), .A2(n13943), .ZN(n13942) );
  AOI21_X2 U11552 ( .B1(n15008), .B2(n15003), .A(n15005), .ZN(n14995) );
  NAND2_X2 U11553 ( .A1(n12167), .A2(n10070), .ZN(n15212) );
  INV_X1 U11554 ( .A(n10881), .ZN(n9724) );
  INV_X2 U11556 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10881) );
  INV_X1 U11557 ( .A(n11016), .ZN(n11005) );
  NAND2_X1 U11558 ( .A1(n11032), .A2(n11101), .ZN(n11117) );
  NAND2_X1 U11559 ( .A1(n11212), .A2(n11213), .ZN(n9727) );
  NAND2_X1 U11560 ( .A1(n11212), .A2(n11213), .ZN(n11237) );
  AND2_X1 U11561 ( .A1(n10950), .A2(n10949), .ZN(n9728) );
  AND2_X1 U11563 ( .A1(n10888), .A2(n13513), .ZN(n9748) );
  NAND2_X1 U11564 ( .A1(n10959), .A2(n10958), .ZN(n9729) );
  NOR2_X2 U11566 ( .A1(n14278), .A2(n10873), .ZN(n15123) );
  AND2_X2 U11567 ( .A1(n14182), .A2(n14192), .ZN(n14190) );
  NAND2_X1 U11568 ( .A1(n11024), .A2(n11548), .ZN(n11572) );
  NAND2_X2 U11569 ( .A1(n10050), .A2(n12720), .ZN(n18642) );
  NOR2_X2 U11570 ( .A1(n17768), .A2(n17986), .ZN(n17657) );
  AOI22_X2 U11571 ( .A1(n17839), .A2(n18061), .B1(n17781), .B2(n16384), .ZN(
        n17768) );
  INV_X4 U11572 ( .A(n15727), .ZN(n17176) );
  OR2_X2 U11573 ( .A1(n11653), .A2(n10100), .ZN(n9810) );
  AND4_X1 U11574 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n11002) );
  INV_X1 U11575 ( .A(n15446), .ZN(n9730) );
  NOR2_X1 U11576 ( .A1(n10075), .A2(n9730), .ZN(n9731) );
  INV_X1 U11577 ( .A(n12146), .ZN(n9733) );
  NAND2_X1 U11578 ( .A1(n10086), .A2(n10085), .ZN(n15445) );
  AND2_X1 U11579 ( .A1(n10218), .A2(n19215), .ZN(n13156) );
  AND2_X2 U11580 ( .A1(n10229), .A2(n13156), .ZN(n9734) );
  XOR2_X1 U11581 ( .A(n10222), .B(n10218), .Z(n12153) );
  NAND2_X1 U11582 ( .A1(n9928), .A2(n9738), .ZN(n9735) );
  AND2_X2 U11583 ( .A1(n9735), .A2(n9736), .ZN(n14769) );
  OR2_X1 U11584 ( .A1(n9737), .A2(n11305), .ZN(n9736) );
  INV_X1 U11585 ( .A(n14770), .ZN(n9737) );
  AND2_X1 U11586 ( .A1(n11301), .A2(n14770), .ZN(n9738) );
  NAND2_X1 U11587 ( .A1(n9932), .A2(n9739), .ZN(n9929) );
  CLKBUF_X1 U11588 ( .A(n11394), .Z(n9740) );
  AND2_X1 U11589 ( .A1(n11298), .A2(n14801), .ZN(n14779) );
  AND2_X2 U11590 ( .A1(n13513), .A2(n13502), .ZN(n11079) );
  AOI21_X1 U11591 ( .B1(n10269), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10268), 
        .ZN(n10271) );
  AND2_X1 U11592 ( .A1(n10888), .A2(n10887), .ZN(n9741) );
  AND2_X4 U11594 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U11595 ( .A1(n12165), .A2(n12185), .ZN(n10266) );
  NAND2_X2 U11596 ( .A1(n10285), .A2(n10284), .ZN(n10721) );
  XOR2_X1 U11597 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12872), .Z(n9742) );
  AND2_X1 U11599 ( .A1(n10250), .A2(n10251), .ZN(n9744) );
  AND2_X1 U11600 ( .A1(n10250), .A2(n10251), .ZN(n10751) );
  AOI21_X2 U11601 ( .B1(n12373), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10239), 
        .ZN(n10240) );
  NAND2_X1 U11602 ( .A1(n10238), .A2(n9795), .ZN(n12373) );
  AND2_X1 U11603 ( .A1(n13503), .A2(n10886), .ZN(n9745) );
  AND2_X1 U11604 ( .A1(n13503), .A2(n10886), .ZN(n9746) );
  AND2_X1 U11605 ( .A1(n13503), .A2(n10886), .ZN(n10969) );
  OR2_X2 U11606 ( .A1(n12170), .A2(n10237), .ZN(n9795) );
  NAND2_X2 U11607 ( .A1(n10241), .A2(n10240), .ZN(n10258) );
  AOI21_X1 U11608 ( .B1(n9726), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11118), .ZN(n11123) );
  NAND2_X1 U11609 ( .A1(n13596), .A2(n11199), .ZN(n20059) );
  AND2_X2 U11610 ( .A1(n10216), .A2(n10218), .ZN(n10181) );
  NAND2_X2 U11611 ( .A1(n11169), .A2(n11125), .ZN(n13519) );
  NAND2_X1 U11612 ( .A1(n9978), .A2(n9975), .ZN(n12217) );
  AND2_X4 U11613 ( .A1(n13432), .A2(n13444), .ZN(n10147) );
  INV_X1 U11614 ( .A(n10147), .ZN(n9756) );
  NAND3_X2 U11616 ( .A1(n10227), .A2(n10181), .A3(n9957), .ZN(n12172) );
  NOR2_X2 U11617 ( .A1(n12611), .A2(n12610), .ZN(n18236) );
  NAND2_X2 U11618 ( .A1(n11368), .A2(n13335), .ZN(n12386) );
  NOR2_X2 U11619 ( .A1(n11013), .A2(n10983), .ZN(n11368) );
  AND2_X2 U11620 ( .A1(n10888), .A2(n13513), .ZN(n12059) );
  INV_X1 U11621 ( .A(n10751), .ZN(n10726) );
  AND2_X1 U11622 ( .A1(n10249), .A2(n12185), .ZN(n10250) );
  XNOR2_X2 U11623 ( .A(n10295), .B(n10294), .ZN(n13180) );
  AND2_X2 U11624 ( .A1(n10307), .A2(n10321), .ZN(n10482) );
  OAI21_X2 U11625 ( .B1(n13797), .B2(n10687), .A(n13647), .ZN(n10448) );
  XNOR2_X1 U11626 ( .A(n11198), .B(n11415), .ZN(n13598) );
  AND2_X2 U11627 ( .A1(n13440), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9751) );
  NAND2_X1 U11628 ( .A1(n13420), .A2(n11165), .ZN(n11198) );
  INV_X4 U11629 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13444) );
  NAND2_X2 U11630 ( .A1(n14079), .A2(n14082), .ZN(n14080) );
  NAND2_X1 U11631 ( .A1(n10248), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9754) );
  AND4_X2 U11632 ( .A1(n12123), .A2(n10246), .A3(n10244), .A4(n10073), .ZN(
        n12165) );
  NOR2_X2 U11633 ( .A1(n18800), .A2(n17798), .ZN(n17687) );
  OAI21_X1 U11634 ( .B1(n10301), .B2(n10299), .A(n10300), .ZN(n13449) );
  INV_X1 U11635 ( .A(n9756), .ZN(n9758) );
  INV_X1 U11636 ( .A(n9756), .ZN(n9759) );
  INV_X1 U11637 ( .A(n9756), .ZN(n9760) );
  AND2_X2 U11638 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10326) );
  AND2_X2 U11639 ( .A1(n13892), .A2(n14105), .ZN(n14079) );
  NOR2_X2 U11640 ( .A1(n13778), .A2(n13893), .ZN(n13892) );
  NOR2_X2 U11641 ( .A1(n15654), .A2(n10236), .ZN(n12185) );
  INV_X2 U11642 ( .A(n10228), .ZN(n10236) );
  NOR2_X2 U11643 ( .A1(n13329), .A2(n13735), .ZN(n13728) );
  XNOR2_X1 U11644 ( .A(n10722), .B(n10724), .ZN(n10720) );
  AOI21_X1 U11645 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10290), .ZN(n10722) );
  NAND2_X2 U11646 ( .A1(n9880), .A2(n10395), .ZN(n13797) );
  XNOR2_X2 U11647 ( .A(n9884), .B(n10258), .ZN(n10296) );
  XNOR2_X2 U11648 ( .A(n11103), .B(n11043), .ZN(n11624) );
  NAND2_X2 U11649 ( .A1(n11120), .A2(n11119), .ZN(n11169) );
  NAND2_X2 U11651 ( .A1(n9873), .A2(n9871), .ZN(n10218) );
  AND2_X1 U11652 ( .A1(n10887), .A2(n13502), .ZN(n9766) );
  AND2_X1 U11653 ( .A1(n10889), .A2(n13502), .ZN(n9767) );
  AND2_X1 U11654 ( .A1(n10889), .A2(n13502), .ZN(n9768) );
  AND2_X1 U11655 ( .A1(n13207), .A2(n13197), .ZN(n10304) );
  AND2_X1 U11656 ( .A1(n13207), .A2(n13181), .ZN(n10307) );
  OR2_X2 U11657 ( .A1(n13207), .A2(n13181), .ZN(n10319) );
  NOR2_X4 U11658 ( .A1(n14567), .A2(n15946), .ZN(n15936) );
  AND2_X1 U11659 ( .A1(n10886), .A2(n10887), .ZN(n11923) );
  NOR2_X2 U11660 ( .A1(n11009), .A2(n12900), .ZN(n11376) );
  OAI21_X2 U11661 ( .B1(n11397), .B2(n11012), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11101) );
  AND2_X4 U11662 ( .A1(n10886), .A2(n13513), .ZN(n11132) );
  OAI21_X2 U11663 ( .B1(n14597), .B2(n14594), .A(n14596), .ZN(n15885) );
  AND2_X1 U11664 ( .A1(n10886), .A2(n10887), .ZN(n9771) );
  AND2_X4 U11665 ( .A1(n10886), .A2(n10887), .ZN(n9772) );
  NAND2_X1 U11666 ( .A1(n9876), .A2(n9804), .ZN(n9874) );
  AND2_X1 U11667 ( .A1(n16380), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13208) );
  NAND4_X1 U11668 ( .A1(n10138), .A2(n10136), .A3(n10135), .A4(n10137), .ZN(
        n9869) );
  INV_X1 U11669 ( .A(n14778), .ZN(n9932) );
  AND2_X1 U11670 ( .A1(n11260), .A2(n11259), .ZN(n11263) );
  INV_X1 U11671 ( .A(n15658), .ZN(n10227) );
  NAND2_X1 U11672 ( .A1(n11021), .A2(n11020), .ZN(n11421) );
  NOR2_X1 U11673 ( .A1(n11536), .A2(n9845), .ZN(n10039) );
  NAND2_X1 U11674 ( .A1(n13909), .A2(n11553), .ZN(n11554) );
  AND2_X2 U11675 ( .A1(n11513), .A2(n11145), .ZN(n11374) );
  NOR2_X1 U11676 ( .A1(n9955), .A2(n10513), .ZN(n9954) );
  NAND2_X1 U11677 ( .A1(n10280), .A2(n10279), .ZN(n10282) );
  NAND2_X1 U11678 ( .A1(n10695), .A2(n10658), .ZN(n10659) );
  AND2_X1 U11679 ( .A1(n10667), .A2(n15026), .ZN(n10657) );
  INV_X1 U11680 ( .A(n13996), .ZN(n9881) );
  OR2_X1 U11681 ( .A1(n10553), .A2(n10552), .ZN(n12257) );
  NAND2_X1 U11682 ( .A1(n12216), .A2(n12236), .ZN(n12222) );
  AND2_X1 U11683 ( .A1(n9710), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13454) );
  NOR2_X1 U11684 ( .A1(n16521), .A2(n12713), .ZN(n16537) );
  OR2_X1 U11685 ( .A1(n17792), .A2(n12528), .ZN(n12529) );
  AOI211_X1 U11686 ( .C1(n18203), .C2(n12666), .A(n12665), .B(n12664), .ZN(
        n12718) );
  AND2_X1 U11687 ( .A1(n16218), .A2(n16217), .ZN(n16220) );
  NAND2_X1 U11688 ( .A1(n12911), .A2(n12910), .ZN(n12913) );
  NOR2_X1 U11689 ( .A1(n10671), .A2(n15164), .ZN(n10672) );
  AOI21_X1 U11690 ( .B1(n13793), .B2(n13208), .A(n13142), .ZN(n13195) );
  AND2_X1 U11691 ( .A1(n19445), .A2(n19444), .ZN(n19414) );
  NAND2_X1 U11692 ( .A1(n10186), .A2(n10334), .ZN(n10193) );
  NOR2_X1 U11693 ( .A1(n19445), .A2(n19444), .ZN(n19661) );
  INV_X1 U11694 ( .A(n17441), .ZN(n16538) );
  INV_X1 U11695 ( .A(n15835), .ZN(n12544) );
  AND2_X1 U11696 ( .A1(n13916), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13917) );
  OR2_X1 U11697 ( .A1(n15361), .A2(n20705), .ZN(n12919) );
  OR2_X1 U11698 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20114), .ZN(
        n11354) );
  AND3_X1 U11699 ( .A1(n11005), .A2(n11006), .A3(n13544), .ZN(n11007) );
  NOR2_X1 U11700 ( .A1(n12828), .A2(n16380), .ZN(n10251) );
  INV_X1 U11701 ( .A(n10201), .ZN(n9976) );
  INV_X1 U11702 ( .A(n10197), .ZN(n9979) );
  NAND2_X1 U11703 ( .A1(n12517), .A2(n12687), .ZN(n12520) );
  AND2_X1 U11704 ( .A1(n14597), .A2(n11990), .ZN(n10106) );
  INV_X1 U11705 ( .A(n14601), .ZN(n11990) );
  INV_X1 U11706 ( .A(n12096), .ZN(n12074) );
  NOR2_X1 U11707 ( .A1(n14257), .A2(n16236), .ZN(n12096) );
  NOR2_X1 U11708 ( .A1(n14207), .A2(n11738), .ZN(n10105) );
  INV_X1 U11709 ( .A(n13901), .ZN(n12099) );
  INV_X1 U11710 ( .A(n11643), .ZN(n11644) );
  INV_X1 U11711 ( .A(n11632), .ZN(n10099) );
  INV_X1 U11712 ( .A(n11669), .ZN(n12046) );
  NAND2_X1 U11713 ( .A1(n9914), .A2(n14598), .ZN(n9913) );
  INV_X1 U11714 ( .A(n11500), .ZN(n9914) );
  INV_X1 U11715 ( .A(n14604), .ZN(n9915) );
  NAND2_X1 U11716 ( .A1(n9929), .A2(n11300), .ZN(n9928) );
  NOR2_X1 U11717 ( .A1(n9818), .A2(n9931), .ZN(n9930) );
  INV_X1 U11718 ( .A(n11263), .ZN(n11261) );
  INV_X1 U11719 ( .A(n11554), .ZN(n11478) );
  INV_X1 U11720 ( .A(n11025), .ZN(n11513) );
  NOR2_X1 U11721 ( .A1(n11096), .A2(n10097), .ZN(n10096) );
  INV_X1 U11722 ( .A(n11077), .ZN(n10097) );
  AND2_X1 U11723 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10915) );
  NAND2_X1 U11724 ( .A1(n10665), .A2(n10669), .ZN(n10662) );
  INV_X1 U11725 ( .A(n10614), .ZN(n9947) );
  OR2_X1 U11726 ( .A1(n10609), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10611) );
  OR2_X1 U11727 ( .A1(n10625), .A2(n9945), .ZN(n9944) );
  NOR2_X1 U11728 ( .A1(n10580), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U11729 ( .A1(n10592), .A2(n10669), .ZN(n10590) );
  OAI21_X1 U11730 ( .B1(n9774), .B2(n14456), .A(n15009), .ZN(n9999) );
  INV_X1 U11731 ( .A(n15047), .ZN(n10005) );
  AND2_X1 U11732 ( .A1(n13143), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13144) );
  NAND2_X1 U11733 ( .A1(n9968), .A2(n12793), .ZN(n9967) );
  INV_X1 U11734 ( .A(n14948), .ZN(n9968) );
  NAND2_X1 U11735 ( .A1(n12956), .A2(n9835), .ZN(n9961) );
  INV_X1 U11736 ( .A(n15036), .ZN(n9958) );
  AND4_X1 U11737 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  INV_X1 U11738 ( .A(n14979), .ZN(n9982) );
  NOR2_X1 U11739 ( .A1(n9993), .A2(n13753), .ZN(n9992) );
  INV_X1 U11740 ( .A(n15565), .ZN(n9993) );
  AND2_X1 U11741 ( .A1(n13307), .A2(n10750), .ZN(n9970) );
  NOR2_X1 U11742 ( .A1(n9989), .A2(n13666), .ZN(n9988) );
  INV_X1 U11743 ( .A(n13620), .ZN(n9989) );
  AND2_X1 U11744 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  INV_X1 U11745 ( .A(n13297), .ZN(n9972) );
  INV_X1 U11746 ( .A(n12810), .ZN(n12838) );
  NAND2_X1 U11747 ( .A1(n9879), .A2(n10849), .ZN(n9862) );
  NAND2_X1 U11748 ( .A1(n10230), .A2(n13494), .ZN(n12369) );
  AND2_X1 U11749 ( .A1(n12214), .A2(n19668), .ZN(n12215) );
  NAND2_X1 U11750 ( .A1(n10228), .A2(n10217), .ZN(n10220) );
  NAND3_X1 U11751 ( .A1(n9747), .A2(n10227), .A3(n19215), .ZN(n10232) );
  OR2_X2 U11752 ( .A1(n13207), .A2(n13197), .ZN(n10316) );
  NAND2_X1 U11753 ( .A1(n10307), .A2(n10306), .ZN(n10374) );
  AND4_X1 U11754 ( .A1(n10228), .A2(n10227), .A3(n10222), .A4(n15654), .ZN(
        n10229) );
  INV_X1 U11755 ( .A(n18209), .ZN(n12657) );
  NOR2_X1 U11756 ( .A1(n12420), .A2(n16910), .ZN(n12461) );
  NOR2_X1 U11757 ( .A1(n18236), .A2(n12707), .ZN(n12721) );
  NAND2_X1 U11758 ( .A1(n10051), .A2(n17770), .ZN(n12533) );
  AND2_X1 U11759 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12524), .ZN(
        n12525) );
  XOR2_X1 U11760 ( .A(n17353), .B(n12523), .Z(n12524) );
  INV_X1 U11761 ( .A(n17359), .ZN(n12687) );
  XNOR2_X1 U11762 ( .A(n12512), .B(n12511), .ZN(n12513) );
  NAND2_X1 U11763 ( .A1(n12719), .A2(n18214), .ZN(n9895) );
  INV_X1 U11764 ( .A(n13537), .ZN(n13134) );
  NOR2_X1 U11765 ( .A1(n13912), .A2(n13911), .ZN(n13919) );
  INV_X1 U11766 ( .A(n14621), .ZN(n9908) );
  NAND2_X1 U11767 ( .A1(n11403), .A2(n11402), .ZN(n11404) );
  INV_X1 U11768 ( .A(n11401), .ZN(n11403) );
  NAND2_X1 U11769 ( .A1(n13287), .A2(n11548), .ZN(n9901) );
  INV_X1 U11770 ( .A(n13565), .ZN(n13564) );
  AND2_X1 U11771 ( .A1(n12055), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12056) );
  NAND2_X1 U11772 ( .A1(n12027), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12054) );
  INV_X1 U11773 ( .A(n11985), .ZN(n11986) );
  NAND2_X1 U11774 ( .A1(n11987), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12026) );
  NAND2_X1 U11775 ( .A1(n10048), .A2(n10047), .ZN(n10046) );
  NOR2_X1 U11776 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U11777 ( .A1(n11848), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11851) );
  NAND2_X1 U11778 ( .A1(n11668), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11677) );
  NAND2_X1 U11779 ( .A1(n11645), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11654) );
  NOR2_X2 U11780 ( .A1(n9788), .A2(n11556), .ZN(n12894) );
  NAND2_X1 U11781 ( .A1(n14186), .A2(n14185), .ZN(n14194) );
  AND2_X1 U11782 ( .A1(n11519), .A2(n11518), .ZN(n13509) );
  NAND2_X1 U11783 ( .A1(n11293), .A2(n10038), .ZN(n10037) );
  INV_X1 U11784 ( .A(n16089), .ZN(n10038) );
  NAND2_X1 U11785 ( .A1(n9707), .A2(n16088), .ZN(n10035) );
  NAND2_X1 U11786 ( .A1(n13765), .A2(n13764), .ZN(n13763) );
  NAND2_X1 U11787 ( .A1(n9900), .A2(n9779), .ZN(n19977) );
  NAND2_X1 U11788 ( .A1(n20115), .A2(n13588), .ZN(n20292) );
  INV_X1 U11789 ( .A(n20187), .ZN(n20354) );
  NOR2_X1 U11790 ( .A1(n14046), .A2(n14045), .ZN(n20494) );
  INV_X1 U11791 ( .A(n13953), .ZN(n14046) );
  OR2_X1 U11792 ( .A1(n13133), .A2(n13134), .ZN(n15821) );
  OR2_X1 U11793 ( .A1(n10032), .A2(n10027), .ZN(n10025) );
  OAI21_X1 U11794 ( .B1(n10642), .B2(n10646), .A(n10641), .ZN(n10645) );
  OR2_X1 U11795 ( .A1(n10032), .A2(n10033), .ZN(n10031) );
  NAND2_X1 U11796 ( .A1(n9952), .A2(n10565), .ZN(n9951) );
  INV_X1 U11797 ( .A(n10570), .ZN(n9952) );
  OR2_X1 U11798 ( .A1(n10574), .A2(n10428), .ZN(n10669) );
  NAND2_X1 U11799 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  NAND2_X1 U11800 ( .A1(n10428), .A2(n10437), .ZN(n9938) );
  NAND2_X1 U11801 ( .A1(n12214), .A2(n12228), .ZN(n9939) );
  AND2_X1 U11802 ( .A1(n13305), .A2(n13304), .ZN(n13553) );
  NOR2_X1 U11803 ( .A1(n9997), .A2(n15013), .ZN(n10002) );
  NAND2_X1 U11804 ( .A1(n9774), .A2(n14456), .ZN(n9997) );
  INV_X1 U11805 ( .A(n10867), .ZN(n9887) );
  INV_X1 U11806 ( .A(n16338), .ZN(n9886) );
  OR3_X1 U11807 ( .A1(n10689), .A2(n10861), .A3(n14289), .ZN(n15124) );
  AOI21_X1 U11808 ( .B1(n15143), .B2(n9846), .A(n10090), .ZN(n10094) );
  NAND2_X1 U11809 ( .A1(n16246), .A2(n10660), .ZN(n10681) );
  NAND2_X1 U11810 ( .A1(n14135), .A2(n12366), .ZN(n14123) );
  NOR2_X1 U11811 ( .A1(n9783), .A2(n14120), .ZN(n9962) );
  INV_X1 U11812 ( .A(n14137), .ZN(n9963) );
  NAND2_X1 U11813 ( .A1(n9868), .A2(n9867), .ZN(n9866) );
  NAND2_X1 U11814 ( .A1(n15629), .A2(n14244), .ZN(n9867) );
  AND2_X1 U11815 ( .A1(n10855), .A2(n10857), .ZN(n10064) );
  CLKBUF_X1 U11816 ( .A(n12367), .Z(n12368) );
  INV_X1 U11817 ( .A(n9985), .ZN(n9987) );
  NOR2_X1 U11818 ( .A1(n13772), .A2(n13192), .ZN(n13193) );
  INV_X1 U11819 ( .A(n9811), .ZN(n13093) );
  INV_X1 U11820 ( .A(n19581), .ZN(n19852) );
  NOR2_X1 U11821 ( .A1(n20708), .A2(n19877), .ZN(n19232) );
  NAND2_X1 U11822 ( .A1(n10072), .A2(n10304), .ZN(n19451) );
  INV_X1 U11823 ( .A(n19232), .ZN(n19479) );
  NAND2_X1 U11824 ( .A1(n19723), .A2(n19668), .ZN(n19581) );
  OR2_X1 U11825 ( .A1(n20708), .A2(n19874), .ZN(n19856) );
  AND2_X1 U11826 ( .A1(n20708), .A2(n19874), .ZN(n19616) );
  INV_X1 U11827 ( .A(n19419), .ZN(n19728) );
  NAND2_X1 U11828 ( .A1(n10825), .A2(n10824), .ZN(n19621) );
  AND2_X1 U11829 ( .A1(n9761), .A2(n10243), .ZN(n13491) );
  NOR3_X1 U11830 ( .A1(n16538), .A2(n16537), .A3(n16536), .ZN(n18631) );
  NOR2_X1 U11831 ( .A1(n15758), .A2(n18833), .ZN(n17380) );
  NOR2_X1 U11832 ( .A1(n17353), .A2(n12523), .ZN(n16416) );
  INV_X1 U11833 ( .A(n12540), .ZN(n12541) );
  XNOR2_X1 U11834 ( .A(n12513), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10059) );
  INV_X1 U11835 ( .A(n18835), .ZN(n18206) );
  AND2_X1 U11836 ( .A1(n20589), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13171) );
  OR2_X1 U11837 ( .A1(n20681), .A2(n13903), .ZN(n20009) );
  INV_X1 U11838 ( .A(n14803), .ZN(n20067) );
  NOR2_X2 U11839 ( .A1(n15821), .A2(n13277), .ZN(n20071) );
  OR2_X1 U11840 ( .A1(n14824), .A2(n14823), .ZN(n9922) );
  OR2_X1 U11841 ( .A1(n9813), .A2(n9923), .ZN(n9918) );
  INV_X1 U11842 ( .A(n9920), .ZN(n9919) );
  AOI211_X1 U11843 ( .C1(n14511), .C2(n11553), .A(n9921), .B(n14515), .ZN(
        n9920) );
  NOR2_X1 U11844 ( .A1(n14511), .A2(n14512), .ZN(n9921) );
  AND2_X1 U11845 ( .A1(n11521), .A2(n11398), .ZN(n20103) );
  CLKBUF_X1 U11846 ( .A(n13948), .Z(n20436) );
  OR2_X1 U11847 ( .A1(n20529), .A2(n20324), .ZN(n20491) );
  INV_X1 U11848 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19723) );
  CLKBUF_X1 U11849 ( .A(n12791), .Z(n19009) );
  AND2_X1 U11850 ( .A1(n13243), .A2(n13242), .ZN(n13244) );
  AND2_X1 U11851 ( .A1(n13555), .A2(n12309), .ZN(n10004) );
  OR2_X1 U11852 ( .A1(n12321), .A2(n12320), .ZN(n13557) );
  NOR2_X1 U11853 ( .A1(n13772), .A2(n13109), .ZN(n19444) );
  OAI21_X1 U11854 ( .B1(n15125), .B2(n15126), .A(n10692), .ZN(n10698) );
  NAND2_X1 U11855 ( .A1(n12860), .A2(n12859), .ZN(n12861) );
  NAND2_X1 U11856 ( .A1(n12845), .A2(n16354), .ZN(n12860) );
  NOR3_X1 U11857 ( .A1(n12858), .A2(n12857), .A3(n12856), .ZN(n12859) );
  NAND2_X1 U11858 ( .A1(n9966), .A2(n12909), .ZN(n15361) );
  NAND2_X1 U11859 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  INV_X1 U11860 ( .A(n12193), .ZN(n9865) );
  AND2_X1 U11861 ( .A1(n12377), .A2(n12213), .ZN(n16359) );
  INV_X1 U11862 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19890) );
  INV_X1 U11863 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19881) );
  INV_X1 U11864 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19871) );
  INV_X1 U11865 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19864) );
  NAND2_X1 U11866 ( .A1(n13224), .A2(n13245), .ZN(n19445) );
  OR2_X1 U11867 ( .A1(n13222), .A2(n13223), .ZN(n13224) );
  AND2_X1 U11868 ( .A1(n19414), .A2(n19868), .ZN(n19344) );
  INV_X1 U11869 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U11870 ( .A1(n18699), .A2(n18632), .ZN(n17443) );
  INV_X1 U11871 ( .A(n17249), .ZN(n17244) );
  AND2_X1 U11872 ( .A1(n17379), .A2(n17280), .ZN(n17295) );
  NAND2_X1 U11873 ( .A1(n17379), .A2(n9896), .ZN(n17323) );
  NOR3_X1 U11874 ( .A1(n17321), .A2(n17233), .A3(n9897), .ZN(n9896) );
  AOI21_X1 U11875 ( .B1(n12880), .B2(n17781), .A(n12879), .ZN(n12881) );
  NAND2_X1 U11876 ( .A1(n17533), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17519) );
  NOR2_X2 U11877 ( .A1(n10049), .A2(n17874), .ZN(n17765) );
  INV_X1 U11878 ( .A(n17863), .ZN(n17874) );
  AOI21_X1 U11879 ( .B1(n12880), .B2(n18107), .A(n12739), .ZN(n12740) );
  NAND2_X1 U11880 ( .A1(n18798), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10055) );
  AOI21_X2 U11881 ( .B1(n12676), .B2(n12675), .A(n18692), .ZN(n18182) );
  AOI211_X1 U11882 ( .C1(n12669), .C2(n18635), .A(n12668), .B(n15759), .ZN(
        n12676) );
  OAI21_X1 U11883 ( .B1(n19480), .B2(n10305), .A(n13143), .ZN(n10310) );
  OAI21_X1 U11884 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18807), .A(
        n12637), .ZN(n12638) );
  INV_X1 U11885 ( .A(n16067), .ZN(n9931) );
  NOR2_X1 U11886 ( .A1(n11236), .A2(n11214), .ZN(n9936) );
  OR2_X1 U11887 ( .A1(n11209), .A2(n11208), .ZN(n11240) );
  AND2_X1 U11888 ( .A1(n11017), .A2(n11008), .ZN(n11371) );
  NAND2_X1 U11889 ( .A1(n13574), .A2(n11328), .ZN(n11175) );
  INV_X1 U11890 ( .A(n11140), .ZN(n11192) );
  OR2_X1 U11891 ( .A1(n11187), .A2(n11186), .ZN(n11241) );
  OAI21_X1 U11892 ( .B1(n10436), .B2(n10428), .A(n10435), .ZN(n10443) );
  NAND2_X1 U11893 ( .A1(n10428), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10435) );
  INV_X1 U11894 ( .A(n10710), .ZN(n10436) );
  INV_X1 U11895 ( .A(n12173), .ZN(n10204) );
  INV_X1 U11896 ( .A(n10654), .ZN(n10076) );
  OR2_X1 U11897 ( .A1(n10366), .A2(n10365), .ZN(n12237) );
  NAND2_X1 U11898 ( .A1(n10297), .A2(n19008), .ZN(n10320) );
  INV_X1 U11899 ( .A(n10320), .ZN(n10321) );
  NAND2_X1 U11900 ( .A1(n18203), .A2(n18835), .ZN(n12713) );
  NAND2_X1 U11901 ( .A1(n12657), .A2(n12713), .ZN(n12660) );
  NOR2_X1 U11902 ( .A1(n11355), .A2(n11354), .ZN(n11384) );
  INV_X1 U11903 ( .A(n15854), .ZN(n10048) );
  NAND2_X1 U11904 ( .A1(n14809), .A2(n11296), .ZN(n14778) );
  OR2_X1 U11905 ( .A1(n11058), .A2(n11057), .ZN(n11286) );
  NAND2_X1 U11906 ( .A1(n11271), .A2(n10045), .ZN(n10043) );
  INV_X1 U11907 ( .A(n11248), .ZN(n10045) );
  OR2_X1 U11908 ( .A1(n11258), .A2(n11257), .ZN(n11279) );
  AND2_X1 U11909 ( .A1(n11144), .A2(n11022), .ZN(n11313) );
  INV_X1 U11910 ( .A(n11286), .ZN(n11290) );
  NAND2_X1 U11911 ( .A1(n9925), .A2(n11100), .ZN(n9924) );
  AND2_X1 U11912 ( .A1(n11103), .A2(n11102), .ZN(n11104) );
  INV_X1 U11913 ( .A(n11287), .ZN(n11107) );
  OR2_X1 U11914 ( .A1(n11093), .A2(n11092), .ZN(n11155) );
  AND2_X1 U11915 ( .A1(n11359), .A2(n11313), .ZN(n11353) );
  INV_X1 U11916 ( .A(n11338), .ZN(n11323) );
  OR2_X1 U11917 ( .A1(n11355), .A2(n11321), .ZN(n11322) );
  INV_X1 U11918 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15810) );
  INV_X1 U11919 ( .A(n12237), .ZN(n10843) );
  NAND2_X1 U11920 ( .A1(n10615), .A2(n9948), .ZN(n10599) );
  NOR2_X1 U11921 ( .A1(n10606), .A2(n9949), .ZN(n9948) );
  NAND2_X1 U11922 ( .A1(n10602), .A2(n10614), .ZN(n9949) );
  NOR2_X1 U11923 ( .A1(n10832), .A2(n10021), .ZN(n10020) );
  INV_X1 U11924 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U11925 ( .A1(n10831), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10832) );
  NAND2_X1 U11926 ( .A1(n10590), .A2(n10591), .ZN(n10627) );
  AND2_X1 U11927 ( .A1(n10428), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10573) );
  NOR2_X1 U11928 ( .A1(n19215), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12226) );
  INV_X1 U11929 ( .A(n12954), .ZN(n9981) );
  NAND2_X1 U11930 ( .A1(n13870), .A2(n10008), .ZN(n10007) );
  INV_X1 U11931 ( .A(n16291), .ZN(n10008) );
  NOR2_X1 U11932 ( .A1(n12941), .A2(n10834), .ZN(n10015) );
  NAND2_X1 U11933 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10017) );
  AND2_X1 U11934 ( .A1(n10020), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10019) );
  NAND2_X1 U11935 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10829) );
  AND2_X1 U11936 ( .A1(n13492), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10239) );
  XNOR2_X1 U11937 ( .A(n10443), .B(n9937), .ZN(n10445) );
  NAND2_X1 U11938 ( .A1(n9744), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10261) );
  OR2_X1 U11939 ( .A1(n10068), .A2(n15406), .ZN(n10067) );
  NAND2_X1 U11940 ( .A1(n10069), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10068) );
  INV_X1 U11941 ( .A(n15430), .ZN(n10069) );
  INV_X1 U11942 ( .A(n15449), .ZN(n9959) );
  AND2_X1 U11943 ( .A1(n10630), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10084) );
  AOI21_X1 U11944 ( .B1(n10082), .B2(n10087), .A(n10081), .ZN(n10080) );
  OAI21_X1 U11945 ( .B1(n10088), .B2(n10633), .A(n10687), .ZN(n10081) );
  NOR2_X1 U11946 ( .A1(n10630), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10082) );
  INV_X1 U11947 ( .A(n12372), .ZN(n9964) );
  NAND2_X1 U11948 ( .A1(n15314), .A2(n10586), .ZN(n12202) );
  NAND2_X1 U11949 ( .A1(n9890), .A2(n9889), .ZN(n10855) );
  AND2_X1 U11950 ( .A1(n10736), .A2(n13249), .ZN(n9973) );
  INV_X1 U11951 ( .A(n13263), .ZN(n10736) );
  NOR2_X1 U11952 ( .A1(n10508), .A2(n10507), .ZN(n12253) );
  OR2_X1 U11953 ( .A1(n10530), .A2(n10519), .ZN(n10518) );
  OAI21_X1 U11954 ( .B1(n9980), .B2(n9979), .A(n10334), .ZN(n9978) );
  OAI21_X1 U11955 ( .B1(n9977), .B2(n9976), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U11956 ( .A1(n10352), .A2(n10351), .ZN(n12228) );
  INV_X1 U11957 ( .A(n12236), .ZN(n12361) );
  OR2_X1 U11958 ( .A1(n10390), .A2(n10389), .ZN(n12243) );
  AND3_X1 U11959 ( .A1(n12138), .A2(n12127), .A3(n12133), .ZN(n10706) );
  NAND2_X1 U11960 ( .A1(n9778), .A2(n9805), .ZN(n9873) );
  NAND2_X1 U11961 ( .A1(n9872), .A2(n9806), .ZN(n9871) );
  AOI21_X1 U11962 ( .B1(n10231), .B2(n10822), .A(n10821), .ZN(n12142) );
  INV_X1 U11963 ( .A(n17159), .ZN(n12410) );
  NOR2_X1 U11964 ( .A1(n12417), .A2(n12420), .ZN(n12549) );
  INV_X1 U11965 ( .A(n17182), .ZN(n17093) );
  INV_X1 U11966 ( .A(n12710), .ZN(n12716) );
  NOR2_X1 U11967 ( .A1(n17505), .A2(n17866), .ZN(n16546) );
  NOR2_X1 U11968 ( .A1(n17691), .A2(n17690), .ZN(n16687) );
  NOR2_X1 U11969 ( .A1(n12686), .A2(n17836), .ZN(n12689) );
  OAI21_X1 U11970 ( .B1(n12650), .B2(n12649), .A(n12648), .ZN(n12673) );
  NOR2_X1 U11971 ( .A1(n12601), .A2(n12600), .ZN(n12711) );
  INV_X1 U11972 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15986) );
  INV_X1 U11973 ( .A(n14627), .ZN(n9906) );
  AND2_X1 U11974 ( .A1(n11692), .A2(n11691), .ZN(n13893) );
  AND2_X1 U11975 ( .A1(n14695), .A2(n12394), .ZN(n13548) );
  NOR2_X1 U11976 ( .A1(n12026), .A2(n15891), .ZN(n12027) );
  AND2_X1 U11977 ( .A1(n12032), .A2(n12031), .ZN(n14588) );
  OR2_X1 U11978 ( .A1(n15875), .A2(n13901), .ZN(n12031) );
  AND2_X1 U11979 ( .A1(n15882), .A2(n12099), .ZN(n12006) );
  NAND2_X1 U11980 ( .A1(n11989), .A2(n11988), .ZN(n14601) );
  NOR2_X1 U11981 ( .A1(n11920), .A2(n15922), .ZN(n11921) );
  NAND2_X1 U11982 ( .A1(n11921), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11985) );
  NOR2_X1 U11983 ( .A1(n11884), .A2(n15933), .ZN(n11885) );
  NAND2_X1 U11984 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11885), .ZN(
        n11920) );
  NOR2_X1 U11985 ( .A1(n11851), .A2(n14772), .ZN(n11852) );
  NAND2_X1 U11986 ( .A1(n11852), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11884) );
  AND2_X1 U11987 ( .A1(n11850), .A2(n11849), .ZN(n14568) );
  OR2_X1 U11988 ( .A1(n11804), .A2(n15966), .ZN(n11805) );
  NOR2_X1 U11989 ( .A1(n20907), .A2(n11805), .ZN(n11848) );
  CLKBUF_X1 U11990 ( .A(n14190), .Z(n14191) );
  NAND2_X1 U11991 ( .A1(n11754), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U11992 ( .A1(n11803), .A2(n10103), .ZN(n10102) );
  INV_X1 U11993 ( .A(n10105), .ZN(n10103) );
  AND2_X1 U11994 ( .A1(n11802), .A2(n14169), .ZN(n11803) );
  NOR2_X1 U11995 ( .A1(n11770), .A2(n15975), .ZN(n11754) );
  OR2_X1 U11996 ( .A1(n11796), .A2(n15986), .ZN(n11770) );
  NAND2_X1 U11997 ( .A1(n11723), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11796) );
  NOR2_X1 U11998 ( .A1(n20950), .A2(n11677), .ZN(n11717) );
  AOI21_X1 U11999 ( .B1(n11674), .B2(n11763), .A(n11673), .ZN(n13781) );
  CLKBUF_X1 U12000 ( .A(n13778), .Z(n13779) );
  INV_X1 U12001 ( .A(n11661), .ZN(n11662) );
  NAND2_X1 U12002 ( .A1(n11662), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11667) );
  INV_X1 U12003 ( .A(n11654), .ZN(n11655) );
  NAND2_X1 U12004 ( .A1(n11655), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11661) );
  NAND2_X1 U12005 ( .A1(n11644), .A2(n11763), .ZN(n11652) );
  NAND2_X1 U12006 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11635) );
  NOR2_X1 U12007 ( .A1(n11635), .A2(n11634), .ZN(n11645) );
  INV_X1 U12008 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11634) );
  CLKBUF_X1 U12009 ( .A(n13329), .Z(n13330) );
  INV_X1 U12010 ( .A(n11613), .ZN(n10101) );
  AOI21_X1 U12011 ( .B1(n11613), .B2(n10100), .A(n10099), .ZN(n10098) );
  INV_X1 U12012 ( .A(n10041), .ZN(n14709) );
  NAND2_X1 U12013 ( .A1(n10041), .A2(n16056), .ZN(n10040) );
  NAND2_X1 U12014 ( .A1(n9912), .A2(n9911), .ZN(n9910) );
  INV_X1 U12015 ( .A(n9913), .ZN(n9912) );
  NOR2_X1 U12016 ( .A1(n9915), .A2(n14590), .ZN(n9911) );
  NOR2_X1 U12017 ( .A1(n11536), .A2(n11535), .ZN(n14740) );
  NOR3_X1 U12018 ( .A1(n14618), .A2(n9915), .A3(n11500), .ZN(n14607) );
  NOR2_X1 U12019 ( .A1(n14618), .A2(n11500), .ZN(n14605) );
  NOR3_X1 U12020 ( .A1(n15959), .A2(n11488), .A3(n11477), .ZN(n15856) );
  NAND2_X1 U12021 ( .A1(n9928), .A2(n11301), .ZN(n9927) );
  INV_X1 U12022 ( .A(n15985), .ZN(n9904) );
  NAND2_X1 U12023 ( .A1(n14209), .A2(n14208), .ZN(n15984) );
  AND2_X1 U12024 ( .A1(n11443), .A2(n11442), .ZN(n14107) );
  AND2_X1 U12025 ( .A1(n11430), .A2(n11429), .ZN(n16217) );
  AND2_X1 U12026 ( .A1(n11426), .A2(n11425), .ZN(n13731) );
  NOR2_X1 U12027 ( .A1(n11409), .A2(n13326), .ZN(n9902) );
  INV_X1 U12028 ( .A(n16172), .ZN(n20097) );
  XNOR2_X1 U12029 ( .A(n11409), .B(n13200), .ZN(n13287) );
  AND2_X1 U12030 ( .A1(n11521), .A2(n11517), .ZN(n16168) );
  NAND2_X1 U12031 ( .A1(n13605), .A2(n11104), .ZN(n11124) );
  NAND2_X1 U12032 ( .A1(n11110), .A2(n11109), .ZN(n11617) );
  NAND2_X1 U12033 ( .A1(n11215), .A2(n11191), .ZN(n20117) );
  CLKBUF_X1 U12034 ( .A(n11368), .Z(n13130) );
  CLKBUF_X1 U12035 ( .A(n11112), .Z(n11113) );
  INV_X1 U12036 ( .A(n13171), .ZN(n13277) );
  INV_X1 U12037 ( .A(n15800), .ZN(n13533) );
  AND3_X1 U12038 ( .A1(n10229), .A2(n13156), .A3(n10243), .ZN(n12819) );
  NAND2_X1 U12039 ( .A1(n9811), .A2(n12828), .ZN(n12123) );
  NAND2_X1 U12040 ( .A1(n10434), .A2(n10433), .ZN(n10710) );
  NAND2_X1 U12041 ( .A1(n12828), .A2(n12128), .ZN(n10433) );
  NAND2_X1 U12042 ( .A1(n10843), .A2(n10429), .ZN(n10434) );
  INV_X1 U12043 ( .A(n12137), .ZN(n10822) );
  NOR2_X1 U12044 ( .A1(n10676), .A2(n10675), .ZN(n10685) );
  AND2_X1 U12045 ( .A1(n15026), .A2(n20956), .ZN(n9956) );
  NAND2_X1 U12046 ( .A1(n10662), .A2(n10663), .ZN(n10676) );
  AND2_X1 U12047 ( .A1(n10025), .A2(n10023), .ZN(n10022) );
  INV_X1 U12048 ( .A(n16259), .ZN(n10023) );
  INV_X1 U12049 ( .A(n15184), .ZN(n10027) );
  OR2_X1 U12050 ( .A1(n16270), .A2(n10032), .ZN(n10028) );
  AND2_X1 U12051 ( .A1(n10031), .A2(n16321), .ZN(n10029) );
  INV_X1 U12052 ( .A(n15211), .ZN(n10033) );
  OR2_X1 U12053 ( .A1(n14983), .A2(n10032), .ZN(n10034) );
  AND2_X1 U12054 ( .A1(n10615), .A2(n9946), .ZN(n10604) );
  NOR2_X1 U12055 ( .A1(n10606), .A2(n9947), .ZN(n9946) );
  NAND2_X1 U12056 ( .A1(n10011), .A2(n10010), .ZN(n10013) );
  INV_X1 U12057 ( .A(n15248), .ZN(n10010) );
  INV_X1 U12058 ( .A(n18900), .ZN(n10011) );
  NOR2_X1 U12059 ( .A1(n9944), .A2(n9821), .ZN(n9943) );
  INV_X1 U12060 ( .A(n9944), .ZN(n9942) );
  OR2_X1 U12061 ( .A1(n9953), .A2(n9950), .ZN(n10571) );
  INV_X1 U12062 ( .A(n10565), .ZN(n9950) );
  NOR2_X1 U12063 ( .A1(n13476), .A2(n13026), .ZN(n12977) );
  BUF_X1 U12064 ( .A(n10286), .Z(n10818) );
  NOR2_X1 U12065 ( .A1(n14137), .A2(n14136), .ZN(n14138) );
  CLKBUF_X1 U12066 ( .A(n13941), .Z(n19025) );
  NAND2_X1 U12067 ( .A1(n10000), .A2(n9998), .ZN(n15008) );
  AOI21_X1 U12068 ( .B1(n15013), .B2(n10003), .A(n9999), .ZN(n9998) );
  OR2_X1 U12069 ( .A1(n16287), .A2(n15044), .ZN(n16280) );
  CLKBUF_X1 U12070 ( .A(n15041), .Z(n15042) );
  NOR2_X1 U12071 ( .A1(n13869), .A2(n10007), .ZN(n16294) );
  NAND2_X1 U12072 ( .A1(n10006), .A2(n13870), .ZN(n16292) );
  INV_X1 U12073 ( .A(n13869), .ZN(n10006) );
  INV_X1 U12074 ( .A(n12933), .ZN(n15651) );
  CLKBUF_X1 U12075 ( .A(n12784), .Z(n12785) );
  INV_X1 U12076 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U12077 ( .A1(n10271), .A2(n10270), .ZN(n10301) );
  NOR2_X1 U12078 ( .A1(n10341), .A2(n10340), .ZN(n13099) );
  NAND2_X1 U12079 ( .A1(n11596), .A2(n10095), .ZN(n10089) );
  OR2_X1 U12080 ( .A1(n12940), .A2(n10861), .ZN(n15139) );
  NOR2_X1 U12081 ( .A1(n10655), .A2(n15422), .ZN(n15178) );
  NAND2_X1 U12082 ( .A1(n12956), .A2(n9833), .ZN(n15451) );
  AND4_X1 U12083 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10419) );
  AND4_X1 U12084 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10420) );
  AND4_X1 U12085 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10421) );
  AND2_X1 U12086 ( .A1(n12850), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10070) );
  INV_X1 U12087 ( .A(n13824), .ZN(n10763) );
  AND2_X1 U12088 ( .A1(n9992), .A2(n15536), .ZN(n9991) );
  NAND2_X1 U12089 ( .A1(n15568), .A2(n15539), .ZN(n9877) );
  INV_X1 U12090 ( .A(n13723), .ZN(n9969) );
  INV_X1 U12091 ( .A(n9861), .ZN(n9860) );
  NAND2_X1 U12092 ( .A1(n10450), .A2(n10449), .ZN(n13800) );
  NAND2_X2 U12093 ( .A1(n10243), .A2(n12217), .ZN(n12828) );
  AND3_X1 U12094 ( .A1(n10228), .A2(n10216), .A3(n15654), .ZN(n10224) );
  CLKBUF_X1 U12095 ( .A(n12373), .Z(n12374) );
  NOR2_X1 U12096 ( .A1(n13216), .A2(n9995), .ZN(n9994) );
  INV_X1 U12097 ( .A(n13213), .ZN(n9995) );
  NAND2_X1 U12099 ( .A1(n19857), .A2(n19444), .ZN(n19609) );
  AND2_X1 U12100 ( .A1(n19621), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19216) );
  NOR2_X1 U12101 ( .A1(n12657), .A2(n18650), .ZN(n12712) );
  NOR2_X1 U12102 ( .A1(n17526), .A2(n16616), .ZN(n16615) );
  NOR2_X1 U12103 ( .A1(n16549), .A2(n16551), .ZN(n17535) );
  NOR2_X1 U12104 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16693), .ZN(n16678) );
  NOR2_X1 U12105 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16855), .ZN(n16846) );
  NOR2_X1 U12106 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16880), .ZN(n16869) );
  NAND2_X1 U12107 ( .A1(n18853), .A2(n16540), .ZN(n16544) );
  NAND2_X1 U12108 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16985), .ZN(n16979) );
  INV_X1 U12109 ( .A(n18203), .ZN(n16540) );
  NOR2_X1 U12110 ( .A1(n17387), .A2(n17389), .ZN(n9893) );
  OR2_X1 U12111 ( .A1(n12457), .A2(n12456), .ZN(n12512) );
  NAND2_X1 U12112 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12458) );
  NOR2_X1 U12113 ( .A1(n18227), .A2(n12711), .ZN(n18664) );
  NAND4_X1 U12114 ( .A1(n16540), .A2(n12721), .A3(n12711), .A4(n12716), .ZN(
        n17441) );
  CLKBUF_X1 U12115 ( .A(n16546), .Z(n16559) );
  NAND2_X1 U12116 ( .A1(n17525), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17505) );
  NOR2_X1 U12117 ( .A1(n17611), .A2(n17587), .ZN(n16552) );
  NAND2_X1 U12118 ( .A1(n16687), .A2(n17667), .ZN(n17652) );
  INV_X1 U12119 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17680) );
  NAND2_X1 U12120 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17709) );
  NAND2_X1 U12121 ( .A1(n16783), .A2(n10118), .ZN(n17734) );
  NOR2_X1 U12122 ( .A1(n12705), .A2(n17779), .ZN(n17739) );
  NOR2_X1 U12123 ( .A1(n12699), .A2(n12703), .ZN(n12705) );
  NOR2_X1 U12124 ( .A1(n17801), .A2(n17808), .ZN(n16783) );
  NOR2_X1 U12125 ( .A1(n16421), .A2(n16400), .ZN(n15772) );
  NAND2_X1 U12126 ( .A1(n16394), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10057) );
  NOR2_X1 U12127 ( .A1(n10054), .A2(n9841), .ZN(n10053) );
  INV_X1 U12128 ( .A(n12548), .ZN(n10054) );
  NOR2_X1 U12129 ( .A1(n17603), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10052) );
  NOR2_X1 U12130 ( .A1(n17512), .A2(n10107), .ZN(n15776) );
  NOR2_X1 U12131 ( .A1(n17538), .A2(n17880), .ZN(n17877) );
  AND2_X1 U12132 ( .A1(n17541), .A2(n10108), .ZN(n12538) );
  NOR2_X1 U12133 ( .A1(n17563), .A2(n12537), .ZN(n17554) );
  INV_X1 U12134 ( .A(n12536), .ZN(n12537) );
  OAI21_X1 U12135 ( .B1(n17661), .B2(n12723), .A(n12535), .ZN(n12536) );
  NOR2_X1 U12136 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17605), .ZN(
        n17583) );
  AND2_X1 U12137 ( .A1(n12533), .A2(n10109), .ZN(n12531) );
  AND2_X1 U12138 ( .A1(n12724), .A2(n12533), .ZN(n17661) );
  NOR2_X1 U12139 ( .A1(n17694), .A2(n17674), .ZN(n17695) );
  OAI21_X1 U12140 ( .B1(n12722), .B2(n12727), .A(n18649), .ZN(n18663) );
  AOI21_X1 U12141 ( .B1(n12704), .B2(n12703), .A(n12702), .ZN(n17780) );
  NOR2_X1 U12142 ( .A1(n12529), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17769) );
  NOR2_X1 U12143 ( .A1(n18124), .A2(n17804), .ZN(n17803) );
  NAND2_X1 U12144 ( .A1(n10062), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10061) );
  NOR2_X1 U12145 ( .A1(n17812), .A2(n17811), .ZN(n17810) );
  OR2_X1 U12146 ( .A1(n17814), .A2(n17815), .ZN(n10063) );
  NOR2_X1 U12147 ( .A1(n17838), .A2(n17837), .ZN(n17836) );
  NAND2_X1 U12148 ( .A1(n17869), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17868) );
  INV_X1 U12149 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12635) );
  INV_X1 U12150 ( .A(n18661), .ZN(n18644) );
  INV_X1 U12151 ( .A(n18650), .ZN(n9894) );
  NAND3_X1 U12152 ( .A1(n12569), .A2(n12568), .A3(n12567), .ZN(n18209) );
  AOI211_X1 U12153 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n12566), .B(n12565), .ZN(n12567) );
  NOR2_X1 U12154 ( .A1(n12591), .A2(n12590), .ZN(n18218) );
  INV_X1 U12155 ( .A(n15651), .ZN(n15653) );
  INV_X1 U12156 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14096) );
  NAND2_X1 U12157 ( .A1(n20009), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19996) );
  INV_X1 U12158 ( .A(n15977), .ZN(n19959) );
  INV_X1 U12159 ( .A(n19932), .ZN(n19964) );
  INV_X1 U12160 ( .A(n19996), .ZN(n20014) );
  AND2_X1 U12161 ( .A1(n13919), .A2(n13915), .ZN(n20006) );
  INV_X1 U12162 ( .A(n19980), .ZN(n20005) );
  AND2_X1 U12163 ( .A1(n13907), .A2(n15977), .ZN(n20017) );
  NAND2_X1 U12164 ( .A1(n9919), .A2(n9918), .ZN(n14818) );
  INV_X1 U12165 ( .A(n14629), .ZN(n20021) );
  AND2_X2 U12166 ( .A1(n12892), .A2(n13171), .ZN(n20023) );
  OAI211_X1 U12167 ( .C1(n12384), .C2(n12888), .A(n13273), .B(n13268), .ZN(
        n12392) );
  INV_X1 U12168 ( .A(n14690), .ZN(n16024) );
  NAND2_X1 U12169 ( .A1(n14695), .A2(n13547), .ZN(n14690) );
  INV_X1 U12170 ( .A(n16029), .ZN(n14692) );
  AND2_X1 U12171 ( .A1(n13548), .A2(n13564), .ZN(n16025) );
  NOR2_X2 U12172 ( .A1(n16024), .A2(n13548), .ZN(n14705) );
  INV_X1 U12173 ( .A(n20035), .ZN(n20045) );
  NOR2_X1 U12174 ( .A1(n13388), .A2(n11022), .ZN(n20054) );
  INV_X2 U12175 ( .A(n20054), .ZN(n13418) );
  XNOR2_X1 U12176 ( .A(n12112), .B(n12111), .ZN(n13916) );
  OR2_X1 U12177 ( .A1(n12110), .A2(n14713), .ZN(n12112) );
  AOI21_X1 U12178 ( .B1(n14547), .B2(n14545), .A(n14546), .ZN(n14724) );
  INV_X1 U12179 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20907) );
  AOI21_X1 U12180 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n16079) );
  CLKBUF_X1 U12181 ( .A(n14080), .Z(n14081) );
  INV_X1 U12182 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20950) );
  AND2_X1 U12183 ( .A1(n16227), .A2(n20538), .ZN(n20062) );
  INV_X1 U12184 ( .A(n20062), .ZN(n20076) );
  OR2_X1 U12185 ( .A1(n20071), .A2(n12108), .ZN(n14803) );
  INV_X1 U12186 ( .A(n20071), .ZN(n19906) );
  XNOR2_X1 U12187 ( .A(n9933), .B(n14820), .ZN(n14835) );
  NAND2_X1 U12188 ( .A1(n9935), .A2(n9934), .ZN(n9933) );
  OAI21_X1 U12189 ( .B1(n14708), .B2(n11604), .A(n9749), .ZN(n9934) );
  NAND2_X1 U12190 ( .A1(n14710), .A2(n16056), .ZN(n9935) );
  AOI21_X1 U12191 ( .B1(n16201), .B2(n16109), .A(n16106), .ZN(n14863) );
  NAND2_X1 U12192 ( .A1(n10035), .A2(n10036), .ZN(n14152) );
  AND2_X1 U12193 ( .A1(n10037), .A2(n11295), .ZN(n10036) );
  NAND2_X1 U12194 ( .A1(n13763), .A2(n11248), .ZN(n16097) );
  OR2_X1 U12195 ( .A1(n12107), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16209) );
  AND2_X1 U12196 ( .A1(n11521), .A2(n15802), .ZN(n16169) );
  INV_X1 U12197 ( .A(n20530), .ZN(n20538) );
  INV_X1 U12198 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20114) );
  INV_X1 U12199 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13534) );
  OAI21_X1 U12200 ( .B1(n20194), .B2(n20190), .A(n20189), .ZN(n20219) );
  OAI21_X1 U12201 ( .B1(n20282), .B2(n20265), .A(n20494), .ZN(n20285) );
  INV_X1 U12202 ( .A(n20279), .ZN(n20284) );
  AOI22_X1 U12203 ( .A1(n14049), .A2(n14047), .B1(n14042), .B2(n20191), .ZN(
        n14092) );
  OR2_X1 U12204 ( .A1(n20292), .A2(n20402), .ZN(n13989) );
  NOR2_X1 U12205 ( .A1(n20390), .A2(n20262), .ZN(n20345) );
  INV_X1 U12206 ( .A(n20357), .ZN(n20386) );
  INV_X1 U12207 ( .A(n20527), .ZN(n20432) );
  INV_X1 U12208 ( .A(n20545), .ZN(n20447) );
  INV_X1 U12209 ( .A(n20556), .ZN(n20457) );
  INV_X1 U12210 ( .A(n20561), .ZN(n20462) );
  INV_X1 U12211 ( .A(n20567), .ZN(n20467) );
  INV_X1 U12212 ( .A(n20572), .ZN(n20472) );
  INV_X1 U12213 ( .A(n20579), .ZN(n20477) );
  OR2_X1 U12214 ( .A1(n20529), .A2(n20262), .ZN(n20479) );
  OAI211_X1 U12215 ( .C1(n20496), .C2(n20513), .A(n20495), .B(n20494), .ZN(
        n20516) );
  AND2_X1 U12216 ( .A1(n11145), .A2(n13701), .ZN(n20556) );
  AND2_X1 U12217 ( .A1(n11144), .A2(n13701), .ZN(n20567) );
  AND2_X1 U12218 ( .A1(n11016), .A2(n13701), .ZN(n20572) );
  INV_X1 U12219 ( .A(n20543), .ZN(n20583) );
  AND2_X1 U12220 ( .A1(n11008), .A2(n13701), .ZN(n20579) );
  NAND2_X1 U12221 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13537), .ZN(n15792) );
  INV_X1 U12222 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16236) );
  CLKBUF_X1 U12223 ( .A(n12123), .Z(n14934) );
  AOI21_X1 U12224 ( .B1(n9794), .B2(n10647), .A(n10646), .ZN(n10648) );
  AND2_X1 U12225 ( .A1(n10028), .A2(n10027), .ZN(n14975) );
  AND2_X1 U12226 ( .A1(n10034), .A2(n10033), .ZN(n12951) );
  OAI22_X1 U12227 ( .A1(n18900), .A2(n10009), .B1(n10012), .B2(n18886), .ZN(
        n18885) );
  OR2_X1 U12228 ( .A1(n18886), .A2(n15248), .ZN(n10009) );
  OR2_X1 U12229 ( .A1(n14267), .A2(n14266), .ZN(n20698) );
  NAND2_X1 U12230 ( .A1(n14932), .A2(n12825), .ZN(n20697) );
  NAND2_X1 U12231 ( .A1(n10441), .A2(n9937), .ZN(n13791) );
  OR2_X1 U12232 ( .A1(n12335), .A2(n12334), .ZN(n19023) );
  OR2_X1 U12233 ( .A1(n12283), .A2(n12282), .ZN(n13305) );
  AND2_X1 U12234 ( .A1(n13874), .A2(n15651), .ZN(n19061) );
  AND2_X1 U12235 ( .A1(n19095), .A2(n13156), .ZN(n19059) );
  NOR2_X1 U12236 ( .A1(n19106), .A2(n19120), .ZN(n19102) );
  OR2_X1 U12237 ( .A1(n19059), .A2(n13874), .ZN(n19096) );
  NAND2_X1 U12238 ( .A1(n19095), .A2(n13165), .ZN(n19124) );
  INV_X1 U12239 ( .A(n19063), .ZN(n19120) );
  INV_X1 U12240 ( .A(n19124), .ZN(n19106) );
  NAND2_X1 U12241 ( .A1(n13030), .A2(n13029), .ZN(n19154) );
  INV_X1 U12242 ( .A(n14267), .ZN(n13048) );
  NAND2_X1 U12243 ( .A1(n19184), .A2(n13101), .ZN(n19172) );
  OAI211_X1 U12244 ( .C1(n15356), .C2(n15355), .A(n15354), .B(n10117), .ZN(
        n15357) );
  NOR2_X1 U12245 ( .A1(n15143), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10092) );
  NAND2_X1 U12246 ( .A1(n10681), .A2(n10661), .ZN(n15156) );
  INV_X1 U12247 ( .A(n15187), .ZN(n15416) );
  NOR2_X1 U12248 ( .A1(n15113), .A2(n15112), .ZN(n14980) );
  INV_X1 U12249 ( .A(n9866), .ZN(n12194) );
  NAND2_X1 U12250 ( .A1(n15312), .A2(n9809), .ZN(n15612) );
  NAND2_X1 U12251 ( .A1(n13621), .A2(n13620), .ZN(n13665) );
  AND2_X1 U12252 ( .A1(n10065), .A2(n10066), .ZN(n14022) );
  CLKBUF_X1 U12253 ( .A(n14000), .Z(n14001) );
  INV_X1 U12254 ( .A(n19444), .ZN(n19884) );
  XNOR2_X1 U12255 ( .A(n13195), .B(n13194), .ZN(n19877) );
  NOR2_X1 U12256 ( .A1(n13311), .A2(n12242), .ZN(n13649) );
  INV_X1 U12257 ( .A(n19877), .ZN(n19874) );
  XNOR2_X1 U12258 ( .A(n13219), .B(n13196), .ZN(n20708) );
  AND2_X1 U12259 ( .A1(n10234), .A2(n10233), .ZN(n9965) );
  OR2_X1 U12260 ( .A1(n19609), .A2(n19419), .ZN(n19218) );
  OAI21_X1 U12261 ( .B1(n19273), .B2(n19272), .A(n19621), .ZN(n19290) );
  INV_X1 U12262 ( .A(n19308), .ZN(n19324) );
  OAI21_X1 U12263 ( .B1(n19335), .B2(n19334), .A(n19333), .ZN(n19353) );
  AND2_X1 U12264 ( .A1(n19414), .A2(n19616), .ZN(n19387) );
  OAI21_X1 U12265 ( .B1(n19456), .B2(n19455), .A(n19454), .ZN(n19474) );
  NOR2_X2 U12266 ( .A1(n19446), .A2(n19479), .ZN(n19503) );
  INV_X1 U12267 ( .A(n19524), .ZN(n19541) );
  OAI21_X1 U12268 ( .B1(n19546), .B2(n19520), .A(n19519), .ZN(n19540) );
  OR3_X1 U12269 ( .A1(n19551), .A2(n19730), .A3(n19550), .ZN(n19573) );
  INV_X1 U12270 ( .A(n19718), .ZN(n19664) );
  OR3_X1 U12271 ( .A1(n19670), .A2(n19730), .A3(n19669), .ZN(n19715) );
  INV_X1 U12272 ( .A(n19686), .ZN(n19744) );
  NAND2_X1 U12273 ( .A1(n19661), .A2(n19728), .ZN(n19781) );
  OR3_X1 U12274 ( .A1(n19731), .A2(n19730), .A3(n19729), .ZN(n19778) );
  OR2_X1 U12275 ( .A1(n13496), .A2(n13495), .ZN(n16367) );
  NOR2_X1 U12276 ( .A1(n16538), .A2(n12712), .ZN(n16521) );
  NOR2_X1 U12277 ( .A1(n18631), .A2(n17443), .ZN(n18853) );
  OR2_X1 U12278 ( .A1(n18639), .A2(n18692), .ZN(n16522) );
  NOR2_X2 U12279 ( .A1(n18686), .A2(n16544), .ZN(n16871) );
  INV_X1 U12280 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17651) );
  NOR2_X1 U12281 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16809), .ZN(n16801) );
  INV_X1 U12282 ( .A(n16928), .ZN(n16915) );
  INV_X1 U12283 ( .A(n16871), .ZN(n16921) );
  INV_X1 U12284 ( .A(n16889), .ZN(n16905) );
  NAND2_X1 U12285 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16922), .ZN(n16913) );
  INV_X1 U12286 ( .A(n16922), .ZN(n16924) );
  NOR3_X1 U12287 ( .A1(n17119), .A2(n17048), .A3(n14221), .ZN(n17050) );
  NOR2_X1 U12288 ( .A1(n16811), .A2(n17194), .ZN(n17149) );
  NOR2_X1 U12289 ( .A1(n17203), .A2(n17208), .ZN(n17207) );
  INV_X1 U12290 ( .A(n17228), .ZN(n17227) );
  NAND2_X1 U12291 ( .A1(n17263), .A2(n9787), .ZN(n17249) );
  NAND2_X1 U12292 ( .A1(n17263), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17259) );
  NOR2_X1 U12293 ( .A1(n17391), .A2(n17268), .ZN(n17263) );
  NOR2_X1 U12294 ( .A1(n17273), .A2(n17280), .ZN(n17269) );
  NAND2_X1 U12295 ( .A1(n17269), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17268) );
  NOR3_X1 U12296 ( .A1(n17313), .A2(n17279), .A3(n17397), .ZN(n17274) );
  NAND2_X1 U12297 ( .A1(n17274), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17273) );
  NOR2_X1 U12298 ( .A1(n17449), .A2(n17301), .ZN(n17296) );
  NAND2_X1 U12299 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17317), .ZN(n17313) );
  NOR2_X1 U12300 ( .A1(n17492), .A2(n17323), .ZN(n17317) );
  NOR2_X1 U12301 ( .A1(n12426), .A2(n12425), .ZN(n17353) );
  NOR2_X1 U12302 ( .A1(n12483), .A2(n12482), .ZN(n17359) );
  AOI21_X1 U12303 ( .B1(n15873), .B2(n15872), .A(n18692), .ZN(n17379) );
  NOR2_X1 U12304 ( .A1(n18664), .A2(n17366), .ZN(n17373) );
  NAND2_X1 U12305 ( .A1(n17381), .A2(n17380), .ZN(n17440) );
  CLKBUF_X1 U12306 ( .A(n17488), .Z(n17483) );
  OR2_X1 U12307 ( .A1(n18687), .A2(n17443), .ZN(n17491) );
  NOR2_X1 U12308 ( .A1(n17596), .A2(n9844), .ZN(n17533) );
  NAND2_X1 U12309 ( .A1(n17697), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17940) );
  NAND2_X1 U12310 ( .A1(n17657), .A2(n17938), .ZN(n17596) );
  INV_X1 U12311 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17665) );
  INV_X1 U12312 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17690) );
  INV_X1 U12313 ( .A(n17765), .ZN(n17784) );
  NAND2_X1 U12314 ( .A1(n17809), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17801) );
  INV_X1 U12315 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17830) );
  INV_X1 U12316 ( .A(n16426), .ZN(n17511) );
  NOR2_X1 U12317 ( .A1(n18661), .A2(n18642), .ZN(n18076) );
  INV_X1 U12318 ( .A(n10059), .ZN(n17851) );
  AND2_X1 U12319 ( .A1(n10059), .A2(n10058), .ZN(n17850) );
  INV_X1 U12320 ( .A(n18642), .ZN(n18665) );
  INV_X1 U12321 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18674) );
  INV_X1 U12322 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18789) );
  AND2_X1 U12323 ( .A1(n12404), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n13565)
         );
  AND2_X1 U12325 ( .A1(n9917), .A2(n9916), .ZN(n14825) );
  NOR2_X1 U12326 ( .A1(n14822), .A2(n9922), .ZN(n9916) );
  NOR2_X1 U12327 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  AND2_X1 U12328 ( .A1(n11531), .A2(n11530), .ZN(n11532) );
  NAND2_X1 U12329 ( .A1(n11399), .A2(n20103), .ZN(n11533) );
  AND2_X1 U12330 ( .A1(n12919), .A2(n12918), .ZN(n12920) );
  AND2_X1 U12331 ( .A1(n9755), .A2(n10004), .ZN(n13558) );
  AOI21_X1 U12332 ( .B1(n12863), .B2(n12862), .A(n12861), .ZN(n12868) );
  NAND2_X1 U12333 ( .A1(n9864), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9863) );
  OAI21_X1 U12334 ( .B1(n12882), .B2(n17875), .A(n12881), .ZN(n12883) );
  OAI21_X1 U12335 ( .B1(n12882), .B2(n18190), .A(n12740), .ZN(n12741) );
  INV_X1 U12336 ( .A(n10945), .ZN(n11006) );
  CLKBUF_X3 U12337 ( .A(n12485), .Z(n17162) );
  NAND2_X1 U12338 ( .A1(n12746), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12747) );
  NAND2_X1 U12339 ( .A1(n14438), .A2(n10121), .ZN(n9774) );
  NAND2_X1 U12340 ( .A1(n10104), .A2(n14207), .ZN(n14206) );
  AND2_X1 U12341 ( .A1(n15936), .A2(n9817), .ZN(n14623) );
  NAND2_X1 U12342 ( .A1(n11405), .A2(n11404), .ZN(n11409) );
  AND2_X1 U12343 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9775) );
  INV_X2 U12344 ( .A(n13659), .ZN(n10032) );
  NOR2_X1 U12345 ( .A1(n10316), .A2(n10320), .ZN(n10493) );
  OR2_X1 U12346 ( .A1(n15113), .A2(n9815), .ZN(n9776) );
  OR2_X1 U12347 ( .A1(n12943), .A2(n12944), .ZN(n9777) );
  AND3_X1 U12348 ( .A1(n10145), .A2(n10144), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9778) );
  INV_X1 U12349 ( .A(n19215), .ZN(n9957) );
  AND2_X1 U12350 ( .A1(n19973), .A2(n19972), .ZN(n9779) );
  AND2_X1 U12351 ( .A1(n9775), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9781) );
  AND2_X1 U12352 ( .A1(n10563), .A2(n9816), .ZN(n9782) );
  NAND2_X1 U12353 ( .A1(n13247), .A2(n13249), .ZN(n13248) );
  NAND2_X1 U12354 ( .A1(n12746), .A2(n10019), .ZN(n12776) );
  NAND2_X1 U12355 ( .A1(n12757), .A2(n9775), .ZN(n12755) );
  AND2_X1 U12356 ( .A1(n15564), .A2(n9992), .ZN(n13752) );
  NAND2_X1 U12357 ( .A1(n12757), .A2(n9825), .ZN(n12751) );
  OR2_X1 U12358 ( .A1(n9964), .A2(n14136), .ZN(n9783) );
  OR2_X1 U12359 ( .A1(n12193), .A2(n9838), .ZN(n9784) );
  OR3_X1 U12360 ( .A1(n12944), .A2(n14955), .A3(n12817), .ZN(n9785) );
  NAND2_X1 U12361 ( .A1(n9901), .A2(n9903), .ZN(n9786) );
  AND2_X1 U12362 ( .A1(n9893), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9787) );
  AND2_X2 U12363 ( .A1(n12217), .A2(n19668), .ZN(n12218) );
  OR2_X1 U12364 ( .A1(n14618), .A2(n9910), .ZN(n9788) );
  OR2_X1 U12365 ( .A1(n9750), .A2(n16193), .ZN(n9789) );
  OR2_X1 U12366 ( .A1(n12522), .A2(n12521), .ZN(n9790) );
  OR2_X1 U12367 ( .A1(n9909), .A2(n9908), .ZN(n9792) );
  OR2_X1 U12368 ( .A1(n12417), .A2(n12418), .ZN(n9793) );
  OR2_X1 U12369 ( .A1(n10645), .A2(n10644), .ZN(n9794) );
  NAND2_X1 U12370 ( .A1(n10078), .A2(n10077), .ZN(n15154) );
  AND2_X1 U12371 ( .A1(n10590), .A2(n9942), .ZN(n10617) );
  NAND2_X1 U12372 ( .A1(n12167), .A2(n12850), .ZN(n15239) );
  NAND2_X1 U12373 ( .A1(n10590), .A2(n9943), .ZN(n10609) );
  NOR2_X1 U12374 ( .A1(n15190), .A2(n15430), .ZN(n15173) );
  NOR2_X1 U12375 ( .A1(n15190), .A2(n10068), .ZN(n15162) );
  INV_X1 U12376 ( .A(n10050), .ZN(n16536) );
  NAND2_X1 U12377 ( .A1(n9801), .A2(n9894), .ZN(n10050) );
  AND2_X1 U12378 ( .A1(n17263), .A2(n9893), .ZN(n9796) );
  NOR2_X1 U12379 ( .A1(n12419), .A2(n12415), .ZN(n12477) );
  INV_X1 U12380 ( .A(n12477), .ZN(n15706) );
  NAND2_X1 U12381 ( .A1(n17695), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12724) );
  AND2_X1 U12382 ( .A1(n10133), .A2(n10132), .ZN(n9797) );
  INV_X1 U12383 ( .A(n12511), .ZN(n12496) );
  NAND2_X1 U12384 ( .A1(n9747), .A2(n10222), .ZN(n10221) );
  OR2_X1 U12385 ( .A1(n12511), .A2(n18799), .ZN(n9798) );
  OR2_X1 U12386 ( .A1(n14723), .A2(n16186), .ZN(n9799) );
  AND2_X1 U12387 ( .A1(n10862), .A2(n10560), .ZN(n10857) );
  AOI211_X1 U12388 ( .C1(n18206), .C2(n12714), .A(n16537), .B(n16538), .ZN(
        n12720) );
  AND4_X1 U12389 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n9800) );
  NOR2_X1 U12390 ( .A1(n14949), .A2(n14948), .ZN(n12792) );
  AND2_X1 U12391 ( .A1(n12720), .A2(n18649), .ZN(n9801) );
  OR3_X1 U12392 ( .A1(n14618), .A2(n9913), .A3(n9915), .ZN(n9802) );
  INV_X1 U12393 ( .A(n15179), .ZN(n10079) );
  NAND2_X1 U12394 ( .A1(n15936), .A2(n11883), .ZN(n9803) );
  NAND2_X1 U12395 ( .A1(n15339), .A2(n10867), .ZN(n16336) );
  AND2_X1 U12396 ( .A1(n13475), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U12397 ( .A1(n10304), .A2(n10306), .ZN(n19513) );
  AND2_X1 U12398 ( .A1(n10146), .A2(n10143), .ZN(n9805) );
  AND2_X1 U12399 ( .A1(n10141), .A2(n10139), .ZN(n9806) );
  AND3_X1 U12400 ( .A1(n10037), .A2(n11295), .A3(n9789), .ZN(n9807) );
  INV_X1 U12401 ( .A(n14080), .ZN(n10104) );
  INV_X1 U12402 ( .A(n14253), .ZN(n15286) );
  NOR2_X1 U12403 ( .A1(n9780), .A2(n15529), .ZN(n14253) );
  AND2_X1 U12404 ( .A1(n10395), .A2(n13798), .ZN(n9808) );
  NAND2_X1 U12405 ( .A1(n10556), .A2(n10555), .ZN(n10854) );
  INV_X1 U12406 ( .A(n10854), .ZN(n10557) );
  INV_X2 U12407 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10334) );
  INV_X1 U12408 ( .A(n9990), .ZN(n14954) );
  NOR3_X1 U12409 ( .A1(n12943), .A2(n12944), .A3(n14955), .ZN(n9990) );
  NAND2_X1 U12410 ( .A1(n10615), .A2(n10614), .ZN(n10605) );
  OR2_X1 U12411 ( .A1(n12167), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9809) );
  NOR2_X1 U12412 ( .A1(n14278), .A2(n15382), .ZN(n15138) );
  INV_X1 U12413 ( .A(n15312), .ZN(n9892) );
  NAND2_X1 U12414 ( .A1(n12167), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15312) );
  INV_X1 U12415 ( .A(n10633), .ZN(n10087) );
  OR2_X1 U12416 ( .A1(n13793), .A2(n19008), .ZN(n10317) );
  INV_X1 U12417 ( .A(n10317), .ZN(n10072) );
  INV_X1 U12418 ( .A(n9868), .ZN(n10119) );
  NAND2_X1 U12419 ( .A1(n14253), .A2(n12199), .ZN(n9868) );
  OR2_X1 U12420 ( .A1(n10243), .A2(n12217), .ZN(n9811) );
  AND2_X1 U12421 ( .A1(n14740), .A2(n9926), .ZN(n9812) );
  AND2_X1 U12422 ( .A1(n14513), .A2(n14512), .ZN(n9813) );
  INV_X1 U12423 ( .A(n9953), .ZN(n10566) );
  AND2_X1 U12424 ( .A1(n10855), .A2(n10852), .ZN(n9814) );
  INV_X1 U12425 ( .A(n13909), .ZN(n14514) );
  NAND2_X1 U12426 ( .A1(n12223), .A2(n12229), .ZN(n12810) );
  NOR2_X1 U12427 ( .A1(n17648), .A2(n17603), .ZN(n17563) );
  AND2_X1 U12428 ( .A1(n12215), .A2(n9761), .ZN(n12236) );
  AND2_X2 U12429 ( .A1(n13530), .A2(n13503), .ZN(n11126) );
  BUF_X1 U12430 ( .A(n11126), .Z(n11050) );
  AND2_X1 U12431 ( .A1(n12529), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16384) );
  AND2_X1 U12432 ( .A1(n12749), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12746) );
  AND2_X1 U12433 ( .A1(n12757), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12754) );
  NAND2_X1 U12434 ( .A1(n9717), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15339) );
  NAND2_X1 U12435 ( .A1(n9712), .A2(n10563), .ZN(n15340) );
  NOR2_X1 U12436 ( .A1(n14080), .A2(n10105), .ZN(n14168) );
  OR3_X1 U12437 ( .A1(n9982), .A2(n15112), .A3(n9981), .ZN(n9815) );
  AND2_X1 U12438 ( .A1(n16332), .A2(n16330), .ZN(n9816) );
  NOR3_X1 U12439 ( .A1(n15113), .A2(n9982), .A3(n15112), .ZN(n12953) );
  AND2_X1 U12440 ( .A1(n13550), .A2(n13551), .ZN(n13549) );
  NOR2_X1 U12441 ( .A1(n12759), .A2(n10829), .ZN(n12758) );
  NOR2_X1 U12442 ( .A1(n13819), .A2(n13820), .ZN(n13821) );
  AND2_X1 U12443 ( .A1(n12748), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12749) );
  AND2_X1 U12444 ( .A1(n12757), .A2(n9781), .ZN(n12752) );
  NOR2_X1 U12445 ( .A1(n12751), .A2(n12766), .ZN(n12748) );
  NOR2_X1 U12446 ( .A1(n11016), .A2(n20525), .ZN(n11763) );
  INV_X1 U12447 ( .A(n11763), .ZN(n10100) );
  AND2_X1 U12448 ( .A1(n11903), .A2(n11883), .ZN(n9817) );
  NAND2_X1 U12449 ( .A1(n11285), .A2(n16089), .ZN(n14112) );
  NAND2_X1 U12450 ( .A1(n13881), .A2(n9859), .ZN(n13994) );
  AND2_X1 U12451 ( .A1(n9749), .A2(n16164), .ZN(n9818) );
  NOR2_X1 U12452 ( .A1(n9961), .A2(n9960), .ZN(n14962) );
  AND2_X1 U12453 ( .A1(n15587), .A2(n15588), .ZN(n15564) );
  AND2_X1 U12454 ( .A1(n15096), .A2(n15097), .ZN(n14966) );
  INV_X1 U12455 ( .A(n9905), .ZN(n9909) );
  NOR3_X1 U12456 ( .A1(n15959), .A2(n11488), .A3(n9823), .ZN(n9905) );
  AND2_X1 U12457 ( .A1(n10439), .A2(n10440), .ZN(n10512) );
  AND2_X1 U12458 ( .A1(n13821), .A2(n15512), .ZN(n14132) );
  XNOR2_X1 U12459 ( .A(n14420), .B(n14422), .ZN(n15021) );
  OR2_X1 U12460 ( .A1(n14137), .A2(n9783), .ZN(n9819) );
  INV_X1 U12461 ( .A(n10028), .ZN(n14974) );
  NAND2_X1 U12462 ( .A1(n10024), .A2(n10025), .ZN(n16257) );
  NAND2_X1 U12463 ( .A1(n13880), .A2(n14006), .ZN(n13881) );
  AND2_X1 U12464 ( .A1(n13728), .A2(n13729), .ZN(n9820) );
  NOR3_X1 U12465 ( .A1(n15113), .A2(n9815), .A3(n15452), .ZN(n15096) );
  AND2_X1 U12466 ( .A1(n10428), .A2(n10597), .ZN(n9821) );
  AND2_X1 U12467 ( .A1(n14208), .A2(n9904), .ZN(n9822) );
  OR2_X1 U12468 ( .A1(n11477), .A2(n9906), .ZN(n9823) );
  INV_X1 U12469 ( .A(n9907), .ZN(n15950) );
  NOR2_X1 U12470 ( .A1(n15959), .A2(n11477), .ZN(n9907) );
  AND2_X1 U12471 ( .A1(n10004), .A2(n13557), .ZN(n9824) );
  AND2_X1 U12472 ( .A1(n9781), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9825) );
  INV_X1 U12473 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15323) );
  NAND2_X1 U12474 ( .A1(n12956), .A2(n12957), .ZN(n12955) );
  AND2_X1 U12475 ( .A1(n15049), .A2(n14986), .ZN(n12956) );
  AND2_X1 U12476 ( .A1(n9988), .A2(n15600), .ZN(n9826) );
  AND2_X1 U12477 ( .A1(n9970), .A2(n9969), .ZN(n9827) );
  AND2_X1 U12478 ( .A1(n10019), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9828) );
  AND2_X1 U12479 ( .A1(n14624), .A2(n9817), .ZN(n9829) );
  AND2_X1 U12480 ( .A1(n10106), .A2(n14588), .ZN(n9830) );
  INV_X1 U12481 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12760) );
  OAI22_X1 U12482 ( .A1(n12745), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16380), 
        .B2(n12744), .ZN(n13659) );
  NAND2_X1 U12483 ( .A1(n20525), .A2(n20321), .ZN(n13901) );
  INV_X1 U12484 ( .A(n10861), .ZN(n10687) );
  NOR2_X1 U12485 ( .A1(n16220), .A2(n16219), .ZN(n9831) );
  NAND2_X1 U12486 ( .A1(n13245), .A2(n13244), .ZN(n13556) );
  NAND2_X1 U12487 ( .A1(n9755), .A2(n13555), .ZN(n13720) );
  NAND2_X1 U12488 ( .A1(n9986), .A2(n9987), .ZN(n13650) );
  NOR2_X1 U12489 ( .A1(n12778), .A2(n10833), .ZN(n12779) );
  NAND2_X1 U12490 ( .A1(n13556), .A2(n9824), .ZN(n13858) );
  AND2_X1 U12491 ( .A1(n12746), .A2(n10020), .ZN(n9832) );
  NAND2_X1 U12492 ( .A1(n13247), .A2(n9973), .ZN(n13261) );
  AND2_X1 U12493 ( .A1(n13621), .A2(n9988), .ZN(n13664) );
  NAND2_X1 U12494 ( .A1(n15564), .A2(n15565), .ZN(n13751) );
  AND2_X1 U12495 ( .A1(n12746), .A2(n9828), .ZN(n12777) );
  AND2_X1 U12496 ( .A1(n9959), .A2(n12957), .ZN(n9833) );
  AND2_X1 U12497 ( .A1(n13656), .A2(n9827), .ZN(n13550) );
  AND2_X1 U12498 ( .A1(n13678), .A2(n13679), .ZN(n13247) );
  NAND2_X1 U12499 ( .A1(n13656), .A2(n13307), .ZN(n13306) );
  NAND2_X1 U12500 ( .A1(n13656), .A2(n9970), .ZN(n13722) );
  NAND2_X1 U12501 ( .A1(n15564), .A2(n9991), .ZN(n13819) );
  NAND2_X1 U12502 ( .A1(n11521), .A2(n11503), .ZN(n16210) );
  INV_X1 U12503 ( .A(n16210), .ZN(n20098) );
  INV_X1 U12504 ( .A(n10591), .ZN(n9945) );
  AND2_X1 U12505 ( .A1(n10013), .A2(n10012), .ZN(n9834) );
  XNOR2_X1 U12506 ( .A(n9924), .B(n11101), .ZN(n13605) );
  AND2_X1 U12507 ( .A1(n10725), .A2(n10126), .ZN(n13678) );
  NOR2_X1 U12508 ( .A1(n10032), .A2(n18885), .ZN(n14982) );
  INV_X1 U12509 ( .A(n10034), .ZN(n12950) );
  NAND2_X1 U12510 ( .A1(n10030), .A2(n10031), .ZN(n15784) );
  AND2_X1 U12511 ( .A1(n13247), .A2(n9971), .ZN(n13296) );
  NAND2_X1 U12512 ( .A1(n10764), .A2(n10763), .ZN(n13823) );
  AND2_X1 U12513 ( .A1(n9833), .A2(n9958), .ZN(n9835) );
  OR2_X1 U12514 ( .A1(n10007), .A2(n10005), .ZN(n9836) );
  OR2_X1 U12515 ( .A1(n19172), .A2(n16321), .ZN(n9837) );
  NOR2_X1 U12516 ( .A1(n15626), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9838) );
  AND2_X1 U12517 ( .A1(n10063), .A2(n9790), .ZN(n9839) );
  AND2_X1 U12518 ( .A1(n9986), .A2(n9984), .ZN(n9840) );
  INV_X1 U12519 ( .A(n16417), .ZN(n10049) );
  NOR2_X1 U12520 ( .A1(n11588), .A2(n12941), .ZN(n11589) );
  NOR3_X1 U12521 ( .A1(n11588), .A2(n12941), .A3(n10018), .ZN(n12786) );
  NAND2_X1 U12522 ( .A1(n9902), .A2(n9901), .ZN(n19976) );
  INV_X1 U12523 ( .A(n19976), .ZN(n9900) );
  AND2_X1 U12524 ( .A1(n18798), .A2(n17770), .ZN(n9841) );
  OR3_X1 U12525 ( .A1(n11588), .A2(n10017), .A3(n12941), .ZN(n9842) );
  AND2_X1 U12526 ( .A1(n10060), .A2(n9798), .ZN(n9843) );
  INV_X1 U12527 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10018) );
  CLKBUF_X3 U12528 ( .A(n11400), .Z(n11553) );
  INV_X1 U12529 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13437) );
  OR2_X1 U12530 ( .A1(n17876), .A2(n17942), .ZN(n9844) );
  OR2_X1 U12531 ( .A1(n11535), .A2(n11583), .ZN(n9845) );
  OR2_X1 U12532 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9846) );
  INV_X1 U12533 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10095) );
  NAND2_X2 U12534 ( .A1(n18851), .A2(n18840), .ZN(n18184) );
  OAI22_X2 U12535 ( .A1(n20807), .A2(n19223), .B1(n19222), .B2(n19221), .ZN(
        n19776) );
  INV_X1 U12536 ( .A(n19213), .ZN(n19221) );
  AOI22_X2 U12537 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19213), .ZN(n19741) );
  AOI22_X2 U12538 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19213), .ZN(n19771) );
  AOI22_X2 U12539 ( .A1(DATAI_19_), .A2(n13699), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n13700), .ZN(n20560) );
  AOI22_X2 U12540 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13700), .B1(DATAI_17_), 
        .B2(n13699), .ZN(n20549) );
  AOI22_X2 U12541 ( .A1(DATAI_21_), .A2(n13699), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13700), .ZN(n20571) );
  AOI22_X2 U12542 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13700), .B1(DATAI_30_), 
        .B2(n13699), .ZN(n20476) );
  AOI22_X2 U12543 ( .A1(DATAI_31_), .A2(n13699), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n13700), .ZN(n20486) );
  AOI22_X2 U12544 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19213), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19214), .ZN(n19753) );
  NOR2_X2 U12545 ( .A1(n15653), .A2(n15652), .ZN(n19214) );
  NOR2_X2 U12546 ( .A1(n15651), .A2(n15652), .ZN(n19213) );
  INV_X1 U12547 ( .A(n19782), .ZN(n9847) );
  INV_X1 U12548 ( .A(n9847), .ZN(n9848) );
  INV_X1 U12549 ( .A(n20588), .ZN(n9849) );
  INV_X1 U12550 ( .A(n9849), .ZN(n9850) );
  INV_X1 U12551 ( .A(n20577), .ZN(n9851) );
  INV_X1 U12552 ( .A(n9851), .ZN(n9852) );
  INV_X1 U12553 ( .A(n20471), .ZN(n9853) );
  INV_X1 U12554 ( .A(n9853), .ZN(n9854) );
  INV_X1 U12555 ( .A(n20461), .ZN(n9855) );
  INV_X1 U12556 ( .A(n9855), .ZN(n9856) );
  INV_X1 U12557 ( .A(n20451), .ZN(n9857) );
  INV_X1 U12558 ( .A(n9857), .ZN(n9858) );
  AOI22_X2 U12559 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n13700), .B1(DATAI_20_), 
        .B2(n13699), .ZN(n20566) );
  AOI22_X2 U12560 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13700), .B1(DATAI_26_), 
        .B2(n13699), .ZN(n20456) );
  OAI22_X2 U12561 ( .A1(n16453), .A2(n19223), .B1(n15118), .B2(n19221), .ZN(
        n19750) );
  INV_X1 U12562 ( .A(n19214), .ZN(n19223) );
  AOI22_X2 U12563 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19213), .ZN(n19747) );
  AOI22_X2 U12564 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13700), .B1(DATAI_24_), 
        .B2(n13699), .ZN(n20544) );
  XNOR2_X2 U12565 ( .A(n9880), .B(n10850), .ZN(n9861) );
  NAND3_X1 U12566 ( .A1(n16319), .A2(n16320), .A3(n9837), .ZN(P2_U2992) );
  NAND3_X1 U12567 ( .A1(n10066), .A2(n10065), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14021) );
  NAND3_X1 U12568 ( .A1(n10220), .A2(n10234), .A3(n10219), .ZN(n9876) );
  NAND3_X1 U12569 ( .A1(n14255), .A2(n14256), .A3(n9863), .ZN(P2_U3030) );
  INV_X2 U12570 ( .A(n10222), .ZN(n10216) );
  NAND2_X2 U12571 ( .A1(n9870), .A2(n9869), .ZN(n10222) );
  OAI211_X2 U12572 ( .C1(n12369), .C2(n12129), .A(n9875), .B(n9874), .ZN(
        n10291) );
  NAND3_X1 U12573 ( .A1(n10206), .A2(n10205), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9875) );
  NAND2_X1 U12574 ( .A1(n9876), .A2(n13475), .ZN(n12184) );
  OAI21_X1 U12575 ( .B1(n9878), .B2(n15551), .A(n15537), .ZN(n15293) );
  XNOR2_X1 U12576 ( .A(n9878), .B(n15551), .ZN(n15559) );
  OAI21_X1 U12577 ( .B1(n15584), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n9878), .ZN(n15577) );
  INV_X2 U12578 ( .A(n19480), .ZN(n10489) );
  XNOR2_X2 U12579 ( .A(n10721), .B(n10720), .ZN(n13207) );
  NAND2_X1 U12580 ( .A1(n9880), .A2(n9808), .ZN(n9879) );
  OR2_X2 U12581 ( .A1(n10475), .A2(n10476), .ZN(n9880) );
  INV_X1 U12582 ( .A(n10856), .ZN(n10853) );
  NAND2_X1 U12583 ( .A1(n9814), .A2(n10856), .ZN(n10065) );
  NAND2_X2 U12584 ( .A1(n9882), .A2(n9881), .ZN(n10856) );
  INV_X1 U12585 ( .A(n13994), .ZN(n9882) );
  NAND2_X1 U12586 ( .A1(n9883), .A2(n9884), .ZN(n10272) );
  INV_X1 U12587 ( .A(n10258), .ZN(n9883) );
  INV_X1 U12588 ( .A(n10257), .ZN(n9884) );
  OAI21_X1 U12589 ( .B1(n9887), .B2(n15338), .A(n9885), .ZN(n16337) );
  NAND2_X1 U12590 ( .A1(n12383), .A2(n9888), .ZN(P2_U3029) );
  INV_X1 U12591 ( .A(n10851), .ZN(n9890) );
  INV_X1 U12592 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9891) );
  NAND3_X1 U12593 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n9897) );
  INV_X2 U12594 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18821) );
  INV_X1 U12595 ( .A(n11409), .ZN(n9903) );
  NAND3_X1 U12596 ( .A1(n9919), .A2(n9918), .A3(n20098), .ZN(n9917) );
  INV_X1 U12597 ( .A(n14515), .ZN(n9923) );
  NAND2_X1 U12598 ( .A1(n11117), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9925) );
  NOR2_X2 U12599 ( .A1(n9926), .A2(n11584), .ZN(n14732) );
  NAND2_X1 U12600 ( .A1(n11212), .A2(n9936), .ZN(n11264) );
  INV_X1 U12601 ( .A(n11264), .ZN(n11262) );
  NAND3_X1 U12602 ( .A1(n11277), .A2(n11660), .A3(n11313), .ZN(n11270) );
  OAI211_X2 U12603 ( .C1(n9941), .C2(n9940), .A(n10661), .B(n10681), .ZN(
        n11597) );
  NOR2_X1 U12604 ( .A1(n10653), .A2(n10079), .ZN(n9941) );
  OAI21_X2 U12605 ( .B1(n11597), .B2(n15164), .A(n11596), .ZN(n15140) );
  NAND2_X1 U12606 ( .A1(n10512), .A2(n10511), .ZN(n10514) );
  NAND2_X1 U12607 ( .A1(n10512), .A2(n9954), .ZN(n9953) );
  INV_X1 U12608 ( .A(n10511), .ZN(n9955) );
  NAND2_X1 U12609 ( .A1(n10667), .A2(n9956), .ZN(n10665) );
  INV_X1 U12610 ( .A(n10662), .ZN(n10695) );
  NOR2_X2 U12611 ( .A1(n10640), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10642) );
  INV_X2 U12612 ( .A(n12214), .ZN(n10428) );
  AND2_X4 U12613 ( .A1(n10326), .A2(n13444), .ZN(n10328) );
  INV_X1 U12614 ( .A(n9961), .ZN(n15037) );
  INV_X1 U12615 ( .A(n14963), .ZN(n9960) );
  NAND2_X1 U12616 ( .A1(n9965), .A2(n13094), .ZN(n13481) );
  AND2_X1 U12617 ( .A1(n9974), .A2(n10218), .ZN(n12223) );
  NAND3_X1 U12618 ( .A1(n10203), .A2(n10200), .A3(n10202), .ZN(n9977) );
  NAND3_X1 U12619 ( .A1(n10199), .A2(n10196), .A3(n10198), .ZN(n9980) );
  NAND3_X1 U12620 ( .A1(n9986), .A2(n9984), .A3(n14008), .ZN(n14007) );
  NAND2_X2 U12621 ( .A1(n14027), .A2(n10110), .ZN(n13621) );
  NOR2_X2 U12622 ( .A1(n12943), .A2(n9785), .ZN(n12911) );
  NAND2_X1 U12623 ( .A1(n13214), .A2(n13213), .ZN(n9996) );
  NAND2_X1 U12624 ( .A1(n13214), .A2(n9994), .ZN(n13217) );
  NAND2_X1 U12625 ( .A1(n9996), .A2(n13216), .ZN(n13243) );
  INV_X1 U12626 ( .A(n15013), .ZN(n10001) );
  NOR2_X1 U12627 ( .A1(n10002), .A2(n14459), .ZN(n15010) );
  INV_X1 U12628 ( .A(n10002), .ZN(n10000) );
  INV_X1 U12629 ( .A(n14456), .ZN(n10003) );
  INV_X1 U12630 ( .A(n10013), .ZN(n14125) );
  NOR2_X2 U12631 ( .A1(n10032), .A2(n12771), .ZN(n18900) );
  NAND2_X1 U12632 ( .A1(n10016), .A2(n10015), .ZN(n10014) );
  INV_X1 U12633 ( .A(n10017), .ZN(n10016) );
  NAND2_X2 U12636 ( .A1(n10035), .A2(n9807), .ZN(n14809) );
  NAND3_X1 U12637 ( .A1(n13765), .A2(n11271), .A3(n13764), .ZN(n10044) );
  XNOR2_X2 U12638 ( .A(n11150), .B(n11151), .ZN(n11622) );
  AND2_X2 U12639 ( .A1(n17863), .A2(n10049), .ZN(n17781) );
  NOR2_X2 U12640 ( .A1(n16522), .A2(n18206), .ZN(n17863) );
  NOR2_X2 U12641 ( .A1(n12420), .A2(n18657), .ZN(n12464) );
  NAND4_X1 U12642 ( .A1(n17769), .A2(n12530), .A3(n18020), .A4(n17755), .ZN(
        n10051) );
  NOR2_X2 U12643 ( .A1(n12419), .A2(n12416), .ZN(n17159) );
  INV_X2 U12644 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12634) );
  NOR2_X2 U12645 ( .A1(n12542), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16426) );
  NOR2_X2 U12646 ( .A1(n17523), .A2(n12541), .ZN(n12542) );
  AOI21_X2 U12647 ( .B1(n10056), .B2(n10055), .A(n10053), .ZN(n12546) );
  NAND3_X1 U12648 ( .A1(n12545), .A2(n15835), .A3(n10057), .ZN(n10056) );
  NAND2_X1 U12649 ( .A1(n10060), .A2(n9798), .ZN(n10058) );
  OR2_X2 U12650 ( .A1(n17860), .A2(n17868), .ZN(n10060) );
  AOI21_X2 U12651 ( .B1(n10059), .B2(n10058), .A(n12514), .ZN(n17841) );
  INV_X1 U12652 ( .A(n10060), .ZN(n17858) );
  INV_X1 U12653 ( .A(n17800), .ZN(n10062) );
  OAI22_X2 U12654 ( .A1(n17814), .A2(n10061), .B1(n9790), .B2(n17800), .ZN(
        n17799) );
  INV_X1 U12655 ( .A(n10063), .ZN(n17813) );
  NOR2_X2 U12656 ( .A1(n17799), .A2(n12525), .ZN(n12527) );
  NAND2_X1 U12657 ( .A1(n10064), .A2(n10853), .ZN(n10066) );
  NOR2_X2 U12658 ( .A1(n15190), .A2(n10067), .ZN(n15152) );
  NAND2_X1 U12659 ( .A1(n10074), .A2(n10245), .ZN(n10073) );
  NAND2_X1 U12660 ( .A1(n12223), .A2(n10222), .ZN(n10074) );
  NAND2_X1 U12661 ( .A1(n15179), .A2(n10076), .ZN(n10075) );
  NAND2_X1 U12662 ( .A1(n15175), .A2(n10653), .ZN(n10077) );
  AOI21_X1 U12663 ( .B1(n10653), .B2(n10654), .A(n10079), .ZN(n10078) );
  NAND2_X1 U12664 ( .A1(n10087), .A2(n15465), .ZN(n10083) );
  INV_X1 U12665 ( .A(n15204), .ZN(n10088) );
  OR2_X1 U12666 ( .A1(n15143), .A2(n10089), .ZN(n10091) );
  INV_X1 U12667 ( .A(n11596), .ZN(n10090) );
  OAI21_X1 U12668 ( .B1(n10678), .B2(n10092), .A(n10094), .ZN(n14275) );
  NAND3_X1 U12669 ( .A1(n10093), .A2(n14274), .A3(n10091), .ZN(n15125) );
  NAND2_X1 U12670 ( .A1(n10678), .A2(n10094), .ZN(n10093) );
  AND3_X2 U12671 ( .A1(n10129), .A2(n13437), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10152) );
  NAND3_X1 U12672 ( .A1(n13728), .A2(n13729), .A3(n13845), .ZN(n13780) );
  INV_X1 U12673 ( .A(n11615), .ZN(n11110) );
  NAND2_X1 U12674 ( .A1(n11098), .A2(n11111), .ZN(n11615) );
  NAND2_X1 U12675 ( .A1(n11078), .A2(n10096), .ZN(n11111) );
  NAND2_X1 U12676 ( .A1(n11078), .A2(n11077), .ZN(n11097) );
  OAI21_X1 U12677 ( .B1(n11609), .B2(n10101), .A(n10098), .ZN(n13325) );
  INV_X1 U12678 ( .A(n13325), .ZN(n11631) );
  NAND2_X1 U12679 ( .A1(n15936), .A2(n9829), .ZN(n14612) );
  INV_X1 U12680 ( .A(n14612), .ZN(n11951) );
  NAND2_X1 U12681 ( .A1(n14556), .A2(n9830), .ZN(n14545) );
  AND2_X1 U12682 ( .A1(n14556), .A2(n10106), .ZN(n14595) );
  AND2_X1 U12683 ( .A1(n14556), .A2(n11990), .ZN(n14594) );
  INV_X1 U12684 ( .A(n14545), .ZN(n12053) );
  XNOR2_X1 U12685 ( .A(n10698), .B(n10697), .ZN(n12865) );
  AOI21_X1 U12686 ( .B1(n14536), .B2(n14534), .A(n14535), .ZN(n14721) );
  NAND2_X1 U12687 ( .A1(n15021), .A2(n15023), .ZN(n15022) );
  NAND2_X1 U12688 ( .A1(n13281), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13282) );
  NOR2_X2 U12689 ( .A1(n14534), .A2(n14536), .ZN(n14535) );
  NAND2_X1 U12690 ( .A1(n11262), .A2(n11261), .ZN(n11277) );
  NOR2_X1 U12691 ( .A1(n10319), .A2(n10318), .ZN(n10479) );
  AND2_X1 U12692 ( .A1(n10147), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U12693 ( .A1(n12172), .A2(n10204), .ZN(n10205) );
  NOR2_X1 U12694 ( .A1(n10316), .A2(n10318), .ZN(n10488) );
  OR2_X1 U12695 ( .A1(n20117), .A2(n20115), .ZN(n20390) );
  NAND2_X1 U12696 ( .A1(n14715), .A2(n12893), .ZN(n12903) );
  AND2_X2 U12697 ( .A1(n10307), .A2(n10072), .ZN(n19580) );
  NAND2_X1 U12698 ( .A1(n10960), .A2(n13911), .ZN(n10983) );
  NAND2_X1 U12699 ( .A1(n11024), .A2(n10960), .ZN(n11514) );
  AND2_X2 U12700 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10889) );
  INV_X1 U12701 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10880) );
  NAND2_X1 U12702 ( .A1(n12865), .A2(n16359), .ZN(n12866) );
  OAI21_X2 U12703 ( .B1(n10297), .B2(n10300), .A(n9709), .ZN(n13793) );
  AOI22_X1 U12704 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U12705 ( .A1(n11145), .A2(n11015), .ZN(n11040) );
  NAND2_X1 U12706 ( .A1(n11005), .A2(n11144), .ZN(n11015) );
  NAND2_X1 U12707 ( .A1(n11601), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11607) );
  NAND2_X1 U12708 ( .A1(n11237), .A2(n11216), .ZN(n11643) );
  OR2_X1 U12709 ( .A1(n11190), .A2(n13587), .ZN(n11191) );
  INV_X1 U12710 ( .A(n10862), .ZN(n10860) );
  XNOR2_X1 U12711 ( .A(n11608), .B(n14821), .ZN(n14826) );
  INV_X1 U12712 ( .A(n13781), .ZN(n11675) );
  INV_X1 U12713 ( .A(n10291), .ZN(n10263) );
  NAND2_X1 U12714 ( .A1(n14516), .A2(n12393), .ZN(n12409) );
  INV_X1 U12715 ( .A(n10448), .ZN(n10450) );
  AND2_X1 U12716 ( .A1(n9764), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10346) );
  AOI22_X1 U12717 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U12718 ( .A1(n12377), .A2(n12376), .ZN(n15614) );
  INV_X1 U12719 ( .A(n15614), .ZN(n12862) );
  NAND2_X1 U12720 ( .A1(n12392), .A2(n13171), .ZN(n16022) );
  INV_X2 U12721 ( .A(n16022), .ZN(n14695) );
  OR2_X1 U12722 ( .A1(n17770), .A2(n17500), .ZN(n10107) );
  OR2_X1 U12723 ( .A1(n17770), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10108) );
  OR2_X1 U12724 ( .A1(n17770), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10109) );
  CLKBUF_X3 U12725 ( .A(n12572), .Z(n17175) );
  OR2_X1 U12726 ( .A1(n10861), .A2(n12361), .ZN(n10110) );
  AND3_X1 U12727 ( .A1(n10149), .A2(n10148), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10111) );
  OR2_X1 U12728 ( .A1(n14731), .A2(n16186), .ZN(n10112) );
  NOR2_X1 U12729 ( .A1(n15212), .A2(n15236), .ZN(n10113) );
  AND3_X1 U12730 ( .A1(n10154), .A2(n10334), .A3(n10153), .ZN(n10114) );
  AND4_X1 U12731 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10115) );
  INV_X1 U12732 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10449) );
  AND2_X1 U12733 ( .A1(n9763), .A2(n10334), .ZN(n10452) );
  INV_X1 U12734 ( .A(n10335), .ZN(n10413) );
  INV_X1 U12735 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11402) );
  NOR2_X1 U12736 ( .A1(n15465), .A2(n15475), .ZN(n10116) );
  NAND2_X1 U12737 ( .A1(n20023), .A2(n11008), .ZN(n14635) );
  INV_X1 U12738 ( .A(n14635), .ZN(n12893) );
  INV_X1 U12739 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10833) );
  INV_X1 U12740 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11604) );
  INV_X1 U12741 ( .A(n10315), .ZN(n10303) );
  INV_X1 U12742 ( .A(n19173), .ZN(n10876) );
  AND3_X1 U12743 ( .A1(n17771), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10118) );
  OR2_X1 U12744 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18705), .ZN(n18849) );
  INV_X1 U12745 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15975) );
  INV_X1 U12746 ( .A(n15853), .ZN(n11306) );
  OR2_X1 U12747 ( .A1(n13429), .A2(n14352), .ZN(n10120) );
  AND2_X1 U12748 ( .A1(n14437), .A2(n14454), .ZN(n10121) );
  INV_X1 U12749 ( .A(n12226), .ZN(n12801) );
  INV_X1 U12750 ( .A(n12801), .ZN(n12325) );
  NAND2_X1 U12751 ( .A1(n12761), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12759) );
  INV_X1 U12752 ( .A(n11589), .ZN(n12787) );
  INV_X1 U12753 ( .A(n17368), .ZN(n17372) );
  INV_X1 U12754 ( .A(n12218), .ZN(n12800) );
  AND3_X1 U12755 ( .A1(n11038), .A2(n13498), .A3(n11037), .ZN(n10122) );
  AND2_X1 U12756 ( .A1(n19023), .A2(n19022), .ZN(n10123) );
  INV_X1 U12757 ( .A(n18488), .ZN(n18575) );
  OR2_X1 U12758 ( .A1(n15001), .A2(n20705), .ZN(n10125) );
  OR2_X1 U12759 ( .A1(n10724), .A2(n10723), .ZN(n10126) );
  AND2_X1 U12760 ( .A1(n11144), .A2(n11016), .ZN(n10127) );
  AND4_X1 U12761 ( .A1(n10885), .A2(n10884), .A3(n10883), .A4(n10882), .ZN(
        n10128) );
  AOI21_X1 U12762 ( .B1(n11359), .B2(n11382), .A(n11330), .ZN(n11340) );
  NOR2_X1 U12763 ( .A1(n11338), .A2(n11381), .ZN(n11344) );
  OAI21_X1 U12764 ( .B1(n10273), .B2(n12971), .A(n10252), .ZN(n10253) );
  INV_X1 U12765 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11318) );
  NOR2_X1 U12766 ( .A1(n12384), .A2(n11010), .ZN(n11011) );
  INV_X1 U12767 ( .A(n15654), .ZN(n10245) );
  AND2_X1 U12768 ( .A1(n20317), .A2(n9724), .ZN(n11331) );
  AND2_X1 U12769 ( .A1(n11235), .A2(n11234), .ZN(n11236) );
  INV_X1 U12770 ( .A(n12828), .ZN(n10429) );
  NAND2_X1 U12771 ( .A1(n10293), .A2(n10292), .ZN(n10724) );
  OR2_X1 U12772 ( .A1(n9754), .A2(n10444), .ZN(n10278) );
  INV_X1 U12773 ( .A(n13324), .ZN(n11630) );
  INV_X1 U12774 ( .A(n14614), .ZN(n11950) );
  INV_X1 U12775 ( .A(n15937), .ZN(n11883) );
  OR2_X1 U12776 ( .A1(n11139), .A2(n11138), .ZN(n11140) );
  NAND2_X1 U12777 ( .A1(n12385), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11287) );
  OR2_X1 U12778 ( .A1(n11233), .A2(n11232), .ZN(n11266) );
  AOI22_X1 U12779 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11126), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10908) );
  INV_X1 U12780 ( .A(n14421), .ZN(n14422) );
  INV_X1 U12781 ( .A(n15586), .ZN(n10750) );
  NAND2_X1 U12782 ( .A1(n10221), .A2(n15658), .ZN(n12148) );
  OR3_X1 U12783 ( .A1(n10701), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n15870), .ZN(n12138) );
  OR2_X1 U12784 ( .A1(n12653), .A2(n12641), .ZN(n12636) );
  INV_X1 U12785 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11581) );
  NOR2_X2 U12786 ( .A1(n11008), .A2(n20525), .ZN(n11669) );
  INV_X1 U12787 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11534) );
  MUX2_X1 U12788 ( .A(n11389), .B(n11388), .S(n11025), .Z(n11390) );
  AND4_X1 U12789 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n10941) );
  AND2_X1 U12790 ( .A1(n11322), .A2(n11354), .ZN(n11386) );
  OR2_X1 U12791 ( .A1(n10701), .A2(n10700), .ZN(n10703) );
  INV_X1 U12792 ( .A(n14378), .ZN(n14380) );
  INV_X1 U12793 ( .A(n13872), .ZN(n13870) );
  INV_X1 U12794 ( .A(n15124), .ZN(n10690) );
  AND2_X1 U12795 ( .A1(n12852), .A2(n15429), .ZN(n15393) );
  OAI21_X1 U12796 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12634), .A(
        n12636), .ZN(n12644) );
  NOR2_X1 U12797 ( .A1(n12697), .A2(n17803), .ZN(n12700) );
  NAND2_X1 U12798 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12504) );
  INV_X1 U12799 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n20874) );
  NAND2_X1 U12800 ( .A1(n13322), .A2(n11632), .ZN(n13328) );
  NAND2_X1 U12801 ( .A1(n12056), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12110) );
  AND2_X1 U12802 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n11986), .ZN(
        n11987) );
  NAND2_X1 U12803 ( .A1(n11717), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11722) );
  INV_X1 U12804 ( .A(n14778), .ZN(n14879) );
  OAI21_X1 U12805 ( .B1(n11614), .B2(n13335), .A(n11159), .ZN(n11161) );
  NAND2_X1 U12806 ( .A1(n11353), .A2(n11386), .ZN(n11367) );
  NAND2_X1 U12807 ( .A1(n10703), .A2(n10702), .ZN(n12137) );
  INV_X1 U12808 ( .A(n11592), .ZN(n10804) );
  NAND2_X1 U12809 ( .A1(n14966), .A2(n14967), .ZN(n14965) );
  AND2_X1 U12810 ( .A1(n13554), .A2(n13553), .ZN(n13555) );
  NOR2_X1 U12811 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  AND2_X1 U12812 ( .A1(n15393), .A2(n15394), .ZN(n15383) );
  AND2_X1 U12813 ( .A1(n10679), .A2(n15406), .ZN(n15164) );
  INV_X1 U12814 ( .A(n13658), .ZN(n10744) );
  AND2_X1 U12815 ( .A1(n12377), .A2(n12187), .ZN(n14242) );
  AOI21_X1 U12816 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18678), .A(
        n12639), .ZN(n12648) );
  NOR2_X1 U12817 ( .A1(n18657), .A2(n12415), .ZN(n12428) );
  INV_X1 U12818 ( .A(n12878), .ZN(n12879) );
  INV_X1 U12819 ( .A(n17709), .ZN(n12870) );
  NOR2_X1 U12820 ( .A1(n17661), .A2(n17645), .ZN(n17602) );
  NAND2_X1 U12821 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17789), .ZN(
        n12703) );
  NOR2_X1 U12822 ( .A1(n12693), .A2(n17810), .ZN(n12695) );
  NOR2_X1 U12823 ( .A1(n11020), .A2(n11022), .ZN(n13114) );
  INV_X1 U12824 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15966) );
  INV_X1 U12825 ( .A(n20006), .ZN(n19984) );
  NAND2_X1 U12826 ( .A1(n13919), .A2(n13918), .ZN(n19980) );
  NAND2_X1 U12827 ( .A1(n20009), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13912) );
  INV_X1 U12828 ( .A(n11022), .ZN(n13335) );
  AND2_X1 U12829 ( .A1(n11801), .A2(n14170), .ZN(n14169) );
  NOR2_X1 U12830 ( .A1(n11722), .A2(n14096), .ZN(n11723) );
  AOI21_X1 U12831 ( .B1(n11605), .B2(n11604), .A(n11603), .ZN(n11606) );
  NAND2_X1 U12832 ( .A1(n11521), .A2(n13509), .ZN(n16172) );
  AND2_X1 U12833 ( .A1(n20226), .A2(n20252), .ZN(n20231) );
  OR2_X1 U12834 ( .A1(n20292), .A2(n20324), .ZN(n14043) );
  OR2_X1 U12835 ( .A1(n20292), .A2(n20487), .ZN(n14089) );
  AOI221_X1 U12836 ( .B1(n20680), .B2(n15792), .C1(n16229), .C2(n15792), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n13953) );
  NOR2_X1 U12837 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20389) );
  INV_X1 U12838 ( .A(n20550), .ZN(n20452) );
  INV_X1 U12839 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20524) );
  AND2_X1 U12840 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13953), .ZN(n13701) );
  INV_X2 U12841 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20525) );
  INV_X1 U12842 ( .A(n10243), .ZN(n13475) );
  INV_X1 U12843 ( .A(n12754), .ZN(n12765) );
  NAND2_X1 U12844 ( .A1(n13221), .A2(n13220), .ZN(n13223) );
  OR2_X1 U12845 ( .A1(n14267), .A2(n14936), .ZN(n13029) );
  OR2_X1 U12846 ( .A1(n15476), .A2(n15504), .ZN(n15493) );
  AND2_X1 U12847 ( .A1(n14242), .A2(n15515), .ZN(n12192) );
  XNOR2_X1 U12848 ( .A(n12232), .B(n12233), .ZN(n12970) );
  OR3_X1 U12849 ( .A1(n19234), .A2(n19417), .A3(n19230), .ZN(n19260) );
  NAND2_X1 U12850 ( .A1(n19445), .A2(n19884), .ZN(n19386) );
  OR2_X1 U12851 ( .A1(n12142), .A2(n13497), .ZN(n10825) );
  OR2_X1 U12852 ( .A1(n19618), .A2(n19612), .ZN(n19655) );
  INV_X1 U12853 ( .A(n19445), .ZN(n19857) );
  NAND2_X1 U12854 ( .A1(n20708), .A2(n19877), .ZN(n19419) );
  INV_X1 U12855 ( .A(n16571), .ZN(n16572) );
  NOR2_X1 U12856 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16765), .ZN(n16750) );
  NOR2_X1 U12857 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16831), .ZN(n16821) );
  INV_X1 U12858 ( .A(n16927), .ZN(n16868) );
  INV_X1 U12859 ( .A(n9696), .ZN(n16887) );
  NOR2_X1 U12860 ( .A1(n17880), .A2(n17540), .ZN(n17883) );
  OAI21_X1 U12861 ( .B1(n17610), .B2(n17866), .A(n18488), .ZN(n17707) );
  INV_X1 U12862 ( .A(n17707), .ZN(n17630) );
  INV_X1 U12863 ( .A(n12724), .ZN(n17579) );
  CLKBUF_X1 U12864 ( .A(n16747), .Z(n17708) );
  INV_X1 U12865 ( .A(n16384), .ZN(n17660) );
  NAND2_X1 U12866 ( .A1(n17705), .A2(n17871), .ZN(n17610) );
  NOR2_X1 U12867 ( .A1(n17823), .A2(n17822), .ZN(n17821) );
  INV_X1 U12868 ( .A(n18663), .ZN(n18082) );
  INV_X1 U12869 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20932) );
  NOR2_X1 U12870 ( .A1(n12621), .A2(n12620), .ZN(n12707) );
  OR3_X1 U12871 ( .A1(n13113), .A2(n13134), .A3(n13277), .ZN(n13336) );
  OAI22_X1 U12872 ( .A1(n14526), .A2(n14629), .B1(n14531), .B2(n20023), .ZN(
        n12901) );
  INV_X1 U12873 ( .A(n11008), .ZN(n12900) );
  AND2_X1 U12874 ( .A1(n13173), .A2(n13172), .ZN(n20035) );
  INV_X1 U12875 ( .A(n13361), .ZN(n20053) );
  NAND2_X1 U12876 ( .A1(n13334), .A2(n13333), .ZN(n13388) );
  AND2_X1 U12877 ( .A1(n11919), .A2(n11918), .ZN(n14624) );
  AND2_X1 U12878 ( .A1(n14699), .A2(n14700), .ZN(n14701) );
  INV_X1 U12879 ( .A(n11667), .ZN(n11668) );
  AND2_X1 U12880 ( .A1(n14803), .A2(n12109), .ZN(n20070) );
  OR2_X1 U12881 ( .A1(n11562), .A2(n11561), .ZN(n14856) );
  NOR2_X1 U12882 ( .A1(n20101), .A2(n13290), .ZN(n20108) );
  INV_X1 U12883 ( .A(n20216), .ZN(n20184) );
  OR2_X1 U12884 ( .A1(n14902), .A2(n11622), .ZN(n20324) );
  NAND2_X1 U12885 ( .A1(n20117), .A2(n20116), .ZN(n20224) );
  OR2_X1 U12886 ( .A1(n14902), .A2(n13609), .ZN(n20262) );
  INV_X1 U12887 ( .A(n14043), .ZN(n20312) );
  OAI211_X1 U12888 ( .C1(n13988), .C2(n20439), .A(n20354), .B(n13956), .ZN(
        n13987) );
  INV_X1 U12889 ( .A(n20383), .ZN(n20339) );
  OAI22_X1 U12890 ( .A1(n20361), .A2(n20360), .B1(n20359), .B2(n20489), .ZN(
        n20385) );
  INV_X1 U12891 ( .A(n20389), .ZN(n20530) );
  OAI22_X1 U12892 ( .A1(n20444), .A2(n20443), .B1(n20490), .B2(n20442), .ZN(
        n20481) );
  INV_X1 U12893 ( .A(n20390), .ZN(n20404) );
  INV_X1 U12894 ( .A(n20491), .ZN(n20515) );
  AND2_X1 U12895 ( .A1(n16233), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20589) );
  INV_X1 U12896 ( .A(n20703), .ZN(n19005) );
  AND2_X1 U12897 ( .A1(n14943), .A2(n12829), .ZN(n20703) );
  INV_X1 U12898 ( .A(n20697), .ZN(n18986) );
  INV_X1 U12899 ( .A(n20705), .ZN(n19007) );
  INV_X1 U12900 ( .A(n19041), .ZN(n19018) );
  AND2_X1 U12901 ( .A1(n13874), .A2(n15653), .ZN(n19060) );
  INV_X1 U12902 ( .A(n19095), .ZN(n19119) );
  INV_X1 U12903 ( .A(n19152), .ZN(n19157) );
  INV_X1 U12904 ( .A(n13051), .ZN(n13038) );
  OAI21_X1 U12905 ( .B1(n16278), .B2(n15652), .A(n10837), .ZN(n10838) );
  INV_X1 U12906 ( .A(n19172), .ZN(n16343) );
  INV_X1 U12907 ( .A(n19184), .ZN(n16322) );
  NOR2_X1 U12908 ( .A1(n15567), .A2(n12198), .ZN(n15516) );
  INV_X1 U12909 ( .A(n15629), .ZN(n16357) );
  AND2_X1 U12910 ( .A1(n12377), .A2(n12371), .ZN(n16354) );
  OAI21_X1 U12911 ( .B1(n15646), .B2(n15649), .A(n15644), .ZN(n19224) );
  NOR2_X2 U12912 ( .A1(n19479), .A2(n19386), .ZN(n19262) );
  NOR2_X1 U12913 ( .A1(n19608), .A2(n19386), .ZN(n19380) );
  OAI21_X1 U12914 ( .B1(n19408), .B2(n19668), .A(n19393), .ZN(n19410) );
  NOR2_X2 U12915 ( .A1(n19419), .A2(n19386), .ZN(n19440) );
  OAI21_X1 U12916 ( .B1(n19473), .B2(n19452), .A(n19621), .ZN(n19475) );
  INV_X1 U12917 ( .A(n19856), .ZN(n19868) );
  INV_X1 U12918 ( .A(n19536), .ZN(n19572) );
  OAI21_X1 U12919 ( .B1(n19579), .B2(n19578), .A(n19577), .ZN(n19603) );
  INV_X1 U12920 ( .A(n19660), .ZN(n19650) );
  OAI21_X1 U12921 ( .B1(n19676), .B2(n19675), .A(n19674), .ZN(n19714) );
  INV_X1 U12922 ( .A(n19616), .ZN(n19608) );
  INV_X1 U12923 ( .A(n19700), .ZN(n19760) );
  INV_X1 U12924 ( .A(n19218), .ZN(n19777) );
  AND3_X1 U12925 ( .A1(n13837), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18862) );
  AOI22_X1 U12926 ( .A1(n18634), .A2(n18630), .B1(n16418), .B2(n18635), .ZN(
        n18639) );
  XNOR2_X1 U12927 ( .A(n16573), .B(n16572), .ZN(n16577) );
  NOR2_X1 U12928 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16653), .ZN(n16637) );
  NOR2_X1 U12929 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16668), .ZN(n16656) );
  NOR2_X1 U12930 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16737), .ZN(n16724) );
  NOR2_X1 U12931 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16789), .ZN(n16769) );
  NAND2_X1 U12932 ( .A1(n16539), .A2(n18184), .ZN(n16922) );
  INV_X1 U12933 ( .A(n16913), .ZN(n16896) );
  NOR2_X1 U12934 ( .A1(n17011), .A2(n17012), .ZN(n16985) );
  NOR2_X1 U12935 ( .A1(n17280), .A2(n17036), .ZN(n17023) );
  NAND2_X1 U12936 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17135), .ZN(n17119) );
  NAND4_X1 U12937 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17227), .A4(n17209), .ZN(n17208) );
  INV_X1 U12938 ( .A(n17243), .ZN(n17239) );
  NOR3_X1 U12939 ( .A1(n17280), .A2(n17313), .A3(n17446), .ZN(n17305) );
  NAND3_X1 U12940 ( .A1(n12495), .A2(n12494), .A3(n12493), .ZN(n16417) );
  INV_X2 U12941 ( .A(n17295), .ZN(n17366) );
  INV_X1 U12942 ( .A(n17438), .ZN(n17436) );
  NAND2_X1 U12943 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17506) );
  NOR2_X1 U12944 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18201), .ZN(n18305) );
  INV_X1 U12945 ( .A(n17770), .ZN(n17603) );
  OR2_X1 U12946 ( .A1(n17556), .A2(n17917), .ZN(n17540) );
  INV_X1 U12947 ( .A(n18182), .ZN(n18176) );
  INV_X1 U12948 ( .A(n18190), .ZN(n18150) );
  INV_X1 U12949 ( .A(n18141), .ZN(n18178) );
  INV_X1 U12950 ( .A(n18636), .ZN(n16418) );
  INV_X1 U12951 ( .A(n18305), .ZN(n18486) );
  INV_X1 U12952 ( .A(n18692), .ZN(n18699) );
  INV_X1 U12953 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18705) );
  NAND2_X1 U12954 ( .A1(n13336), .A2(n13147), .ZN(n20681) );
  INV_X1 U12955 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20321) );
  INV_X1 U12956 ( .A(n19993), .ZN(n20010) );
  NAND2_X1 U12957 ( .A1(n20009), .A2(n13906), .ZN(n15977) );
  NAND2_X1 U12958 ( .A1(n20009), .A2(n13917), .ZN(n19991) );
  INV_X1 U12959 ( .A(n14715), .ZN(n14648) );
  NAND2_X1 U12960 ( .A1(n13548), .A2(n13565), .ZN(n16029) );
  INV_X1 U12961 ( .A(n20038), .ZN(n20044) );
  INV_X1 U12962 ( .A(n13351), .ZN(n13387) );
  INV_X1 U12963 ( .A(n12114), .ZN(n12115) );
  XNOR2_X1 U12964 ( .A(n11312), .B(n14746), .ZN(n14760) );
  OAI21_X1 U12965 ( .B1(n14701), .B2(n14639), .A(n14638), .ZN(n15978) );
  INV_X1 U12966 ( .A(n20070), .ZN(n20066) );
  INV_X1 U12967 ( .A(n20103), .ZN(n16186) );
  INV_X1 U12968 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20317) );
  NAND2_X1 U12969 ( .A1(n20119), .A2(n20118), .ZN(n20182) );
  OR2_X1 U12970 ( .A1(n20224), .A2(n20324), .ZN(n20216) );
  OR2_X1 U12971 ( .A1(n20224), .A2(n20487), .ZN(n20253) );
  OR2_X1 U12972 ( .A1(n20224), .A2(n20402), .ZN(n20279) );
  OR2_X1 U12973 ( .A1(n20292), .A2(n20262), .ZN(n20316) );
  INV_X1 U12974 ( .A(n20345), .ZN(n20342) );
  NAND2_X1 U12975 ( .A1(n20404), .A2(n20325), .ZN(n20383) );
  NAND2_X1 U12976 ( .A1(n20404), .A2(n20349), .ZN(n20430) );
  NAND2_X1 U12977 ( .A1(n20404), .A2(n20403), .ZN(n20485) );
  OR2_X1 U12978 ( .A1(n20529), .A2(n20487), .ZN(n20543) );
  OR2_X1 U12979 ( .A1(n20529), .A2(n20402), .ZN(n20587) );
  INV_X1 U12980 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16233) );
  INV_X1 U12981 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19666) );
  OR2_X1 U12982 ( .A1(n14932), .A2(n12794), .ZN(n20705) );
  AND2_X1 U12983 ( .A1(n13111), .A2(n18862), .ZN(n19048) );
  NAND2_X1 U12984 ( .A1(n13155), .A2(n13154), .ZN(n19095) );
  INV_X1 U12985 ( .A(n19096), .ZN(n19128) );
  INV_X1 U12986 ( .A(n19166), .ZN(n19152) );
  INV_X1 U12987 ( .A(n19154), .ZN(n19170) );
  OR2_X1 U12988 ( .A1(n12981), .A2(n13143), .ZN(n14267) );
  INV_X1 U12989 ( .A(n10838), .ZN(n10878) );
  INV_X1 U12990 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16342) );
  NAND2_X1 U12991 ( .A1(n18864), .A2(n10826), .ZN(n19184) );
  NOR2_X1 U12992 ( .A1(n12382), .A2(n12381), .ZN(n12383) );
  INV_X1 U12993 ( .A(n16359), .ZN(n15623) );
  INV_X1 U12994 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15870) );
  NAND2_X1 U12995 ( .A1(n19232), .A2(n19414), .ZN(n19293) );
  AND2_X1 U12996 ( .A1(n19300), .A2(n19299), .ZN(n19308) );
  INV_X1 U12997 ( .A(n19317), .ZN(n19327) );
  INV_X1 U12998 ( .A(n19344), .ZN(n19356) );
  INV_X1 U12999 ( .A(n19380), .ZN(n19378) );
  INV_X1 U13000 ( .A(n19387), .ZN(n19413) );
  NAND2_X1 U13001 ( .A1(n19414), .A2(n19728), .ZN(n19478) );
  INV_X1 U13002 ( .A(n19503), .ZN(n19511) );
  AND2_X1 U13003 ( .A1(n19518), .A2(n19621), .ZN(n19524) );
  OR2_X1 U13004 ( .A1(n19609), .A2(n19479), .ZN(n19544) );
  OR2_X1 U13005 ( .A1(n19609), .A2(n19856), .ZN(n19607) );
  OR2_X1 U13006 ( .A1(n19609), .A2(n19608), .ZN(n19718) );
  INV_X1 U13007 ( .A(n19565), .ZN(n19765) );
  INV_X1 U13008 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13837) );
  INV_X1 U13009 ( .A(n19851), .ZN(n19783) );
  NOR2_X1 U13010 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16718), .ZN(n16709) );
  INV_X1 U13011 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17737) );
  INV_X1 U13012 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17203) );
  NOR2_X1 U13013 ( .A1(n16979), .A2(n15664), .ZN(n16969) );
  NOR2_X1 U13014 ( .A1(n16966), .A2(n16979), .ZN(n16984) );
  NOR2_X1 U13015 ( .A1(n16790), .A2(n17121), .ZN(n17135) );
  AND2_X1 U13016 ( .A1(n17227), .A2(n17280), .ZN(n17229) );
  NOR2_X1 U13017 ( .A1(n17420), .A2(n17341), .ZN(n17344) );
  INV_X1 U13018 ( .A(n12677), .ZN(n17356) );
  INV_X1 U13019 ( .A(n17373), .ZN(n17371) );
  INV_X1 U13020 ( .A(n17407), .ZN(n17406) );
  NAND2_X1 U13021 ( .A1(n17438), .A2(n17440), .ZN(n17439) );
  INV_X1 U13022 ( .A(n17489), .ZN(n17481) );
  INV_X1 U13023 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17808) );
  OAI21_X2 U13024 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18842), .A(n16522), 
        .ZN(n17871) );
  INV_X1 U13025 ( .A(n17839), .ZN(n17875) );
  NAND2_X1 U13026 ( .A1(n18184), .A2(n18176), .ZN(n18141) );
  INV_X1 U13027 ( .A(n18089), .ZN(n18110) );
  INV_X1 U13028 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18668) );
  INV_X1 U13029 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18678) );
  INV_X1 U13030 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18800) );
  INV_X1 U13031 ( .A(n18786), .ZN(n18783) );
  INV_X1 U13032 ( .A(n16476), .ZN(n16475) );
  NAND2_X1 U13033 ( .A1(n12903), .A2(n12902), .ZN(P1_U2842) );
  NAND2_X1 U13034 ( .A1(n12409), .A2(n12408), .ZN(P1_U2873) );
  NAND2_X1 U13035 ( .A1(n10112), .A2(n11569), .ZN(P1_U3003) );
  OAI211_X1 U13036 ( .C1(n15138), .C2(n11600), .A(n11599), .B(n11598), .ZN(
        P2_U2987) );
  AOI22_X1 U13037 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10133) );
  AND3_X4 U13038 ( .A1(n13437), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10327) );
  AND3_X4 U13039 ( .A1(n13444), .A2(n10129), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U13040 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U13041 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U13042 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10134) );
  AND2_X1 U13043 ( .A1(n10134), .A2(n10334), .ZN(n10138) );
  AOI22_X1 U13044 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9693), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13045 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13046 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U13047 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U13048 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13049 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U13050 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U13051 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U13052 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13053 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U13054 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U13055 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13056 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9751), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13057 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13058 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10148) );
  NAND3_X1 U13059 ( .A1(n10151), .A2(n10150), .A3(n10111), .ZN(n10158) );
  AOI22_X1 U13060 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13061 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U13062 ( .A1(n10328), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9693), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10155) );
  NAND3_X1 U13063 ( .A1(n10156), .A2(n10114), .A3(n10155), .ZN(n10157) );
  NAND2_X1 U13064 ( .A1(n12153), .A2(n10227), .ZN(n12152) );
  AOI22_X1 U13065 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13066 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13067 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13068 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10159) );
  NAND4_X1 U13069 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10163) );
  NAND2_X1 U13070 ( .A1(n10163), .A2(n10334), .ZN(n10170) );
  AOI22_X1 U13071 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13072 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U13073 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9751), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13074 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10164) );
  NAND4_X1 U13075 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10168) );
  NAND2_X1 U13076 ( .A1(n10168), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10169) );
  NAND3_X1 U13077 ( .A1(n12152), .A2(n12148), .A3(n19215), .ZN(n12179) );
  AOI22_X1 U13078 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13079 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13080 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13081 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10171) );
  NAND4_X1 U13082 ( .A1(n10174), .A2(n10173), .A3(n10172), .A4(n10171), .ZN(
        n10180) );
  AOI22_X1 U13083 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9763), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13084 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U13085 ( .A1(n10328), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9751), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13086 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10175) );
  NAND4_X1 U13087 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10179) );
  NAND2_X1 U13088 ( .A1(n12179), .A2(n15654), .ZN(n10195) );
  AOI22_X1 U13089 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13090 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9693), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13091 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13092 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10182) );
  NAND4_X1 U13093 ( .A1(n10185), .A2(n10184), .A3(n10183), .A4(n10182), .ZN(
        n10186) );
  AOI22_X1 U13094 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9751), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13095 ( .A1(n9758), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13096 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13097 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10187) );
  NAND4_X1 U13098 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10191) );
  NAND2_X1 U13099 ( .A1(n10191), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10192) );
  AOI21_X1 U13100 ( .B1(n12172), .B2(n10245), .A(n13475), .ZN(n10194) );
  NAND2_X1 U13101 ( .A1(n10195), .A2(n10194), .ZN(n10206) );
  AOI22_X1 U13102 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9693), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U13103 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13104 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13105 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13106 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13107 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13108 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13109 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U13110 ( .A1(n10221), .A2(n9761), .ZN(n12173) );
  AOI22_X1 U13111 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9753), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13112 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13113 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9693), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13114 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13115 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9752), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13116 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13117 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9751), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13118 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10211) );
  MUX2_X2 U13119 ( .A(n10115), .B(n10215), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10228) );
  AND2_X1 U13120 ( .A1(n12214), .A2(n10216), .ZN(n10217) );
  NAND2_X1 U13121 ( .A1(n10232), .A2(n10236), .ZN(n10219) );
  NAND2_X1 U13122 ( .A1(n10221), .A2(n15654), .ZN(n10246) );
  NAND2_X1 U13123 ( .A1(n15658), .A2(n19215), .ZN(n10242) );
  OAI21_X1 U13124 ( .B1(n10222), .B2(n15658), .A(n10242), .ZN(n10223) );
  INV_X1 U13125 ( .A(n10232), .ZN(n10225) );
  NOR2_X1 U13126 ( .A1(n9761), .A2(n10236), .ZN(n10226) );
  NAND2_X1 U13127 ( .A1(n10717), .A2(n10226), .ZN(n10230) );
  NAND2_X1 U13128 ( .A1(n10243), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12129) );
  INV_X1 U13129 ( .A(n12129), .ZN(n10231) );
  NAND2_X1 U13130 ( .A1(n10291), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10241) );
  NOR2_X1 U13131 ( .A1(n10232), .A2(n10228), .ZN(n10233) );
  INV_X1 U13132 ( .A(n12819), .ZN(n10235) );
  NAND2_X1 U13133 ( .A1(n12145), .A2(n10235), .ZN(n12367) );
  INV_X1 U13134 ( .A(n12367), .ZN(n10238) );
  NAND2_X1 U13135 ( .A1(n12185), .A2(n13093), .ZN(n12170) );
  AND2_X1 U13136 ( .A1(n19215), .A2(n10216), .ZN(n13157) );
  NAND2_X1 U13137 ( .A1(n13157), .A2(n10218), .ZN(n10237) );
  NOR2_X1 U13138 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13492) );
  INV_X1 U13139 ( .A(n10242), .ZN(n10244) );
  NAND2_X1 U13140 ( .A1(n9734), .A2(n13491), .ZN(n10247) );
  NAND2_X2 U13141 ( .A1(n10248), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10286) );
  INV_X1 U13142 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10256) );
  INV_X1 U13143 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U13144 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10252) );
  INV_X1 U13145 ( .A(n10286), .ZN(n10259) );
  INV_X1 U13146 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13097) );
  NAND2_X1 U13147 ( .A1(n10259), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10265) );
  NAND2_X1 U13148 ( .A1(n10815), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10262) );
  INV_X1 U13149 ( .A(n13492), .ZN(n10267) );
  NAND2_X1 U13150 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10260) );
  INV_X1 U13151 ( .A(n10266), .ZN(n10269) );
  NAND2_X1 U13152 ( .A1(n10291), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10270) );
  NAND2_X2 U13153 ( .A1(n10299), .A2(n10301), .ZN(n10300) );
  INV_X1 U13154 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10444) );
  INV_X1 U13155 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20696) );
  NAND2_X1 U13156 ( .A1(n9744), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U13157 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10274) );
  OAI211_X1 U13158 ( .C1(n20696), .C2(n10273), .A(n10275), .B(n10274), .ZN(
        n10276) );
  INV_X1 U13159 ( .A(n10276), .ZN(n10277) );
  NAND2_X1 U13160 ( .A1(n10278), .A2(n10277), .ZN(n10281) );
  NAND2_X1 U13161 ( .A1(n10291), .A2(n14352), .ZN(n10280) );
  AOI21_X1 U13162 ( .B1(n16380), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U13163 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  INV_X1 U13164 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U13165 ( .A1(n10751), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U13166 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10287) );
  OAI211_X1 U13167 ( .C1(n10289), .C2(n10273), .A(n10288), .B(n10287), .ZN(
        n10290) );
  NAND2_X1 U13168 ( .A1(n10291), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10293) );
  NAND2_X1 U13169 ( .A1(n13492), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U13170 ( .A1(n13793), .A2(n13449), .ZN(n10318) );
  AOI22_X1 U13171 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9701), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10314) );
  INV_X1 U13172 ( .A(n10297), .ZN(n10302) );
  INV_X1 U13173 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10305) );
  INV_X1 U13174 ( .A(n10318), .ZN(n10306) );
  INV_X1 U13175 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10308) );
  NOR2_X1 U13176 ( .A1(n10374), .A2(n10308), .ZN(n10309) );
  NOR2_X1 U13177 ( .A1(n10310), .A2(n10309), .ZN(n10313) );
  AOI22_X1 U13178 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10483), .B1(
        n19580), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10312) );
  AND2_X2 U13179 ( .A1(n10307), .A2(n10303), .ZN(n10480) );
  AOI22_X1 U13180 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10493), .B1(
        n10480), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U13181 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10369) );
  AOI22_X1 U13182 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10492), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10325) );
  NOR2_X2 U13183 ( .A1(n10316), .A2(n10315), .ZN(n10537) );
  NOR2_X1 U13184 ( .A1(n10319), .A2(n10317), .ZN(n10481) );
  AOI22_X1 U13185 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10537), .B1(
        n10481), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10324) );
  NOR2_X1 U13186 ( .A1(n10319), .A2(n10320), .ZN(n10490) );
  AOI22_X1 U13187 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10479), .B1(
        n10490), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10323) );
  AND2_X2 U13188 ( .A1(n10304), .A2(n10321), .ZN(n10491) );
  AOI22_X1 U13189 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10482), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13190 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10368) );
  AND2_X2 U13191 ( .A1(n13454), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14368) );
  AOI22_X1 U13192 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13193 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10331) );
  AND2_X2 U13194 ( .A1(n10327), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10384) );
  AOI22_X1 U13195 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10330) );
  AND2_X2 U13196 ( .A1(n13454), .A2(n13444), .ZN(n14369) );
  AOI22_X1 U13197 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13198 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10341) );
  AND2_X2 U13199 ( .A1(n14467), .A2(n10334), .ZN(n10459) );
  AOI22_X1 U13200 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10339) );
  AND2_X1 U13201 ( .A1(n10147), .A2(n10334), .ZN(n10396) );
  AOI22_X1 U13202 ( .A1(n10396), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10338) );
  INV_X1 U13203 ( .A(n10333), .ZN(n13430) );
  AOI22_X1 U13204 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10337) );
  AND2_X1 U13205 ( .A1(n14400), .A2(n10334), .ZN(n10335) );
  AOI22_X1 U13206 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10336) );
  NAND4_X1 U13207 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10340) );
  AOI22_X1 U13208 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13209 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13210 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13211 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10342) );
  NAND4_X1 U13212 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10342), .ZN(
        n10352) );
  AOI22_X1 U13213 ( .A1(n10396), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13214 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13215 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13216 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U13217 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  NOR2_X1 U13218 ( .A1(n13099), .A2(n12228), .ZN(n10353) );
  NAND2_X1 U13219 ( .A1(n9761), .A2(n10353), .ZN(n10844) );
  AOI22_X1 U13220 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10452), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13221 ( .A1(n10396), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13222 ( .A1(n10379), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13223 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10355) );
  NAND4_X1 U13224 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10366) );
  AOI22_X1 U13225 ( .A1(n10359), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13226 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13227 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13228 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10361) );
  NAND4_X1 U13229 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10365) );
  NAND2_X1 U13230 ( .A1(n10844), .A2(n10843), .ZN(n10367) );
  OAI21_X2 U13231 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(n10475) );
  AOI22_X1 U13232 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10488), .B1(
        n10489), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13233 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19580), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13234 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10493), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13235 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10492), .B1(
        n10479), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10370) );
  NAND4_X1 U13236 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10394) );
  INV_X2 U13237 ( .A(n10374), .ZN(n19673) );
  AOI22_X1 U13238 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19673), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13239 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9701), .B1(
        n10480), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13240 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10490), .B1(
        n10481), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13241 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10483), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13242 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10393) );
  AOI22_X1 U13243 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10452), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13244 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13245 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13246 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10380) );
  NAND4_X1 U13247 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10390) );
  AOI22_X1 U13248 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13249 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13250 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13251 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U13252 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  INV_X1 U13253 ( .A(n12243), .ZN(n10391) );
  NAND2_X1 U13254 ( .A1(n10391), .A2(n9761), .ZN(n10392) );
  OAI21_X2 U13255 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(n10476) );
  NAND2_X1 U13256 ( .A1(n10475), .A2(n10476), .ZN(n10395) );
  NAND2_X1 U13257 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10400) );
  NAND2_X1 U13258 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13259 ( .A1(n10396), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10398) );
  NAND2_X1 U13260 ( .A1(n10379), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10397) );
  NAND2_X1 U13261 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13262 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13263 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10402) );
  NAND2_X1 U13264 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10401) );
  NAND2_X1 U13265 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10411) );
  NAND2_X1 U13266 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13267 ( .A1(n10359), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10409) );
  INV_X1 U13268 ( .A(n10405), .ZN(n10407) );
  INV_X1 U13269 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10406) );
  OR2_X1 U13270 ( .A1(n10407), .A2(n10406), .ZN(n10408) );
  NAND2_X1 U13271 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10417) );
  NAND2_X1 U13272 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10416) );
  NAND2_X1 U13273 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10415) );
  INV_X1 U13274 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10412) );
  OR2_X1 U13275 ( .A1(n10413), .A2(n10412), .ZN(n10414) );
  AND4_X2 U13276 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10861) );
  XNOR2_X1 U13277 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U13278 ( .A1(n19890), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10704) );
  INV_X1 U13279 ( .A(n10704), .ZN(n10422) );
  NAND2_X1 U13280 ( .A1(n12125), .A2(n10422), .ZN(n10424) );
  NAND2_X1 U13281 ( .A1(n19881), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U13282 ( .A1(n10424), .A2(n10423), .ZN(n10432) );
  XNOR2_X1 U13283 ( .A(n14352), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13284 ( .A1(n10432), .A2(n10430), .ZN(n10426) );
  NAND2_X1 U13285 ( .A1(n19871), .A2(n14352), .ZN(n10425) );
  NAND2_X1 U13286 ( .A1(n10426), .A2(n10425), .ZN(n10471) );
  XNOR2_X1 U13287 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10470) );
  INV_X1 U13288 ( .A(n10470), .ZN(n10427) );
  XNOR2_X1 U13289 ( .A(n10471), .B(n10427), .ZN(n12133) );
  MUX2_X1 U13290 ( .A(n12243), .B(n12133), .S(n12828), .Z(n10713) );
  INV_X1 U13291 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13644) );
  MUX2_X1 U13292 ( .A(n10713), .B(n13644), .S(n10428), .Z(n10440) );
  INV_X1 U13293 ( .A(n10430), .ZN(n10431) );
  XNOR2_X1 U13294 ( .A(n10432), .B(n10431), .ZN(n12127) );
  INV_X1 U13295 ( .A(n12127), .ZN(n12128) );
  INV_X1 U13296 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13145) );
  INV_X1 U13297 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n18998) );
  NAND2_X1 U13298 ( .A1(n13145), .A2(n18998), .ZN(n10437) );
  INV_X1 U13299 ( .A(n10512), .ZN(n10438) );
  OAI21_X1 U13300 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(n13647) );
  OAI21_X1 U13301 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19890), .A(
        n10704), .ZN(n10699) );
  MUX2_X1 U13302 ( .A(n10699), .B(n13099), .S(n10429), .Z(n10712) );
  MUX2_X1 U13303 ( .A(n10712), .B(n18998), .S(n10428), .Z(n19004) );
  NOR2_X1 U13304 ( .A1(n19004), .A2(n13097), .ZN(n13096) );
  INV_X1 U13305 ( .A(n13096), .ZN(n12967) );
  NAND3_X1 U13306 ( .A1(n10428), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10441) );
  NOR2_X1 U13307 ( .A1(n12967), .A2(n13791), .ZN(n10442) );
  NAND2_X1 U13308 ( .A1(n12967), .A2(n13791), .ZN(n12966) );
  OAI21_X1 U13309 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10442), .A(
        n12966), .ZN(n14233) );
  XNOR2_X1 U13310 ( .A(n10445), .B(n10444), .ZN(n14232) );
  OR2_X1 U13311 ( .A1(n14233), .A2(n14232), .ZN(n14235) );
  INV_X1 U13312 ( .A(n10445), .ZN(n20702) );
  NAND2_X1 U13313 ( .A1(n20702), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10446) );
  NAND2_X1 U13314 ( .A1(n14235), .A2(n10446), .ZN(n13801) );
  INV_X1 U13315 ( .A(n13801), .ZN(n10447) );
  NAND2_X1 U13316 ( .A1(n13799), .A2(n10447), .ZN(n10451) );
  INV_X1 U13317 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19047) );
  AOI22_X1 U13318 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10452), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13319 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10462) );
  INV_X1 U13320 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n20853) );
  INV_X1 U13321 ( .A(n10453), .ZN(n10457) );
  INV_X1 U13322 ( .A(n10454), .ZN(n10456) );
  INV_X1 U13323 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10455) );
  OAI22_X1 U13324 ( .A1(n20853), .A2(n10457), .B1(n10456), .B2(n10455), .ZN(
        n10458) );
  INV_X1 U13325 ( .A(n10458), .ZN(n10461) );
  AOI22_X1 U13326 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10460) );
  NAND4_X1 U13327 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10469) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13329 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13330 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13331 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10464) );
  NAND4_X1 U13332 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10468) );
  NAND2_X1 U13333 ( .A1(n10471), .A2(n10470), .ZN(n10473) );
  NAND2_X1 U13334 ( .A1(n19864), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13335 ( .A1(n10473), .A2(n10472), .ZN(n10701) );
  MUX2_X1 U13336 ( .A(n12248), .B(n12138), .S(n12828), .Z(n12121) );
  MUX2_X1 U13337 ( .A(n19047), .B(n12121), .S(n12214), .Z(n10511) );
  XNOR2_X1 U13338 ( .A(n10512), .B(n9955), .ZN(n10474) );
  XNOR2_X1 U13339 ( .A(n10474), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13884) );
  INV_X1 U13340 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14006) );
  INV_X1 U13341 ( .A(n10474), .ZN(n13688) );
  INV_X1 U13342 ( .A(n10475), .ZN(n10478) );
  INV_X1 U13343 ( .A(n10476), .ZN(n10477) );
  AOI22_X1 U13344 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19269), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13345 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19580), .B1(
        n10480), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13346 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n15647), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13347 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10483), .B1(
        n19673), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13348 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10488), .B1(
        n10489), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13349 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19302), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13350 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n9701), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13351 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10492), .B1(
        n10493), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10494) );
  AND4_X1 U13352 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10498) );
  NAND2_X1 U13353 ( .A1(n9800), .A2(n10498), .ZN(n10510) );
  AOI22_X1 U13354 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13355 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13356 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13357 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10499) );
  NAND4_X1 U13358 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10508) );
  AOI22_X1 U13359 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13360 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13361 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13362 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10503) );
  NAND4_X1 U13363 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10507) );
  NAND2_X1 U13364 ( .A1(n12253), .A2(n9761), .ZN(n10509) );
  NAND2_X1 U13365 ( .A1(n10510), .A2(n10509), .ZN(n10530) );
  MUX2_X1 U13366 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12253), .S(n12214), .Z(
        n10513) );
  AND2_X1 U13367 ( .A1(n10514), .A2(n10513), .ZN(n10515) );
  OR2_X1 U13368 ( .A1(n10515), .A2(n10566), .ZN(n18983) );
  AND2_X1 U13369 ( .A1(n18983), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10519) );
  AND2_X1 U13370 ( .A1(n10861), .A2(n9891), .ZN(n10520) );
  INV_X1 U13371 ( .A(n10520), .ZN(n10516) );
  NAND2_X1 U13372 ( .A1(n10530), .A2(n10516), .ZN(n10517) );
  NAND2_X1 U13373 ( .A1(n10518), .A2(n10517), .ZN(n10525) );
  MUX2_X1 U13374 ( .A(n10520), .B(n10519), .S(n10530), .Z(n10521) );
  NAND2_X1 U13375 ( .A1(n10526), .A2(n10521), .ZN(n10524) );
  OAI21_X1 U13376 ( .B1(n10861), .B2(n9891), .A(n18983), .ZN(n10522) );
  OAI21_X1 U13377 ( .B1(n18983), .B2(n9891), .A(n10522), .ZN(n10523) );
  OAI211_X1 U13378 ( .C1(n10526), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n13999) );
  NAND2_X1 U13379 ( .A1(n14000), .A2(n13999), .ZN(n10529) );
  OAI21_X1 U13380 ( .B1(n10851), .B2(n10687), .A(n18983), .ZN(n10527) );
  NAND2_X1 U13381 ( .A1(n10527), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10528) );
  NAND2_X1 U13382 ( .A1(n10529), .A2(n10528), .ZN(n14036) );
  INV_X1 U13383 ( .A(n10530), .ZN(n10532) );
  INV_X1 U13384 ( .A(n10559), .ZN(n10558) );
  AOI22_X1 U13385 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10492), .B1(
        n10489), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13386 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19269), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19302), .B1(
        n9701), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13388 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10483), .B1(
        n19673), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10533) );
  NAND4_X1 U13389 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10543) );
  AOI22_X1 U13390 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10493), .B1(
        n10488), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10541) );
  INV_X1 U13391 ( .A(n10537), .ZN(n19358) );
  AOI22_X1 U13392 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10537), .B1(
        n19580), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13393 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n15647), .B1(
        n10480), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10482), .B1(
        n9699), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10538) );
  NAND4_X1 U13395 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10542) );
  AOI22_X1 U13396 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10452), .B1(
        n10346), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13397 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10396), .B1(
        n10453), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13398 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10379), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U13400 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10553) );
  AOI22_X1 U13401 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12265), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13402 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n14369), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13403 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13404 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14368), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10548) );
  NAND4_X1 U13405 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10552) );
  INV_X1 U13406 ( .A(n12257), .ZN(n10554) );
  NAND2_X1 U13407 ( .A1(n10554), .A2(n9761), .ZN(n10555) );
  NAND2_X1 U13408 ( .A1(n10559), .A2(n10854), .ZN(n10560) );
  INV_X1 U13409 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13266) );
  MUX2_X1 U13410 ( .A(n12257), .B(n13266), .S(n10428), .Z(n10565) );
  XNOR2_X1 U13411 ( .A(n10566), .B(n10565), .ZN(n18971) );
  INV_X1 U13412 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14033) );
  NAND2_X1 U13413 ( .A1(n10562), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10563) );
  MUX2_X1 U13414 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n10861), .S(n12214), .Z(
        n10570) );
  NAND3_X1 U13415 ( .A1(n10574), .A2(P2_EBX_REG_8__SCAN_IN), .A3(n10428), .ZN(
        n10568) );
  OR2_X1 U13416 ( .A1(n10574), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10567) );
  AND3_X1 U13417 ( .A1(n10669), .A2(n10568), .A3(n10567), .ZN(n13670) );
  INV_X1 U13418 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20760) );
  NOR2_X1 U13419 ( .A1(n10861), .A2(n20760), .ZN(n10569) );
  NAND2_X1 U13420 ( .A1(n13670), .A2(n10569), .ZN(n16332) );
  NAND2_X1 U13421 ( .A1(n10571), .A2(n10570), .ZN(n10572) );
  NAND2_X1 U13422 ( .A1(n10574), .A2(n10572), .ZN(n13622) );
  INV_X1 U13423 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15618) );
  OR2_X1 U13424 ( .A1(n13622), .A2(n15618), .ZN(n16330) );
  NOR2_X2 U13425 ( .A1(n10574), .A2(n10573), .ZN(n10585) );
  INV_X1 U13426 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U13427 ( .A1(n10585), .A2(n10575), .ZN(n10580) );
  NAND2_X1 U13428 ( .A1(n10428), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10576) );
  OR2_X1 U13429 ( .A1(n10577), .A2(n10576), .ZN(n10579) );
  INV_X1 U13430 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U13431 ( .A1(n10577), .A2(n13725), .ZN(n10592) );
  INV_X1 U13432 ( .A(n10590), .ZN(n10578) );
  NAND2_X1 U13433 ( .A1(n10579), .A2(n10578), .ZN(n18938) );
  OR2_X1 U13434 ( .A1(n18938), .A2(n10861), .ZN(n10587) );
  INV_X1 U13435 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U13436 ( .A1(n10587), .A2(n15572), .ZN(n15319) );
  NAND2_X1 U13437 ( .A1(n10428), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10581) );
  MUX2_X1 U13438 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n10581), .S(n10580), .Z(
        n10582) );
  NAND2_X1 U13439 ( .A1(n10582), .A2(n10669), .ZN(n18951) );
  OR2_X1 U13440 ( .A1(n18951), .A2(n10861), .ZN(n10589) );
  INV_X1 U13441 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15594) );
  NAND2_X1 U13442 ( .A1(n10589), .A2(n15594), .ZN(n15316) );
  INV_X1 U13443 ( .A(n13670), .ZN(n10583) );
  OAI21_X1 U13444 ( .B1(n10583), .B2(n10861), .A(n20760), .ZN(n16333) );
  NAND2_X1 U13445 ( .A1(n13622), .A2(n15618), .ZN(n15341) );
  AND2_X1 U13446 ( .A1(n16333), .A2(n15341), .ZN(n15313) );
  AND2_X1 U13447 ( .A1(n10428), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10584) );
  XNOR2_X1 U13448 ( .A(n10585), .B(n10584), .ZN(n18962) );
  NAND2_X1 U13449 ( .A1(n18962), .A2(n10687), .ZN(n10588) );
  INV_X1 U13450 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15560) );
  NAND2_X1 U13451 ( .A1(n10588), .A2(n15560), .ZN(n15315) );
  AND4_X1 U13452 ( .A1(n15319), .A2(n15316), .A3(n15313), .A4(n15315), .ZN(
        n10586) );
  OR2_X1 U13453 ( .A1(n10587), .A2(n15572), .ZN(n15320) );
  NOR2_X1 U13454 ( .A1(n10588), .A2(n15560), .ZN(n15580) );
  NOR2_X1 U13455 ( .A1(n15594), .A2(n10589), .ZN(n15578) );
  NOR2_X1 U13456 ( .A1(n15580), .A2(n15578), .ZN(n15317) );
  AND2_X1 U13457 ( .A1(n15320), .A2(n15317), .ZN(n12204) );
  NAND2_X1 U13458 ( .A1(n12202), .A2(n12204), .ZN(n15303) );
  NAND2_X1 U13459 ( .A1(n10428), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U13460 ( .A1(n9945), .A2(n10592), .ZN(n10593) );
  AND2_X1 U13461 ( .A1(n10627), .A2(n10593), .ZN(n13747) );
  INV_X1 U13462 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15551) );
  NOR2_X1 U13463 ( .A1(n10861), .A2(n15551), .ZN(n10594) );
  AND2_X1 U13464 ( .A1(n13747), .A2(n10594), .ZN(n12203) );
  NAND2_X1 U13465 ( .A1(n13747), .A2(n10687), .ZN(n10595) );
  NAND2_X1 U13466 ( .A1(n10595), .A2(n15551), .ZN(n15304) );
  OAI21_X1 U13467 ( .B1(n15303), .B2(n12203), .A(n15304), .ZN(n10596) );
  INV_X1 U13468 ( .A(n10596), .ZN(n15294) );
  NAND2_X1 U13469 ( .A1(n10428), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10598) );
  INV_X1 U13470 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n20871) );
  NOR2_X1 U13471 ( .A1(n12214), .A2(n20871), .ZN(n10625) );
  INV_X1 U13472 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10619) );
  INV_X1 U13473 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18917) );
  NAND2_X1 U13474 ( .A1(n10619), .A2(n18917), .ZN(n10597) );
  NAND2_X1 U13475 ( .A1(n10428), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10614) );
  AND2_X1 U13476 ( .A1(n10428), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13477 ( .A1(n10428), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10602) );
  MUX2_X1 U13478 ( .A(n10428), .B(n10598), .S(n10599), .Z(n10600) );
  OR2_X2 U13479 ( .A1(n10599), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13480 ( .A1(n10600), .A2(n10640), .ZN(n14991) );
  OR2_X1 U13481 ( .A1(n14991), .A2(n10861), .ZN(n10601) );
  INV_X1 U13482 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13483 ( .A1(n10601), .A2(n10780), .ZN(n15218) );
  INV_X1 U13484 ( .A(n10602), .ZN(n10603) );
  XNOR2_X1 U13485 ( .A(n10604), .B(n10603), .ZN(n18887) );
  NAND2_X1 U13486 ( .A1(n18887), .A2(n10687), .ZN(n10634) );
  INV_X1 U13487 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15236) );
  NAND2_X1 U13488 ( .A1(n10634), .A2(n15236), .ZN(n15228) );
  INV_X1 U13489 ( .A(n10606), .ZN(n10607) );
  XNOR2_X1 U13490 ( .A(n10605), .B(n10607), .ZN(n14126) );
  NAND2_X1 U13491 ( .A1(n14126), .A2(n10687), .ZN(n10608) );
  INV_X1 U13492 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15504) );
  NAND2_X1 U13493 ( .A1(n10608), .A2(n15504), .ZN(n15242) );
  AND2_X1 U13494 ( .A1(n15228), .A2(n15242), .ZN(n15219) );
  AND2_X1 U13495 ( .A1(n10428), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10610) );
  INV_X1 U13496 ( .A(n10669), .ZN(n10646) );
  AOI21_X1 U13497 ( .B1(n10609), .B2(n10610), .A(n10646), .ZN(n10612) );
  NAND2_X1 U13498 ( .A1(n10612), .A2(n10611), .ZN(n14140) );
  OR2_X1 U13499 ( .A1(n14140), .A2(n10861), .ZN(n10613) );
  XNOR2_X1 U13500 ( .A(n10613), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14249) );
  OR2_X1 U13501 ( .A1(n10615), .A2(n10614), .ZN(n10616) );
  NAND2_X1 U13502 ( .A1(n10605), .A2(n10616), .ZN(n18897) );
  INV_X1 U13503 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10771) );
  OAI21_X1 U13504 ( .B1(n18897), .B2(n10861), .A(n10771), .ZN(n15199) );
  NAND2_X1 U13505 ( .A1(n10428), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10618) );
  MUX2_X1 U13506 ( .A(n10618), .B(n10428), .S(n10617), .Z(n10620) );
  NAND2_X1 U13507 ( .A1(n10617), .A2(n10619), .ZN(n10622) );
  NAND2_X1 U13508 ( .A1(n10620), .A2(n10622), .ZN(n13832) );
  OR2_X1 U13509 ( .A1(n13832), .A2(n10861), .ZN(n10636) );
  INV_X1 U13510 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15529) );
  NAND2_X1 U13511 ( .A1(n10636), .A2(n15529), .ZN(n15282) );
  AND2_X1 U13512 ( .A1(n10428), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U13513 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  NAND2_X1 U13514 ( .A1(n10623), .A2(n10609), .ZN(n18907) );
  OR2_X1 U13515 ( .A1(n18907), .A2(n10861), .ZN(n10624) );
  INV_X1 U13516 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U13517 ( .A1(n10624), .A2(n15515), .ZN(n15272) );
  INV_X1 U13518 ( .A(n10625), .ZN(n10626) );
  XNOR2_X1 U13519 ( .A(n10627), .B(n10626), .ZN(n18919) );
  NAND2_X1 U13520 ( .A1(n18919), .A2(n10687), .ZN(n10628) );
  INV_X1 U13521 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15537) );
  NAND2_X1 U13522 ( .A1(n10628), .A2(n15537), .ZN(n15296) );
  AND4_X1 U13523 ( .A1(n15199), .A2(n15282), .A3(n15272), .A4(n15296), .ZN(
        n10629) );
  AND4_X1 U13524 ( .A1(n15218), .A2(n15219), .A3(n14249), .A4(n10629), .ZN(
        n10630) );
  INV_X1 U13525 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15465) );
  NAND3_X1 U13526 ( .A1(n10640), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10428), 
        .ZN(n10631) );
  OAI211_X1 U13527 ( .C1(n10640), .C2(P2_EBX_REG_21__SCAN_IN), .A(n10631), .B(
        n10669), .ZN(n15204) );
  INV_X1 U13528 ( .A(n18897), .ZN(n10632) );
  NAND2_X1 U13529 ( .A1(n10632), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12212) );
  INV_X1 U13530 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15261) );
  OR2_X1 U13531 ( .A1(n14140), .A2(n15261), .ZN(n12210) );
  NAND2_X1 U13532 ( .A1(n12212), .A2(n12210), .ZN(n10633) );
  OR2_X1 U13533 ( .A1(n10634), .A2(n15236), .ZN(n15229) );
  NOR2_X1 U13534 ( .A1(n10861), .A2(n15504), .ZN(n10635) );
  NAND2_X1 U13535 ( .A1(n14126), .A2(n10635), .ZN(n15241) );
  AND2_X1 U13536 ( .A1(n15229), .A2(n15241), .ZN(n15202) );
  INV_X1 U13537 ( .A(n10636), .ZN(n10637) );
  NAND2_X1 U13538 ( .A1(n10637), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15283) );
  OR3_X1 U13539 ( .A1(n18907), .A2(n10861), .A3(n15515), .ZN(n15271) );
  AND2_X1 U13540 ( .A1(n15283), .A2(n15271), .ZN(n12208) );
  NOR2_X1 U13541 ( .A1(n10861), .A2(n15537), .ZN(n10638) );
  NAND2_X1 U13542 ( .A1(n18919), .A2(n10638), .ZN(n15295) );
  OR3_X1 U13543 ( .A1(n14991), .A2(n10861), .A3(n10780), .ZN(n15217) );
  NAND4_X1 U13544 ( .A1(n15202), .A2(n12208), .A3(n15295), .A4(n15217), .ZN(
        n10639) );
  NAND2_X1 U13545 ( .A1(n10428), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10641) );
  OAI21_X1 U13546 ( .B1(n10642), .B2(n10641), .A(n10645), .ZN(n15780) );
  OR2_X1 U13547 ( .A1(n15780), .A2(n10861), .ZN(n10650) );
  INV_X1 U13548 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20823) );
  NAND2_X1 U13549 ( .A1(n10650), .A2(n20823), .ZN(n15446) );
  AND2_X1 U13550 ( .A1(n10428), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10644) );
  INV_X1 U13551 ( .A(n10644), .ZN(n10643) );
  XNOR2_X1 U13552 ( .A(n10645), .B(n10643), .ZN(n16265) );
  NAND2_X1 U13553 ( .A1(n16265), .A2(n10687), .ZN(n15177) );
  INV_X1 U13554 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15176) );
  AND2_X1 U13555 ( .A1(n15177), .A2(n15176), .ZN(n10654) );
  INV_X1 U13556 ( .A(n10667), .ZN(n10649) );
  AND2_X1 U13557 ( .A1(n10428), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U13558 ( .A1(n10649), .A2(n10648), .ZN(n14973) );
  OR2_X1 U13559 ( .A1(n14973), .A2(n10861), .ZN(n10655) );
  INV_X1 U13560 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15422) );
  INV_X1 U13561 ( .A(n10650), .ZN(n10651) );
  NAND2_X1 U13562 ( .A1(n10651), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15447) );
  AOI21_X1 U13563 ( .B1(n15447), .B2(n15176), .A(n15177), .ZN(n10652) );
  NOR2_X1 U13564 ( .A1(n15178), .A2(n10652), .ZN(n10653) );
  NAND2_X1 U13565 ( .A1(n10655), .A2(n15422), .ZN(n15179) );
  INV_X1 U13566 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15026) );
  INV_X1 U13567 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n20956) );
  NAND2_X1 U13568 ( .A1(n10428), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10656) );
  OR2_X1 U13569 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  INV_X1 U13570 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15399) );
  OAI21_X1 U13571 ( .B1(n10659), .B2(n10861), .A(n15399), .ZN(n10661) );
  INV_X1 U13572 ( .A(n10659), .ZN(n16246) );
  NOR2_X1 U13573 ( .A1(n10861), .A2(n15399), .ZN(n10660) );
  INV_X1 U13574 ( .A(n11597), .ZN(n10673) );
  NAND2_X1 U13575 ( .A1(n10428), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10663) );
  INV_X1 U13576 ( .A(n10663), .ZN(n10664) );
  NAND2_X1 U13577 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  NAND2_X1 U13578 ( .A1(n10676), .A2(n10666), .ZN(n12940) );
  INV_X1 U13579 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15382) );
  AND2_X1 U13580 ( .A1(n15139), .A2(n15382), .ZN(n10671) );
  NAND2_X1 U13581 ( .A1(n10428), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10668) );
  MUX2_X1 U13582 ( .A(n10668), .B(P2_EBX_REG_25__SCAN_IN), .S(n10667), .Z(
        n10670) );
  AND2_X1 U13583 ( .A1(n10670), .A2(n10669), .ZN(n16253) );
  NAND2_X1 U13584 ( .A1(n16253), .A2(n10687), .ZN(n10679) );
  INV_X1 U13585 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15406) );
  NAND2_X1 U13586 ( .A1(n10673), .A2(n10672), .ZN(n10678) );
  INV_X1 U13587 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10674) );
  NOR2_X1 U13588 ( .A1(n12214), .A2(n10674), .ZN(n10675) );
  AND2_X1 U13589 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NOR2_X1 U13590 ( .A1(n10685), .A2(n10677), .ZN(n14959) );
  AND2_X1 U13591 ( .A1(n14959), .A2(n10687), .ZN(n15143) );
  INV_X1 U13592 ( .A(n10679), .ZN(n10680) );
  NAND2_X1 U13593 ( .A1(n10680), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15165) );
  NAND2_X1 U13594 ( .A1(n10428), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10684) );
  INV_X1 U13595 ( .A(n10684), .ZN(n10682) );
  XNOR2_X1 U13596 ( .A(n10685), .B(n10682), .ZN(n12830) );
  NAND2_X1 U13597 ( .A1(n12830), .A2(n10687), .ZN(n10683) );
  INV_X1 U13598 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14289) );
  NAND2_X1 U13599 ( .A1(n10683), .A2(n14289), .ZN(n14274) );
  NAND2_X1 U13600 ( .A1(n10685), .A2(n10684), .ZN(n10693) );
  NAND2_X1 U13601 ( .A1(n10428), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10686) );
  XNOR2_X1 U13602 ( .A(n10693), .B(n10686), .ZN(n12917) );
  AOI21_X1 U13603 ( .B1(n12917), .B2(n10687), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15126) );
  INV_X1 U13604 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12847) );
  NOR2_X1 U13605 ( .A1(n10861), .A2(n12847), .ZN(n10688) );
  NAND2_X1 U13606 ( .A1(n12917), .A2(n10688), .ZN(n15127) );
  INV_X1 U13607 ( .A(n15127), .ZN(n10691) );
  INV_X1 U13608 ( .A(n12830), .ZN(n10689) );
  NOR2_X1 U13609 ( .A1(n10693), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10694) );
  MUX2_X1 U13610 ( .A(n10695), .B(n10694), .S(n10428), .Z(n14271) );
  NAND2_X1 U13611 ( .A1(n14271), .A2(n10687), .ZN(n10696) );
  INV_X1 U13612 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12744) );
  XNOR2_X1 U13613 ( .A(n10696), .B(n12744), .ZN(n10697) );
  INV_X1 U13614 ( .A(n10699), .ZN(n12124) );
  AND2_X1 U13615 ( .A1(n15870), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10700) );
  INV_X1 U13616 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13486) );
  NAND2_X1 U13617 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13486), .ZN(
        n10702) );
  XNOR2_X1 U13618 ( .A(n12125), .B(n10704), .ZN(n12118) );
  NAND2_X1 U13619 ( .A1(n12118), .A2(n10706), .ZN(n10705) );
  NAND2_X1 U13620 ( .A1(n12137), .A2(n10705), .ZN(n13476) );
  AOI21_X1 U13621 ( .B1(n12124), .B2(n10706), .A(n13476), .ZN(n10709) );
  INV_X1 U13622 ( .A(n10384), .ZN(n10707) );
  NOR2_X1 U13623 ( .A1(n13454), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13091) );
  NAND2_X1 U13624 ( .A1(n10707), .A2(n13091), .ZN(n10708) );
  INV_X1 U13625 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18865) );
  NAND2_X1 U13626 ( .A1(n10708), .A2(n18865), .ZN(n19886) );
  MUX2_X1 U13627 ( .A(n10709), .B(n19886), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n15866) );
  INV_X1 U13628 ( .A(n12125), .ZN(n10711) );
  OAI21_X1 U13629 ( .B1(n10712), .B2(n10711), .A(n10710), .ZN(n10715) );
  AND2_X1 U13630 ( .A1(n12121), .A2(n10713), .ZN(n10714) );
  AOI21_X1 U13631 ( .B1(n10715), .B2(n10714), .A(n10822), .ZN(n10716) );
  MUX2_X1 U13632 ( .A(n15866), .B(n10716), .S(n9761), .Z(n19895) );
  NAND2_X1 U13633 ( .A1(n10243), .A2(n18862), .ZN(n10718) );
  NOR2_X1 U13634 ( .A1(n10717), .A2(n10718), .ZN(n10719) );
  NAND2_X1 U13635 ( .A1(n19895), .A2(n10719), .ZN(n18864) );
  NOR2_X1 U13636 ( .A1(n18864), .A2(n9761), .ZN(n15335) );
  NAND2_X1 U13637 ( .A1(n12865), .A2(n16346), .ZN(n10879) );
  NAND2_X1 U13638 ( .A1(n10721), .A2(n10720), .ZN(n10725) );
  INV_X1 U13639 ( .A(n10722), .ZN(n10723) );
  INV_X1 U13640 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12251) );
  OR2_X1 U13641 ( .A1(n10286), .A2(n14006), .ZN(n10728) );
  INV_X2 U13642 ( .A(n10726), .ZN(n10814) );
  AOI22_X1 U13643 ( .A1(n10814), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10727) );
  OAI211_X1 U13644 ( .C1(n10785), .C2(n12251), .A(n10728), .B(n10727), .ZN(
        n13679) );
  INV_X1 U13645 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10731) );
  OR2_X1 U13646 ( .A1(n10286), .A2(n9891), .ZN(n10730) );
  AOI22_X1 U13647 ( .A1(n10814), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10729) );
  OAI211_X1 U13648 ( .C1(n10785), .C2(n10731), .A(n10730), .B(n10729), .ZN(
        n13249) );
  INV_X1 U13649 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U13650 ( .A1(n10814), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10733) );
  NAND2_X1 U13651 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10732) );
  OAI211_X1 U13652 ( .C1(n10734), .C2(n10785), .A(n10733), .B(n10732), .ZN(
        n10735) );
  AOI21_X1 U13653 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10735), .ZN(n13263) );
  INV_X1 U13654 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13655 ( .A1(n10814), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13656 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10737) );
  OAI211_X1 U13657 ( .C1(n10739), .C2(n10785), .A(n10738), .B(n10737), .ZN(
        n10740) );
  AOI21_X1 U13658 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10740), .ZN(n13297) );
  INV_X1 U13659 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U13660 ( .A1(n10814), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13661 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10741) );
  OAI211_X1 U13662 ( .C1(n13663), .C2(n10785), .A(n10742), .B(n10741), .ZN(
        n10743) );
  AOI21_X1 U13663 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10743), .ZN(n13658) );
  INV_X1 U13664 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15329) );
  OR2_X1 U13665 ( .A1(n10818), .A2(n15560), .ZN(n10746) );
  AOI22_X1 U13666 ( .A1(n10814), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10745) );
  OAI211_X1 U13667 ( .C1(n10785), .C2(n15329), .A(n10746), .B(n10745), .ZN(
        n13307) );
  INV_X1 U13668 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U13669 ( .A1(n10814), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10747) );
  OAI211_X1 U13671 ( .C1(n12298), .C2(n10785), .A(n10748), .B(n10747), .ZN(
        n10749) );
  AOI21_X1 U13672 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10749), .ZN(n15586) );
  INV_X1 U13673 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19811) );
  NAND2_X1 U13674 ( .A1(n10814), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13675 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10752) );
  OAI211_X1 U13676 ( .C1(n19811), .C2(n10785), .A(n10753), .B(n10752), .ZN(
        n10754) );
  AOI21_X1 U13677 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10754), .ZN(n13723) );
  INV_X1 U13678 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10757) );
  OR2_X1 U13679 ( .A1(n10818), .A2(n15551), .ZN(n10756) );
  AOI22_X1 U13680 ( .A1(n10814), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10755) );
  OAI211_X1 U13681 ( .C1(n10785), .C2(n10757), .A(n10756), .B(n10755), .ZN(
        n13551) );
  INV_X1 U13682 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15298) );
  OR2_X1 U13683 ( .A1(n10818), .A2(n15537), .ZN(n10759) );
  AOI22_X1 U13684 ( .A1(n10814), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10758) );
  OAI211_X1 U13685 ( .C1(n10785), .C2(n15298), .A(n10759), .B(n10758), .ZN(
        n13760) );
  NAND2_X1 U13686 ( .A1(n13549), .A2(n13760), .ZN(n13759) );
  INV_X1 U13687 ( .A(n13759), .ZN(n10764) );
  INV_X1 U13688 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19815) );
  NAND2_X1 U13689 ( .A1(n10814), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10761) );
  NAND2_X1 U13690 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10760) );
  OAI211_X1 U13691 ( .C1(n19815), .C2(n10785), .A(n10761), .B(n10760), .ZN(
        n10762) );
  AOI21_X1 U13692 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10762), .ZN(n13824) );
  INV_X1 U13693 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19817) );
  NAND2_X1 U13694 ( .A1(n10814), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U13695 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10765) );
  OAI211_X1 U13696 ( .C1(n19817), .C2(n10785), .A(n10766), .B(n10765), .ZN(
        n10767) );
  AOI21_X1 U13697 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10767), .ZN(n13939) );
  INV_X1 U13698 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U13699 ( .A1(n10814), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U13700 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10768) );
  OAI211_X1 U13701 ( .C1(n14142), .C2(n10785), .A(n10769), .B(n10768), .ZN(
        n10770) );
  AOI21_X1 U13702 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10770), .ZN(n14136) );
  INV_X1 U13703 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19819) );
  OR2_X1 U13704 ( .A1(n10818), .A2(n10771), .ZN(n10773) );
  AOI22_X1 U13705 ( .A1(n10814), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10772) );
  OAI211_X1 U13706 ( .C1(n10785), .C2(n19819), .A(n10773), .B(n10772), .ZN(
        n12372) );
  INV_X1 U13707 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U13708 ( .A1(n10814), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10775) );
  NAND2_X1 U13709 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10774) );
  OAI211_X1 U13710 ( .C1(n15245), .C2(n10785), .A(n10775), .B(n10774), .ZN(
        n10776) );
  AOI21_X1 U13711 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10776), .ZN(n14120) );
  INV_X1 U13712 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19822) );
  NAND2_X1 U13713 ( .A1(n10814), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U13714 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10777) );
  OAI211_X1 U13715 ( .C1(n19822), .C2(n10785), .A(n10778), .B(n10777), .ZN(
        n10779) );
  AOI21_X1 U13716 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10779), .ZN(n15051) );
  INV_X1 U13717 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19824) );
  OR2_X1 U13718 ( .A1(n10818), .A2(n10780), .ZN(n10782) );
  AOI22_X1 U13719 ( .A1(n10814), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10781) );
  OAI211_X1 U13720 ( .C1(n10785), .C2(n19824), .A(n10782), .B(n10781), .ZN(
        n14986) );
  INV_X1 U13721 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19826) );
  OR2_X1 U13722 ( .A1(n10818), .A2(n15465), .ZN(n10784) );
  AOI22_X1 U13723 ( .A1(n10814), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10783) );
  OAI211_X1 U13724 ( .C1(n10785), .C2(n19826), .A(n10784), .B(n10783), .ZN(
        n12957) );
  INV_X1 U13725 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U13726 ( .A1(n10814), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13727 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10786) );
  OAI211_X1 U13728 ( .C1(n10788), .C2(n10785), .A(n10787), .B(n10786), .ZN(
        n10789) );
  AOI21_X1 U13729 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10789), .ZN(n15449) );
  INV_X1 U13730 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n10792) );
  NAND2_X1 U13731 ( .A1(n10814), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10791) );
  NAND2_X1 U13732 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10790) );
  OAI211_X1 U13733 ( .C1(n10792), .C2(n10785), .A(n10791), .B(n10790), .ZN(
        n10793) );
  AOI21_X1 U13734 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10793), .ZN(n15036) );
  INV_X1 U13735 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15183) );
  OR2_X1 U13736 ( .A1(n10818), .A2(n15422), .ZN(n10795) );
  AOI22_X1 U13737 ( .A1(n10814), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10794) );
  OAI211_X1 U13738 ( .C1(n10785), .C2(n15183), .A(n10795), .B(n10794), .ZN(
        n14963) );
  INV_X1 U13739 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19831) );
  OR2_X1 U13740 ( .A1(n10818), .A2(n15406), .ZN(n10797) );
  AOI22_X1 U13741 ( .A1(n10814), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10796) );
  OAI211_X1 U13742 ( .C1(n10785), .C2(n19831), .A(n10797), .B(n10796), .ZN(
        n15024) );
  NAND2_X1 U13743 ( .A1(n14962), .A2(n15024), .ZN(n15016) );
  INV_X1 U13744 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19833) );
  NAND2_X1 U13745 ( .A1(n10814), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13746 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10798) );
  OAI211_X1 U13747 ( .C1(n19833), .C2(n10785), .A(n10799), .B(n10798), .ZN(
        n10800) );
  AOI21_X1 U13748 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10800), .ZN(n15018) );
  INV_X1 U13749 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19836) );
  NAND2_X1 U13750 ( .A1(n10814), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U13751 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10801) );
  OAI211_X1 U13752 ( .C1(n19836), .C2(n10785), .A(n10802), .B(n10801), .ZN(
        n10803) );
  AOI21_X1 U13753 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10803), .ZN(n11592) );
  INV_X1 U13754 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15146) );
  NAND2_X1 U13755 ( .A1(n10814), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10806) );
  NAND2_X1 U13756 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10805) );
  OAI211_X1 U13757 ( .C1(n15146), .C2(n10785), .A(n10806), .B(n10805), .ZN(
        n10807) );
  AOI21_X1 U13758 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10807), .ZN(n14948) );
  INV_X1 U13759 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19838) );
  OR2_X1 U13760 ( .A1(n10818), .A2(n14289), .ZN(n10809) );
  AOI22_X1 U13761 ( .A1(n10814), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10808) );
  OAI211_X1 U13762 ( .C1(n10785), .C2(n19838), .A(n10809), .B(n10808), .ZN(
        n12793) );
  INV_X1 U13763 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15131) );
  NAND2_X1 U13764 ( .A1(n10814), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10811) );
  NAND2_X1 U13765 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10810) );
  OAI211_X1 U13766 ( .C1(n15131), .C2(n10785), .A(n10811), .B(n10810), .ZN(
        n10812) );
  AOI21_X1 U13767 ( .B1(n10813), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10812), .ZN(n12907) );
  AOI22_X1 U13768 ( .A1(n10814), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10817) );
  NAND2_X1 U13769 ( .A1(n10815), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10816) );
  OAI211_X1 U13770 ( .C1(n10818), .C2(n12744), .A(n10817), .B(n10816), .ZN(
        n10819) );
  INV_X1 U13771 ( .A(n10819), .ZN(n10820) );
  XNOR2_X1 U13772 ( .A(n9966), .B(n10820), .ZN(n16278) );
  NOR2_X1 U13773 ( .A1(n19581), .A2(n19666), .ZN(n19869) );
  NOR2_X1 U13774 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n10821) );
  NAND2_X1 U13775 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n16380), .ZN(n13497) );
  NOR2_X1 U13776 ( .A1(n13837), .A2(n19723), .ZN(n19887) );
  INV_X1 U13777 ( .A(n19887), .ZN(n16368) );
  NAND2_X1 U13778 ( .A1(n13837), .A2(n19723), .ZN(n16377) );
  NAND2_X1 U13779 ( .A1(n16380), .A2(n16377), .ZN(n14939) );
  INV_X1 U13780 ( .A(n14939), .ZN(n10823) );
  NAND2_X1 U13781 ( .A1(n16368), .A2(n10823), .ZN(n10824) );
  INV_X1 U13782 ( .A(n15652), .ZN(n19176) );
  NOR2_X1 U13783 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13840) );
  INV_X1 U13784 ( .A(n13840), .ZN(n19854) );
  NAND2_X1 U13785 ( .A1(n19581), .A2(n19854), .ZN(n19872) );
  NAND2_X1 U13786 ( .A1(n19872), .A2(n16380), .ZN(n10826) );
  NAND2_X1 U13787 ( .A1(n13840), .A2(n19723), .ZN(n14930) );
  INV_X1 U13788 ( .A(n14930), .ZN(n10827) );
  NAND2_X1 U13789 ( .A1(n16380), .A2(n10827), .ZN(n18933) );
  INV_X1 U13790 ( .A(n18985), .ZN(n18970) );
  INV_X1 U13791 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12842) );
  NOR2_X1 U13792 ( .A1(n18970), .A2(n12842), .ZN(n12857) );
  INV_X1 U13793 ( .A(n13208), .ZN(n13104) );
  NAND2_X1 U13794 ( .A1(n19666), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13795 ( .A1(n13104), .A2(n10828), .ZN(n13101) );
  AND2_X1 U13796 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U13797 ( .A1(n12758), .A2(n10830), .ZN(n12756) );
  INV_X1 U13798 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12766) );
  INV_X1 U13799 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15287) );
  INV_X1 U13800 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15234) );
  INV_X1 U13801 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15246) );
  NOR2_X1 U13802 ( .A1(n15234), .A2(n15246), .ZN(n10831) );
  INV_X1 U13803 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20983) );
  INV_X1 U13804 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U13805 ( .A1(n12777), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12778) );
  NAND2_X1 U13806 ( .A1(n12779), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12782) );
  INV_X1 U13807 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15168) );
  NAND2_X1 U13808 ( .A1(n12784), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11588) );
  INV_X1 U13809 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12941) );
  INV_X1 U13810 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10834) );
  XNOR2_X1 U13811 ( .A(n10835), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12745) );
  NOR2_X1 U13812 ( .A1(n19172), .A2(n12745), .ZN(n10836) );
  AOI211_X1 U13813 ( .C1(n16322), .C2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12857), .B(n10836), .ZN(n10837) );
  NAND2_X1 U13814 ( .A1(n13099), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13098) );
  INV_X1 U13815 ( .A(n13098), .ZN(n10840) );
  INV_X1 U13816 ( .A(n12228), .ZN(n10839) );
  NAND2_X1 U13817 ( .A1(n10840), .A2(n10839), .ZN(n10842) );
  AND2_X1 U13818 ( .A1(n13097), .A2(n13099), .ZN(n10841) );
  XOR2_X1 U13819 ( .A(n12228), .B(n10841), .Z(n12973) );
  NAND2_X1 U13820 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12973), .ZN(
        n12972) );
  NAND2_X1 U13821 ( .A1(n10842), .A2(n12972), .ZN(n10845) );
  XOR2_X1 U13822 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10845), .Z(
        n14231) );
  XNOR2_X1 U13823 ( .A(n10844), .B(n10843), .ZN(n14230) );
  NAND2_X1 U13824 ( .A1(n14231), .A2(n14230), .ZN(n10847) );
  NAND2_X1 U13825 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10845), .ZN(
        n10846) );
  NAND2_X1 U13826 ( .A1(n10847), .A2(n10846), .ZN(n10848) );
  XNOR2_X1 U13827 ( .A(n10848), .B(n10449), .ZN(n13798) );
  NAND2_X1 U13828 ( .A1(n10848), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10849) );
  INV_X1 U13829 ( .A(n12248), .ZN(n10850) );
  NAND2_X1 U13830 ( .A1(n10857), .A2(n13995), .ZN(n10852) );
  NAND2_X1 U13831 ( .A1(n10856), .A2(n13995), .ZN(n10858) );
  NAND2_X1 U13832 ( .A1(n10858), .A2(n10857), .ZN(n10859) );
  NAND2_X1 U13833 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  NAND2_X1 U13834 ( .A1(n10868), .A2(n10863), .ZN(n10864) );
  INV_X1 U13835 ( .A(n10864), .ZN(n10865) );
  INV_X1 U13836 ( .A(n10868), .ZN(n10869) );
  NAND2_X1 U13837 ( .A1(n10869), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10870) );
  NAND2_X2 U13838 ( .A1(n16337), .A2(n10870), .ZN(n12167) );
  AND2_X1 U13839 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15568) );
  AND2_X1 U13840 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15539) );
  AND2_X1 U13841 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10871) );
  NAND3_X1 U13842 ( .A1(n15568), .A2(n15539), .A3(n10871), .ZN(n12189) );
  AND2_X1 U13843 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U13844 ( .A1(n12199), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12846) );
  NOR2_X1 U13845 ( .A1(n12189), .A2(n12846), .ZN(n12850) );
  NAND2_X1 U13846 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U13847 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15430) );
  NAND2_X1 U13848 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14277) );
  OR2_X1 U13849 ( .A1(n14277), .A2(n14289), .ZN(n10873) );
  NAND2_X1 U13850 ( .A1(n15123), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10874) );
  XNOR2_X2 U13851 ( .A(n10874), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12864) );
  INV_X1 U13852 ( .A(n18864), .ZN(n10875) );
  NAND2_X1 U13853 ( .A1(n10875), .A2(n9761), .ZN(n19173) );
  NAND2_X1 U13854 ( .A1(n12864), .A2(n10876), .ZN(n10877) );
  NAND3_X1 U13855 ( .A1(n10879), .A2(n10878), .A3(n10877), .ZN(P2_U2983) );
  NOR2_X4 U13856 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13530) );
  NOR2_X4 U13857 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10887) );
  AND2_X2 U13858 ( .A1(n13530), .A2(n10887), .ZN(n11133) );
  AOI22_X1 U13859 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10885) );
  INV_X1 U13860 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11112) );
  AND2_X4 U13861 ( .A1(n13508), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13513) );
  AND2_X4 U13862 ( .A1(n10880), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13503) );
  AND2_X4 U13863 ( .A1(n13503), .A2(n13502), .ZN(n11080) );
  AOI22_X1 U13864 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10884) );
  AND2_X4 U13865 ( .A1(n10881), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10888) );
  AND2_X4 U13866 ( .A1(n10886), .A2(n10889), .ZN(n11131) );
  AOI22_X1 U13867 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10883) );
  AND2_X4 U13868 ( .A1(n13530), .A2(n10889), .ZN(n11181) );
  AOI22_X1 U13869 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13870 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13871 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13872 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13873 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13874 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9766), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13875 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13876 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13877 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10895) );
  AND4_X2 U13878 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10904) );
  AOI22_X1 U13879 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13880 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11923), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13881 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9741), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13882 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U13883 ( .A1(n10945), .A2(n11008), .ZN(n11027) );
  AOI22_X1 U13884 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9691), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13885 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13886 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13887 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13888 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13889 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11133), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13890 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11079), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10909) );
  NAND2_X1 U13891 ( .A1(n11027), .A2(n11010), .ZN(n10944) );
  AOI22_X1 U13892 ( .A1(n9772), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9741), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13893 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13894 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13895 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13896 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13897 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U13898 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10927) );
  NAND2_X1 U13899 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10926) );
  NAND2_X1 U13900 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10925) );
  NAND2_X1 U13901 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10924) );
  NAND2_X1 U13902 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10931) );
  NAND2_X1 U13903 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10930) );
  NAND2_X1 U13904 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10929) );
  NAND2_X1 U13905 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10928) );
  NAND2_X1 U13906 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U13907 ( .A1(n9772), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10934) );
  NAND2_X1 U13908 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10933) );
  NAND2_X1 U13909 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10932) );
  NAND2_X1 U13910 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10939) );
  NAND2_X1 U13911 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10938) );
  NAND2_X1 U13912 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10937) );
  NAND2_X1 U13913 ( .A1(n11081), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10936) );
  AND2_X2 U13914 ( .A1(n11144), .A2(n11006), .ZN(n10960) );
  AOI22_X1 U13915 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13916 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13917 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13918 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10946) );
  AND2_X1 U13919 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  AOI22_X1 U13920 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12059), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U13921 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U13922 ( .A1(n9772), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9741), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U13923 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U13924 ( .A1(n10127), .A2(n11513), .ZN(n10956) );
  OAI21_X1 U13925 ( .B1(n10960), .B2(n11513), .A(n10956), .ZN(n10957) );
  INV_X1 U13926 ( .A(n10957), .ZN(n10958) );
  NAND2_X1 U13927 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10964) );
  NAND2_X1 U13928 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10963) );
  NAND2_X1 U13929 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10962) );
  NAND2_X1 U13930 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10961) );
  NAND2_X1 U13931 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10968) );
  NAND2_X1 U13932 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10967) );
  NAND2_X1 U13933 ( .A1(n9772), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10966) );
  NAND2_X1 U13934 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10965) );
  NAND2_X1 U13935 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10974) );
  NAND2_X1 U13936 ( .A1(n11771), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10973) );
  NAND2_X1 U13937 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10972) );
  NAND2_X1 U13938 ( .A1(n11087), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U13939 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10978) );
  NAND2_X1 U13940 ( .A1(n9766), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10977) );
  NAND2_X1 U13941 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10976) );
  NAND2_X1 U13942 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10975) );
  NAND2_X1 U13943 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10987) );
  NAND2_X1 U13944 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10986) );
  NAND2_X1 U13945 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10985) );
  NAND2_X1 U13946 ( .A1(n9772), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U13947 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10991) );
  NAND2_X1 U13948 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10990) );
  NAND2_X1 U13949 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10989) );
  NAND3_X1 U13950 ( .A1(n10989), .A2(n10990), .A3(n10991), .ZN(n10992) );
  AOI21_X2 U13951 ( .B1(n11771), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n10992), .ZN(n11003) );
  NAND2_X1 U13952 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10996) );
  NAND2_X1 U13953 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10995) );
  NAND2_X1 U13954 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10994) );
  NAND2_X1 U13955 ( .A1(n9766), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10993) );
  NAND2_X1 U13956 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11000) );
  NAND2_X1 U13957 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10999) );
  NAND2_X1 U13958 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10998) );
  NAND2_X1 U13959 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10997) );
  NAND4_X4 U13960 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11022) );
  INV_X2 U13961 ( .A(n11144), .ZN(n13544) );
  BUF_X4 U13962 ( .A(n11020), .Z(n11328) );
  NAND2_X1 U13963 ( .A1(n11376), .A2(n13909), .ZN(n12389) );
  NAND2_X1 U13964 ( .A1(n12386), .A2(n12389), .ZN(n11397) );
  NAND2_X1 U13965 ( .A1(n13131), .A2(n11008), .ZN(n13113) );
  NAND2_X1 U13966 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20607) );
  OAI21_X1 U13967 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20607), .ZN(n11377) );
  AND2_X2 U13968 ( .A1(n11014), .A2(n13544), .ZN(n12890) );
  INV_X1 U13969 ( .A(n11011), .ZN(n11394) );
  OAI21_X1 U13970 ( .B1(n9729), .B2(n11014), .A(n13911), .ZN(n11030) );
  NAND2_X1 U13971 ( .A1(n13544), .A2(n11016), .ZN(n11017) );
  NAND2_X1 U13972 ( .A1(n11369), .A2(n11035), .ZN(n11039) );
  NAND2_X1 U13973 ( .A1(n11369), .A2(n11328), .ZN(n11018) );
  NAND2_X1 U13974 ( .A1(n11018), .A2(n20677), .ZN(n11019) );
  NAND2_X1 U13975 ( .A1(n11039), .A2(n11019), .ZN(n11512) );
  INV_X1 U13976 ( .A(n11145), .ZN(n11021) );
  INV_X1 U13977 ( .A(n11374), .ZN(n11023) );
  NAND2_X1 U13978 ( .A1(n11401), .A2(n11023), .ZN(n11506) );
  INV_X1 U13979 ( .A(n11400), .ZN(n11024) );
  NAND2_X1 U13980 ( .A1(n11025), .A2(n11328), .ZN(n11026) );
  AND2_X2 U13981 ( .A1(n11514), .A2(n11026), .ZN(n13498) );
  NAND2_X1 U13982 ( .A1(n13911), .A2(n11022), .ZN(n13908) );
  NAND2_X1 U13983 ( .A1(n11039), .A2(n14257), .ZN(n11028) );
  NAND4_X1 U13984 ( .A1(n11030), .A2(n11512), .A3(n11029), .A4(n11028), .ZN(
        n11031) );
  NAND2_X1 U13985 ( .A1(n11031), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U13986 ( .A1(n11117), .A2(n9724), .ZN(n11034) );
  NOR2_X1 U13987 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U13988 ( .A1(n14262), .A2(n16236), .ZN(n12107) );
  MUX2_X1 U13989 ( .A(n12107), .B(n20589), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11033) );
  NAND2_X1 U13990 ( .A1(n11014), .A2(n9725), .ZN(n11516) );
  AND4_X1 U13991 ( .A1(n11516), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14262), 
        .A4(n13908), .ZN(n11038) );
  INV_X1 U13992 ( .A(n11035), .ZN(n11036) );
  NAND2_X1 U13993 ( .A1(n11036), .A2(n11502), .ZN(n11037) );
  NAND3_X1 U13994 ( .A1(n11039), .A2(n11022), .A3(n14257), .ZN(n11042) );
  OAI21_X1 U13995 ( .B1(n13904), .B2(n11040), .A(n9729), .ZN(n11041) );
  NAND3_X1 U13996 ( .A1(n10122), .A2(n11042), .A3(n11041), .ZN(n11102) );
  INV_X1 U13997 ( .A(n11102), .ZN(n11043) );
  NAND2_X1 U13998 ( .A1(n11624), .A2(n16236), .ZN(n11072) );
  AOI22_X1 U13999 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11180), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U14000 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14001 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11047) );
  BUF_X1 U14002 ( .A(n11181), .Z(n11045) );
  AOI22_X1 U14003 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11046) );
  NAND4_X1 U14004 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n11058) );
  AOI22_X1 U14005 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U14006 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14007 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14008 ( .A1(n9770), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11053) );
  NAND4_X1 U14009 ( .A1(n11056), .A2(n11055), .A3(n11054), .A4(n11053), .ZN(
        n11057) );
  AOI22_X1 U14010 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U14011 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U14012 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14013 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11087), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11059) );
  NAND4_X1 U14014 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11069) );
  AOI22_X1 U14015 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9770), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14017 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14018 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14019 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11064) );
  NAND4_X1 U14020 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11068) );
  XNOR2_X1 U14021 ( .A(n11290), .B(n11156), .ZN(n11070) );
  NAND2_X1 U14022 ( .A1(n11070), .A2(n11107), .ZN(n11071) );
  NAND2_X1 U14023 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11076) );
  NAND2_X1 U14024 ( .A1(n13911), .A2(n11156), .ZN(n11073) );
  OAI211_X1 U14025 ( .C1(n11290), .C2(n13574), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n11073), .ZN(n11074) );
  INV_X1 U14026 ( .A(n11074), .ZN(n11075) );
  NAND2_X1 U14027 ( .A1(n11150), .A2(n11151), .ZN(n11078) );
  NAND2_X1 U14028 ( .A1(n11107), .A2(n11286), .ZN(n11077) );
  NAND2_X1 U14029 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11095) );
  NOR2_X1 U14030 ( .A1(n11328), .A2(n16236), .ZN(n11141) );
  AOI22_X1 U14031 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14032 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14033 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14034 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11082) );
  NAND4_X1 U14035 ( .A1(n11085), .A2(n11084), .A3(n11083), .A4(n11082), .ZN(
        n11093) );
  AOI22_X1 U14036 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14037 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14038 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9703), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14039 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11088) );
  NAND4_X1 U14040 ( .A1(n11091), .A2(n11090), .A3(n11089), .A4(n11088), .ZN(
        n11092) );
  NAND2_X1 U14041 ( .A1(n11141), .A2(n11155), .ZN(n11094) );
  OAI211_X1 U14042 ( .C1(n11287), .C2(n11286), .A(n11095), .B(n11094), .ZN(
        n11096) );
  NAND2_X1 U14043 ( .A1(n11097), .A2(n11096), .ZN(n11098) );
  NAND2_X1 U14044 ( .A1(n20524), .A2(n20317), .ZN(n20431) );
  NAND2_X1 U14045 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20520) );
  NAND2_X1 U14046 ( .A1(n20431), .A2(n20520), .ZN(n20353) );
  OR2_X1 U14047 ( .A1(n20589), .A2(n20524), .ZN(n11114) );
  OAI21_X1 U14048 ( .B1(n12107), .B2(n20353), .A(n11114), .ZN(n11099) );
  INV_X1 U14049 ( .A(n11099), .ZN(n11100) );
  INV_X1 U14050 ( .A(n13605), .ZN(n11106) );
  INV_X1 U14051 ( .A(n11104), .ZN(n11105) );
  NAND2_X1 U14052 ( .A1(n11124), .A2(n13562), .ZN(n13948) );
  NAND2_X1 U14053 ( .A1(n11107), .A2(n11155), .ZN(n11108) );
  INV_X1 U14054 ( .A(n11614), .ZN(n11109) );
  NAND2_X1 U14055 ( .A1(n11617), .A2(n11111), .ZN(n11168) );
  INV_X1 U14056 ( .A(n11101), .ZN(n11116) );
  NAND2_X1 U14057 ( .A1(n11114), .A2(n11113), .ZN(n11115) );
  NAND2_X1 U14058 ( .A1(n11116), .A2(n11115), .ZN(n11122) );
  NAND2_X1 U14059 ( .A1(n11124), .A2(n11122), .ZN(n11120) );
  NOR2_X1 U14060 ( .A1(n20589), .A2(n15810), .ZN(n11118) );
  INV_X1 U14061 ( .A(n12107), .ZN(n11172) );
  XNOR2_X1 U14062 ( .A(n20520), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13952) );
  NAND2_X1 U14063 ( .A1(n11172), .A2(n13952), .ZN(n11121) );
  NAND2_X1 U14064 ( .A1(n11123), .A2(n11121), .ZN(n11119) );
  NAND4_X1 U14065 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .ZN(
        n11125) );
  AOI22_X1 U14066 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14067 ( .A1(n11050), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14068 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14069 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11127) );
  NAND4_X1 U14070 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11139) );
  AOI22_X1 U14071 ( .A1(n12059), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U14072 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11136) );
  AOI22_X1 U14073 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11135) );
  AOI22_X1 U14074 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11134) );
  NAND4_X1 U14075 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11138) );
  OAI22_X2 U14076 ( .A1(n13519), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11192), 
        .B2(n11287), .ZN(n11143) );
  AOI22_X1 U14077 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11141), .B2(n11140), .ZN(n11142) );
  XNOR2_X2 U14078 ( .A(n11143), .B(n11142), .ZN(n11166) );
  XNOR2_X1 U14079 ( .A(n11168), .B(n11166), .ZN(n11609) );
  NAND2_X1 U14080 ( .A1(n11609), .A2(n11313), .ZN(n11149) );
  NAND2_X1 U14081 ( .A1(n11155), .A2(n11156), .ZN(n11193) );
  XNOR2_X1 U14082 ( .A(n11193), .B(n11192), .ZN(n11147) );
  NAND2_X1 U14083 ( .A1(n13911), .A2(n11145), .ZN(n11152) );
  INV_X1 U14084 ( .A(n11152), .ZN(n11146) );
  AOI21_X1 U14085 ( .B1(n11147), .B2(n11502), .A(n11146), .ZN(n11148) );
  NAND2_X1 U14086 ( .A1(n11149), .A2(n11148), .ZN(n13421) );
  INV_X1 U14087 ( .A(n11313), .ZN(n11239) );
  OAI21_X1 U14088 ( .B1(n20677), .B2(n11156), .A(n11152), .ZN(n11153) );
  INV_X1 U14089 ( .A(n11153), .ZN(n11154) );
  OAI21_X1 U14090 ( .B1(n11156), .B2(n11155), .A(n11193), .ZN(n11157) );
  OAI211_X1 U14091 ( .C1(n11157), .C2(n20677), .A(n11374), .B(n11144), .ZN(
        n11158) );
  INV_X1 U14092 ( .A(n11158), .ZN(n11159) );
  INV_X1 U14093 ( .A(n11160), .ZN(n11162) );
  NAND2_X1 U14094 ( .A1(n11162), .A2(n11161), .ZN(n11163) );
  INV_X1 U14095 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20107) );
  NAND2_X1 U14096 ( .A1(n13421), .A2(n13422), .ZN(n13420) );
  NAND2_X1 U14097 ( .A1(n11164), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11165) );
  INV_X1 U14098 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11415) );
  INV_X1 U14099 ( .A(n11166), .ZN(n11167) );
  NOR2_X2 U14100 ( .A1(n11168), .A2(n11167), .ZN(n11190) );
  NAND2_X1 U14101 ( .A1(n9726), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11174) );
  NOR2_X1 U14102 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15810), .ZN(
        n20288) );
  INV_X1 U14103 ( .A(n20520), .ZN(n20391) );
  NAND2_X1 U14104 ( .A1(n20288), .A2(n20391), .ZN(n13702) );
  OAI21_X1 U14105 ( .B1(n20520), .B2(n15810), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U14106 ( .A1(n13702), .A2(n11170), .ZN(n20127) );
  INV_X1 U14107 ( .A(n20589), .ZN(n11171) );
  AOI22_X1 U14108 ( .A1(n20127), .A2(n11172), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11171), .ZN(n11173) );
  AOI22_X1 U14109 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14110 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14111 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14112 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11176) );
  NAND4_X1 U14113 ( .A1(n11179), .A2(n11178), .A3(n11177), .A4(n11176), .ZN(
        n11187) );
  AOI22_X1 U14114 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14115 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14116 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14117 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11182) );
  NAND4_X1 U14118 ( .A1(n11185), .A2(n11184), .A3(n11183), .A4(n11182), .ZN(
        n11186) );
  AOI22_X1 U14119 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11323), .B2(n11241), .ZN(n11188) );
  NAND2_X1 U14120 ( .A1(n11190), .A2(n13587), .ZN(n11215) );
  OR2_X1 U14121 ( .A1(n20117), .A2(n11239), .ZN(n11197) );
  NAND2_X1 U14122 ( .A1(n11193), .A2(n11192), .ZN(n11243) );
  INV_X1 U14123 ( .A(n11241), .ZN(n11194) );
  XNOR2_X1 U14124 ( .A(n11243), .B(n11194), .ZN(n11195) );
  NAND2_X1 U14125 ( .A1(n11195), .A2(n11502), .ZN(n11196) );
  NAND2_X1 U14126 ( .A1(n11197), .A2(n11196), .ZN(n13597) );
  NAND2_X1 U14127 ( .A1(n13598), .A2(n13597), .ZN(n13596) );
  NAND2_X1 U14128 ( .A1(n11198), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11199) );
  INV_X1 U14129 ( .A(n11215), .ZN(n11212) );
  NAND2_X1 U14130 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11211) );
  AOI22_X1 U14131 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14132 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14133 ( .A1(n9772), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14134 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11200) );
  NAND4_X1 U14135 ( .A1(n11203), .A2(n11202), .A3(n11201), .A4(n11200), .ZN(
        n11209) );
  AOI22_X1 U14136 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14137 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14138 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14139 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11204) );
  NAND4_X1 U14140 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11208) );
  NAND2_X1 U14141 ( .A1(n11323), .A2(n11240), .ZN(n11210) );
  NAND2_X1 U14142 ( .A1(n11211), .A2(n11210), .ZN(n11213) );
  INV_X1 U14143 ( .A(n11213), .ZN(n11214) );
  NAND2_X1 U14144 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  OR2_X1 U14145 ( .A1(n11643), .A2(n11239), .ZN(n11220) );
  NAND2_X1 U14146 ( .A1(n11243), .A2(n11241), .ZN(n11217) );
  XNOR2_X1 U14147 ( .A(n11217), .B(n11240), .ZN(n11218) );
  NAND2_X1 U14148 ( .A1(n11218), .A2(n11502), .ZN(n11219) );
  NAND2_X1 U14149 ( .A1(n11220), .A2(n11219), .ZN(n11222) );
  INV_X1 U14150 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11221) );
  XNOR2_X1 U14151 ( .A(n11222), .B(n11221), .ZN(n20058) );
  NAND2_X1 U14152 ( .A1(n20059), .A2(n20058), .ZN(n20057) );
  NAND2_X1 U14153 ( .A1(n11222), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14154 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11235) );
  AOI22_X1 U14155 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14156 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11226) );
  INV_X1 U14157 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U14158 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14159 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11224) );
  NAND4_X1 U14160 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(
        n11233) );
  AOI22_X1 U14161 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14162 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14163 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14164 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14165 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11232) );
  NAND2_X1 U14166 ( .A1(n11323), .A2(n11266), .ZN(n11234) );
  NAND2_X1 U14167 ( .A1(n9727), .A2(n11236), .ZN(n11238) );
  NAND2_X1 U14168 ( .A1(n11264), .A2(n11238), .ZN(n11653) );
  OR2_X1 U14169 ( .A1(n11653), .A2(n11239), .ZN(n11246) );
  AND2_X1 U14170 ( .A1(n11241), .A2(n11240), .ZN(n11242) );
  NAND2_X1 U14171 ( .A1(n11243), .A2(n11242), .ZN(n11265) );
  XNOR2_X1 U14172 ( .A(n11265), .B(n11266), .ZN(n11244) );
  NAND2_X1 U14173 ( .A1(n11244), .A2(n11502), .ZN(n11245) );
  NAND2_X1 U14174 ( .A1(n11246), .A2(n11245), .ZN(n11247) );
  INV_X1 U14175 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20890) );
  XNOR2_X1 U14176 ( .A(n11247), .B(n20890), .ZN(n13764) );
  NAND2_X1 U14177 ( .A1(n11247), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14178 ( .A1(n11359), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11260) );
  AOI22_X1 U14179 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14180 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14181 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14182 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11249) );
  NAND4_X1 U14183 ( .A1(n11252), .A2(n11251), .A3(n11250), .A4(n11249), .ZN(
        n11258) );
  AOI22_X1 U14184 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14185 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14186 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14187 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11253) );
  NAND4_X1 U14188 ( .A1(n11256), .A2(n11255), .A3(n11254), .A4(n11253), .ZN(
        n11257) );
  NAND2_X1 U14189 ( .A1(n11323), .A2(n11279), .ZN(n11259) );
  NAND2_X1 U14190 ( .A1(n11264), .A2(n11263), .ZN(n11660) );
  INV_X1 U14191 ( .A(n11265), .ZN(n11267) );
  NAND2_X1 U14192 ( .A1(n11267), .A2(n11266), .ZN(n11278) );
  XNOR2_X1 U14193 ( .A(n11278), .B(n11279), .ZN(n11268) );
  NAND2_X1 U14194 ( .A1(n11268), .A2(n11502), .ZN(n11269) );
  INV_X1 U14195 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16094) );
  NAND2_X1 U14196 ( .A1(n16095), .A2(n16094), .ZN(n11271) );
  INV_X1 U14197 ( .A(n16095), .ZN(n11272) );
  NAND2_X1 U14198 ( .A1(n11272), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11273) );
  INV_X1 U14199 ( .A(n11359), .ZN(n11350) );
  INV_X1 U14200 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U14201 ( .A1(n11323), .A2(n11286), .ZN(n11274) );
  OAI21_X1 U14202 ( .B1(n11350), .B2(n11275), .A(n11274), .ZN(n11276) );
  INV_X1 U14203 ( .A(n11278), .ZN(n11280) );
  NAND2_X1 U14204 ( .A1(n11280), .A2(n11279), .ZN(n11291) );
  XNOR2_X1 U14205 ( .A(n11291), .B(n11286), .ZN(n11281) );
  AND2_X1 U14206 ( .A1(n11281), .A2(n11502), .ZN(n11282) );
  AOI21_X1 U14207 ( .B1(n11674), .B2(n11313), .A(n11282), .ZN(n11283) );
  INV_X1 U14208 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16215) );
  NAND2_X1 U14209 ( .A1(n11283), .A2(n16215), .ZN(n16090) );
  NAND2_X1 U14210 ( .A1(n16088), .A2(n16090), .ZN(n11285) );
  INV_X1 U14211 ( .A(n11283), .ZN(n11284) );
  NAND2_X1 U14212 ( .A1(n11284), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16089) );
  NAND2_X1 U14213 ( .A1(n11313), .A2(n11286), .ZN(n11288) );
  NOR2_X1 U14214 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  OR3_X1 U14215 ( .A1(n11291), .A2(n11290), .A3(n20677), .ZN(n11292) );
  INV_X1 U14216 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U14217 ( .A1(n14114), .A2(n14113), .ZN(n11293) );
  INV_X1 U14218 ( .A(n14114), .ZN(n11294) );
  NAND2_X1 U14219 ( .A1(n11294), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11295) );
  INV_X1 U14220 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16193) );
  NAND2_X1 U14221 ( .A1(n9750), .A2(n16193), .ZN(n11296) );
  INV_X1 U14222 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U14223 ( .A1(n9750), .A2(n11303), .ZN(n14800) );
  NAND2_X1 U14224 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11297) );
  NAND2_X1 U14225 ( .A1(n9750), .A2(n11297), .ZN(n14798) );
  AND2_X1 U14226 ( .A1(n14800), .A2(n14798), .ZN(n11298) );
  XNOR2_X1 U14227 ( .A(n9749), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14801) );
  INV_X1 U14228 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16142) );
  NAND2_X1 U14229 ( .A1(n9750), .A2(n16142), .ZN(n16067) );
  INV_X1 U14230 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16164) );
  OAI21_X1 U14231 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n16056), .ZN(n11300) );
  INV_X1 U14232 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14233 ( .A1(n9749), .A2(n11472), .ZN(n11301) );
  INV_X1 U14234 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14788) );
  NAND2_X1 U14235 ( .A1(n14788), .A2(n16164), .ZN(n11302) );
  NAND2_X1 U14236 ( .A1(n16056), .A2(n11302), .ZN(n16064) );
  NAND2_X1 U14237 ( .A1(n16056), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16068) );
  NAND2_X1 U14238 ( .A1(n16064), .A2(n16068), .ZN(n14781) );
  NOR2_X1 U14239 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14796) );
  AND2_X1 U14240 ( .A1(n14796), .A2(n11303), .ZN(n11304) );
  NOR2_X1 U14241 ( .A1(n9750), .A2(n11304), .ZN(n14780) );
  NOR2_X1 U14242 ( .A1(n14781), .A2(n14780), .ZN(n11305) );
  XNOR2_X1 U14243 ( .A(n9749), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14770) );
  NAND2_X1 U14244 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15853) );
  INV_X1 U14245 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14878) );
  NAND2_X1 U14246 ( .A1(n11306), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11307) );
  OAI21_X2 U14247 ( .B1(n14769), .B2(n11307), .A(n9749), .ZN(n14763) );
  NAND2_X1 U14248 ( .A1(n14763), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14249 ( .A1(n11310), .A2(n9750), .ZN(n11580) );
  NAND2_X1 U14250 ( .A1(n11580), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14747) );
  INV_X1 U14251 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11308) );
  INV_X1 U14252 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11483) );
  NAND2_X1 U14253 ( .A1(n11308), .A2(n11483), .ZN(n15854) );
  NAND2_X1 U14254 ( .A1(n11309), .A2(n16056), .ZN(n14764) );
  NAND2_X1 U14255 ( .A1(n11310), .A2(n14764), .ZN(n11536) );
  INV_X1 U14256 ( .A(n11536), .ZN(n14737) );
  NAND2_X1 U14257 ( .A1(n14737), .A2(n14747), .ZN(n11311) );
  MUX2_X1 U14258 ( .A(n14747), .B(n11311), .S(n16056), .Z(n11312) );
  INV_X1 U14259 ( .A(n14760), .ZN(n11399) );
  XNOR2_X1 U14260 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U14261 ( .A1(n11331), .A2(n11329), .ZN(n11315) );
  NAND2_X1 U14262 ( .A1(n20524), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U14263 ( .A1(n11315), .A2(n11314), .ZN(n11327) );
  XNOR2_X1 U14264 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11326) );
  NAND2_X1 U14265 ( .A1(n11327), .A2(n11326), .ZN(n11317) );
  NAND2_X1 U14266 ( .A1(n15810), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11316) );
  NAND2_X1 U14267 ( .A1(n11317), .A2(n11316), .ZN(n11325) );
  MUX2_X1 U14268 ( .A(n11318), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11324) );
  NAND2_X1 U14269 ( .A1(n11325), .A2(n11324), .ZN(n11320) );
  NAND2_X1 U14270 ( .A1(n11318), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11319) );
  NAND2_X1 U14271 ( .A1(n11320), .A2(n11319), .ZN(n11355) );
  NOR2_X1 U14272 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13534), .ZN(
        n11321) );
  NAND2_X1 U14273 ( .A1(n11386), .A2(n11323), .ZN(n11365) );
  XNOR2_X1 U14274 ( .A(n11325), .B(n11324), .ZN(n11383) );
  XNOR2_X1 U14275 ( .A(n11327), .B(n11326), .ZN(n11381) );
  AOI21_X1 U14276 ( .B1(n13544), .B2(n11328), .A(n11022), .ZN(n11345) );
  AOI211_X1 U14277 ( .C1(n11359), .C2(n11381), .A(n11344), .B(n11345), .ZN(
        n11349) );
  XNOR2_X1 U14278 ( .A(n11329), .B(n11331), .ZN(n11382) );
  NAND2_X1 U14279 ( .A1(n13544), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11337) );
  OAI21_X1 U14280 ( .B1(n13335), .B2(n11338), .A(n11337), .ZN(n11330) );
  INV_X1 U14281 ( .A(n11340), .ZN(n11343) );
  INV_X1 U14282 ( .A(n11331), .ZN(n11333) );
  NAND2_X1 U14283 ( .A1(n10881), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11332) );
  NAND2_X1 U14284 ( .A1(n11333), .A2(n11332), .ZN(n11336) );
  AOI21_X1 U14285 ( .B1(n10960), .B2(n11328), .A(n11345), .ZN(n11334) );
  NOR3_X1 U14286 ( .A1(n11334), .A2(n11338), .A3(n11336), .ZN(n11335) );
  AOI21_X1 U14287 ( .B1(n11353), .B2(n11336), .A(n11335), .ZN(n11339) );
  INV_X1 U14288 ( .A(n11339), .ZN(n11342) );
  NAND3_X1 U14289 ( .A1(n11338), .A2(n11022), .A3(n11337), .ZN(n11357) );
  AOI22_X1 U14290 ( .A1(n11382), .A2(n11357), .B1(n11340), .B2(n11339), .ZN(
        n11341) );
  AOI21_X1 U14291 ( .B1(n11343), .B2(n11342), .A(n11341), .ZN(n11348) );
  INV_X1 U14292 ( .A(n11344), .ZN(n11347) );
  INV_X1 U14293 ( .A(n11345), .ZN(n11346) );
  OAI22_X1 U14294 ( .A1(n11349), .A2(n11348), .B1(n11347), .B2(n11346), .ZN(
        n11352) );
  NAND2_X1 U14295 ( .A1(n11350), .A2(n11383), .ZN(n11351) );
  AOI22_X1 U14296 ( .A1(n11353), .A2(n11383), .B1(n11352), .B2(n11351), .ZN(
        n11362) );
  INV_X1 U14297 ( .A(n11384), .ZN(n11356) );
  NOR2_X1 U14298 ( .A1(n11359), .A2(n11356), .ZN(n11361) );
  INV_X1 U14299 ( .A(n11357), .ZN(n11358) );
  NAND3_X1 U14300 ( .A1(n11359), .A2(n11358), .A3(n11384), .ZN(n11360) );
  OAI21_X1 U14301 ( .B1(n11362), .B2(n11361), .A(n11360), .ZN(n11363) );
  AOI21_X1 U14302 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16236), .A(
        n11363), .ZN(n11364) );
  NAND2_X1 U14303 ( .A1(n11365), .A2(n11364), .ZN(n11366) );
  NOR2_X1 U14304 ( .A1(n14257), .A2(n13335), .ZN(n11518) );
  INV_X1 U14305 ( .A(n11518), .ZN(n11392) );
  INV_X1 U14306 ( .A(n11369), .ZN(n11370) );
  NAND2_X1 U14307 ( .A1(n11370), .A2(n12385), .ZN(n11372) );
  AND2_X1 U14308 ( .A1(n11372), .A2(n11371), .ZN(n11508) );
  NAND2_X1 U14309 ( .A1(n14257), .A2(n13911), .ZN(n11373) );
  AND3_X1 U14310 ( .A1(n11508), .A2(n11374), .A3(n11373), .ZN(n12388) );
  OR2_X1 U14311 ( .A1(n13130), .A2(n12388), .ZN(n11375) );
  NAND2_X1 U14312 ( .A1(n11375), .A2(n11512), .ZN(n13270) );
  INV_X1 U14313 ( .A(n13270), .ZN(n11391) );
  OR2_X1 U14314 ( .A1(n11377), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15843) );
  INV_X1 U14315 ( .A(n15843), .ZN(n15795) );
  NAND2_X1 U14316 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20603) );
  OAI21_X1 U14317 ( .B1(n11022), .B2(n15795), .A(n20603), .ZN(n13913) );
  INV_X1 U14318 ( .A(n13913), .ZN(n11378) );
  NAND2_X1 U14319 ( .A1(n11376), .A2(n11378), .ZN(n11379) );
  NAND3_X1 U14320 ( .A1(n11379), .A2(n11328), .A3(n11010), .ZN(n11380) );
  NAND2_X1 U14321 ( .A1(n11380), .A2(n13537), .ZN(n11389) );
  NOR4_X1 U14322 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11385) );
  NOR2_X1 U14323 ( .A1(n11386), .A2(n11385), .ZN(n13128) );
  NAND2_X1 U14324 ( .A1(n13128), .A2(n20603), .ZN(n12387) );
  AND2_X1 U14325 ( .A1(n11022), .A2(n15843), .ZN(n11387) );
  OR2_X1 U14326 ( .A1(n12387), .A2(n11387), .ZN(n11388) );
  OAI211_X1 U14327 ( .C1(n13537), .C2(n11392), .A(n11391), .B(n11390), .ZN(
        n11393) );
  OAI21_X1 U14328 ( .B1(n10960), .B2(n13904), .A(n12388), .ZN(n11395) );
  OAI21_X1 U14329 ( .B1(n12385), .B2(n9740), .A(n11395), .ZN(n11396) );
  OR2_X1 U14330 ( .A1(n11397), .A2(n11396), .ZN(n11398) );
  MUX2_X1 U14331 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11405) );
  INV_X1 U14332 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11406) );
  OR2_X1 U14333 ( .A1(n11446), .A2(n11406), .ZN(n11408) );
  NAND2_X1 U14334 ( .A1(n11024), .A2(n11406), .ZN(n11407) );
  NAND2_X1 U14335 ( .A1(n11408), .A2(n11407), .ZN(n13200) );
  MUX2_X1 U14336 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11410) );
  OAI21_X1 U14337 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n11401), .A(
        n11410), .ZN(n13326) );
  INV_X1 U14338 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20846) );
  NAND2_X1 U14339 ( .A1(n11478), .A2(n20846), .ZN(n11414) );
  NAND2_X1 U14340 ( .A1(n13909), .A2(n20846), .ZN(n11412) );
  NAND2_X1 U14341 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11411) );
  NAND3_X1 U14342 ( .A1(n11412), .A2(n11446), .A3(n11411), .ZN(n11413) );
  AND2_X1 U14343 ( .A1(n11414), .A2(n11413), .ZN(n19973) );
  OR2_X1 U14344 ( .A1(n11572), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U14345 ( .A1(n11446), .A2(n11415), .ZN(n11418) );
  INV_X1 U14346 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U14347 ( .A1(n13909), .A2(n11416), .ZN(n11417) );
  NAND3_X1 U14348 ( .A1(n11418), .A2(n11553), .A3(n11417), .ZN(n11419) );
  NAND2_X1 U14349 ( .A1(n11420), .A2(n11419), .ZN(n19972) );
  OR2_X1 U14350 ( .A1(n11572), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11426) );
  NAND2_X1 U14351 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11422) );
  NAND2_X1 U14352 ( .A1(n11446), .A2(n11422), .ZN(n11424) );
  INV_X1 U14353 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U14354 ( .A1(n11548), .A2(n13733), .ZN(n11423) );
  NAND2_X1 U14355 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  INV_X1 U14356 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20020) );
  NAND2_X1 U14357 ( .A1(n11478), .A2(n20020), .ZN(n11430) );
  NAND2_X1 U14358 ( .A1(n11548), .A2(n20020), .ZN(n11428) );
  NAND2_X1 U14359 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11427) );
  NAND3_X1 U14360 ( .A1(n11428), .A2(n11446), .A3(n11427), .ZN(n11429) );
  OR2_X1 U14361 ( .A1(n11572), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U14362 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11431) );
  NAND2_X1 U14363 ( .A1(n11446), .A2(n11431), .ZN(n11433) );
  INV_X1 U14364 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13784) );
  NAND2_X1 U14365 ( .A1(n11548), .A2(n13784), .ZN(n11432) );
  NAND2_X1 U14366 ( .A1(n11433), .A2(n11432), .ZN(n11434) );
  NAND2_X1 U14367 ( .A1(n11435), .A2(n11434), .ZN(n13783) );
  INV_X1 U14368 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13897) );
  NAND2_X1 U14369 ( .A1(n11548), .A2(n13897), .ZN(n11437) );
  NAND2_X1 U14370 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11436) );
  NAND3_X1 U14371 ( .A1(n11437), .A2(n11446), .A3(n11436), .ZN(n11438) );
  OAI21_X1 U14372 ( .B1(n11554), .B2(P1_EBX_REG_8__SCAN_IN), .A(n11438), .ZN(
        n13894) );
  OR2_X1 U14373 ( .A1(n11572), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11443) );
  NAND2_X1 U14374 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11439) );
  NAND2_X1 U14375 ( .A1(n11446), .A2(n11439), .ZN(n11441) );
  INV_X1 U14376 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U14377 ( .A1(n11548), .A2(n14111), .ZN(n11440) );
  NAND2_X1 U14378 ( .A1(n11441), .A2(n11440), .ZN(n11442) );
  MUX2_X1 U14379 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11444) );
  OAI21_X1 U14380 ( .B1(n11401), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11444), .ZN(n14084) );
  INV_X1 U14381 ( .A(n14084), .ZN(n11445) );
  OR2_X1 U14382 ( .A1(n11572), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n11451) );
  NAND2_X1 U14383 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11447) );
  NAND2_X1 U14384 ( .A1(n11446), .A2(n11447), .ZN(n11449) );
  INV_X1 U14385 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14211) );
  NAND2_X1 U14386 ( .A1(n11548), .A2(n14211), .ZN(n11448) );
  NAND2_X1 U14387 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NAND2_X1 U14388 ( .A1(n11451), .A2(n11450), .ZN(n14208) );
  INV_X1 U14389 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16007) );
  NAND2_X1 U14390 ( .A1(n11548), .A2(n16007), .ZN(n11453) );
  NAND2_X1 U14391 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11452) );
  NAND3_X1 U14392 ( .A1(n11453), .A2(n11446), .A3(n11452), .ZN(n11454) );
  OAI21_X1 U14393 ( .B1(n11554), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11454), .ZN(
        n15985) );
  MUX2_X1 U14394 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11455) );
  OAI21_X1 U14395 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n11401), .A(
        n11455), .ZN(n11456) );
  INV_X1 U14396 ( .A(n11456), .ZN(n14174) );
  OR2_X1 U14397 ( .A1(n11572), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U14398 ( .A1(n11446), .A2(n14788), .ZN(n11459) );
  INV_X1 U14399 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14400 ( .A1(n11548), .A2(n11457), .ZN(n11458) );
  NAND3_X1 U14401 ( .A1(n11459), .A2(n11553), .A3(n11458), .ZN(n11460) );
  NAND2_X1 U14402 ( .A1(n11461), .A2(n11460), .ZN(n14640) );
  NAND2_X1 U14403 ( .A1(n14174), .A2(n14640), .ZN(n11462) );
  OR2_X1 U14404 ( .A1(n11572), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14405 ( .A1(n11446), .A2(n16142), .ZN(n11464) );
  INV_X1 U14406 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15965) );
  NAND2_X1 U14407 ( .A1(n11548), .A2(n15965), .ZN(n11463) );
  NAND3_X1 U14408 ( .A1(n11464), .A2(n11553), .A3(n11463), .ZN(n11465) );
  NAND2_X1 U14409 ( .A1(n11466), .A2(n11465), .ZN(n14185) );
  MUX2_X1 U14410 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11467) );
  OAI21_X1 U14411 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n11401), .A(
        n11467), .ZN(n14195) );
  INV_X1 U14412 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U14413 ( .A1(n11478), .A2(n14632), .ZN(n11471) );
  NAND2_X1 U14414 ( .A1(n11548), .A2(n14632), .ZN(n11469) );
  NAND2_X1 U14415 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11468) );
  NAND3_X1 U14416 ( .A1(n11469), .A2(n11446), .A3(n11468), .ZN(n11470) );
  AND2_X1 U14417 ( .A1(n11471), .A2(n11470), .ZN(n14574) );
  OR2_X1 U14418 ( .A1(n11572), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U14419 ( .A1(n11446), .A2(n11472), .ZN(n11474) );
  INV_X1 U14420 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16005) );
  NAND2_X1 U14421 ( .A1(n11548), .A2(n16005), .ZN(n11473) );
  NAND3_X1 U14422 ( .A1(n11474), .A2(n11553), .A3(n11473), .ZN(n11475) );
  NAND2_X1 U14423 ( .A1(n11476), .A2(n11475), .ZN(n15958) );
  NAND2_X1 U14424 ( .A1(n14574), .A2(n15958), .ZN(n11477) );
  INV_X1 U14425 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n16001) );
  NAND2_X1 U14426 ( .A1(n11478), .A2(n16001), .ZN(n11482) );
  NAND2_X1 U14427 ( .A1(n11548), .A2(n16001), .ZN(n11480) );
  NAND2_X1 U14428 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11479) );
  NAND3_X1 U14429 ( .A1(n11480), .A2(n11446), .A3(n11479), .ZN(n11481) );
  AND2_X1 U14430 ( .A1(n11482), .A2(n11481), .ZN(n15855) );
  OR2_X1 U14431 ( .A1(n11572), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U14432 ( .A1(n11446), .A2(n11483), .ZN(n11485) );
  INV_X1 U14433 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16003) );
  NAND2_X1 U14434 ( .A1(n11548), .A2(n16003), .ZN(n11484) );
  NAND3_X1 U14435 ( .A1(n11485), .A2(n11553), .A3(n11484), .ZN(n11486) );
  NAND2_X1 U14436 ( .A1(n11487), .A2(n11486), .ZN(n15949) );
  NAND2_X1 U14437 ( .A1(n15855), .A2(n15949), .ZN(n11488) );
  OR2_X1 U14438 ( .A1(n11572), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U14439 ( .A1(n11446), .A2(n14878), .ZN(n11490) );
  INV_X1 U14440 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15924) );
  NAND2_X1 U14441 ( .A1(n11548), .A2(n15924), .ZN(n11489) );
  NAND3_X1 U14442 ( .A1(n11490), .A2(n11553), .A3(n11489), .ZN(n11491) );
  NAND2_X1 U14443 ( .A1(n11492), .A2(n11491), .ZN(n14627) );
  MUX2_X1 U14444 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11494) );
  OR2_X1 U14445 ( .A1(n11401), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11493) );
  AND2_X1 U14446 ( .A1(n11494), .A2(n11493), .ZN(n14621) );
  OR2_X1 U14447 ( .A1(n11572), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n11498) );
  INV_X1 U14448 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14862) );
  NAND2_X1 U14449 ( .A1(n11446), .A2(n14862), .ZN(n11496) );
  INV_X1 U14450 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15905) );
  NAND2_X1 U14451 ( .A1(n11548), .A2(n15905), .ZN(n11495) );
  NAND3_X1 U14452 ( .A1(n11496), .A2(n11553), .A3(n11495), .ZN(n11497) );
  AND2_X1 U14453 ( .A1(n11498), .A2(n11497), .ZN(n14616) );
  MUX2_X1 U14454 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11499) );
  OAI21_X1 U14455 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n11401), .A(
        n11499), .ZN(n11500) );
  AND2_X1 U14456 ( .A1(n14618), .A2(n11500), .ZN(n11501) );
  OR2_X1 U14457 ( .A1(n11501), .A2(n14605), .ZN(n14610) );
  INV_X1 U14458 ( .A(n14610), .ZN(n11504) );
  NAND2_X1 U14459 ( .A1(n11376), .A2(n11502), .ZN(n15797) );
  OAI21_X1 U14460 ( .B1(n9740), .B2(n13574), .A(n15797), .ZN(n11503) );
  NAND2_X1 U14461 ( .A1(n11504), .A2(n20098), .ZN(n11531) );
  AND2_X1 U14462 ( .A1(n13130), .A2(n11022), .ZN(n15802) );
  OR2_X1 U14463 ( .A1(n10960), .A2(n13908), .ZN(n11505) );
  AND2_X1 U14464 ( .A1(n11506), .A2(n11505), .ZN(n11519) );
  NAND2_X1 U14465 ( .A1(n9729), .A2(n13904), .ZN(n11511) );
  INV_X1 U14466 ( .A(n11014), .ZN(n11507) );
  NAND2_X1 U14467 ( .A1(n11508), .A2(n11507), .ZN(n11509) );
  NAND2_X1 U14468 ( .A1(n11509), .A2(n11022), .ZN(n11510) );
  AND4_X1 U14469 ( .A1(n11512), .A2(n11519), .A3(n11511), .A4(n11510), .ZN(
        n13500) );
  MUX2_X1 U14470 ( .A(n11514), .B(n11513), .S(n11328), .Z(n11515) );
  NAND3_X1 U14471 ( .A1(n13500), .A2(n11516), .A3(n11515), .ZN(n11517) );
  NOR2_X1 U14472 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16169), .ZN(
        n13290) );
  NAND2_X1 U14473 ( .A1(n20101), .A2(n16172), .ZN(n16201) );
  NAND2_X1 U14474 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16109) );
  INV_X1 U14475 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16194) );
  NAND3_X1 U14476 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14156) );
  NOR3_X1 U14477 ( .A1(n16194), .A2(n16193), .A3(n14156), .ZN(n14886) );
  NAND2_X1 U14478 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14886), .ZN(
        n16181) );
  NOR2_X1 U14479 ( .A1(n11303), .A2(n16181), .ZN(n11520) );
  NAND2_X1 U14480 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20079) );
  INV_X1 U14481 ( .A(n20079), .ZN(n14161) );
  NOR2_X1 U14482 ( .A1(n20107), .A2(n11402), .ZN(n14155) );
  NAND2_X1 U14483 ( .A1(n14161), .A2(n14155), .ZN(n13767) );
  NOR2_X1 U14484 ( .A1(n20890), .A2(n13767), .ZN(n14883) );
  AND2_X1 U14485 ( .A1(n11520), .A2(n14883), .ZN(n16167) );
  NAND2_X1 U14486 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16167), .ZN(
        n16125) );
  INV_X1 U14487 ( .A(n20101), .ZN(n16126) );
  NAND4_X1 U14488 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11524) );
  INV_X1 U14489 ( .A(n11524), .ZN(n16127) );
  NAND2_X1 U14490 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16127), .ZN(
        n15850) );
  AOI21_X1 U14491 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20093) );
  NOR3_X1 U14492 ( .A1(n20093), .A2(n20890), .A3(n20079), .ZN(n14158) );
  NAND2_X1 U14493 ( .A1(n14158), .A2(n11520), .ZN(n16171) );
  NOR2_X1 U14494 ( .A1(n14788), .A2(n16171), .ZN(n16161) );
  INV_X1 U14495 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13284) );
  INV_X2 U14496 ( .A(n16209), .ZN(n20106) );
  NOR2_X1 U14497 ( .A1(n20106), .A2(n11521), .ZN(n14895) );
  OAI21_X1 U14498 ( .B1(n16161), .B2(n16172), .A(n20100), .ZN(n16124) );
  AOI221_X1 U14499 ( .B1(n16125), .B2(n16126), .C1(n15850), .C2(n16126), .A(
        n16124), .ZN(n15851) );
  NOR2_X1 U14500 ( .A1(n15853), .A2(n15850), .ZN(n14871) );
  INV_X1 U14501 ( .A(n20100), .ZN(n14153) );
  NOR2_X1 U14502 ( .A1(n16201), .A2(n14153), .ZN(n14157) );
  AOI21_X1 U14503 ( .B1(n9692), .B2(n14871), .A(n14157), .ZN(n16106) );
  OAI21_X1 U14504 ( .B1(n16172), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14863), .ZN(n11561) );
  AOI21_X1 U14505 ( .B1(n20108), .B2(n14862), .A(n11561), .ZN(n11522) );
  OR2_X1 U14506 ( .A1(n11522), .A2(n14746), .ZN(n11529) );
  INV_X1 U14507 ( .A(n16125), .ZN(n11523) );
  AOI22_X1 U14508 ( .A1(n20097), .A2(n16161), .B1(n11523), .B2(n20108), .ZN(
        n16134) );
  NOR2_X1 U14509 ( .A1(n16134), .A2(n11524), .ZN(n16130) );
  NAND2_X1 U14510 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16130), .ZN(
        n16120) );
  INV_X1 U14511 ( .A(n16120), .ZN(n11526) );
  NOR2_X1 U14512 ( .A1(n15853), .A2(n16109), .ZN(n11525) );
  NAND2_X1 U14513 ( .A1(n11526), .A2(n11525), .ZN(n14868) );
  NOR2_X1 U14514 ( .A1(n14862), .A2(n14868), .ZN(n11527) );
  AOI22_X1 U14515 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20106), .B1(n11527), 
        .B2(n14746), .ZN(n11528) );
  AND2_X1 U14516 ( .A1(n11529), .A2(n11528), .ZN(n11530) );
  NAND2_X1 U14517 ( .A1(n11533), .A2(n11532), .ZN(P1_U3007) );
  NAND3_X1 U14518 ( .A1(n14746), .A2(n11534), .A3(n14862), .ZN(n11535) );
  INV_X1 U14519 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14844) );
  NAND2_X1 U14520 ( .A1(n14740), .A2(n14844), .ZN(n11539) );
  NAND3_X1 U14521 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14522 ( .A1(n9749), .A2(n11584), .ZN(n14738) );
  NAND3_X1 U14523 ( .A1(n11536), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14738), .ZN(n11538) );
  MUX2_X1 U14524 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14844), .S(
        n9749), .Z(n11537) );
  AOI21_X1 U14525 ( .B1(n11539), .B2(n11538), .A(n11537), .ZN(n11540) );
  XNOR2_X1 U14526 ( .A(n11540), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14731) );
  OR2_X1 U14527 ( .A1(n11572), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n11544) );
  NAND2_X1 U14528 ( .A1(n11446), .A2(n11534), .ZN(n11542) );
  INV_X1 U14529 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15893) );
  NAND2_X1 U14530 ( .A1(n11548), .A2(n15893), .ZN(n11541) );
  NAND3_X1 U14531 ( .A1(n11542), .A2(n11553), .A3(n11541), .ZN(n11543) );
  NAND2_X1 U14532 ( .A1(n11544), .A2(n11543), .ZN(n14604) );
  MUX2_X1 U14533 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11546) );
  OR2_X1 U14534 ( .A1(n11401), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11545) );
  AND2_X1 U14535 ( .A1(n11546), .A2(n11545), .ZN(n14598) );
  OR2_X1 U14536 ( .A1(n11572), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U14537 ( .A1(n11553), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14538 ( .A1(n11446), .A2(n11547), .ZN(n11550) );
  INV_X1 U14539 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U14540 ( .A1(n11548), .A2(n14592), .ZN(n11549) );
  NAND2_X1 U14541 ( .A1(n11550), .A2(n11549), .ZN(n11551) );
  AND2_X1 U14542 ( .A1(n11552), .A2(n11551), .ZN(n14590) );
  MUX2_X1 U14543 ( .A(n11554), .B(n11553), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11555) );
  OAI21_X1 U14544 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11401), .A(
        n11555), .ZN(n11556) );
  AND2_X1 U14545 ( .A1(n9788), .A2(n11556), .ZN(n11557) );
  OR2_X1 U14546 ( .A1(n11557), .A2(n12894), .ZN(n14586) );
  NAND2_X1 U14547 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14548 ( .A1(n16169), .A2(n11584), .ZN(n11560) );
  OR2_X1 U14549 ( .A1(n14746), .A2(n14862), .ZN(n11558) );
  NAND2_X1 U14550 ( .A1(n16168), .A2(n11558), .ZN(n11559) );
  OAI211_X1 U14551 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16172), .A(
        n11560), .B(n11559), .ZN(n11562) );
  INV_X1 U14552 ( .A(n11577), .ZN(n14837) );
  INV_X1 U14553 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14548) );
  NOR2_X1 U14554 ( .A1(n16209), .A2(n14548), .ZN(n14727) );
  AOI21_X1 U14555 ( .B1(n14837), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14727), .ZN(n11564) );
  OAI21_X1 U14556 ( .B1(n14586), .B2(n16210), .A(n11564), .ZN(n11568) );
  INV_X1 U14557 ( .A(n11584), .ZN(n14845) );
  NAND2_X1 U14558 ( .A1(n14845), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11565) );
  NOR2_X1 U14559 ( .A1(n14868), .A2(n11565), .ZN(n14840) );
  XNOR2_X1 U14560 ( .A(n11581), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11566) );
  AND2_X1 U14561 ( .A1(n14840), .A2(n11566), .ZN(n11567) );
  AND2_X1 U14562 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U14563 ( .A1(n14840), .A2(n11585), .ZN(n14827) );
  OR2_X1 U14564 ( .A1(n11401), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11571) );
  INV_X1 U14565 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14585) );
  NAND2_X1 U14566 ( .A1(n11548), .A2(n14585), .ZN(n11570) );
  NAND2_X1 U14567 ( .A1(n11571), .A2(n11570), .ZN(n12896) );
  OAI22_X1 U14568 ( .A1(n12896), .A2(n11024), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11572), .ZN(n11573) );
  NAND2_X1 U14569 ( .A1(n12894), .A2(n11573), .ZN(n14511) );
  OR2_X1 U14570 ( .A1(n12894), .A2(n11573), .ZN(n11574) );
  NAND2_X1 U14571 ( .A1(n14511), .A2(n11574), .ZN(n14584) );
  INV_X1 U14572 ( .A(n11585), .ZN(n11575) );
  NAND2_X1 U14573 ( .A1(n16201), .A2(n11575), .ZN(n11576) );
  NAND2_X1 U14574 ( .A1(n11577), .A2(n11576), .ZN(n14819) );
  INV_X1 U14575 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20652) );
  NOR2_X1 U14576 ( .A1(n16209), .A2(n20652), .ZN(n14717) );
  AOI21_X1 U14577 ( .B1(n14819), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14717), .ZN(n11578) );
  OAI21_X1 U14578 ( .B1(n14584), .B2(n16210), .A(n11578), .ZN(n11579) );
  INV_X1 U14579 ( .A(n11579), .ZN(n11587) );
  INV_X1 U14580 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U14581 ( .A1(n11582), .A2(n11581), .ZN(n11583) );
  NAND2_X1 U14582 ( .A1(n14732), .A2(n11585), .ZN(n14708) );
  XNOR2_X1 U14583 ( .A(n9750), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11586) );
  XNOR2_X1 U14584 ( .A(n11605), .B(n11586), .ZN(n14723) );
  OAI211_X1 U14585 ( .C1(n14827), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11587), .B(n9799), .ZN(P1_U3002) );
  INV_X1 U14586 ( .A(n15138), .ZN(n15380) );
  NAND2_X1 U14587 ( .A1(n14278), .A2(n15382), .ZN(n15379) );
  NAND2_X1 U14588 ( .A1(n15379), .A2(n10876), .ZN(n11600) );
  AOI21_X1 U14589 ( .B1(n12941), .B2(n11588), .A(n11589), .ZN(n12939) );
  NOR2_X1 U14590 ( .A1(n18970), .A2(n19836), .ZN(n15381) );
  INV_X1 U14591 ( .A(n15381), .ZN(n11590) );
  OAI21_X1 U14592 ( .B1(n19184), .B2(n12941), .A(n11590), .ZN(n11595) );
  INV_X1 U14593 ( .A(n11591), .ZN(n15017) );
  NAND2_X1 U14594 ( .A1(n15017), .A2(n11592), .ZN(n11593) );
  NAND2_X1 U14595 ( .A1(n14949), .A2(n11593), .ZN(n15386) );
  NOR2_X1 U14596 ( .A1(n15386), .A2(n15652), .ZN(n11594) );
  AOI211_X1 U14597 ( .C1(n16343), .C2(n12939), .A(n11595), .B(n11594), .ZN(
        n11599) );
  XNOR2_X1 U14598 ( .A(n15140), .B(n15139), .ZN(n15142) );
  XNOR2_X1 U14599 ( .A(n15142), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15392) );
  INV_X1 U14600 ( .A(n15335), .ZN(n19179) );
  INV_X1 U14601 ( .A(n11605), .ZN(n11601) );
  MUX2_X1 U14602 ( .A(n11604), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .S(
        n9749), .Z(n11602) );
  INV_X1 U14603 ( .A(n11602), .ZN(n11603) );
  NAND2_X1 U14604 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  NAND2_X1 U14605 ( .A1(n12388), .A2(n10960), .ZN(n13133) );
  INV_X1 U14606 ( .A(n11010), .ZN(n12394) );
  AND2_X1 U14607 ( .A1(n12394), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11640) );
  NAND2_X1 U14608 ( .A1(n11640), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11612) );
  INV_X1 U14609 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19995) );
  XNOR2_X1 U14610 ( .A(n19995), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20001) );
  NAND2_X1 U14611 ( .A1(n20525), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11831) );
  OAI21_X1 U14612 ( .B1(n20001), .B2(n13901), .A(n11831), .ZN(n11610) );
  AOI21_X1 U14613 ( .B1(n11669), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11610), .ZN(
        n11611) );
  AND2_X1 U14614 ( .A1(n11612), .A2(n11611), .ZN(n11613) );
  INV_X1 U14615 ( .A(n11831), .ZN(n12103) );
  NAND2_X1 U14616 ( .A1(n12103), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11632) );
  NAND2_X1 U14617 ( .A1(n11615), .A2(n11614), .ZN(n11616) );
  NAND2_X1 U14618 ( .A1(n14902), .A2(n11763), .ZN(n11621) );
  INV_X1 U14619 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13397) );
  NAND2_X1 U14620 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20525), .ZN(
        n11618) );
  OAI21_X1 U14621 ( .B1(n12046), .B2(n13397), .A(n11618), .ZN(n11619) );
  AOI21_X1 U14622 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11640), .A(
        n11619), .ZN(n11620) );
  NAND2_X1 U14623 ( .A1(n11621), .A2(n11620), .ZN(n13294) );
  NAND2_X1 U14624 ( .A1(n11622), .A2(n9725), .ZN(n11623) );
  NAND2_X1 U14625 ( .A1(n11623), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13203) );
  INV_X1 U14626 ( .A(n11640), .ZN(n11649) );
  NAND2_X1 U14627 ( .A1(n11669), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11626) );
  NAND2_X1 U14628 ( .A1(n20525), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11625) );
  OAI211_X1 U14629 ( .C1(n11649), .C2(n10881), .A(n11626), .B(n11625), .ZN(
        n11627) );
  AOI21_X1 U14630 ( .B1(n11624), .B2(n11763), .A(n11627), .ZN(n11628) );
  OR2_X1 U14631 ( .A1(n13203), .A2(n11628), .ZN(n13204) );
  INV_X1 U14632 ( .A(n11628), .ZN(n13205) );
  OR2_X1 U14633 ( .A1(n13205), .A2(n13901), .ZN(n11629) );
  NAND2_X1 U14634 ( .A1(n13204), .A2(n11629), .ZN(n13293) );
  NAND2_X1 U14635 ( .A1(n13294), .A2(n13293), .ZN(n13324) );
  NAND2_X1 U14636 ( .A1(n11631), .A2(n11630), .ZN(n13322) );
  INV_X1 U14637 ( .A(n20117), .ZN(n11633) );
  NAND2_X1 U14638 ( .A1(n11633), .A2(n11763), .ZN(n11642) );
  INV_X1 U14639 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13411) );
  INV_X1 U14640 ( .A(n11635), .ZN(n11637) );
  INV_X1 U14641 ( .A(n11645), .ZN(n11636) );
  OAI21_X1 U14642 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11637), .A(
        n11636), .ZN(n13923) );
  AOI22_X1 U14643 ( .A1(n12099), .A2(n13923), .B1(n12103), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11638) );
  OAI21_X1 U14644 ( .B1(n12046), .B2(n13411), .A(n11638), .ZN(n11639) );
  AOI21_X1 U14645 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11640), .A(
        n11639), .ZN(n11641) );
  NAND2_X1 U14646 ( .A1(n11642), .A2(n11641), .ZN(n13331) );
  NAND2_X1 U14647 ( .A1(n13328), .A2(n13331), .ZN(n13329) );
  OAI21_X1 U14648 ( .B1(n11645), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11654), .ZN(n20065) );
  INV_X1 U14649 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11646) );
  AOI21_X1 U14650 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n11646), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11647) );
  AOI21_X1 U14651 ( .B1(n11669), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11647), .ZN(
        n11648) );
  OAI21_X1 U14652 ( .B1(n13534), .B2(n11649), .A(n11648), .ZN(n11650) );
  OAI21_X1 U14653 ( .B1(n20065), .B2(n13901), .A(n11650), .ZN(n11651) );
  AND2_X2 U14654 ( .A1(n11652), .A2(n11651), .ZN(n13735) );
  INV_X1 U14655 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13734) );
  OAI21_X1 U14656 ( .B1(n11655), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n11661), .ZN(n19971) );
  NAND2_X1 U14657 ( .A1(n19971), .A2(n12099), .ZN(n11657) );
  NAND2_X1 U14658 ( .A1(n12103), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11656) );
  OAI211_X1 U14659 ( .C1(n12046), .C2(n13734), .A(n11657), .B(n11656), .ZN(
        n11658) );
  INV_X1 U14660 ( .A(n11658), .ZN(n11659) );
  NAND2_X1 U14661 ( .A1(n11660), .A2(n11763), .ZN(n11666) );
  OAI21_X1 U14662 ( .B1(n11662), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11667), .ZN(n19962) );
  INV_X1 U14663 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13846) );
  INV_X1 U14664 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11663) );
  OAI22_X1 U14665 ( .A1(n12046), .A2(n13846), .B1(n11831), .B2(n11663), .ZN(
        n11664) );
  AOI21_X1 U14666 ( .B1(n12099), .B2(n19962), .A(n11664), .ZN(n11665) );
  INV_X1 U14667 ( .A(n13780), .ZN(n11676) );
  INV_X1 U14668 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11672) );
  OAI21_X1 U14669 ( .B1(n11668), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11677), .ZN(n19953) );
  NAND2_X1 U14670 ( .A1(n19953), .A2(n12099), .ZN(n11671) );
  NAND2_X1 U14671 ( .A1(n11669), .A2(P1_EAX_REG_7__SCAN_IN), .ZN(n11670) );
  OAI211_X1 U14672 ( .C1(n11831), .C2(n11672), .A(n11671), .B(n11670), .ZN(
        n11673) );
  NAND2_X1 U14673 ( .A1(n11676), .A2(n11675), .ZN(n13778) );
  AOI21_X1 U14674 ( .B1(n11677), .B2(n20950), .A(n11717), .ZN(n19942) );
  OR2_X1 U14675 ( .A1(n19942), .A2(n13901), .ZN(n11692) );
  AOI22_X1 U14676 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14677 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14678 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14679 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U14680 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11687) );
  AOI22_X1 U14681 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14682 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11923), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14683 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14684 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U14685 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11686) );
  NOR2_X1 U14686 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  OAI22_X1 U14687 ( .A1(n10100), .A2(n11688), .B1(n11831), .B2(n20950), .ZN(
        n11690) );
  INV_X1 U14688 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13938) );
  NOR2_X1 U14689 ( .A1(n12046), .A2(n13938), .ZN(n11689) );
  NOR2_X1 U14690 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  INV_X1 U14691 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19922) );
  XNOR2_X1 U14692 ( .A(n19922), .B(n11717), .ZN(n19928) );
  AOI22_X1 U14693 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14694 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14695 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14696 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14697 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11702) );
  AOI22_X1 U14698 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14699 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14700 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14701 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14702 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  NOR2_X1 U14703 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  OAI22_X1 U14704 ( .A1(n10100), .A2(n11703), .B1(n11831), .B2(n19922), .ZN(
        n11705) );
  INV_X1 U14705 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14106) );
  NOR2_X1 U14706 ( .A1(n12046), .A2(n14106), .ZN(n11704) );
  NOR2_X1 U14707 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  OAI21_X1 U14708 ( .B1(n19928), .B2(n13901), .A(n11706), .ZN(n14105) );
  AOI22_X1 U14709 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14710 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14711 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14712 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11707) );
  NAND4_X1 U14713 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11716) );
  AOI22_X1 U14714 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14715 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14716 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14717 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11711) );
  NAND4_X1 U14718 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11715) );
  NOR2_X1 U14719 ( .A1(n11716), .A2(n11715), .ZN(n11721) );
  NAND2_X1 U14720 ( .A1(n11669), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11720) );
  INV_X1 U14721 ( .A(n11722), .ZN(n11718) );
  XNOR2_X1 U14722 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n11718), .ZN(
        n14813) );
  AOI22_X1 U14723 ( .A1(n12099), .A2(n14813), .B1(n12103), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11719) );
  OAI211_X1 U14724 ( .C1(n11721), .C2(n10100), .A(n11720), .B(n11719), .ZN(
        n14082) );
  OR2_X1 U14725 ( .A1(n11723), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14726 ( .A1(n11724), .A2(n11796), .ZN(n16087) );
  INV_X1 U14727 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14216) );
  INV_X1 U14728 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11725) );
  OAI22_X1 U14729 ( .A1(n12046), .A2(n14216), .B1(n11831), .B2(n11725), .ZN(
        n11726) );
  AOI21_X1 U14730 ( .B1(n16087), .B2(n12099), .A(n11726), .ZN(n14205) );
  AOI22_X1 U14731 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14732 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14733 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14734 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11727) );
  NAND4_X1 U14735 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11736) );
  AOI22_X1 U14736 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14737 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14738 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14739 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11731) );
  NAND4_X1 U14740 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11735) );
  OR2_X1 U14741 ( .A1(n11736), .A2(n11735), .ZN(n11737) );
  NAND2_X1 U14742 ( .A1(n11763), .A2(n11737), .ZN(n14636) );
  INV_X1 U14743 ( .A(n14636), .ZN(n11738) );
  XNOR2_X1 U14744 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11804), .ZN(
        n16071) );
  INV_X1 U14745 ( .A(n16071), .ZN(n11753) );
  AOI22_X1 U14746 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14747 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14748 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14749 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11739) );
  NAND4_X1 U14750 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11748) );
  AOI22_X1 U14751 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14752 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14753 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14754 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11743) );
  NAND4_X1 U14755 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11747) );
  OAI21_X1 U14756 ( .B1(n11748), .B2(n11747), .A(n11763), .ZN(n11751) );
  NAND2_X1 U14757 ( .A1(n11669), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U14758 ( .A1(n12103), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11749) );
  NAND3_X1 U14759 ( .A1(n11751), .A2(n11750), .A3(n11749), .ZN(n11752) );
  AOI21_X1 U14760 ( .B1(n11753), .B2(n12099), .A(n11752), .ZN(n14184) );
  INV_X1 U14761 ( .A(n14184), .ZN(n11802) );
  XNOR2_X1 U14762 ( .A(n11754), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14791) );
  AOI22_X1 U14763 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11180), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14764 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14765 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12087), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14766 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14767 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11765) );
  AOI22_X1 U14768 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12082), .B1(
        n9773), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14769 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14770 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12079), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14771 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11759) );
  NAND4_X1 U14772 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11764) );
  OAI21_X1 U14773 ( .B1(n11765), .B2(n11764), .A(n11763), .ZN(n11768) );
  NAND2_X1 U14774 ( .A1(n11669), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U14775 ( .A1(n12103), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11766) );
  NAND3_X1 U14776 ( .A1(n11768), .A2(n11767), .A3(n11766), .ZN(n11769) );
  AOI21_X1 U14777 ( .B1(n14791), .B2(n12099), .A(n11769), .ZN(n14171) );
  INV_X1 U14778 ( .A(n14171), .ZN(n11801) );
  XNOR2_X1 U14779 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11770), .ZN(
        n15981) );
  AOI22_X1 U14780 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14781 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9772), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14782 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14783 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U14784 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11781) );
  AOI22_X1 U14785 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14786 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14787 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14788 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U14789 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  NOR2_X1 U14790 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  OAI22_X1 U14791 ( .A1(n10100), .A2(n11782), .B1(n11831), .B2(n15975), .ZN(
        n11784) );
  INV_X1 U14792 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13403) );
  NOR2_X1 U14793 ( .A1(n12046), .A2(n13403), .ZN(n11783) );
  NOR2_X1 U14794 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  OAI21_X1 U14795 ( .B1(n15981), .B2(n13901), .A(n11785), .ZN(n14639) );
  AOI22_X1 U14796 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14797 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14798 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14799 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U14800 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11795) );
  AOI22_X1 U14801 ( .A1(n9771), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14802 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14803 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14804 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11790) );
  NAND4_X1 U14805 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11794) );
  NOR2_X1 U14806 ( .A1(n11795), .A2(n11794), .ZN(n11800) );
  NAND2_X1 U14807 ( .A1(n11669), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11799) );
  XNOR2_X1 U14808 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11796), .ZN(
        n16080) );
  INV_X1 U14809 ( .A(n16080), .ZN(n11797) );
  AOI22_X1 U14810 ( .A1(n12103), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12099), .B2(n11797), .ZN(n11798) );
  OAI211_X1 U14811 ( .C1(n11800), .C2(n10100), .A(n11799), .B(n11798), .ZN(
        n14700) );
  AND2_X1 U14812 ( .A1(n14639), .A2(n14700), .ZN(n14170) );
  AOI21_X1 U14813 ( .B1(n11805), .B2(n20907), .A(n11848), .ZN(n14783) );
  OAI21_X1 U14814 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20907), .A(n13901), 
        .ZN(n11806) );
  AOI21_X1 U14815 ( .B1(n11669), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11806), .ZN(
        n11818) );
  AOI22_X1 U14816 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14817 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14818 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14819 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11807) );
  NAND4_X1 U14820 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11816) );
  AOI22_X1 U14821 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14822 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14823 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14824 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11811) );
  NAND4_X1 U14825 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11815) );
  OAI21_X1 U14826 ( .B1(n11816), .B2(n11815), .A(n12096), .ZN(n11817) );
  AOI22_X1 U14827 ( .A1(n14783), .A2(n12099), .B1(n11818), .B2(n11817), .ZN(
        n14192) );
  AOI22_X1 U14828 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14829 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14830 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14831 ( .A1(n9771), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11819) );
  NAND4_X1 U14832 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11828) );
  AOI22_X1 U14833 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14834 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14835 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14836 ( .A1(n9770), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11823) );
  NAND4_X1 U14837 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11827) );
  OR2_X1 U14838 ( .A1(n11828), .A2(n11827), .ZN(n11829) );
  NAND2_X1 U14839 ( .A1(n12096), .A2(n11829), .ZN(n11834) );
  XOR2_X1 U14840 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11848), .Z(
        n16060) );
  INV_X1 U14841 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11830) );
  OAI22_X1 U14842 ( .A1(n16060), .A2(n13901), .B1(n11831), .B2(n11830), .ZN(
        n11832) );
  AOI21_X1 U14843 ( .B1(n11669), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11832), .ZN(
        n11833) );
  NAND2_X1 U14844 ( .A1(n11834), .A2(n11833), .ZN(n15955) );
  AOI22_X1 U14845 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14846 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9770), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14847 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14848 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U14849 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11844) );
  AOI22_X1 U14850 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14851 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U14852 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14853 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11839) );
  NAND4_X1 U14854 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11843) );
  NOR2_X1 U14855 ( .A1(n11844), .A2(n11843), .ZN(n11847) );
  AOI21_X1 U14856 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14772), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11845) );
  AOI21_X1 U14857 ( .B1(n11669), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11845), .ZN(
        n11846) );
  OAI21_X1 U14858 ( .B1(n12074), .B2(n11847), .A(n11846), .ZN(n11850) );
  XNOR2_X1 U14859 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B(n11851), .ZN(
        n14776) );
  NAND2_X1 U14860 ( .A1(n12099), .A2(n14776), .ZN(n11849) );
  OR2_X1 U14861 ( .A1(n11852), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11853) );
  NAND2_X1 U14862 ( .A1(n11853), .A2(n11884), .ZN(n16052) );
  AOI22_X1 U14863 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11132), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14864 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14865 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14866 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11854) );
  NAND4_X1 U14867 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11863) );
  AOI22_X1 U14868 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14869 ( .A1(n9770), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14870 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14871 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11858) );
  NAND4_X1 U14872 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11862) );
  OAI21_X1 U14873 ( .B1(n11863), .B2(n11862), .A(n12096), .ZN(n11866) );
  NAND2_X1 U14874 ( .A1(n11669), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14875 ( .A1(n20525), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11864) );
  NAND4_X1 U14876 ( .A1(n11866), .A2(n13901), .A3(n11865), .A4(n11864), .ZN(
        n11867) );
  OAI21_X1 U14877 ( .B1(n16052), .B2(n13901), .A(n11867), .ZN(n15946) );
  AOI22_X1 U14878 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14879 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14880 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14881 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U14882 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11877) );
  AOI22_X1 U14883 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14884 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14885 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14886 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U14887 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11876) );
  NOR2_X1 U14888 ( .A1(n11877), .A2(n11876), .ZN(n11880) );
  INV_X1 U14889 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15933) );
  AOI21_X1 U14890 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15933), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11878) );
  AOI21_X1 U14891 ( .B1(n11669), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11878), .ZN(
        n11879) );
  OAI21_X1 U14892 ( .B1(n12074), .B2(n11880), .A(n11879), .ZN(n11882) );
  XNOR2_X1 U14893 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11884), .ZN(
        n16040) );
  NAND2_X1 U14894 ( .A1(n16040), .A2(n12099), .ZN(n11881) );
  NAND2_X1 U14895 ( .A1(n11882), .A2(n11881), .ZN(n15937) );
  OR2_X1 U14896 ( .A1(n11885), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11886) );
  NAND2_X1 U14897 ( .A1(n11886), .A2(n11920), .ZN(n16039) );
  AOI22_X1 U14898 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14899 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14900 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14901 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U14902 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11897) );
  AOI22_X1 U14903 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14904 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14905 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14906 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U14907 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11896) );
  NOR2_X1 U14908 ( .A1(n11897), .A2(n11896), .ZN(n11901) );
  INV_X1 U14909 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11898) );
  OAI21_X1 U14910 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n11898), .A(n13901), 
        .ZN(n11899) );
  AOI21_X1 U14911 ( .B1(n11669), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11899), .ZN(
        n11900) );
  OAI21_X1 U14912 ( .B1(n12074), .B2(n11901), .A(n11900), .ZN(n11902) );
  OAI21_X1 U14913 ( .B1(n16039), .B2(n13901), .A(n11902), .ZN(n14626) );
  INV_X1 U14914 ( .A(n14626), .ZN(n11903) );
  AOI22_X1 U14915 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11180), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14916 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11929), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14917 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n9773), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14918 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U14919 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11913) );
  AOI22_X1 U14920 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14921 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12082), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14922 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14923 ( .A1(n9771), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14924 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11912) );
  NOR2_X1 U14925 ( .A1(n11913), .A2(n11912), .ZN(n11917) );
  INV_X1 U14926 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14679) );
  NAND2_X1 U14927 ( .A1(n20525), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11914) );
  OAI211_X1 U14928 ( .C1(n12046), .C2(n14679), .A(n13901), .B(n11914), .ZN(
        n11915) );
  INV_X1 U14929 ( .A(n11915), .ZN(n11916) );
  OAI21_X1 U14930 ( .B1(n12074), .B2(n11917), .A(n11916), .ZN(n11919) );
  XNOR2_X1 U14931 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n11920), .ZN(
        n15913) );
  NAND2_X1 U14932 ( .A1(n15913), .A2(n12099), .ZN(n11918) );
  INV_X1 U14933 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15922) );
  OR2_X1 U14934 ( .A1(n11921), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U14935 ( .A1(n11922), .A2(n11985), .ZN(n16034) );
  AOI22_X1 U14936 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U14937 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14938 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14939 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11924) );
  NAND4_X1 U14940 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11935) );
  AOI22_X1 U14941 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14942 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14943 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14944 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11930) );
  NAND4_X1 U14945 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11934) );
  NOR2_X1 U14946 ( .A1(n11935), .A2(n11934), .ZN(n11953) );
  AOI22_X1 U14947 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U14948 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U14949 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U14950 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11936) );
  NAND4_X1 U14951 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11945) );
  AOI22_X1 U14952 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14953 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U14954 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U14955 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U14956 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11944) );
  NOR2_X1 U14957 ( .A1(n11945), .A2(n11944), .ZN(n11952) );
  XNOR2_X1 U14958 ( .A(n11953), .B(n11952), .ZN(n11948) );
  OAI21_X1 U14959 ( .B1(n20321), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n20525), .ZN(n11947) );
  NAND2_X1 U14960 ( .A1(n11669), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n11946) );
  OAI211_X1 U14961 ( .C1(n12074), .C2(n11948), .A(n11947), .B(n11946), .ZN(
        n11949) );
  OAI21_X1 U14962 ( .B1(n16034), .B2(n13901), .A(n11949), .ZN(n14614) );
  NAND2_X1 U14963 ( .A1(n11951), .A2(n11950), .ZN(n14555) );
  NOR2_X1 U14964 ( .A1(n11953), .A2(n11952), .ZN(n11980) );
  AOI22_X1 U14965 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U14966 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U14967 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U14968 ( .A1(n9770), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11954) );
  NAND4_X1 U14969 ( .A1(n11957), .A2(n11956), .A3(n11955), .A4(n11954), .ZN(
        n11963) );
  AOI22_X1 U14970 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U14971 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U14972 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U14973 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11958) );
  NAND4_X1 U14974 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n11962) );
  OR2_X1 U14975 ( .A1(n11963), .A2(n11962), .ZN(n11979) );
  XNOR2_X1 U14976 ( .A(n11980), .B(n11979), .ZN(n11966) );
  INV_X1 U14977 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14755) );
  OAI21_X1 U14978 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14755), .A(n13901), 
        .ZN(n11964) );
  AOI21_X1 U14979 ( .B1(n11669), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11964), .ZN(
        n11965) );
  OAI21_X1 U14980 ( .B1(n11966), .B2(n12074), .A(n11965), .ZN(n11968) );
  XNOR2_X1 U14981 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n11985), .ZN(
        n14757) );
  NAND2_X1 U14982 ( .A1(n12099), .A2(n14757), .ZN(n11967) );
  NAND2_X1 U14983 ( .A1(n11968), .A2(n11967), .ZN(n14558) );
  NOR2_X2 U14984 ( .A1(n14555), .A2(n14558), .ZN(n14556) );
  AOI22_X1 U14985 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U14986 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U14987 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U14988 ( .A1(n9770), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U14989 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11978) );
  AOI22_X1 U14990 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U14991 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U14992 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U14993 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U14994 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11977) );
  NOR2_X1 U14995 ( .A1(n11978), .A2(n11977), .ZN(n11992) );
  NAND2_X1 U14996 ( .A1(n11980), .A2(n11979), .ZN(n11991) );
  XNOR2_X1 U14997 ( .A(n11992), .B(n11991), .ZN(n11984) );
  INV_X1 U14998 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14663) );
  NAND2_X1 U14999 ( .A1(n20525), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11981) );
  OAI211_X1 U15000 ( .C1(n12046), .C2(n14663), .A(n13901), .B(n11981), .ZN(
        n11982) );
  INV_X1 U15001 ( .A(n11982), .ZN(n11983) );
  OAI21_X1 U15002 ( .B1(n11984), .B2(n12074), .A(n11983), .ZN(n11989) );
  OAI21_X1 U15003 ( .B1(n11987), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n12026), .ZN(n15896) );
  OR2_X1 U15004 ( .A1(n15896), .A2(n13901), .ZN(n11988) );
  NOR2_X1 U15005 ( .A1(n11992), .A2(n11991), .ZN(n12020) );
  AOI22_X1 U15006 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15007 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15008 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15009 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11993) );
  NAND4_X1 U15010 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n12002) );
  AOI22_X1 U15011 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15012 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15013 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15014 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U15015 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  OR2_X1 U15016 ( .A1(n12002), .A2(n12001), .ZN(n12019) );
  INV_X1 U15017 ( .A(n12019), .ZN(n12003) );
  XNOR2_X1 U15018 ( .A(n12020), .B(n12003), .ZN(n12004) );
  NAND2_X1 U15019 ( .A1(n12004), .A2(n12096), .ZN(n12008) );
  INV_X1 U15020 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15891) );
  OAI21_X1 U15021 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15891), .A(n13901), 
        .ZN(n12005) );
  AOI21_X1 U15022 ( .B1(n11669), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12005), .ZN(
        n12007) );
  XNOR2_X1 U15023 ( .A(n12026), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15882) );
  AOI21_X1 U15024 ( .B1(n12008), .B2(n12007), .A(n12006), .ZN(n14597) );
  AOI22_X1 U15025 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15026 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15027 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15028 ( .A1(n9770), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12009) );
  NAND4_X1 U15029 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12018) );
  AOI22_X1 U15030 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15031 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11132), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15032 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15033 ( .A1(n11045), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12013) );
  NAND4_X1 U15034 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12017) );
  NOR2_X1 U15035 ( .A1(n12018), .A2(n12017), .ZN(n12034) );
  NAND2_X1 U15036 ( .A1(n12020), .A2(n12019), .ZN(n12033) );
  XNOR2_X1 U15037 ( .A(n12034), .B(n12033), .ZN(n12025) );
  INV_X1 U15038 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12022) );
  NAND2_X1 U15039 ( .A1(n20525), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12021) );
  OAI211_X1 U15040 ( .C1(n12046), .C2(n12022), .A(n13901), .B(n12021), .ZN(
        n12023) );
  INV_X1 U15041 ( .A(n12023), .ZN(n12024) );
  OAI21_X1 U15042 ( .B1(n12025), .B2(n12074), .A(n12024), .ZN(n12032) );
  INV_X1 U15043 ( .A(n12027), .ZN(n12029) );
  INV_X1 U15044 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U15045 ( .A1(n12029), .A2(n12028), .ZN(n12030) );
  NAND2_X1 U15046 ( .A1(n12054), .A2(n12030), .ZN(n15875) );
  NOR2_X1 U15047 ( .A1(n12034), .A2(n12033), .ZN(n12071) );
  AOI22_X1 U15048 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15049 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15050 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15051 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U15052 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12044) );
  AOI22_X1 U15053 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15054 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15055 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15056 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11045), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15057 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12043) );
  OR2_X1 U15058 ( .A1(n12044), .A2(n12043), .ZN(n12070) );
  XNOR2_X1 U15059 ( .A(n12071), .B(n12070), .ZN(n12049) );
  INV_X1 U15060 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U15061 ( .A1(n20525), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12045) );
  OAI211_X1 U15062 ( .C1(n12046), .C2(n14654), .A(n13901), .B(n12045), .ZN(
        n12047) );
  INV_X1 U15063 ( .A(n12047), .ZN(n12048) );
  OAI21_X1 U15064 ( .B1(n12049), .B2(n12074), .A(n12048), .ZN(n12051) );
  XNOR2_X1 U15065 ( .A(n12054), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14728) );
  NAND2_X1 U15066 ( .A1(n14728), .A2(n12099), .ZN(n12050) );
  NAND2_X1 U15067 ( .A1(n12051), .A2(n12050), .ZN(n14547) );
  INV_X1 U15068 ( .A(n14547), .ZN(n12052) );
  NAND2_X1 U15069 ( .A1(n12053), .A2(n12052), .ZN(n14534) );
  INV_X1 U15070 ( .A(n12054), .ZN(n12055) );
  INV_X1 U15071 ( .A(n12056), .ZN(n12057) );
  INV_X1 U15072 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U15073 ( .A1(n12057), .A2(n14538), .ZN(n12058) );
  NAND2_X1 U15074 ( .A1(n12110), .A2(n12058), .ZN(n14719) );
  AOI22_X1 U15075 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15076 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n9770), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15077 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n9773), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15078 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12082), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12060) );
  NAND4_X1 U15079 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12069) );
  AOI22_X1 U15080 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12081), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15081 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9703), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15082 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15083 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12064) );
  NAND4_X1 U15084 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12068) );
  NOR2_X1 U15085 ( .A1(n12069), .A2(n12068), .ZN(n12078) );
  NAND2_X1 U15086 ( .A1(n12071), .A2(n12070), .ZN(n12077) );
  XNOR2_X1 U15087 ( .A(n12078), .B(n12077), .ZN(n12075) );
  AOI21_X1 U15088 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20525), .A(
        n12099), .ZN(n12073) );
  NAND2_X1 U15089 ( .A1(n11669), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12072) );
  OAI211_X1 U15090 ( .C1(n12075), .C2(n12074), .A(n12073), .B(n12072), .ZN(
        n12076) );
  OAI21_X1 U15091 ( .B1(n13901), .B2(n14719), .A(n12076), .ZN(n14536) );
  NOR2_X1 U15092 ( .A1(n12078), .A2(n12077), .ZN(n12095) );
  AOI22_X1 U15093 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15094 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9771), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15095 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15096 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12083) );
  NAND4_X1 U15097 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12093) );
  AOI22_X1 U15098 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15099 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12087), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15100 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15101 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11052), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12088) );
  NAND4_X1 U15102 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n12092) );
  NOR2_X1 U15103 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  XNOR2_X1 U15104 ( .A(n12095), .B(n12094), .ZN(n12097) );
  NAND2_X1 U15105 ( .A1(n12097), .A2(n12096), .ZN(n12102) );
  INV_X1 U15106 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14713) );
  AOI21_X1 U15107 ( .B1(n14713), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12098) );
  AOI21_X1 U15108 ( .B1(n11669), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12098), .ZN(
        n12101) );
  XNOR2_X1 U15109 ( .A(n12110), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14711) );
  AND2_X1 U15110 ( .A1(n14711), .A2(n12099), .ZN(n12100) );
  AOI21_X1 U15111 ( .B1(n12102), .B2(n12101), .A(n12100), .ZN(n12886) );
  NAND2_X1 U15112 ( .A1(n14535), .A2(n12886), .ZN(n12106) );
  AOI22_X1 U15113 ( .A1(n11669), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12103), .ZN(n12104) );
  INV_X1 U15114 ( .A(n12104), .ZN(n12105) );
  XNOR2_X2 U15115 ( .A(n12106), .B(n12105), .ZN(n14516) );
  AND3_X1 U15116 ( .A1(n16236), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16227) );
  NAND2_X1 U15117 ( .A1(n14516), .A2(n20062), .ZN(n12116) );
  NAND2_X1 U15118 ( .A1(n20530), .A2(n12107), .ZN(n20682) );
  AND2_X1 U15119 ( .A1(n20682), .A2(n16236), .ZN(n12108) );
  NOR2_X1 U15120 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20525), .ZN(n20684) );
  AOI21_X1 U15121 ( .B1(n20321), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n20684), 
        .ZN(n13253) );
  INV_X1 U15122 ( .A(n13253), .ZN(n12109) );
  INV_X1 U15123 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12111) );
  INV_X1 U15124 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20656) );
  NOR2_X1 U15125 ( .A1(n16209), .A2(n20656), .ZN(n14823) );
  AOI21_X1 U15126 ( .B1(n20067), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14823), .ZN(n12113) );
  OAI21_X1 U15127 ( .B1(n20066), .B2(n13916), .A(n12113), .ZN(n12114) );
  OAI211_X1 U15128 ( .C1(n14826), .C2(n19906), .A(n12116), .B(n12115), .ZN(
        P1_U2968) );
  INV_X1 U15129 ( .A(n10717), .ZN(n12117) );
  NAND2_X1 U15130 ( .A1(n19895), .A2(n12117), .ZN(n12162) );
  OAI211_X1 U15131 ( .C1(n13143), .C2(n12124), .A(n13475), .B(n12118), .ZN(
        n12134) );
  INV_X1 U15132 ( .A(n12133), .ZN(n12119) );
  AOI21_X1 U15133 ( .B1(n12134), .B2(n12128), .A(n12119), .ZN(n12120) );
  NAND2_X1 U15134 ( .A1(n12121), .A2(n12120), .ZN(n12122) );
  NAND2_X1 U15135 ( .A1(n12122), .A2(n12828), .ZN(n12136) );
  INV_X1 U15136 ( .A(n14934), .ZN(n14935) );
  AND2_X1 U15137 ( .A1(n12125), .A2(n12124), .ZN(n12126) );
  NOR2_X1 U15138 ( .A1(n12127), .A2(n12126), .ZN(n12131) );
  NAND3_X1 U15139 ( .A1(n12129), .A2(n13143), .A3(n12128), .ZN(n12130) );
  OAI21_X1 U15140 ( .B1(n12828), .B2(n12131), .A(n12130), .ZN(n12132) );
  AOI22_X1 U15141 ( .A1(n14935), .A2(n12134), .B1(n12133), .B2(n12132), .ZN(
        n12135) );
  NAND2_X1 U15142 ( .A1(n12136), .A2(n12135), .ZN(n12141) );
  OAI211_X1 U15143 ( .C1(n12828), .C2(n12138), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n12137), .ZN(n12139) );
  INV_X1 U15144 ( .A(n12139), .ZN(n12140) );
  NAND2_X1 U15145 ( .A1(n12141), .A2(n12140), .ZN(n12143) );
  NOR2_X1 U15146 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19795) );
  AOI211_X1 U15147 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19795), .ZN(n19787) );
  AND2_X1 U15148 ( .A1(n19787), .A2(n13143), .ZN(n12144) );
  NAND2_X1 U15149 ( .A1(n13773), .A2(n12144), .ZN(n13027) );
  NAND2_X1 U15150 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n15862) );
  INV_X1 U15151 ( .A(n15862), .ZN(n19793) );
  INV_X1 U15152 ( .A(n12145), .ZN(n12146) );
  NAND2_X1 U15153 ( .A1(n12147), .A2(n12146), .ZN(n13079) );
  INV_X1 U15154 ( .A(n12185), .ZN(n12151) );
  NAND2_X1 U15155 ( .A1(n10243), .A2(n19215), .ZN(n12149) );
  OAI211_X1 U15156 ( .C1(n13143), .C2(n10242), .A(n12149), .B(n10228), .ZN(
        n12150) );
  AND3_X1 U15157 ( .A1(n12152), .A2(n12151), .A3(n12150), .ZN(n12154) );
  OAI21_X1 U15158 ( .B1(n12153), .B2(n9957), .A(n13491), .ZN(n12180) );
  AND2_X1 U15159 ( .A1(n12154), .A2(n12180), .ZN(n13085) );
  NAND2_X1 U15160 ( .A1(n13773), .A2(n13143), .ZN(n12155) );
  OAI211_X1 U15161 ( .C1(n13773), .C2(n10243), .A(n12155), .B(n15658), .ZN(
        n12159) );
  NOR2_X1 U15162 ( .A1(n13143), .A2(n19787), .ZN(n12156) );
  OAI22_X1 U15163 ( .A1(n13494), .A2(n12156), .B1(n10228), .B2(n13143), .ZN(
        n12157) );
  NOR2_X1 U15164 ( .A1(n19793), .A2(n13476), .ZN(n13082) );
  NAND2_X1 U15165 ( .A1(n12157), .A2(n13082), .ZN(n12158) );
  NAND4_X1 U15166 ( .A1(n12148), .A2(n13085), .A3(n12159), .A4(n12158), .ZN(
        n12160) );
  AOI21_X1 U15167 ( .B1(n10236), .B2(n13079), .A(n12160), .ZN(n12161) );
  INV_X1 U15168 ( .A(n18862), .ZN(n13026) );
  INV_X1 U15169 ( .A(n13491), .ZN(n12163) );
  NOR2_X1 U15170 ( .A1(n10717), .A2(n12163), .ZN(n12164) );
  AND3_X1 U15171 ( .A1(n12214), .A2(n9761), .A3(n10228), .ZN(n12166) );
  AND2_X1 U15172 ( .A1(n12165), .A2(n12166), .ZN(n13470) );
  NAND2_X1 U15173 ( .A1(n12377), .A2(n13470), .ZN(n14244) );
  INV_X1 U15174 ( .A(n15568), .ZN(n15538) );
  INV_X1 U15175 ( .A(n12377), .ZN(n12168) );
  NAND2_X1 U15176 ( .A1(n12168), .A2(n18933), .ZN(n15625) );
  INV_X1 U15177 ( .A(n14244), .ZN(n12169) );
  NOR2_X1 U15178 ( .A1(n10256), .A2(n13097), .ZN(n14241) );
  NOR2_X1 U15179 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14241), .ZN(
        n12195) );
  NAND2_X1 U15180 ( .A1(n12169), .A2(n12195), .ZN(n14236) );
  NAND2_X1 U15181 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14241), .ZN(
        n12196) );
  INV_X1 U15182 ( .A(n12170), .ZN(n12171) );
  NAND2_X1 U15183 ( .A1(n12171), .A2(n10249), .ZN(n13150) );
  NAND2_X1 U15184 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  NAND2_X1 U15185 ( .A1(n12174), .A2(n14934), .ZN(n12175) );
  NAND2_X1 U15186 ( .A1(n12175), .A2(n12185), .ZN(n12178) );
  NAND2_X1 U15187 ( .A1(n14935), .A2(n15658), .ZN(n12177) );
  NAND2_X1 U15188 ( .A1(n10243), .A2(n10236), .ZN(n12176) );
  AND4_X1 U15189 ( .A1(n13150), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12183) );
  NAND2_X1 U15190 ( .A1(n12179), .A2(n13143), .ZN(n13438) );
  NAND2_X1 U15191 ( .A1(n13438), .A2(n12180), .ZN(n12181) );
  NAND2_X1 U15192 ( .A1(n12181), .A2(n15654), .ZN(n12182) );
  AND3_X1 U15193 ( .A1(n12184), .A2(n12183), .A3(n12182), .ZN(n13448) );
  AND2_X1 U15194 ( .A1(n12185), .A2(n10429), .ZN(n12186) );
  NAND2_X1 U15195 ( .A1(n12186), .A2(n10249), .ZN(n13428) );
  NAND2_X1 U15196 ( .A1(n13448), .A2(n13428), .ZN(n12187) );
  AOI21_X1 U15197 ( .B1(n12196), .B2(n14242), .A(n10449), .ZN(n12188) );
  NAND3_X1 U15198 ( .A1(n15625), .A2(n14236), .A3(n12188), .ZN(n14030) );
  NAND2_X1 U15199 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14031) );
  NOR3_X1 U15200 ( .A1(n14033), .A2(n15618), .A3(n14031), .ZN(n16361) );
  NAND2_X1 U15201 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16361), .ZN(
        n12197) );
  NOR2_X1 U15202 ( .A1(n14030), .A2(n12197), .ZN(n15607) );
  INV_X1 U15203 ( .A(n12189), .ZN(n12191) );
  INV_X1 U15204 ( .A(n14242), .ZN(n14240) );
  NAND2_X1 U15205 ( .A1(n15626), .A2(n15625), .ZN(n15599) );
  INV_X1 U15206 ( .A(n15599), .ZN(n12190) );
  AOI21_X1 U15207 ( .B1(n15607), .B2(n12191), .A(n12190), .ZN(n15514) );
  OR2_X1 U15208 ( .A1(n15514), .A2(n12192), .ZN(n12193) );
  AOI211_X1 U15209 ( .C1(n14244), .C2(n12196), .A(n12195), .B(n15626), .ZN(
        n13810) );
  NAND2_X1 U15210 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13810), .ZN(
        n14028) );
  NOR2_X1 U15211 ( .A1(n14028), .A2(n12197), .ZN(n15561) );
  NAND2_X1 U15212 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15561), .ZN(
        n15567) );
  NAND3_X1 U15213 ( .A1(n15568), .A2(n15539), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15214 ( .A1(n10119), .A2(n16357), .B1(n12199), .B2(n15516), .ZN(
        n12200) );
  INV_X1 U15215 ( .A(n15304), .ZN(n12201) );
  NOR2_X1 U15216 ( .A1(n9711), .A2(n12201), .ZN(n12206) );
  INV_X1 U15217 ( .A(n12203), .ZN(n15305) );
  NAND3_X1 U15218 ( .A1(n12204), .A2(n15305), .A3(n15295), .ZN(n12205) );
  OAI21_X1 U15219 ( .B1(n12206), .B2(n12205), .A(n15296), .ZN(n15285) );
  INV_X1 U15220 ( .A(n15282), .ZN(n12207) );
  NOR2_X1 U15221 ( .A1(n15285), .A2(n12207), .ZN(n15274) );
  INV_X1 U15222 ( .A(n12208), .ZN(n12209) );
  OAI21_X1 U15223 ( .B1(n15274), .B2(n12209), .A(n15272), .ZN(n14250) );
  INV_X1 U15224 ( .A(n14249), .ZN(n12211) );
  OAI22_X1 U15225 ( .A1(n14250), .A2(n12211), .B1(n10861), .B2(n12210), .ZN(
        n15201) );
  OAI21_X1 U15226 ( .B1(n12212), .B2(n10861), .A(n15199), .ZN(n15200) );
  XNOR2_X1 U15227 ( .A(n15201), .B(n15200), .ZN(n15252) );
  NOR2_X1 U15228 ( .A1(n10717), .A2(n12828), .ZN(n12213) );
  INV_X1 U15229 ( .A(n13099), .ZN(n12216) );
  INV_X1 U15230 ( .A(n10221), .ZN(n13165) );
  NAND2_X1 U15231 ( .A1(n13165), .A2(n12218), .ZN(n12238) );
  INV_X1 U15232 ( .A(n12229), .ZN(n12219) );
  NAND2_X1 U15233 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19890), .ZN(n19882) );
  NAND2_X1 U15234 ( .A1(n12219), .A2(n19882), .ZN(n12220) );
  AND2_X1 U15235 ( .A1(n12238), .A2(n12220), .ZN(n12221) );
  INV_X1 U15236 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18997) );
  AOI21_X1 U15237 ( .B1(n13143), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U15238 ( .A1(n9957), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12224) );
  OAI211_X1 U15239 ( .C1(n12810), .C2(n18997), .A(n12225), .B(n12224), .ZN(
        n13159) );
  AOI22_X1 U15240 ( .A1(n12226), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12227) );
  OAI21_X1 U15241 ( .B1(n12810), .B2(n12971), .A(n12227), .ZN(n12233) );
  OR2_X1 U15242 ( .A1(n12228), .A2(n12361), .ZN(n12231) );
  AOI22_X1 U15243 ( .A1(n10221), .A2(n12229), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U15244 ( .A1(n12231), .A2(n12230), .ZN(n12969) );
  NOR2_X1 U15245 ( .A1(n12970), .A2(n12969), .ZN(n12235) );
  NOR2_X1 U15246 ( .A1(n12232), .A2(n12233), .ZN(n12234) );
  NOR2_X2 U15247 ( .A1(n12235), .A2(n12234), .ZN(n12241) );
  NAND2_X1 U15248 ( .A1(n12236), .A2(n12237), .ZN(n12239) );
  OAI211_X1 U15249 ( .C1(n19668), .C2(n19871), .A(n12239), .B(n12238), .ZN(
        n12240) );
  XNOR2_X1 U15250 ( .A(n12241), .B(n12240), .ZN(n13313) );
  INV_X1 U15251 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19163) );
  OAI222_X1 U15252 ( .A1(n12800), .A2(n10444), .B1(n12801), .B2(n19163), .C1(
        n12810), .C2(n20696), .ZN(n13312) );
  NOR2_X1 U15253 ( .A1(n13313), .A2(n13312), .ZN(n13311) );
  NOR2_X1 U15254 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  NAND2_X1 U15255 ( .A1(n12838), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15256 ( .A1(n12218), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12246) );
  NAND2_X1 U15257 ( .A1(n12236), .A2(n12243), .ZN(n12245) );
  NAND2_X1 U15258 ( .A1(n12325), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15259 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n13648) );
  AOI22_X1 U15260 ( .A1(n12325), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U15261 ( .A1(n12236), .A2(n12248), .ZN(n12249) );
  OAI211_X1 U15262 ( .C1(n12810), .C2(n12251), .A(n12250), .B(n12249), .ZN(
        n13682) );
  INV_X1 U15263 ( .A(n13682), .ZN(n12252) );
  AOI22_X1 U15264 ( .A1(n12838), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12325), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12256) );
  INV_X1 U15265 ( .A(n12253), .ZN(n12254) );
  AOI22_X1 U15266 ( .A1(n12236), .A2(n12254), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12218), .ZN(n12255) );
  NAND2_X1 U15267 ( .A1(n12256), .A2(n12255), .ZN(n14008) );
  NAND2_X1 U15268 ( .A1(n12236), .A2(n12257), .ZN(n14024) );
  NAND2_X1 U15269 ( .A1(n14007), .A2(n14024), .ZN(n12259) );
  AOI22_X1 U15270 ( .A1(n12325), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12258) );
  OAI21_X1 U15271 ( .B1(n12810), .B2(n10734), .A(n12258), .ZN(n14023) );
  NAND2_X1 U15272 ( .A1(n12259), .A2(n14023), .ZN(n14027) );
  AOI22_X1 U15273 ( .A1(n12325), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12260) );
  OAI21_X1 U15274 ( .B1(n12810), .B2(n10739), .A(n12260), .ZN(n13620) );
  AOI22_X1 U15275 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15276 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15277 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15278 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12261) );
  NAND4_X1 U15279 ( .A1(n12264), .A2(n12263), .A3(n12262), .A4(n12261), .ZN(
        n12271) );
  AOI22_X1 U15280 ( .A1(n12265), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15281 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15282 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15283 ( .A1(n10359), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12266) );
  NAND4_X1 U15284 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12270) );
  OR2_X1 U15285 ( .A1(n12271), .A2(n12270), .ZN(n13302) );
  INV_X1 U15286 ( .A(n13302), .ZN(n19043) );
  AOI22_X1 U15287 ( .A1(n12325), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12272) );
  OAI21_X1 U15288 ( .B1(n12361), .B2(n19043), .A(n12272), .ZN(n12273) );
  AOI21_X1 U15289 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(n12838), .A(n12273), .ZN(
        n13666) );
  AOI22_X1 U15290 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15291 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15292 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15293 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15294 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12283) );
  AOI22_X1 U15295 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15296 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15297 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15298 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15299 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  NAND2_X1 U15300 ( .A1(n12236), .A2(n13305), .ZN(n12285) );
  AOI22_X1 U15301 ( .A1(n12325), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12284) );
  OAI211_X1 U15302 ( .C1(n12810), .C2(n15329), .A(n12285), .B(n12284), .ZN(
        n15600) );
  AOI22_X1 U15303 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15304 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15305 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15306 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12286) );
  NAND4_X1 U15307 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n12286), .ZN(
        n12295) );
  AOI22_X1 U15308 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15309 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15310 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15311 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15312 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12294) );
  NOR2_X1 U15313 ( .A1(n12295), .A2(n12294), .ZN(n19031) );
  INV_X1 U15314 ( .A(n19031), .ZN(n13554) );
  NAND2_X1 U15315 ( .A1(n12236), .A2(n13554), .ZN(n12297) );
  AOI22_X1 U15316 ( .A1(n12325), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12296) );
  OAI211_X1 U15317 ( .C1(n12810), .C2(n12298), .A(n12297), .B(n12296), .ZN(
        n15588) );
  AOI22_X1 U15318 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10396), .B1(
        n10452), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15319 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15320 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15321 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12299) );
  NAND4_X1 U15322 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n12308) );
  AOI22_X1 U15323 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15324 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15325 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15326 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15327 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12307) );
  NOR2_X1 U15328 ( .A1(n12308), .A2(n12307), .ZN(n13721) );
  INV_X1 U15329 ( .A(n13721), .ZN(n12309) );
  NAND2_X1 U15330 ( .A1(n12236), .A2(n12309), .ZN(n12311) );
  AOI22_X1 U15331 ( .A1(n12325), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12310) );
  OAI211_X1 U15332 ( .C1(n12810), .C2(n19811), .A(n12311), .B(n12310), .ZN(
        n15565) );
  AOI22_X1 U15333 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10396), .B1(
        n10452), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15334 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15335 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15336 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12312) );
  NAND4_X1 U15337 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n12321) );
  AOI22_X1 U15338 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15339 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15340 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15341 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U15342 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12320) );
  INV_X1 U15343 ( .A(n13557), .ZN(n12323) );
  AOI22_X1 U15344 ( .A1(n12325), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12322) );
  OAI21_X1 U15345 ( .B1(n12361), .B2(n12323), .A(n12322), .ZN(n12324) );
  AOI21_X1 U15346 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n12838), .A(n12324), 
        .ZN(n13753) );
  AOI22_X1 U15347 ( .A1(n12838), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n12325), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15348 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15349 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15350 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15351 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U15352 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12335) );
  AOI22_X1 U15353 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15354 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15355 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15356 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12330) );
  NAND4_X1 U15357 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12334) );
  AOI22_X1 U15358 ( .A1(n12236), .A2(n19023), .B1(n12218), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U15359 ( .A1(n12337), .A2(n12336), .ZN(n15536) );
  AOI22_X1 U15360 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10396), .B1(
        n10452), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15361 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15362 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15363 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10354), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12338) );
  NAND4_X1 U15364 ( .A1(n12341), .A2(n12340), .A3(n12339), .A4(n12338), .ZN(
        n12347) );
  AOI22_X1 U15365 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n14368), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15366 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10335), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15367 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12265), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15368 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14369), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12342) );
  NAND4_X1 U15369 ( .A1(n12345), .A2(n12344), .A3(n12343), .A4(n12342), .ZN(
        n12346) );
  OR2_X1 U15370 ( .A1(n12347), .A2(n12346), .ZN(n19022) );
  NAND2_X1 U15371 ( .A1(n12236), .A2(n19022), .ZN(n12349) );
  AOI22_X1 U15372 ( .A1(n12325), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12348) );
  OAI211_X1 U15373 ( .C1(n12810), .C2(n19815), .A(n12349), .B(n12348), .ZN(
        n12350) );
  INV_X1 U15374 ( .A(n12350), .ZN(n13820) );
  AOI22_X1 U15375 ( .A1(n12325), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15376 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10396), .B1(
        n10452), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15377 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15378 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15379 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12351) );
  NAND4_X1 U15380 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n12360) );
  AOI22_X1 U15381 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15382 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15383 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15384 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U15385 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12359) );
  NOR2_X1 U15386 ( .A1(n12360), .A2(n12359), .ZN(n13943) );
  OR2_X1 U15387 ( .A1(n12361), .A2(n13943), .ZN(n12362) );
  OAI211_X1 U15388 ( .C1(n12810), .C2(n19817), .A(n12363), .B(n12362), .ZN(
        n15512) );
  AOI22_X1 U15389 ( .A1(n12325), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12364) );
  OAI21_X1 U15390 ( .B1(n12810), .B2(n14142), .A(n12364), .ZN(n14133) );
  AOI22_X1 U15391 ( .A1(n12325), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12365) );
  OAI21_X1 U15392 ( .B1(n12810), .B2(n19819), .A(n12365), .ZN(n12366) );
  OAI21_X1 U15393 ( .B1(n14135), .B2(n12366), .A(n14123), .ZN(n18905) );
  NAND2_X1 U15394 ( .A1(n12368), .A2(n13143), .ZN(n12370) );
  NAND2_X1 U15395 ( .A1(n12165), .A2(n12369), .ZN(n13431) );
  NAND2_X1 U15396 ( .A1(n12370), .A2(n13431), .ZN(n12371) );
  NOR2_X1 U15397 ( .A1(n18905), .A2(n15355), .ZN(n12379) );
  OAI21_X1 U15398 ( .B1(n14138), .B2(n12372), .A(n9819), .ZN(n15253) );
  NAND2_X1 U15399 ( .A1(n12374), .A2(n9761), .ZN(n12375) );
  NAND2_X1 U15400 ( .A1(n12375), .A2(n10266), .ZN(n12376) );
  NAND2_X1 U15401 ( .A1(n18985), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15255) );
  OAI21_X1 U15402 ( .B1(n15253), .B2(n15614), .A(n15255), .ZN(n12378) );
  AOI211_X1 U15403 ( .C1(n15252), .C2(n16359), .A(n12379), .B(n12378), .ZN(
        n12380) );
  INV_X1 U15404 ( .A(n12380), .ZN(n12381) );
  NAND3_X1 U15405 ( .A1(n12385), .A2(n12900), .A3(n11016), .ZN(n12888) );
  OR2_X1 U15406 ( .A1(n12386), .A2(n12387), .ZN(n13273) );
  NAND2_X1 U15407 ( .A1(n12388), .A2(n13904), .ZN(n13510) );
  INV_X1 U15408 ( .A(n20603), .ZN(n20593) );
  OR2_X1 U15409 ( .A1(n12389), .A2(n20593), .ZN(n12390) );
  NAND2_X1 U15410 ( .A1(n13510), .A2(n12390), .ZN(n12391) );
  NAND2_X1 U15411 ( .A1(n12391), .A2(n13537), .ZN(n13268) );
  AND2_X1 U15412 ( .A1(n14695), .A2(n12900), .ZN(n12393) );
  NOR4_X1 U15413 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12398) );
  NOR4_X1 U15414 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12397) );
  NOR4_X1 U15415 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12396) );
  NOR4_X1 U15416 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12395) );
  AND4_X1 U15417 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12403) );
  NOR4_X1 U15418 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12401) );
  NOR4_X1 U15419 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12400) );
  NOR4_X1 U15420 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12399) );
  INV_X1 U15421 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20613) );
  AND4_X1 U15422 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n20613), .ZN(
        n12402) );
  NAND2_X1 U15423 ( .A1(n12403), .A2(n12402), .ZN(n12404) );
  INV_X1 U15424 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19054) );
  NOR2_X1 U15425 ( .A1(n16029), .A2(n19054), .ZN(n12407) );
  AOI22_X1 U15426 ( .A1(n16025), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16022), .ZN(n12405) );
  INV_X1 U15427 ( .A(n12405), .ZN(n12406) );
  NOR2_X1 U15428 ( .A1(n12407), .A2(n12406), .ZN(n12408) );
  NOR2_X2 U15429 ( .A1(n16910), .A2(n12415), .ZN(n12485) );
  INV_X2 U15430 ( .A(n9793), .ZN(n15746) );
  AOI22_X1 U15431 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15433 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12413) );
  NOR2_X2 U15434 ( .A1(n12417), .A2(n12416), .ZN(n17182) );
  NOR2_X2 U15435 ( .A1(n16910), .A2(n12418), .ZN(n12484) );
  AOI22_X1 U15436 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12484), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15437 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12411) );
  NAND4_X1 U15438 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n12426) );
  OR2_X2 U15439 ( .A1(n18657), .A2(n12418), .ZN(n12571) );
  INV_X2 U15440 ( .A(n12571), .ZN(n17108) );
  AOI22_X1 U15441 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12424) );
  INV_X2 U15442 ( .A(n15706), .ZN(n17123) );
  AOI22_X1 U15443 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12423) );
  INV_X2 U15444 ( .A(n9791), .ZN(n17152) );
  AOI22_X1 U15445 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12422) );
  NOR2_X2 U15446 ( .A1(n12418), .A2(n12419), .ZN(n12462) );
  BUF_X4 U15447 ( .A(n9697), .Z(n17181) );
  AOI22_X1 U15448 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12421) );
  NAND4_X1 U15449 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12425) );
  AOI22_X1 U15450 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15451 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12436) );
  INV_X1 U15452 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n20736) );
  AOI22_X1 U15453 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12427) );
  OAI21_X1 U15454 ( .B1(n17093), .B2(n20736), .A(n12427), .ZN(n12434) );
  AOI22_X1 U15455 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12432) );
  INV_X2 U15456 ( .A(n16878), .ZN(n17173) );
  AOI22_X1 U15457 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15458 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12430) );
  INV_X1 U15459 ( .A(n12461), .ZN(n15727) );
  AOI22_X1 U15460 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12429) );
  NAND4_X1 U15461 ( .A1(n12432), .A2(n12431), .A3(n12430), .A4(n12429), .ZN(
        n12433) );
  AOI211_X1 U15462 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n12434), .B(n12433), .ZN(n12435) );
  NAND3_X1 U15463 ( .A1(n12437), .A2(n12436), .A3(n12435), .ZN(n12677) );
  INV_X2 U15464 ( .A(n9791), .ZN(n17185) );
  AOI22_X1 U15465 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15466 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12446) );
  BUF_X4 U15467 ( .A(n12462), .Z(n17151) );
  INV_X1 U15468 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U15469 ( .A1(n12484), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12438) );
  OAI21_X1 U15470 ( .B1(n12410), .B2(n20884), .A(n12438), .ZN(n12444) );
  AOI22_X1 U15471 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15472 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15473 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12464), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15474 ( .A1(n9697), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12572), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12439) );
  NAND4_X1 U15475 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12443) );
  AOI211_X1 U15476 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n12444), .B(n12443), .ZN(n12445) );
  NAND3_X1 U15477 ( .A1(n12447), .A2(n12446), .A3(n12445), .ZN(n17362) );
  AOI22_X1 U15478 ( .A1(n12485), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15479 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15480 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15481 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12448) );
  NAND4_X1 U15482 ( .A1(n12451), .A2(n12450), .A3(n12449), .A4(n12448), .ZN(
        n12457) );
  AOI22_X1 U15483 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15484 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12461), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15485 ( .A1(n12503), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12464), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15486 ( .A1(n12484), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12572), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15487 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12456) );
  AOI22_X1 U15488 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12484), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n12485), .ZN(n12460) );
  AOI22_X1 U15489 ( .A1(n12503), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12477), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12459) );
  NAND3_X1 U15490 ( .A1(n12460), .A2(n12459), .A3(n12458), .ZN(n12472) );
  AOI22_X1 U15491 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17159), .ZN(n12468) );
  AOI22_X1 U15492 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12461), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15493 ( .A1(n12463), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12572), .ZN(n12466) );
  AOI22_X1 U15494 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n12549), .ZN(n12465) );
  NAND4_X1 U15495 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(
        n12471) );
  INV_X1 U15496 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U15497 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12428), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12469) );
  OAI21_X1 U15498 ( .B1(n20719), .B2(n9793), .A(n12469), .ZN(n12470) );
  AOI22_X1 U15499 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15500 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15501 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15502 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12473) );
  NAND4_X1 U15503 ( .A1(n12476), .A2(n12475), .A3(n12474), .A4(n12473), .ZN(
        n12483) );
  AOI22_X1 U15504 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12481) );
  INV_X2 U15505 ( .A(n15706), .ZN(n17183) );
  AOI22_X1 U15506 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15507 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15508 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12478) );
  NAND4_X1 U15509 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12482) );
  INV_X2 U15510 ( .A(n12571), .ZN(n17172) );
  AOI22_X1 U15511 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15512 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12494) );
  INV_X1 U15513 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U15514 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12486) );
  OAI21_X1 U15515 ( .B1(n16878), .B2(n17198), .A(n12486), .ZN(n12492) );
  AOI22_X1 U15516 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15517 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15518 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15519 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12487) );
  NAND4_X1 U15520 ( .A1(n12490), .A2(n12489), .A3(n12488), .A4(n12487), .ZN(
        n12491) );
  AOI211_X1 U15521 ( .C1(n17161), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12492), .B(n12491), .ZN(n12493) );
  NAND2_X1 U15522 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17603), .ZN(
        n12548) );
  OAI21_X1 U15523 ( .B1(n16416), .B2(n16417), .A(n17770), .ZN(n12526) );
  INV_X1 U15524 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U15525 ( .A1(n12461), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12497) );
  OAI21_X1 U15526 ( .B1(n17093), .B2(n20872), .A(n12497), .ZN(n12498) );
  INV_X1 U15527 ( .A(n12498), .ZN(n12510) );
  AOI22_X1 U15528 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U15529 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15530 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15531 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15532 ( .A1(n12484), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12572), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15533 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12507) );
  AOI22_X1 U15534 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U15535 ( .A1(n12505), .A2(n12504), .ZN(n12506) );
  NOR2_X1 U15536 ( .A1(n12507), .A2(n12506), .ZN(n12508) );
  NAND3_X1 U15537 ( .A1(n12510), .A2(n12509), .A3(n12508), .ZN(n17869) );
  INV_X1 U15538 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18799) );
  INV_X1 U15539 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18156) );
  NOR2_X1 U15540 ( .A1(n18156), .A2(n12513), .ZN(n12514) );
  XNOR2_X1 U15541 ( .A(n17362), .B(n12515), .ZN(n17842) );
  NOR2_X1 U15542 ( .A1(n17841), .A2(n17842), .ZN(n12516) );
  NAND2_X1 U15543 ( .A1(n17841), .A2(n17842), .ZN(n17840) );
  OAI21_X1 U15544 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n12516), .A(
        n17840), .ZN(n17825) );
  XNOR2_X1 U15545 ( .A(n17359), .B(n12517), .ZN(n12518) );
  XNOR2_X1 U15546 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12518), .ZN(
        n17826) );
  NOR2_X1 U15547 ( .A1(n17825), .A2(n17826), .ZN(n17824) );
  NOR2_X2 U15548 ( .A1(n17824), .A2(n12519), .ZN(n12522) );
  XOR2_X1 U15549 ( .A(n12677), .B(n12520), .Z(n12521) );
  INV_X1 U15550 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17815) );
  XNOR2_X1 U15551 ( .A(n12522), .B(n12521), .ZN(n17814) );
  XNOR2_X1 U15552 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12524), .ZN(
        n17800) );
  XNOR2_X1 U15553 ( .A(n12526), .B(n12527), .ZN(n17793) );
  INV_X1 U15554 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17794) );
  NOR2_X1 U15555 ( .A1(n17793), .A2(n17794), .ZN(n17792) );
  NOR2_X1 U15556 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  INV_X1 U15557 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18092) );
  INV_X1 U15558 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18074) );
  NOR2_X1 U15559 ( .A1(n18092), .A2(n18074), .ZN(n17740) );
  NAND2_X1 U15560 ( .A1(n17740), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18039) );
  INV_X1 U15561 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18059) );
  NOR2_X1 U15562 ( .A1(n18039), .A2(n18059), .ZN(n18022) );
  NAND2_X1 U15563 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17674) );
  INV_X1 U15564 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18003) );
  NAND2_X1 U15565 ( .A1(n12724), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12532) );
  NOR2_X1 U15566 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17755) );
  NOR4_X1 U15567 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12530) );
  INV_X1 U15568 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18020) );
  NAND2_X1 U15569 ( .A1(n12532), .A2(n12531), .ZN(n17649) );
  NAND2_X1 U15570 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17645) );
  NOR2_X1 U15571 ( .A1(n17563), .A2(n17602), .ZN(n17604) );
  INV_X1 U15572 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17636) );
  INV_X1 U15573 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17945) );
  NAND2_X1 U15574 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17939) );
  NOR3_X1 U15575 ( .A1(n17636), .A2(n17945), .A3(n17939), .ZN(n17582) );
  NAND2_X1 U15576 ( .A1(n17582), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12729) );
  NOR2_X1 U15577 ( .A1(n17645), .A2(n12729), .ZN(n16412) );
  NAND2_X1 U15578 ( .A1(n16412), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12723) );
  NAND2_X1 U15579 ( .A1(n17636), .A2(n17770), .ZN(n17635) );
  NOR2_X1 U15580 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17635), .ZN(
        n12534) );
  INV_X1 U15581 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17936) );
  NAND2_X1 U15582 ( .A1(n12534), .A2(n17936), .ZN(n17605) );
  INV_X1 U15583 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17942) );
  INV_X1 U15584 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17922) );
  NAND3_X1 U15585 ( .A1(n17583), .A2(n17942), .A3(n17922), .ZN(n12535) );
  INV_X1 U15586 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17556) );
  NAND2_X1 U15587 ( .A1(n17554), .A2(n17556), .ZN(n17553) );
  NAND3_X1 U15588 ( .A1(n17562), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17553), .ZN(n12539) );
  INV_X1 U15589 ( .A(n12539), .ZN(n17542) );
  INV_X1 U15590 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20775) );
  NAND2_X1 U15591 ( .A1(n17770), .A2(n17553), .ZN(n17541) );
  OAI21_X1 U15592 ( .B1(n17542), .B2(n20775), .A(n12538), .ZN(n17524) );
  NOR2_X2 U15593 ( .A1(n17524), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17523) );
  NAND2_X1 U15594 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17880) );
  OAI21_X1 U15595 ( .B1(n12539), .B2(n17880), .A(n17603), .ZN(n12540) );
  INV_X1 U15596 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16400) );
  NAND2_X1 U15597 ( .A1(n15775), .A2(n16400), .ZN(n15835) );
  AOI21_X1 U15598 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12544), .A(
        n17603), .ZN(n12543) );
  NAND2_X1 U15599 ( .A1(n12542), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17512) );
  INV_X1 U15600 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17500) );
  NAND2_X1 U15601 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15776), .ZN(
        n15834) );
  NAND2_X1 U15602 ( .A1(n17603), .A2(n15834), .ZN(n12545) );
  OAI21_X1 U15603 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12543), .A(
        n12545), .ZN(n12547) );
  INV_X1 U15604 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18798) );
  INV_X1 U15605 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16394) );
  AOI21_X2 U15606 ( .B1(n12548), .B2(n12547), .A(n12546), .ZN(n12869) );
  AOI22_X1 U15607 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15608 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15609 ( .A1(n15746), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12551) );
  BUF_X2 U15610 ( .A(n12549), .Z(n17154) );
  AOI22_X1 U15611 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17154), .ZN(n12550) );
  NAND4_X1 U15612 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12559) );
  BUF_X4 U15613 ( .A(n12464), .Z(n17153) );
  AOI22_X1 U15614 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15615 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15616 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17176), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17172), .ZN(n12555) );
  AOI22_X1 U15617 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12484), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12554) );
  NAND4_X1 U15618 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12558) );
  AOI22_X1 U15619 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15620 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12568) );
  INV_X1 U15621 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U15622 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12560) );
  OAI21_X1 U15623 ( .B1(n12571), .B2(n20827), .A(n12560), .ZN(n12566) );
  AOI22_X1 U15624 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15625 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15626 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15627 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U15628 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12565) );
  NOR2_X1 U15629 ( .A1(n18206), .A2(n18209), .ZN(n12670) );
  AOI22_X1 U15630 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15631 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15632 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12570) );
  OAI21_X1 U15633 ( .B1(n15727), .B2(n20874), .A(n12570), .ZN(n12578) );
  AOI22_X1 U15634 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15635 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15636 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15637 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12573) );
  NAND4_X1 U15638 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12577) );
  AOI211_X1 U15639 ( .C1(n17161), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12578), .B(n12577), .ZN(n12579) );
  NAND3_X1 U15640 ( .A1(n12581), .A2(n12580), .A3(n12579), .ZN(n18227) );
  AND2_X1 U15641 ( .A1(n12670), .A2(n18227), .ZN(n12669) );
  AOI22_X1 U15642 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15643 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15644 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15645 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12582) );
  NAND4_X1 U15646 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12591) );
  AOI22_X1 U15647 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15648 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15649 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15650 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U15651 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12590) );
  AOI22_X1 U15652 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15653 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15654 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15655 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15656 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12601) );
  AOI22_X1 U15657 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15658 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15659 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15660 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12596) );
  NAND4_X1 U15661 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  AOI22_X1 U15662 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15663 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15664 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15665 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12602) );
  NAND4_X1 U15666 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n12602), .ZN(
        n12611) );
  AOI22_X1 U15667 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15668 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15669 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15670 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12606) );
  NAND4_X1 U15671 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12610) );
  AOI22_X1 U15672 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15673 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15674 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15675 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12612) );
  NAND4_X1 U15676 ( .A1(n12615), .A2(n12614), .A3(n12613), .A4(n12612), .ZN(
        n12621) );
  AOI22_X1 U15677 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15678 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12484), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15679 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15680 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12616) );
  NAND4_X1 U15681 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        n12620) );
  INV_X1 U15682 ( .A(n12711), .ZN(n18223) );
  NOR2_X1 U15683 ( .A1(n17235), .A2(n18223), .ZN(n12708) );
  AOI22_X1 U15684 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15685 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15686 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15687 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12622) );
  NAND4_X1 U15688 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12631) );
  AOI22_X1 U15689 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15690 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U15691 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15692 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12626) );
  NAND4_X1 U15693 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12626), .ZN(
        n12630) );
  NOR2_X1 U15694 ( .A1(n12708), .A2(n12660), .ZN(n12632) );
  OAI211_X1 U15695 ( .C1(n18218), .C2(n18664), .A(n12721), .B(n12632), .ZN(
        n12633) );
  INV_X1 U15696 ( .A(n12633), .ZN(n12667) );
  NAND2_X1 U15697 ( .A1(n12669), .A2(n12667), .ZN(n18636) );
  NAND2_X1 U15698 ( .A1(n18668), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12641) );
  OAI21_X1 U15699 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18668), .A(
        n12641), .ZN(n12652) );
  INV_X1 U15700 ( .A(n12652), .ZN(n12651) );
  AOI22_X1 U15701 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20932), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12634), .ZN(n12642) );
  AOI22_X1 U15702 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18674), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18807), .ZN(n12643) );
  INV_X1 U15703 ( .A(n12642), .ZN(n12653) );
  NAND2_X1 U15704 ( .A1(n12643), .A2(n12644), .ZN(n12637) );
  NAND2_X1 U15705 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12638), .ZN(
        n12645) );
  OAI22_X1 U15706 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18678), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12638), .ZN(n12647) );
  AOI21_X1 U15707 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12645), .A(
        n12647), .ZN(n12639) );
  NAND2_X1 U15708 ( .A1(n12642), .A2(n12641), .ZN(n12640) );
  OAI211_X1 U15709 ( .C1(n12642), .C2(n12641), .A(n12648), .B(n12640), .ZN(
        n12672) );
  XNOR2_X1 U15710 ( .A(n12644), .B(n12643), .ZN(n12650) );
  NOR2_X1 U15711 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18678), .ZN(
        n12646) );
  AOI22_X1 U15712 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12647), .B1(
        n12646), .B2(n12645), .ZN(n12655) );
  INV_X1 U15713 ( .A(n12655), .ZN(n12649) );
  OAI21_X1 U15714 ( .B1(n12651), .B2(n12672), .A(n12673), .ZN(n18635) );
  NOR2_X2 U15715 ( .A1(n12711), .A2(n17235), .ZN(n12662) );
  NAND2_X1 U15716 ( .A1(n12657), .A2(n12662), .ZN(n12658) );
  NOR2_X1 U15717 ( .A1(n12653), .A2(n12652), .ZN(n12654) );
  AOI21_X1 U15718 ( .B1(n12655), .B2(n12654), .A(n12673), .ZN(n18634) );
  INV_X1 U15719 ( .A(n18634), .ZN(n15763) );
  AOI21_X1 U15720 ( .B1(n18218), .B2(n12658), .A(n15763), .ZN(n12668) );
  NAND2_X1 U15721 ( .A1(n18203), .A2(n17280), .ZN(n12709) );
  INV_X1 U15722 ( .A(n12709), .ZN(n12656) );
  NAND3_X1 U15723 ( .A1(n12657), .A2(n18218), .A3(n17235), .ZN(n12710) );
  NAND2_X1 U15724 ( .A1(n12710), .A2(n12658), .ZN(n12666) );
  AOI22_X1 U15725 ( .A1(n12709), .A2(n12707), .B1(n18218), .B2(n18664), .ZN(
        n12659) );
  INV_X1 U15726 ( .A(n12659), .ZN(n12665) );
  NOR2_X1 U15727 ( .A1(n18236), .A2(n12662), .ZN(n12663) );
  INV_X1 U15728 ( .A(n12660), .ZN(n12661) );
  OAI22_X1 U15729 ( .A1(n18218), .A2(n12663), .B1(n12662), .B2(n12661), .ZN(
        n12664) );
  OAI211_X1 U15730 ( .C1(n18236), .C2(n18664), .A(n16540), .B(n18206), .ZN(
        n12715) );
  OAI211_X1 U15731 ( .C1(n12712), .C2(n12667), .A(n12718), .B(n12715), .ZN(
        n15759) );
  AOI21_X1 U15732 ( .B1(n18206), .B2(n18209), .A(n12670), .ZN(n12671) );
  INV_X1 U15733 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18719) );
  INV_X2 U15734 ( .A(n18849), .ZN(n18848) );
  OAI211_X1 U15735 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18719), .B(n18776), .ZN(n18833) );
  NAND2_X1 U15736 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18844) );
  INV_X1 U15737 ( .A(n18844), .ZN(n18837) );
  AOI21_X1 U15738 ( .B1(n12671), .B2(n18833), .A(n18837), .ZN(n16519) );
  NOR2_X1 U15739 ( .A1(n12711), .A2(n18209), .ZN(n12717) );
  INV_X1 U15740 ( .A(n12717), .ZN(n12674) );
  NAND2_X1 U15741 ( .A1(n12673), .A2(n12672), .ZN(n18632) );
  NAND3_X1 U15742 ( .A1(n16519), .A2(n12674), .A3(n18632), .ZN(n12675) );
  NAND3_X1 U15743 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(n18800), .ZN(n18692) );
  NAND2_X1 U15744 ( .A1(n16418), .A2(n18182), .ZN(n18188) );
  NOR2_X2 U15745 ( .A1(n10049), .A2(n18188), .ZN(n18089) );
  NAND2_X1 U15746 ( .A1(n12869), .A2(n18089), .ZN(n12743) );
  NAND2_X1 U15747 ( .A1(n17869), .A2(n12511), .ZN(n12679) );
  NAND2_X1 U15748 ( .A1(n17367), .A2(n12679), .ZN(n12678) );
  NAND2_X1 U15749 ( .A1(n12678), .A2(n17362), .ZN(n12688) );
  NOR2_X1 U15750 ( .A1(n17359), .A2(n12688), .ZN(n12692) );
  NAND2_X1 U15751 ( .A1(n12692), .A2(n12677), .ZN(n12694) );
  NOR2_X1 U15752 ( .A1(n17353), .A2(n12694), .ZN(n12698) );
  NAND2_X1 U15753 ( .A1(n12698), .A2(n16417), .ZN(n12699) );
  INV_X1 U15754 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18140) );
  XNOR2_X1 U15755 ( .A(n12678), .B(n17362), .ZN(n12685) );
  NOR2_X1 U15756 ( .A1(n18140), .A2(n12685), .ZN(n12686) );
  XOR2_X1 U15757 ( .A(n17367), .B(n12679), .Z(n12682) );
  NOR2_X1 U15758 ( .A1(n12682), .A2(n18156), .ZN(n12684) );
  INV_X1 U15759 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18818) );
  NOR2_X1 U15760 ( .A1(n12496), .A2(n18818), .ZN(n12681) );
  INV_X1 U15761 ( .A(n17869), .ZN(n17859) );
  NAND3_X1 U15762 ( .A1(n17859), .A2(n12496), .A3(n18818), .ZN(n12680) );
  OAI221_X1 U15763 ( .B1(n12681), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17859), .C2(n12496), .A(n12680), .ZN(n17853) );
  XNOR2_X1 U15764 ( .A(n18156), .B(n12682), .ZN(n17852) );
  NOR2_X1 U15765 ( .A1(n17853), .A2(n17852), .ZN(n12683) );
  NOR2_X1 U15766 ( .A1(n12684), .A2(n12683), .ZN(n17838) );
  XNOR2_X1 U15767 ( .A(n18140), .B(n12685), .ZN(n17837) );
  INV_X1 U15768 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12726) );
  NOR2_X1 U15769 ( .A1(n12689), .A2(n12726), .ZN(n12690) );
  XOR2_X1 U15770 ( .A(n12688), .B(n12687), .Z(n17823) );
  XNOR2_X1 U15771 ( .A(n12726), .B(n12689), .ZN(n17822) );
  NOR2_X2 U15772 ( .A1(n12690), .A2(n17821), .ZN(n12691) );
  NOR2_X1 U15773 ( .A1(n12691), .A2(n17815), .ZN(n12693) );
  XNOR2_X1 U15774 ( .A(n17815), .B(n12691), .ZN(n17812) );
  XOR2_X1 U15775 ( .A(n12692), .B(n17356), .Z(n17811) );
  XNOR2_X1 U15776 ( .A(n12694), .B(n17353), .ZN(n12696) );
  NOR2_X1 U15777 ( .A1(n12695), .A2(n12696), .ZN(n12697) );
  INV_X1 U15778 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18124) );
  XNOR2_X1 U15779 ( .A(n12696), .B(n12695), .ZN(n17804) );
  XNOR2_X1 U15780 ( .A(n12698), .B(n16417), .ZN(n12701) );
  NAND2_X1 U15781 ( .A1(n12700), .A2(n12701), .ZN(n17789) );
  INV_X1 U15782 ( .A(n12699), .ZN(n12704) );
  OR2_X1 U15783 ( .A1(n12701), .A2(n12700), .ZN(n17790) );
  OAI21_X1 U15784 ( .B1(n12704), .B2(n12703), .A(n17790), .ZN(n12702) );
  INV_X1 U15785 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18103) );
  NAND3_X1 U15786 ( .A1(n18022), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17998) );
  NAND2_X1 U15787 ( .A1(n17920), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17538) );
  NAND3_X1 U15788 ( .A1(n17877), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16421) );
  NAND2_X1 U15789 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15772), .ZN(
        n12706) );
  XOR2_X1 U15790 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12706), .Z(
        n12882) );
  XOR2_X1 U15791 ( .A(n18206), .B(n18203), .Z(n18854) );
  NOR2_X1 U15792 ( .A1(n18218), .A2(n18227), .ZN(n18648) );
  NAND3_X1 U15793 ( .A1(n12721), .A2(n12717), .A3(n18648), .ZN(n15764) );
  INV_X1 U15794 ( .A(n12707), .ZN(n18214) );
  NOR2_X1 U15795 ( .A1(n18214), .A2(n18209), .ZN(n18647) );
  NAND2_X1 U15796 ( .A1(n18647), .A2(n12708), .ZN(n14220) );
  NOR2_X1 U15797 ( .A1(n12709), .A2(n14220), .ZN(n12714) );
  INV_X1 U15798 ( .A(n12720), .ZN(n12722) );
  OAI21_X1 U15799 ( .B1(n12717), .B2(n12716), .A(n12715), .ZN(n12719) );
  NOR2_X1 U15800 ( .A1(n18206), .A2(n12721), .ZN(n18646) );
  NOR2_X1 U15801 ( .A1(n18647), .A2(n18646), .ZN(n12727) );
  NOR2_X4 U15802 ( .A1(n18835), .A2(n18100), .ZN(n18630) );
  NAND2_X1 U15803 ( .A1(n18630), .A2(n18182), .ZN(n18190) );
  INV_X1 U15804 ( .A(n12723), .ZN(n17555) );
  NAND2_X1 U15805 ( .A1(n17555), .A2(n17579), .ZN(n17917) );
  NAND3_X1 U15806 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n17883), .ZN(n16420) );
  NOR2_X1 U15807 ( .A1(n16400), .A2(n16420), .ZN(n15771) );
  NAND2_X1 U15808 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15771), .ZN(
        n12725) );
  XNOR2_X1 U15809 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12725), .ZN(
        n12880) );
  NOR2_X1 U15810 ( .A1(n16417), .A2(n18188), .ZN(n18107) );
  NOR2_X1 U15811 ( .A1(n17998), .A2(n18020), .ZN(n17662) );
  NAND2_X1 U15812 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18099) );
  OR2_X1 U15813 ( .A1(n18103), .A2(n18099), .ZN(n18010) );
  NOR3_X1 U15814 ( .A1(n17815), .A2(n18140), .A3(n12726), .ZN(n17984) );
  OAI21_X1 U15815 ( .B1(n18818), .B2(n18799), .A(n18156), .ZN(n18137) );
  NAND2_X1 U15816 ( .A1(n17984), .A2(n18137), .ZN(n18096) );
  NOR2_X1 U15817 ( .A1(n18010), .A2(n18096), .ZN(n18085) );
  NAND2_X1 U15818 ( .A1(n17662), .A2(n18085), .ZN(n12728) );
  NAND3_X1 U15819 ( .A1(n9801), .A2(n12727), .A3(n18650), .ZN(n18095) );
  OAI21_X1 U15820 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18642), .A(
        n18095), .ZN(n18165) );
  NOR2_X1 U15821 ( .A1(n18156), .A2(n18799), .ZN(n18138) );
  NAND2_X1 U15822 ( .A1(n18138), .A2(n17984), .ZN(n18094) );
  NOR2_X1 U15823 ( .A1(n18094), .A2(n18010), .ZN(n17997) );
  NAND2_X1 U15824 ( .A1(n17997), .A2(n17662), .ZN(n17977) );
  OAI22_X1 U15825 ( .A1(n18644), .A2(n12728), .B1(n18165), .B2(n17977), .ZN(
        n16410) );
  NAND2_X1 U15826 ( .A1(n16412), .A2(n16410), .ZN(n17904) );
  INV_X1 U15827 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17887) );
  NOR2_X1 U15828 ( .A1(n17922), .A2(n17556), .ZN(n17879) );
  NAND2_X1 U15829 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17879), .ZN(
        n17876) );
  INV_X1 U15830 ( .A(n17876), .ZN(n17893) );
  NAND2_X1 U15831 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17893), .ZN(
        n12733) );
  NOR2_X1 U15832 ( .A1(n17887), .A2(n12733), .ZN(n12730) );
  NAND2_X1 U15833 ( .A1(n18182), .A2(n12730), .ZN(n16413) );
  NOR3_X1 U15834 ( .A1(n17500), .A2(n17904), .A3(n16413), .ZN(n15769) );
  NOR3_X1 U15835 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16394), .A3(
        n16400), .ZN(n12737) );
  INV_X1 U15836 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18773) );
  NAND2_X1 U15837 ( .A1(n18800), .A2(n18789), .ZN(n18803) );
  NOR2_X1 U15838 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18803), .ZN(n18851) );
  INV_X1 U15839 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18840) );
  NOR2_X1 U15840 ( .A1(n18773), .A2(n18184), .ZN(n12877) );
  NAND2_X1 U15841 ( .A1(n18100), .A2(n18182), .ZN(n18171) );
  INV_X1 U15842 ( .A(n18171), .ZN(n15774) );
  NAND3_X1 U15843 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16385) );
  INV_X1 U15844 ( .A(n17645), .ZN(n17980) );
  INV_X1 U15845 ( .A(n12728), .ZN(n17935) );
  NAND2_X1 U15846 ( .A1(n17980), .A2(n17935), .ZN(n17982) );
  NOR2_X1 U15847 ( .A1(n12729), .A2(n17982), .ZN(n17921) );
  AOI21_X1 U15848 ( .B1(n17879), .B2(n17921), .A(n18644), .ZN(n17902) );
  AOI21_X1 U15849 ( .B1(n18661), .B2(n17880), .A(n17902), .ZN(n17881) );
  INV_X1 U15850 ( .A(n12730), .ZN(n12731) );
  INV_X1 U15851 ( .A(n16412), .ZN(n17566) );
  NOR2_X1 U15852 ( .A1(n17566), .A2(n17977), .ZN(n12732) );
  NAND2_X1 U15853 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12732), .ZN(
        n17941) );
  OAI21_X1 U15854 ( .B1(n12731), .B2(n17941), .A(n18663), .ZN(n12735) );
  INV_X1 U15855 ( .A(n12732), .ZN(n17878) );
  OAI21_X1 U15856 ( .B1(n12733), .B2(n17878), .A(n18642), .ZN(n12734) );
  NAND4_X1 U15857 ( .A1(n17881), .A2(n18141), .A3(n12735), .A4(n12734), .ZN(
        n15770) );
  AOI22_X1 U15858 ( .A1(n15774), .A2(n16385), .B1(n18184), .B2(n15770), .ZN(
        n15841) );
  AOI221_X1 U15859 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15841), 
        .C1(n18171), .C2(n15841), .A(n18798), .ZN(n12736) );
  AOI211_X1 U15860 ( .C1(n15769), .C2(n12737), .A(n12877), .B(n12736), .ZN(
        n12738) );
  INV_X1 U15861 ( .A(n12738), .ZN(n12739) );
  INV_X1 U15862 ( .A(n12741), .ZN(n12742) );
  NAND2_X1 U15863 ( .A1(n12743), .A2(n12742), .ZN(P3_U2831) );
  OAI21_X1 U15864 ( .B1(n12746), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n12747), .ZN(n15265) );
  INV_X1 U15865 ( .A(n15265), .ZN(n14147) );
  INV_X1 U15866 ( .A(n12748), .ZN(n12768) );
  AND2_X1 U15867 ( .A1(n12768), .A2(n15287), .ZN(n12750) );
  OR2_X1 U15868 ( .A1(n12750), .A2(n12749), .ZN(n13830) );
  INV_X1 U15869 ( .A(n13830), .ZN(n15290) );
  OR2_X1 U15870 ( .A1(n12752), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12753) );
  AND2_X1 U15871 ( .A1(n12751), .A2(n12753), .ZN(n15307) );
  OAI21_X1 U15872 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12754), .A(
        n12755), .ZN(n16328) );
  INV_X1 U15873 ( .A(n16328), .ZN(n18949) );
  AOI21_X1 U15874 ( .B1(n16342), .B2(n12756), .A(n12757), .ZN(n16329) );
  INV_X1 U15875 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16350) );
  INV_X1 U15876 ( .A(n12758), .ZN(n12762) );
  AND2_X1 U15877 ( .A1(n12758), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12764) );
  AOI21_X1 U15878 ( .B1(n16350), .B2(n12762), .A(n12764), .ZN(n18976) );
  INV_X1 U15879 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20984) );
  NOR2_X1 U15880 ( .A1(n20984), .A2(n12759), .ZN(n12763) );
  AOI21_X1 U15881 ( .B1(n20984), .B2(n12759), .A(n12763), .ZN(n13932) );
  AOI21_X1 U15882 ( .B1(n13071), .B2(n12760), .A(n12761), .ZN(n20693) );
  AOI22_X1 U15883 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16380), .ZN(n13786) );
  AOI22_X1 U15884 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13071), .B2(n16380), .ZN(
        n13785) );
  NAND2_X1 U15885 ( .A1(n13786), .A2(n13785), .ZN(n20691) );
  NOR2_X1 U15886 ( .A1(n20693), .A2(n20691), .ZN(n13641) );
  OAI21_X1 U15887 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12761), .A(
        n12759), .ZN(n13803) );
  NAND2_X1 U15888 ( .A1(n13641), .A2(n13803), .ZN(n13675) );
  NOR2_X1 U15889 ( .A1(n13932), .A2(n13675), .ZN(n18987) );
  OAI21_X1 U15890 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12763), .A(
        n12762), .ZN(n18990) );
  NAND2_X1 U15891 ( .A1(n18987), .A2(n18990), .ZN(n18974) );
  NOR2_X1 U15892 ( .A1(n18976), .A2(n18974), .ZN(n13618) );
  OAI21_X1 U15893 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12764), .A(
        n12756), .ZN(n15344) );
  NAND2_X1 U15894 ( .A1(n13618), .A2(n15344), .ZN(n13660) );
  NOR2_X1 U15895 ( .A1(n16329), .A2(n13660), .ZN(n18959) );
  OAI21_X1 U15896 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n12757), .A(
        n12765), .ZN(n18961) );
  NAND2_X1 U15897 ( .A1(n18959), .A2(n18961), .ZN(n18948) );
  NOR2_X1 U15898 ( .A1(n18949), .A2(n18948), .ZN(n18943) );
  AOI21_X1 U15899 ( .B1(n12755), .B2(n15323), .A(n12752), .ZN(n15325) );
  INV_X1 U15900 ( .A(n15325), .ZN(n18946) );
  NAND2_X1 U15901 ( .A1(n18943), .A2(n18946), .ZN(n18941) );
  NOR2_X1 U15902 ( .A1(n15307), .A2(n18941), .ZN(n18929) );
  NAND2_X1 U15903 ( .A1(n12751), .A2(n12766), .ZN(n12767) );
  NAND2_X1 U15904 ( .A1(n12768), .A2(n12767), .ZN(n18928) );
  NAND2_X1 U15905 ( .A1(n18929), .A2(n18928), .ZN(n13826) );
  NOR2_X1 U15906 ( .A1(n15290), .A2(n13826), .ZN(n18909) );
  INV_X1 U15907 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18906) );
  INV_X1 U15908 ( .A(n12749), .ZN(n12769) );
  AOI21_X1 U15909 ( .B1(n18906), .B2(n12769), .A(n12746), .ZN(n15277) );
  INV_X1 U15910 ( .A(n15277), .ZN(n18911) );
  NAND2_X1 U15911 ( .A1(n18909), .A2(n18911), .ZN(n14145) );
  NOR2_X1 U15912 ( .A1(n14147), .A2(n14145), .ZN(n18902) );
  OR2_X1 U15913 ( .A1(n12747), .A2(n20983), .ZN(n12772) );
  NAND2_X1 U15914 ( .A1(n12747), .A2(n20983), .ZN(n12770) );
  NAND2_X1 U15915 ( .A1(n12772), .A2(n12770), .ZN(n18901) );
  AND2_X1 U15916 ( .A1(n18902), .A2(n18901), .ZN(n12771) );
  OR2_X1 U15917 ( .A1(n12772), .A2(n15246), .ZN(n12774) );
  NAND2_X1 U15918 ( .A1(n12772), .A2(n15246), .ZN(n12773) );
  AND2_X1 U15919 ( .A1(n12774), .A2(n12773), .ZN(n15248) );
  AND2_X1 U15920 ( .A1(n12774), .A2(n15234), .ZN(n12775) );
  NOR2_X1 U15921 ( .A1(n9832), .A2(n12775), .ZN(n18886) );
  OAI21_X1 U15922 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9832), .A(
        n12776), .ZN(n15223) );
  INV_X1 U15923 ( .A(n15223), .ZN(n14984) );
  NOR2_X1 U15924 ( .A1(n14982), .A2(n14984), .ZN(n14983) );
  AOI21_X1 U15925 ( .B1(n15208), .B2(n12776), .A(n12777), .ZN(n15211) );
  OAI21_X1 U15926 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12777), .A(
        n12778), .ZN(n16321) );
  INV_X1 U15927 ( .A(n16321), .ZN(n15786) );
  NOR2_X1 U15928 ( .A1(n10032), .A2(n15785), .ZN(n16269) );
  AOI21_X1 U15929 ( .B1(n10833), .B2(n12778), .A(n12779), .ZN(n16271) );
  NOR2_X1 U15930 ( .A1(n16269), .A2(n16271), .ZN(n16270) );
  INV_X1 U15931 ( .A(n12779), .ZN(n12781) );
  INV_X1 U15932 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12780) );
  NAND2_X1 U15933 ( .A1(n12781), .A2(n12780), .ZN(n12783) );
  AND2_X1 U15934 ( .A1(n12783), .A2(n12782), .ZN(n15184) );
  AOI21_X1 U15935 ( .B1(n15168), .B2(n12782), .A(n12785), .ZN(n16259) );
  NOR2_X1 U15936 ( .A1(n10032), .A2(n16258), .ZN(n16240) );
  OAI21_X1 U15937 ( .B1(n12785), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11588), .ZN(n15159) );
  INV_X1 U15938 ( .A(n15159), .ZN(n16242) );
  NOR2_X1 U15939 ( .A1(n16240), .A2(n16242), .ZN(n16241) );
  NOR2_X1 U15940 ( .A1(n10032), .A2(n16241), .ZN(n12937) );
  NOR2_X1 U15941 ( .A1(n12937), .A2(n12939), .ZN(n12938) );
  NOR2_X1 U15942 ( .A1(n10032), .A2(n12938), .ZN(n14951) );
  AOI21_X1 U15943 ( .B1(n10018), .B2(n12787), .A(n12786), .ZN(n15148) );
  NOR2_X1 U15944 ( .A1(n14951), .A2(n15148), .ZN(n14952) );
  NOR2_X1 U15945 ( .A1(n10032), .A2(n14952), .ZN(n12789) );
  OR2_X1 U15946 ( .A1(n12786), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12788) );
  AND2_X1 U15947 ( .A1(n9842), .A2(n12788), .ZN(n14284) );
  NOR2_X1 U15948 ( .A1(n14284), .A2(n12789), .ZN(n12904) );
  AOI21_X1 U15949 ( .B1(n12789), .B2(n14284), .A(n12904), .ZN(n12790) );
  INV_X1 U15950 ( .A(n12790), .ZN(n12837) );
  NOR4_X1 U15951 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n13837), .ZN(n12791) );
  INV_X1 U15952 ( .A(n19009), .ZN(n12836) );
  NAND2_X1 U15953 ( .A1(n12368), .A2(n12977), .ZN(n14932) );
  NOR2_X1 U15954 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19793), .ZN(n12820) );
  NAND2_X1 U15955 ( .A1(n10429), .A2(n12820), .ZN(n12794) );
  AOI22_X1 U15956 ( .A1(n12325), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U15957 ( .B1(n12810), .B2(n15245), .A(n12795), .ZN(n12796) );
  INV_X1 U15958 ( .A(n12796), .ZN(n14124) );
  OR2_X2 U15959 ( .A1(n14123), .A2(n14124), .ZN(n15113) );
  AOI22_X1 U15960 ( .A1(n12325), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12797) );
  OAI21_X1 U15961 ( .B1(n12810), .B2(n19822), .A(n12797), .ZN(n12798) );
  INV_X1 U15962 ( .A(n12798), .ZN(n15112) );
  AOI22_X1 U15963 ( .A1(n12325), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12799) );
  OAI21_X1 U15964 ( .B1(n12810), .B2(n19824), .A(n12799), .ZN(n14979) );
  INV_X1 U15965 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15105) );
  OAI222_X1 U15966 ( .A1(n12810), .A2(n19826), .B1(n12801), .B2(n15105), .C1(
        n15465), .C2(n12800), .ZN(n12954) );
  NAND2_X1 U15967 ( .A1(n12838), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15968 ( .A1(n12325), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12802) );
  AND2_X1 U15969 ( .A1(n12803), .A2(n12802), .ZN(n15452) );
  AOI22_X1 U15970 ( .A1(n12325), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12804) );
  OAI21_X1 U15971 ( .B1(n12810), .B2(n10792), .A(n12804), .ZN(n15097) );
  NAND2_X1 U15972 ( .A1(n12838), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U15973 ( .A1(n12325), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U15974 ( .A1(n12806), .A2(n12805), .ZN(n14967) );
  NAND2_X1 U15975 ( .A1(n12838), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U15976 ( .A1(n12325), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12807) );
  AND2_X1 U15977 ( .A1(n12808), .A2(n12807), .ZN(n15082) );
  NOR2_X2 U15978 ( .A1(n14965), .A2(n15082), .ZN(n15075) );
  AOI22_X1 U15979 ( .A1(n12325), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12809) );
  OAI21_X1 U15980 ( .B1(n12810), .B2(n19833), .A(n12809), .ZN(n15074) );
  NAND2_X1 U15981 ( .A1(n15075), .A2(n15074), .ZN(n12943) );
  NAND2_X1 U15982 ( .A1(n12838), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15983 ( .A1(n12226), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12811) );
  AND2_X1 U15984 ( .A1(n12812), .A2(n12811), .ZN(n12944) );
  NAND2_X1 U15985 ( .A1(n12838), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U15986 ( .A1(n12226), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12813) );
  AND2_X1 U15987 ( .A1(n12814), .A2(n12813), .ZN(n14955) );
  NAND2_X1 U15988 ( .A1(n12838), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U15989 ( .A1(n12226), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12815) );
  AND2_X1 U15990 ( .A1(n12816), .A2(n12815), .ZN(n12817) );
  AND2_X1 U15991 ( .A1(n14954), .A2(n12817), .ZN(n12818) );
  NAND2_X1 U15992 ( .A1(n12819), .A2(n12977), .ZN(n12981) );
  INV_X1 U15993 ( .A(n19787), .ZN(n14936) );
  INV_X1 U15994 ( .A(n12820), .ZN(n12826) );
  NOR2_X1 U15995 ( .A1(n14936), .A2(n12826), .ZN(n13490) );
  INV_X1 U15996 ( .A(n13490), .ZN(n14266) );
  OR2_X1 U15997 ( .A1(n14267), .A2(n13490), .ZN(n12822) );
  OR3_X1 U15998 ( .A1(n12981), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12820), .ZN(
        n12821) );
  NAND2_X1 U15999 ( .A1(n12822), .A2(n12821), .ZN(n20694) );
  AND2_X1 U16000 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19723), .ZN(n19417) );
  NAND2_X1 U16001 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19417), .ZN(n12823) );
  NOR2_X1 U16002 ( .A1(n12823), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16373) );
  NAND2_X1 U16003 ( .A1(n18970), .A2(n12836), .ZN(n12824) );
  NOR2_X1 U16004 ( .A1(n16373), .A2(n12824), .ZN(n12825) );
  INV_X1 U16005 ( .A(n14932), .ZN(n14943) );
  NAND2_X1 U16006 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12826), .ZN(n12827) );
  NOR2_X1 U16007 ( .A1(n12828), .A2(n12827), .ZN(n12829) );
  AND2_X2 U16008 ( .A1(n20697), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19012) );
  AOI22_X1 U16009 ( .A1(n12830), .A2(n20703), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19012), .ZN(n12831) );
  OAI21_X1 U16010 ( .B1(n19838), .B2(n20697), .A(n12831), .ZN(n12832) );
  AOI21_X1 U16011 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n20694), .A(n12832), .ZN(
        n12833) );
  OAI21_X1 U16012 ( .B1(n15059), .B2(n20698), .A(n12833), .ZN(n12834) );
  INV_X1 U16013 ( .A(n12834), .ZN(n12835) );
  OAI211_X1 U16014 ( .C1(n12837), .C2(n12836), .A(n10125), .B(n12835), .ZN(
        P2_U2826) );
  INV_X1 U16015 ( .A(n16278), .ZN(n12863) );
  NAND2_X1 U16016 ( .A1(n12838), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U16017 ( .A1(n12226), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12839) );
  NAND2_X1 U16018 ( .A1(n12840), .A2(n12839), .ZN(n12910) );
  AOI22_X1 U16019 ( .A1(n12325), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12218), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12841) );
  OAI21_X1 U16020 ( .B1(n12810), .B2(n12842), .A(n12841), .ZN(n12843) );
  INV_X1 U16021 ( .A(n12843), .ZN(n12844) );
  XNOR2_X2 U16022 ( .A(n12913), .B(n12844), .ZN(n19053) );
  INV_X1 U16023 ( .A(n19053), .ZN(n12845) );
  NOR2_X1 U16024 ( .A1(n15430), .A2(n15422), .ZN(n12852) );
  INV_X1 U16025 ( .A(n12846), .ZN(n15477) );
  NAND2_X1 U16026 ( .A1(n15516), .A2(n15477), .ZN(n15476) );
  NOR2_X1 U16027 ( .A1(n15475), .A2(n15493), .ZN(n12848) );
  NAND2_X1 U16028 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n12848), .ZN(
        n15455) );
  INV_X1 U16029 ( .A(n15455), .ZN(n15429) );
  NOR2_X1 U16030 ( .A1(n15399), .A2(n15406), .ZN(n15394) );
  INV_X1 U16031 ( .A(n14277), .ZN(n14290) );
  NAND3_X1 U16032 ( .A1(n15383), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14290), .ZN(n15353) );
  NOR3_X1 U16033 ( .A1(n15353), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12847), .ZN(n12858) );
  NAND2_X1 U16034 ( .A1(n12848), .A2(n15465), .ZN(n15464) );
  AND3_X1 U16035 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12849) );
  NAND3_X1 U16036 ( .A1(n15607), .A2(n12850), .A3(n12849), .ZN(n12851) );
  NAND2_X1 U16037 ( .A1(n12851), .A2(n15599), .ZN(n15466) );
  NAND2_X1 U16038 ( .A1(n15464), .A2(n15466), .ZN(n15457) );
  NOR2_X1 U16039 ( .A1(n15626), .A2(n12852), .ZN(n12853) );
  NOR2_X1 U16040 ( .A1(n15457), .A2(n12853), .ZN(n15407) );
  OAI21_X1 U16041 ( .B1(n15394), .B2(n15626), .A(n15407), .ZN(n15389) );
  NOR2_X1 U16042 ( .A1(n15389), .A2(n14277), .ZN(n15367) );
  INV_X1 U16043 ( .A(n15389), .ZN(n14288) );
  AOI22_X1 U16044 ( .A1(n15367), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n15626), .B2(n14288), .ZN(n15358) );
  NOR2_X1 U16045 ( .A1(n15626), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12854) );
  OAI21_X1 U16046 ( .B1(n15358), .B2(n12854), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12855) );
  INV_X1 U16047 ( .A(n12855), .ZN(n12856) );
  NAND2_X1 U16048 ( .A1(n12864), .A2(n16357), .ZN(n12867) );
  NAND3_X1 U16049 ( .A1(n12868), .A2(n12867), .A3(n12866), .ZN(P2_U3015) );
  NAND2_X1 U16050 ( .A1(n12869), .A2(n17765), .ZN(n12885) );
  NAND2_X1 U16051 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17773) );
  NAND2_X1 U16052 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18192) );
  NAND2_X1 U16053 ( .A1(n18789), .A2(n18192), .ZN(n18842) );
  INV_X1 U16054 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17787) );
  INV_X1 U16055 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17774) );
  NOR2_X1 U16056 ( .A1(n17787), .A2(n17774), .ZN(n17771) );
  NOR2_X1 U16057 ( .A1(n17680), .A2(n17665), .ZN(n17667) );
  INV_X1 U16058 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17611) );
  NAND2_X1 U16059 ( .A1(n17589), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17585) );
  INV_X1 U16060 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16549) );
  NOR2_X2 U16061 ( .A1(n17585), .A2(n16549), .ZN(n17567) );
  NAND2_X1 U16062 ( .A1(n17567), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17545) );
  NAND2_X1 U16063 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17546) );
  INV_X1 U16064 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17866) );
  INV_X1 U16065 ( .A(n17506), .ZN(n12871) );
  NAND2_X1 U16066 ( .A1(n16546), .A2(n12871), .ZN(n16405) );
  INV_X1 U16067 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16584) );
  NAND2_X1 U16069 ( .A1(n16404), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12872) );
  INV_X1 U16070 ( .A(n17505), .ZN(n17493) );
  NAND3_X1 U16071 ( .A1(n17493), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16395) );
  NOR2_X1 U16072 ( .A1(n16584), .A2(n16395), .ZN(n12873) );
  INV_X1 U16073 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18836) );
  NOR2_X1 U16074 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18836), .ZN(n17705) );
  NAND2_X1 U16075 ( .A1(n18800), .A2(n18836), .ZN(n18839) );
  NOR2_X1 U16076 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18789), .ZN(
        n18815) );
  AOI21_X1 U16077 ( .B1(n18192), .B2(n18839), .A(n18815), .ZN(n18201) );
  INV_X1 U16078 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16545) );
  NOR3_X2 U16079 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16545), .ZN(n18541) );
  NAND2_X2 U16080 ( .A1(n18305), .A2(n18541), .ZN(n18488) );
  NAND2_X1 U16081 ( .A1(n12873), .A2(n17707), .ZN(n16389) );
  INV_X1 U16082 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16569) );
  XOR2_X1 U16083 ( .A(n16569), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12875) );
  NOR2_X1 U16084 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17610), .ZN(
        n16406) );
  INV_X1 U16085 ( .A(n16405), .ZN(n16547) );
  INV_X1 U16086 ( .A(n17705), .ZN(n17870) );
  OR2_X1 U16087 ( .A1(n18488), .A2(n12873), .ZN(n12874) );
  OAI211_X1 U16088 ( .C1(n16547), .C2(n17870), .A(n17871), .B(n12874), .ZN(
        n16397) );
  NOR2_X1 U16089 ( .A1(n16406), .A2(n16397), .ZN(n16388) );
  OAI22_X1 U16090 ( .A1(n16389), .A2(n12875), .B1(n16388), .B2(n16569), .ZN(
        n12876) );
  AOI211_X1 U16091 ( .C1(n17687), .C2(n16887), .A(n12877), .B(n12876), .ZN(
        n12878) );
  INV_X1 U16092 ( .A(n12883), .ZN(n12884) );
  NAND2_X1 U16093 ( .A1(n12885), .A2(n12884), .ZN(P3_U2799) );
  INV_X1 U16094 ( .A(n12886), .ZN(n12887) );
  XNOR2_X1 U16095 ( .A(n14535), .B(n12887), .ZN(n14715) );
  NAND2_X1 U16096 ( .A1(n13134), .A2(n13509), .ZN(n13269) );
  NOR2_X1 U16097 ( .A1(n12888), .A2(n14514), .ZN(n12889) );
  NAND2_X1 U16098 ( .A1(n12890), .A2(n12889), .ZN(n12891) );
  NAND2_X1 U16099 ( .A1(n13269), .A2(n12891), .ZN(n12892) );
  INV_X1 U16100 ( .A(n14511), .ZN(n14513) );
  INV_X1 U16101 ( .A(n12894), .ZN(n12895) );
  OAI22_X1 U16102 ( .A1(n14513), .A2(n11553), .B1(n12896), .B2(n12895), .ZN(
        n12899) );
  NAND2_X1 U16103 ( .A1(n11401), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12898) );
  NAND2_X1 U16104 ( .A1(n14514), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12897) );
  NAND2_X1 U16105 ( .A1(n12898), .A2(n12897), .ZN(n14512) );
  XNOR2_X1 U16106 ( .A(n12899), .B(n14512), .ZN(n14526) );
  NAND2_X1 U16107 ( .A1(n20023), .A2(n12900), .ZN(n14629) );
  INV_X1 U16108 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14531) );
  INV_X1 U16109 ( .A(n12901), .ZN(n12902) );
  NOR2_X1 U16110 ( .A1(n10032), .A2(n12904), .ZN(n12905) );
  XOR2_X1 U16111 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9842), .Z(n15132) );
  XNOR2_X1 U16112 ( .A(n12905), .B(n15132), .ZN(n12906) );
  NAND2_X1 U16113 ( .A1(n12906), .A2(n19009), .ZN(n12921) );
  NAND2_X1 U16114 ( .A1(n12908), .A2(n12907), .ZN(n12909) );
  OR2_X1 U16115 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  AOI22_X1 U16116 ( .A1(n18986), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n20694), .ZN(n12915) );
  NAND2_X1 U16117 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12914) );
  OAI211_X1 U16118 ( .C1(n15356), .C2(n20698), .A(n12915), .B(n12914), .ZN(
        n12916) );
  AOI21_X1 U16119 ( .B1(n12917), .B2(n20703), .A(n12916), .ZN(n12918) );
  NAND2_X1 U16120 ( .A1(n12921), .A2(n12920), .ZN(P2_U2825) );
  INV_X1 U16121 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20746) );
  NOR3_X1 U16122 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20746), .ZN(n12923) );
  NOR4_X1 U16123 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12922) );
  NAND4_X1 U16124 ( .A1(n13565), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12923), .A4(
        n12922), .ZN(U214) );
  NOR4_X1 U16125 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n12927) );
  NOR4_X1 U16126 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n12926) );
  NOR4_X1 U16127 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n12925) );
  NOR4_X1 U16128 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n12924) );
  NAND4_X1 U16129 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12932) );
  NOR4_X1 U16130 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .A3(P2_ADDRESS_REG_1__SCAN_IN), .A4(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n12930) );
  NOR4_X1 U16131 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n12929) );
  NOR4_X1 U16132 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12928) );
  INV_X1 U16133 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19805) );
  NAND4_X1 U16134 ( .A1(n12930), .A2(n12929), .A3(n12928), .A4(n19805), .ZN(
        n12931) );
  OAI21_X1 U16135 ( .B1(n12932), .B2(n12931), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12933) );
  NOR2_X1 U16136 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12935) );
  NOR4_X1 U16137 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12934) );
  NAND4_X1 U16138 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12935), .A4(n12934), .ZN(n12936) );
  NOR2_X1 U16139 ( .A1(n15653), .A2(n12936), .ZN(n16432) );
  NAND2_X1 U16140 ( .A1(n16432), .A2(U214), .ZN(U212) );
  NOR2_X1 U16141 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12936), .ZN(n16494)
         );
  AOI211_X1 U16142 ( .C1(n12939), .C2(n12937), .A(n12938), .B(n12836), .ZN(
        n12949) );
  OAI22_X1 U16143 ( .A1(n12940), .A2(n19005), .B1(n19836), .B2(n20697), .ZN(
        n12948) );
  INV_X1 U16144 ( .A(n20694), .ZN(n18999) );
  INV_X1 U16145 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12942) );
  INV_X1 U16146 ( .A(n19012), .ZN(n18981) );
  OAI22_X1 U16147 ( .A1(n18999), .A2(n12942), .B1(n12941), .B2(n18981), .ZN(
        n12947) );
  NAND2_X1 U16148 ( .A1(n12943), .A2(n12944), .ZN(n12945) );
  NAND2_X1 U16149 ( .A1(n9777), .A2(n12945), .ZN(n15385) );
  OAI22_X1 U16150 ( .A1(n15386), .A2(n20705), .B1(n20698), .B2(n15385), .ZN(
        n12946) );
  OR4_X1 U16151 ( .A1(n12949), .A2(n12948), .A3(n12947), .A4(n12946), .ZN(
        P2_U2828) );
  AOI211_X1 U16152 ( .C1(n15211), .C2(n12950), .A(n12951), .B(n12836), .ZN(
        n12962) );
  OAI22_X1 U16153 ( .A1(n15208), .A2(n18981), .B1(n19826), .B2(n20697), .ZN(
        n12961) );
  INV_X1 U16154 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12952) );
  OAI22_X1 U16155 ( .A1(n15204), .A2(n19005), .B1(n18999), .B2(n12952), .ZN(
        n12960) );
  OAI21_X1 U16156 ( .B1(n12953), .B2(n12954), .A(n9776), .ZN(n15467) );
  OR2_X1 U16157 ( .A1(n12956), .A2(n12957), .ZN(n12958) );
  NAND2_X1 U16158 ( .A1(n12955), .A2(n12958), .ZN(n15462) );
  OAI22_X1 U16159 ( .A1(n15467), .A2(n20698), .B1(n20705), .B2(n15462), .ZN(
        n12959) );
  OR4_X1 U16160 ( .A1(n12962), .A2(n12961), .A3(n12960), .A4(n12959), .ZN(
        P2_U2834) );
  INV_X1 U16161 ( .A(n15626), .ZN(n15415) );
  INV_X1 U16162 ( .A(n14241), .ZN(n12963) );
  OAI211_X1 U16163 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15415), .B(n12963), .ZN(n12965) );
  NAND2_X1 U16164 ( .A1(n12862), .A2(n13793), .ZN(n12964) );
  OAI211_X1 U16165 ( .C1(n10256), .C2(n15625), .A(n12965), .B(n12964), .ZN(
        n12976) );
  OAI21_X1 U16166 ( .B1(n12967), .B2(n13791), .A(n12966), .ZN(n12968) );
  XNOR2_X1 U16167 ( .A(n12968), .B(n10256), .ZN(n13072) );
  XNOR2_X1 U16168 ( .A(n12970), .B(n12969), .ZN(n19879) );
  INV_X1 U16169 ( .A(n19879), .ZN(n13314) );
  OAI22_X1 U16170 ( .A1(n13072), .A2(n15623), .B1(n15355), .B2(n13314), .ZN(
        n12975) );
  NOR2_X1 U16171 ( .A1(n18933), .A2(n12971), .ZN(n13074) );
  OAI21_X1 U16172 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12973), .A(
        n12972), .ZN(n13070) );
  NOR2_X1 U16173 ( .A1(n15629), .A2(n13070), .ZN(n12974) );
  OR4_X1 U16174 ( .A1(n12976), .A2(n12975), .A3(n13074), .A4(n12974), .ZN(
        P2_U3045) );
  INV_X1 U16175 ( .A(n12977), .ZN(n12978) );
  NOR2_X1 U16176 ( .A1(n9733), .A2(n12978), .ZN(n20707) );
  INV_X1 U16177 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19900) );
  OAI211_X1 U16178 ( .C1(n20707), .C2(n19900), .A(n14930), .B(n12981), .ZN(
        P2_U2814) );
  INV_X1 U16179 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n12980) );
  NAND2_X1 U16180 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19668), .ZN(n12979) );
  OAI22_X1 U16181 ( .A1(n14943), .A2(n12980), .B1(n12979), .B2(n16377), .ZN(
        P2_U2816) );
  INV_X1 U16182 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19141) );
  INV_X1 U16183 ( .A(n12981), .ZN(n12984) );
  NAND3_X1 U16184 ( .A1(n12984), .A2(n15862), .A3(n13143), .ZN(n13051) );
  NAND2_X1 U16185 ( .A1(n15653), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12983) );
  INV_X1 U16186 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16458) );
  OR2_X1 U16187 ( .A1(n15653), .A2(n16458), .ZN(n12982) );
  NAND2_X1 U16188 ( .A1(n12983), .A2(n12982), .ZN(n19077) );
  NAND2_X1 U16189 ( .A1(n13038), .A2(n19077), .ZN(n13043) );
  OAI21_X1 U16190 ( .B1(n9761), .B2(n15862), .A(n12984), .ZN(n12991) );
  NAND2_X1 U16191 ( .A1(n12991), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12985) );
  OAI211_X1 U16192 ( .C1(n19141), .C2(n14267), .A(n13043), .B(n12985), .ZN(
        P2_U2979) );
  AOI22_X1 U16193 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12991), .B1(n13048), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16194 ( .A1(n15651), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15653), .ZN(n19129) );
  INV_X1 U16195 ( .A(n19129), .ZN(n19191) );
  NAND2_X1 U16196 ( .A1(n13038), .A2(n19191), .ZN(n12992) );
  NAND2_X1 U16197 ( .A1(n12986), .A2(n12992), .ZN(P2_U2953) );
  AOI22_X1 U16198 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12991), .B1(n13048), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16199 ( .A1(n15651), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15653), .ZN(n19118) );
  INV_X1 U16200 ( .A(n19118), .ZN(n15645) );
  NAND2_X1 U16201 ( .A1(n13038), .A2(n15645), .ZN(n13013) );
  NAND2_X1 U16202 ( .A1(n12987), .A2(n13013), .ZN(P2_U2955) );
  AOI22_X1 U16203 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12991), .B1(n13048), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12988) );
  OAI22_X1 U16204 ( .A1(n15653), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15651), .ZN(n19110) );
  INV_X1 U16205 ( .A(n19110), .ZN(n16303) );
  NAND2_X1 U16206 ( .A1(n13038), .A2(n16303), .ZN(n13000) );
  NAND2_X1 U16207 ( .A1(n12988), .A2(n13000), .ZN(P2_U2956) );
  AOI22_X1 U16208 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12991), .B1(n13048), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U16209 ( .A1(n15651), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15653), .ZN(n19092) );
  INV_X1 U16210 ( .A(n19092), .ZN(n19220) );
  NAND2_X1 U16211 ( .A1(n13038), .A2(n19220), .ZN(n13016) );
  NAND2_X1 U16212 ( .A1(n12989), .A2(n13016), .ZN(P2_U2959) );
  AOI22_X1 U16213 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12991), .B1(n13048), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16214 ( .A1(n15651), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15653), .ZN(n15106) );
  INV_X1 U16215 ( .A(n15106), .ZN(n19203) );
  NAND2_X1 U16216 ( .A1(n13038), .A2(n19203), .ZN(n13024) );
  NAND2_X1 U16217 ( .A1(n12990), .A2(n13024), .ZN(P2_U2957) );
  CLKBUF_X2 U16218 ( .A(n12991), .Z(n13049) );
  AOI22_X1 U16219 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U16220 ( .A1(n12993), .A2(n12992), .ZN(P2_U2968) );
  AOI22_X1 U16221 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12996) );
  INV_X1 U16222 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13337) );
  OR2_X1 U16223 ( .A1(n15653), .A2(n13337), .ZN(n12995) );
  NAND2_X1 U16224 ( .A1(n15653), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12994) );
  AND2_X1 U16225 ( .A1(n12995), .A2(n12994), .ZN(n19081) );
  INV_X1 U16226 ( .A(n19081), .ZN(n15067) );
  NAND2_X1 U16227 ( .A1(n13038), .A2(n15067), .ZN(n13009) );
  NAND2_X1 U16228 ( .A1(n12996), .A2(n13009), .ZN(P2_U2963) );
  AOI22_X1 U16229 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16230 ( .A1(n15653), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12998) );
  INV_X1 U16231 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16463) );
  OR2_X1 U16232 ( .A1(n15653), .A2(n16463), .ZN(n12997) );
  NAND2_X1 U16233 ( .A1(n12998), .A2(n12997), .ZN(n19085) );
  NAND2_X1 U16234 ( .A1(n13038), .A2(n19085), .ZN(n13045) );
  NAND2_X1 U16235 ( .A1(n12999), .A2(n13045), .ZN(P2_U2961) );
  AOI22_X1 U16236 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13001) );
  NAND2_X1 U16237 ( .A1(n13001), .A2(n13000), .ZN(P2_U2971) );
  AOI22_X1 U16238 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13002) );
  INV_X1 U16239 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20904) );
  INV_X1 U16240 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U16241 ( .A1(n15651), .A2(n20904), .B1(n18210), .B2(n15653), .ZN(
        n19197) );
  NAND2_X1 U16242 ( .A1(n13038), .A2(n19197), .ZN(n13018) );
  NAND2_X1 U16243 ( .A1(n13002), .A2(n13018), .ZN(P2_U2969) );
  AOI22_X1 U16244 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13004) );
  INV_X1 U16245 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13373) );
  NOR2_X1 U16246 ( .A1(n15653), .A2(n13373), .ZN(n13003) );
  AOI21_X1 U16247 ( .B1(n15653), .B2(BUF2_REG_13__SCAN_IN), .A(n13003), .ZN(
        n19075) );
  INV_X1 U16248 ( .A(n19075), .ZN(n15056) );
  NAND2_X1 U16249 ( .A1(n13038), .A2(n15056), .ZN(n13007) );
  NAND2_X1 U16250 ( .A1(n13004), .A2(n13007), .ZN(P2_U2980) );
  AOI22_X1 U16251 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13005) );
  INV_X1 U16252 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16478) );
  INV_X1 U16253 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U16254 ( .A1(n15651), .A2(n16478), .B1(n18200), .B2(n15653), .ZN(
        n19185) );
  NAND2_X1 U16255 ( .A1(n13038), .A2(n19185), .ZN(n13022) );
  NAND2_X1 U16256 ( .A1(n13005), .A2(n13022), .ZN(P2_U2952) );
  AOI22_X1 U16257 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13006) );
  OAI22_X1 U16258 ( .A1(n15653), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15651), .ZN(n19094) );
  INV_X1 U16259 ( .A(n19094), .ZN(n19207) );
  NAND2_X1 U16260 ( .A1(n13038), .A2(n19207), .ZN(n13011) );
  NAND2_X1 U16261 ( .A1(n13006), .A2(n13011), .ZN(P2_U2973) );
  AOI22_X1 U16262 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U16263 ( .A1(n13008), .A2(n13007), .ZN(P2_U2965) );
  AOI22_X1 U16264 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13010) );
  NAND2_X1 U16265 ( .A1(n13010), .A2(n13009), .ZN(P2_U2978) );
  AOI22_X1 U16266 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U16267 ( .A1(n13012), .A2(n13011), .ZN(P2_U2958) );
  AOI22_X1 U16268 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13014) );
  NAND2_X1 U16269 ( .A1(n13014), .A2(n13013), .ZN(P2_U2970) );
  AOI22_X1 U16270 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U16271 ( .A1(n15651), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15653), .ZN(n19089) );
  INV_X1 U16272 ( .A(n19089), .ZN(n15090) );
  NAND2_X1 U16273 ( .A1(n13038), .A2(n15090), .ZN(n13020) );
  NAND2_X1 U16274 ( .A1(n13015), .A2(n13020), .ZN(P2_U2975) );
  AOI22_X1 U16275 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U16276 ( .A1(n13017), .A2(n13016), .ZN(P2_U2974) );
  AOI22_X1 U16277 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16278 ( .A1(n13019), .A2(n13018), .ZN(P2_U2954) );
  AOI22_X1 U16279 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13021) );
  NAND2_X1 U16280 ( .A1(n13021), .A2(n13020), .ZN(P2_U2960) );
  AOI22_X1 U16281 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13023) );
  NAND2_X1 U16282 ( .A1(n13023), .A2(n13022), .ZN(P2_U2967) );
  AOI22_X1 U16283 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U16284 ( .A1(n13025), .A2(n13024), .ZN(P2_U2972) );
  INV_X1 U16285 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13032) );
  OR2_X1 U16286 ( .A1(n9733), .A2(n13026), .ZN(n13028) );
  OR2_X1 U16287 ( .A1(n13028), .A2(n13027), .ZN(n13030) );
  NAND2_X1 U16288 ( .A1(n19154), .A2(n10231), .ZN(n19131) );
  OR2_X1 U16289 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16368), .ZN(n19156) );
  INV_X2 U16290 ( .A(n19156), .ZN(n19167) );
  NOR2_X2 U16291 ( .A1(n19154), .A2(n19167), .ZN(n19166) );
  AOI22_X1 U16292 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n19166), .B1(n19167), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13031) );
  OAI21_X1 U16293 ( .B1(n13032), .B2(n19131), .A(n13031), .ZN(P2_U2924) );
  INV_X1 U16294 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19137) );
  NAND2_X1 U16295 ( .A1(n15653), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13034) );
  INV_X1 U16296 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13346) );
  OR2_X1 U16297 ( .A1(n15653), .A2(n13346), .ZN(n13033) );
  NAND2_X1 U16298 ( .A1(n13034), .A2(n13033), .ZN(n19071) );
  NAND2_X1 U16299 ( .A1(n13038), .A2(n19071), .ZN(n13041) );
  NAND2_X1 U16300 ( .A1(n13049), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13035) );
  OAI211_X1 U16301 ( .C1(n19137), .C2(n14267), .A(n13041), .B(n13035), .ZN(
        P2_U2981) );
  INV_X1 U16302 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13055) );
  NAND2_X1 U16303 ( .A1(n15653), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13037) );
  INV_X1 U16304 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16461) );
  OR2_X1 U16305 ( .A1(n15653), .A2(n16461), .ZN(n13036) );
  NAND2_X1 U16306 ( .A1(n13037), .A2(n13036), .ZN(n19082) );
  NAND2_X1 U16307 ( .A1(n13038), .A2(n19082), .ZN(n13047) );
  NAND2_X1 U16308 ( .A1(n13049), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13039) );
  OAI211_X1 U16309 ( .C1(n13055), .C2(n14267), .A(n13047), .B(n13039), .ZN(
        P2_U2962) );
  INV_X1 U16310 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U16311 ( .A1(n13049), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13040) );
  OAI211_X1 U16312 ( .C1(n13120), .C2(n14267), .A(n13041), .B(n13040), .ZN(
        P2_U2966) );
  INV_X1 U16313 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13059) );
  NAND2_X1 U16314 ( .A1(n13049), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13042) );
  OAI211_X1 U16315 ( .C1(n13059), .C2(n14267), .A(n13043), .B(n13042), .ZN(
        P2_U2964) );
  INV_X1 U16316 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19147) );
  NAND2_X1 U16317 ( .A1(n13049), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13044) );
  OAI211_X1 U16318 ( .C1(n19147), .C2(n14267), .A(n13045), .B(n13044), .ZN(
        P2_U2976) );
  INV_X1 U16319 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19145) );
  NAND2_X1 U16320 ( .A1(n13049), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13046) );
  OAI211_X1 U16321 ( .C1(n19145), .C2(n14267), .A(n13047), .B(n13046), .ZN(
        P2_U2977) );
  AOI22_X1 U16322 ( .A1(n15651), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15653), .ZN(n19070) );
  AOI22_X1 U16323 ( .A1(P2_LWORD_REG_15__SCAN_IN), .A2(n13049), .B1(n13048), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n13050) );
  OAI21_X1 U16324 ( .B1(n19070), .B2(n13051), .A(n13050), .ZN(P2_U2982) );
  INV_X1 U16325 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16326 ( .A1(n19167), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13052) );
  OAI21_X1 U16327 ( .B1(n13053), .B2(n19131), .A(n13052), .ZN(P2_U2922) );
  AOI22_X1 U16328 ( .A1(n19167), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13054) );
  OAI21_X1 U16329 ( .B1(n13055), .B2(n19131), .A(n13054), .ZN(P2_U2925) );
  INV_X1 U16330 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16331 ( .A1(n19167), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13056) );
  OAI21_X1 U16332 ( .B1(n13057), .B2(n19131), .A(n13056), .ZN(P2_U2926) );
  AOI22_X1 U16333 ( .A1(n19167), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13058) );
  OAI21_X1 U16334 ( .B1(n13059), .B2(n19131), .A(n13058), .ZN(P2_U2923) );
  INV_X1 U16335 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U16336 ( .A1(n19167), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13060) );
  OAI21_X1 U16337 ( .B1(n13873), .B2(n19131), .A(n13060), .ZN(P2_U2934) );
  INV_X1 U16338 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U16339 ( .A1(n19167), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13061) );
  OAI21_X1 U16340 ( .B1(n15114), .B2(n19131), .A(n13061), .ZN(P2_U2932) );
  INV_X1 U16341 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16342 ( .A1(n19167), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13062) );
  OAI21_X1 U16343 ( .B1(n13063), .B2(n19131), .A(n13062), .ZN(P2_U2931) );
  AOI22_X1 U16344 ( .A1(n19167), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13064) );
  OAI21_X1 U16345 ( .B1(n15105), .B2(n19131), .A(n13064), .ZN(P2_U2930) );
  INV_X1 U16346 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16347 ( .A1(n19167), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13065) );
  OAI21_X1 U16348 ( .B1(n13066), .B2(n19131), .A(n13065), .ZN(P2_U2929) );
  INV_X1 U16349 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16350 ( .A1(n19167), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13067) );
  OAI21_X1 U16351 ( .B1(n13068), .B2(n19131), .A(n13067), .ZN(P2_U2927) );
  INV_X1 U16352 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13069) );
  INV_X1 U16353 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16502) );
  INV_X1 U16354 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n20734) );
  OAI222_X1 U16355 ( .A1(n19131), .A2(n13069), .B1(n19152), .B2(n16502), .C1(
        n19156), .C2(n20734), .ZN(P2_U2928) );
  INV_X1 U16356 ( .A(n13070), .ZN(n13075) );
  OAI22_X1 U16357 ( .A1(n13072), .A2(n19179), .B1(n13071), .B2(n19184), .ZN(
        n13073) );
  AOI211_X1 U16358 ( .C1(n10876), .C2(n13075), .A(n13074), .B(n13073), .ZN(
        n13077) );
  NAND2_X1 U16359 ( .A1(n13793), .A2(n19176), .ZN(n13076) );
  OAI211_X1 U16360 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19172), .A(
        n13077), .B(n13076), .ZN(P2_U3013) );
  NAND2_X1 U16361 ( .A1(n12148), .A2(n10228), .ZN(n13078) );
  NAND2_X1 U16362 ( .A1(n13079), .A2(n13078), .ZN(n13087) );
  OR2_X1 U16363 ( .A1(n13773), .A2(n13431), .ZN(n13110) );
  NAND2_X1 U16364 ( .A1(n13470), .A2(n13773), .ZN(n13151) );
  NAND2_X1 U16365 ( .A1(n12368), .A2(n14934), .ZN(n13081) );
  NAND2_X1 U16366 ( .A1(n9734), .A2(n19787), .ZN(n13080) );
  NAND2_X1 U16367 ( .A1(n13081), .A2(n13080), .ZN(n13083) );
  NAND2_X1 U16368 ( .A1(n13083), .A2(n13082), .ZN(n13084) );
  AND4_X1 U16369 ( .A1(n13110), .A2(n13085), .A3(n13151), .A4(n13084), .ZN(
        n13086) );
  NAND2_X1 U16370 ( .A1(n13087), .A2(n13086), .ZN(n13485) );
  NAND2_X1 U16371 ( .A1(n13485), .A2(n18862), .ZN(n13090) );
  NAND2_X1 U16372 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19887), .ZN(n15863) );
  NOR2_X1 U16373 ( .A1(n18865), .A2(n15863), .ZN(n15867) );
  INV_X1 U16374 ( .A(n13497), .ZN(n13088) );
  NOR2_X1 U16375 ( .A1(n15867), .A2(n13088), .ZN(n13089) );
  NAND2_X1 U16376 ( .A1(n13090), .A2(n13089), .ZN(n15641) );
  INV_X1 U16377 ( .A(n15641), .ZN(n13843) );
  INV_X1 U16378 ( .A(n13091), .ZN(n13092) );
  AND2_X1 U16379 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  OR3_X1 U16380 ( .A1(n13843), .A2(n19854), .A3(n13481), .ZN(n13095) );
  OAI21_X1 U16381 ( .B1(n13486), .B2(n15641), .A(n13095), .ZN(P2_U3595) );
  AOI21_X1 U16382 ( .B1(n13097), .B2(n19004), .A(n13096), .ZN(n15627) );
  NOR2_X1 U16383 ( .A1(n18933), .A2(n18997), .ZN(n15631) );
  OAI21_X1 U16384 ( .B1(n13099), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13098), .ZN(n15628) );
  NOR2_X1 U16385 ( .A1(n19173), .A2(n15628), .ZN(n13100) );
  AOI211_X1 U16386 ( .C1(n15627), .C2(n16346), .A(n15631), .B(n13100), .ZN(
        n13103) );
  OAI21_X1 U16387 ( .B1(n16322), .B2(n13101), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13102) );
  OAI211_X1 U16388 ( .C1(n15652), .C2(n13449), .A(n13103), .B(n13102), .ZN(
        P2_U3014) );
  OAI21_X1 U16389 ( .B1(n9706), .B2(n16380), .A(n19668), .ZN(n13212) );
  NOR2_X1 U16390 ( .A1(n19581), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13105) );
  AOI21_X1 U16391 ( .B1(n13212), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13105), .ZN(n13106) );
  INV_X1 U16392 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20885) );
  NAND2_X1 U16393 ( .A1(n13143), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13108) );
  AND4_X1 U16394 ( .A1(n9706), .A2(n13108), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19668), .ZN(n13109) );
  NAND2_X1 U16395 ( .A1(n13110), .A2(n13428), .ZN(n13111) );
  NAND2_X1 U16396 ( .A1(n19048), .A2(n19215), .ZN(n19041) );
  MUX2_X1 U16397 ( .A(n13449), .B(n18998), .S(n19052), .Z(n13112) );
  OAI21_X1 U16398 ( .B1(n19884), .B2(n19041), .A(n13112), .ZN(P2_U2887) );
  NAND2_X1 U16399 ( .A1(n13130), .A2(n13128), .ZN(n13115) );
  INV_X1 U16400 ( .A(n13114), .ZN(n13125) );
  AOI22_X1 U16401 ( .A1(n13115), .A2(n13113), .B1(n13134), .B2(n13125), .ZN(
        n13127) );
  AND2_X1 U16402 ( .A1(n13127), .A2(n13171), .ZN(n13118) );
  INV_X1 U16403 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n13117) );
  INV_X1 U16404 ( .A(n14262), .ZN(n14926) );
  NOR2_X1 U16405 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n16236), .ZN(n16228) );
  INV_X1 U16406 ( .A(n16228), .ZN(n13116) );
  OAI22_X1 U16407 ( .A1(n13118), .A2(n13117), .B1(n14926), .B2(n13116), .ZN(
        P1_U2803) );
  AOI22_X1 U16408 ( .A1(n19167), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13119) );
  OAI21_X1 U16409 ( .B1(n13120), .B2(n19131), .A(n13119), .ZN(P2_U2921) );
  INV_X1 U16410 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16411 ( .A1(n19167), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U16412 ( .B1(n13122), .B2(n19131), .A(n13121), .ZN(P2_U2935) );
  AND2_X1 U16413 ( .A1(n13128), .A2(n13171), .ZN(n13123) );
  NAND2_X1 U16414 ( .A1(n13130), .A2(n13123), .ZN(n13147) );
  AND2_X1 U16415 ( .A1(n20538), .A2(n16233), .ZN(n14094) );
  INV_X1 U16416 ( .A(n13336), .ZN(n13334) );
  AOI211_X1 U16417 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13147), .A(n14094), 
        .B(n13334), .ZN(n13124) );
  INV_X1 U16418 ( .A(n13124), .ZN(P1_U2801) );
  NAND3_X1 U16419 ( .A1(n13125), .A2(n14514), .A3(n15843), .ZN(n13126) );
  NAND2_X1 U16420 ( .A1(n13126), .A2(n20603), .ZN(n20678) );
  AND2_X1 U16421 ( .A1(n13127), .A2(n20678), .ZN(n15818) );
  NOR2_X1 U16422 ( .A1(n15818), .A2(n13277), .ZN(n19908) );
  INV_X1 U16423 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15816) );
  INV_X1 U16424 ( .A(n13128), .ZN(n13129) );
  AOI22_X1 U16425 ( .A1(n13130), .A2(n13129), .B1(n13509), .B2(n13537), .ZN(
        n13137) );
  INV_X1 U16426 ( .A(n13131), .ZN(n13132) );
  NAND3_X1 U16427 ( .A1(n13510), .A2(n13133), .A3(n13132), .ZN(n13135) );
  NAND2_X1 U16428 ( .A1(n13135), .A2(n13134), .ZN(n13136) );
  NAND2_X1 U16429 ( .A1(n13137), .A2(n13136), .ZN(n13138) );
  NAND2_X1 U16430 ( .A1(n13138), .A2(n11008), .ZN(n15819) );
  INV_X1 U16431 ( .A(n15819), .ZN(n13139) );
  NAND2_X1 U16432 ( .A1(n19908), .A2(n13139), .ZN(n13140) );
  OAI21_X1 U16433 ( .B1(n19908), .B2(n15816), .A(n13140), .ZN(P1_U3484) );
  NAND2_X1 U16434 ( .A1(n13212), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13141) );
  NAND2_X1 U16435 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19547) );
  NAND2_X1 U16436 ( .A1(n19881), .A2(n19890), .ZN(n19447) );
  AND2_X1 U16437 ( .A1(n19547), .A2(n19447), .ZN(n19389) );
  NAND2_X1 U16438 ( .A1(n19389), .A2(n19852), .ZN(n19520) );
  NAND2_X1 U16439 ( .A1(n13141), .A2(n19520), .ZN(n13142) );
  NAND2_X1 U16440 ( .A1(n13144), .A2(n9706), .ZN(n14397) );
  INV_X1 U16441 ( .A(n14397), .ZN(n14454) );
  NAND2_X1 U16442 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13191) );
  INV_X1 U16443 ( .A(n13793), .ZN(n13441) );
  MUX2_X1 U16444 ( .A(n13145), .B(n13441), .S(n19048), .Z(n13146) );
  OAI21_X1 U16445 ( .B1(n19874), .B2(n19041), .A(n13146), .ZN(P2_U2886) );
  NOR2_X1 U16446 ( .A1(n14094), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13149)
         );
  OAI21_X1 U16447 ( .B1(n11024), .B2(n13904), .A(n20681), .ZN(n13148) );
  OAI21_X1 U16448 ( .B1(n13149), .B2(n20681), .A(n13148), .ZN(P1_U3487) );
  NAND2_X1 U16449 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U16450 ( .A1(n13152), .A2(n18862), .ZN(n13155) );
  NAND2_X1 U16451 ( .A1(n14934), .A2(n15862), .ZN(n13153) );
  OR2_X1 U16452 ( .A1(n14932), .A2(n13153), .ZN(n13154) );
  AND2_X1 U16453 ( .A1(n19095), .A2(n13157), .ZN(n13874) );
  INV_X1 U16454 ( .A(n19185), .ZN(n13169) );
  INV_X1 U16455 ( .A(n12232), .ZN(n13163) );
  INV_X1 U16456 ( .A(n13158), .ZN(n13161) );
  INV_X1 U16457 ( .A(n13159), .ZN(n13160) );
  NAND2_X1 U16458 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  NAND2_X1 U16459 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  INV_X1 U16460 ( .A(n13164), .ZN(n19001) );
  NOR2_X1 U16461 ( .A1(n19884), .A2(n13164), .ZN(n19123) );
  INV_X1 U16462 ( .A(n19123), .ZN(n13166) );
  OAI211_X1 U16463 ( .C1(n19444), .C2(n19001), .A(n13166), .B(n19106), .ZN(
        n13168) );
  NAND2_X1 U16464 ( .A1(n19095), .A2(n9957), .ZN(n19063) );
  AOI22_X1 U16465 ( .A1(n19120), .A2(n19001), .B1(n19119), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13167) );
  OAI211_X1 U16466 ( .C1(n19128), .C2(n13169), .A(n13168), .B(n13167), .ZN(
        P2_U2919) );
  INV_X1 U16467 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13175) );
  INV_X1 U16468 ( .A(n15797), .ZN(n13170) );
  OR2_X1 U16469 ( .A1(n15802), .A2(n13170), .ZN(n13173) );
  AND3_X1 U16470 ( .A1(n13537), .A2(n15795), .A3(n13171), .ZN(n13172) );
  NAND2_X1 U16471 ( .A1(n20035), .A2(n11328), .ZN(n13241) );
  NOR2_X1 U16472 ( .A1(n20525), .A2(n16233), .ZN(n16229) );
  NAND2_X1 U16473 ( .A1(n16229), .A2(n16236), .ZN(n20046) );
  INV_X2 U16474 ( .A(n20046), .ZN(n20036) );
  NOR2_X4 U16475 ( .A1(n20035), .A2(n20036), .ZN(n20038) );
  AOI22_X1 U16476 ( .A1(n20036), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13174) );
  OAI21_X1 U16477 ( .B1(n13175), .B2(n13241), .A(n13174), .ZN(P1_U2920) );
  INV_X1 U16478 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16479 ( .A1(n20036), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13176) );
  OAI21_X1 U16480 ( .B1(n13350), .B2(n13241), .A(n13176), .ZN(P1_U2906) );
  INV_X1 U16481 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16482 ( .A1(n20036), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13177) );
  OAI21_X1 U16483 ( .B1(n13178), .B2(n13241), .A(n13177), .ZN(P1_U2918) );
  INV_X1 U16484 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n20804) );
  INV_X1 U16485 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13179) );
  INV_X1 U16486 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n20840) );
  OAI222_X1 U16487 ( .A1(n20044), .A2(n20804), .B1(n13241), .B2(n13179), .C1(
        n20840), .C2(n20046), .ZN(P1_U2919) );
  NAND2_X1 U16488 ( .A1(n13181), .A2(n13208), .ZN(n13186) );
  NAND2_X1 U16489 ( .A1(n19547), .A2(n19871), .ZN(n13183) );
  NAND2_X1 U16490 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19719) );
  INV_X1 U16491 ( .A(n19719), .ZN(n13182) );
  NAND2_X1 U16492 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13182), .ZN(
        n13210) );
  NAND2_X1 U16493 ( .A1(n13183), .A2(n13210), .ZN(n19328) );
  NOR2_X1 U16494 ( .A1(n19328), .A2(n19581), .ZN(n13184) );
  AOI21_X1 U16495 ( .B1(n13212), .B2(n14352), .A(n13184), .ZN(n13185) );
  NAND2_X1 U16496 ( .A1(n13186), .A2(n13185), .ZN(n13189) );
  INV_X1 U16497 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13187) );
  NOR2_X1 U16498 ( .A1(n14397), .A2(n13187), .ZN(n13188) );
  OR2_X1 U16499 ( .A1(n13189), .A2(n13188), .ZN(n13190) );
  NAND2_X1 U16500 ( .A1(n13189), .A2(n13188), .ZN(n13220) );
  INV_X1 U16501 ( .A(n13191), .ZN(n13192) );
  INV_X1 U16502 ( .A(n13218), .ZN(n13196) );
  INV_X1 U16503 ( .A(n20708), .ZN(n19866) );
  INV_X1 U16504 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13198) );
  MUX2_X1 U16505 ( .A(n13197), .B(n13198), .S(n19052), .Z(n13199) );
  OAI21_X1 U16506 ( .B1(n19866), .B2(n19041), .A(n13199), .ZN(P2_U2885) );
  INV_X1 U16507 ( .A(n13200), .ZN(n13202) );
  OR2_X1 U16508 ( .A1(n11401), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13201) );
  NAND2_X1 U16509 ( .A1(n13202), .A2(n13201), .ZN(n13978) );
  INV_X1 U16510 ( .A(n13203), .ZN(n13206) );
  OAI21_X1 U16511 ( .B1(n13206), .B2(n13205), .A(n13204), .ZN(n13983) );
  OAI222_X1 U16512 ( .A1(n13978), .A2(n14629), .B1(n11406), .B2(n20023), .C1(
        n13983), .C2(n14635), .ZN(P1_U2872) );
  NAND2_X1 U16513 ( .A1(n13207), .A2(n13208), .ZN(n13214) );
  INV_X1 U16514 ( .A(n13210), .ZN(n13209) );
  NAND2_X1 U16515 ( .A1(n13209), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19721) );
  NAND2_X1 U16516 ( .A1(n19864), .A2(n13210), .ZN(n13211) );
  AND3_X1 U16517 ( .A1(n19721), .A2(n19852), .A3(n13211), .ZN(n19576) );
  AOI21_X1 U16518 ( .B1(n13212), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19576), .ZN(n13213) );
  INV_X1 U16519 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13215) );
  NOR2_X1 U16520 ( .A1(n14397), .A2(n13215), .ZN(n13216) );
  NAND2_X1 U16521 ( .A1(n13219), .A2(n13218), .ZN(n13221) );
  NAND2_X1 U16522 ( .A1(n13223), .A2(n13222), .ZN(n13245) );
  NAND2_X1 U16523 ( .A1(n19052), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U16524 ( .A1(n13207), .A2(n19048), .ZN(n13225) );
  OAI211_X1 U16525 ( .C1(n19445), .C2(n19041), .A(n13226), .B(n13225), .ZN(
        P2_U2884) );
  INV_X1 U16526 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13360) );
  AOI22_X1 U16527 ( .A1(n20036), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U16528 ( .B1(n13360), .B2(n13241), .A(n13227), .ZN(P1_U2912) );
  INV_X1 U16529 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U16530 ( .A1(n20036), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13228) );
  OAI21_X1 U16531 ( .B1(n14673), .B2(n13241), .A(n13228), .ZN(P1_U2913) );
  INV_X1 U16532 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U16533 ( .A1(n20036), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13229) );
  OAI21_X1 U16534 ( .B1(n13230), .B2(n13241), .A(n13229), .ZN(P1_U2917) );
  AOI22_X1 U16535 ( .A1(n20036), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16536 ( .B1(n14654), .B2(n13241), .A(n13231), .ZN(P1_U2908) );
  AOI22_X1 U16537 ( .A1(n20036), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13232) );
  OAI21_X1 U16538 ( .B1(n14679), .B2(n13241), .A(n13232), .ZN(P1_U2914) );
  INV_X1 U16539 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U16540 ( .A1(n20036), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16541 ( .B1(n13234), .B2(n13241), .A(n13233), .ZN(P1_U2910) );
  INV_X1 U16542 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16543 ( .A1(n20036), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16544 ( .B1(n13236), .B2(n13241), .A(n13235), .ZN(P1_U2916) );
  AOI22_X1 U16545 ( .A1(n20036), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13237) );
  OAI21_X1 U16546 ( .B1(n14663), .B2(n13241), .A(n13237), .ZN(P1_U2911) );
  AOI22_X1 U16547 ( .A1(n20036), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U16548 ( .B1(n12022), .B2(n13241), .A(n13238), .ZN(P1_U2909) );
  AOI22_X1 U16549 ( .A1(n20036), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U16550 ( .B1(n14649), .B2(n13241), .A(n13239), .ZN(P1_U2907) );
  INV_X1 U16551 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n20858) );
  AOI22_X1 U16552 ( .A1(n20036), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16553 ( .B1(n20858), .B2(n13241), .A(n13240), .ZN(P1_U2915) );
  NAND2_X1 U16554 ( .A1(n10216), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13242) );
  INV_X1 U16555 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13246) );
  NOR2_X1 U16556 ( .A1(n14397), .A2(n13246), .ZN(n19037) );
  NAND2_X1 U16557 ( .A1(n9755), .A2(n19037), .ZN(n13674) );
  XOR2_X1 U16558 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13674), .Z(n13252)
         );
  OAI21_X1 U16559 ( .B1(n13247), .B2(n13249), .A(n13248), .ZN(n18991) );
  NOR2_X1 U16560 ( .A1(n18991), .A2(n19052), .ZN(n13250) );
  AOI21_X1 U16561 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n19052), .A(n13250), .ZN(
        n13251) );
  OAI21_X1 U16562 ( .B1(n13252), .B2(n19041), .A(n13251), .ZN(P2_U2882) );
  NAND2_X1 U16563 ( .A1(n13253), .A2(n14803), .ZN(n13257) );
  INV_X1 U16564 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13254) );
  NOR2_X1 U16565 ( .A1(n16209), .A2(n13254), .ZN(n14893) );
  OAI21_X1 U16566 ( .B1(n13255), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11160), .ZN(n14892) );
  NOR2_X1 U16567 ( .A1(n14892), .A2(n19906), .ZN(n13256) );
  AOI211_X1 U16568 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13257), .A(
        n14893), .B(n13256), .ZN(n13258) );
  OAI21_X1 U16569 ( .B1(n20076), .B2(n13983), .A(n13258), .ZN(P1_U2999) );
  INV_X1 U16570 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13259) );
  NOR2_X1 U16571 ( .A1(n13674), .A2(n13259), .ZN(n13260) );
  NAND2_X1 U16572 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13301) );
  OR2_X1 U16573 ( .A1(n13674), .A2(n13301), .ZN(n13295) );
  OAI211_X1 U16574 ( .C1(n13260), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19018), .B(n13295), .ZN(n13265) );
  INV_X1 U16575 ( .A(n13261), .ZN(n13262) );
  AOI21_X1 U16576 ( .B1(n13263), .B2(n13248), .A(n13262), .ZN(n18977) );
  NAND2_X1 U16577 ( .A1(n18977), .A2(n19048), .ZN(n13264) );
  OAI211_X1 U16578 ( .C1(n19048), .C2(n13266), .A(n13265), .B(n13264), .ZN(
        P2_U2881) );
  OR2_X1 U16579 ( .A1(n13908), .A2(n11025), .ZN(n13267) );
  AND2_X1 U16580 ( .A1(n13268), .A2(n13267), .ZN(n13276) );
  INV_X1 U16581 ( .A(n13269), .ZN(n13271) );
  NOR2_X1 U16582 ( .A1(n13271), .A2(n13270), .ZN(n13275) );
  NOR2_X1 U16583 ( .A1(n15843), .A2(n20593), .ZN(n13272) );
  OAI211_X1 U16584 ( .C1(n15802), .C2(n11376), .A(n13272), .B(n13537), .ZN(
        n13274) );
  NAND4_X1 U16585 ( .A1(n13276), .A2(n13275), .A3(n13274), .A4(n13273), .ZN(
        n15800) );
  NAND2_X1 U16586 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16229), .ZN(n16239) );
  INV_X1 U16587 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19907) );
  OAI22_X1 U16588 ( .A1(n13533), .A2(n13277), .B1(n16239), .B2(n19907), .ZN(
        n13279) );
  AOI21_X1 U16589 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n16236), .A(n13279), 
        .ZN(n14928) );
  INV_X1 U16590 ( .A(n14928), .ZN(n14916) );
  INV_X1 U16591 ( .A(n13604), .ZN(n13561) );
  NOR2_X1 U16592 ( .A1(n11169), .A2(n13561), .ZN(n13278) );
  XNOR2_X1 U16593 ( .A(n13278), .B(n13534), .ZN(n19981) );
  INV_X1 U16594 ( .A(n12386), .ZN(n13531) );
  NAND4_X1 U16595 ( .A1(n19981), .A2(n14262), .A3(n13531), .A4(n13279), .ZN(
        n13280) );
  OAI21_X1 U16596 ( .B1(n13534), .B2(n14916), .A(n13280), .ZN(P1_U3468) );
  OAI21_X1 U16597 ( .B1(n13281), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13282), .ZN(n20068) );
  INV_X1 U16598 ( .A(n14895), .ZN(n13286) );
  INV_X1 U16599 ( .A(n16168), .ZN(n13283) );
  NAND2_X1 U16600 ( .A1(n13283), .A2(n16172), .ZN(n13285) );
  NAND2_X1 U16601 ( .A1(n13285), .A2(n13284), .ZN(n14897) );
  AOI21_X1 U16602 ( .B1(n13286), .B2(n14897), .A(n11402), .ZN(n13289) );
  XNOR2_X1 U16603 ( .A(n13287), .B(n14514), .ZN(n20011) );
  NOR2_X1 U16604 ( .A1(n16210), .A2(n20011), .ZN(n13288) );
  AOI211_X1 U16605 ( .C1(P1_REIP_REG_1__SCAN_IN), .C2(n20106), .A(n13289), .B(
        n13288), .ZN(n13292) );
  INV_X1 U16606 ( .A(n16201), .ZN(n16143) );
  OR3_X1 U16607 ( .A1(n16143), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13290), .ZN(n13291) );
  OAI211_X1 U16608 ( .C1(n20068), .C2(n16186), .A(n13292), .B(n13291), .ZN(
        P1_U3030) );
  OAI21_X1 U16609 ( .B1(n13294), .B2(n13293), .A(n13324), .ZN(n20075) );
  INV_X1 U16610 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20776) );
  OAI222_X1 U16611 ( .A1(n20075), .A2(n14635), .B1(n20023), .B2(n20776), .C1(
        n20011), .C2(n14629), .ZN(P1_U2871) );
  XOR2_X1 U16612 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13295), .Z(n13300)
         );
  INV_X1 U16613 ( .A(n13296), .ZN(n13657) );
  NAND2_X1 U16614 ( .A1(n13261), .A2(n13297), .ZN(n13298) );
  NAND2_X1 U16615 ( .A1(n13657), .A2(n13298), .ZN(n15615) );
  INV_X1 U16616 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13623) );
  MUX2_X1 U16617 ( .A(n15615), .B(n13623), .S(n19052), .Z(n13299) );
  OAI21_X1 U16618 ( .B1(n13300), .B2(n19041), .A(n13299), .ZN(P2_U2880) );
  INV_X1 U16619 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19227) );
  NOR2_X1 U16620 ( .A1(n19227), .A2(n13301), .ZN(n19038) );
  AND2_X1 U16621 ( .A1(n13302), .A2(n19038), .ZN(n13303) );
  AND2_X1 U16622 ( .A1(n13303), .A2(n19037), .ZN(n13304) );
  AND2_X1 U16623 ( .A1(n9755), .A2(n13304), .ZN(n19040) );
  NAND2_X1 U16624 ( .A1(n9755), .A2(n13553), .ZN(n19032) );
  OAI211_X1 U16625 ( .C1(n19040), .C2(n13305), .A(n19018), .B(n19032), .ZN(
        n13310) );
  OR2_X1 U16626 ( .A1(n13656), .A2(n13307), .ZN(n13308) );
  AND2_X1 U16627 ( .A1(n13306), .A2(n13308), .ZN(n18964) );
  NAND2_X1 U16628 ( .A1(n18964), .A2(n19048), .ZN(n13309) );
  OAI211_X1 U16629 ( .C1(n19048), .C2(n10575), .A(n13310), .B(n13309), .ZN(
        P2_U2878) );
  AOI21_X1 U16630 ( .B1(n13313), .B2(n13312), .A(n13311), .ZN(n20699) );
  XOR2_X1 U16631 ( .A(n20699), .B(n20708), .Z(n13318) );
  NAND2_X1 U16632 ( .A1(n19874), .A2(n13314), .ZN(n13315) );
  OAI21_X1 U16633 ( .B1(n19874), .B2(n13314), .A(n13315), .ZN(n19122) );
  NOR2_X1 U16634 ( .A1(n19122), .A2(n19123), .ZN(n19121) );
  INV_X1 U16635 ( .A(n13315), .ZN(n13316) );
  NOR2_X1 U16636 ( .A1(n19121), .A2(n13316), .ZN(n13317) );
  NOR2_X1 U16637 ( .A1(n13318), .A2(n13317), .ZN(n19097) );
  AOI21_X1 U16638 ( .B1(n13318), .B2(n13317), .A(n19097), .ZN(n13321) );
  AOI22_X1 U16639 ( .A1(n19096), .A2(n19197), .B1(n19119), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13320) );
  INV_X1 U16640 ( .A(n20699), .ZN(n14239) );
  NAND2_X1 U16641 ( .A1(n14239), .A2(n19120), .ZN(n13319) );
  OAI211_X1 U16642 ( .C1(n13321), .C2(n19124), .A(n13320), .B(n13319), .ZN(
        P2_U2917) );
  INV_X1 U16643 ( .A(n13322), .ZN(n13323) );
  AOI21_X1 U16644 ( .B1(n13325), .B2(n13324), .A(n13323), .ZN(n13426) );
  INV_X1 U16645 ( .A(n13426), .ZN(n19999) );
  AOI21_X1 U16646 ( .B1(n9786), .B2(n13326), .A(n9900), .ZN(n20099) );
  INV_X1 U16647 ( .A(n20023), .ZN(n14642) );
  AOI22_X1 U16648 ( .A1(n20099), .A2(n20021), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14642), .ZN(n13327) );
  OAI21_X1 U16649 ( .B1(n19999), .B2(n14635), .A(n13327), .ZN(P1_U2870) );
  OAI21_X1 U16650 ( .B1(n13328), .B2(n13331), .A(n13330), .ZN(n13930) );
  XNOR2_X1 U16651 ( .A(n19976), .B(n19972), .ZN(n20086) );
  AOI22_X1 U16652 ( .A1(n20086), .A2(n20021), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14642), .ZN(n13332) );
  OAI21_X1 U16653 ( .B1(n13930), .B2(n14635), .A(n13332), .ZN(P1_U2869) );
  NAND2_X1 U16654 ( .A1(n20677), .A2(n20593), .ZN(n13333) );
  NOR3_X1 U16655 ( .A1(n13336), .A2(n13335), .A3(n20593), .ZN(n13351) );
  NOR2_X1 U16656 ( .A1(n13564), .A2(n13337), .ZN(n13338) );
  AOI21_X1 U16657 ( .B1(DATAI_11_), .B2(n13564), .A(n13338), .ZN(n14217) );
  INV_X1 U16658 ( .A(n14217), .ZN(n16008) );
  NAND2_X1 U16659 ( .A1(n13351), .A2(n16008), .ZN(n20049) );
  NAND2_X1 U16660 ( .A1(n13388), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13339) );
  OAI211_X1 U16661 ( .C1(n13418), .C2(n12022), .A(n20049), .B(n13339), .ZN(
        P1_U2948) );
  INV_X1 U16662 ( .A(DATAI_12_), .ZN(n13340) );
  MUX2_X1 U16663 ( .A(n13340), .B(n16458), .S(n13565), .Z(n14706) );
  INV_X1 U16664 ( .A(n14706), .ZN(n13341) );
  NAND2_X1 U16665 ( .A1(n13351), .A2(n13341), .ZN(n20051) );
  NAND2_X1 U16666 ( .A1(n13388), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13342) );
  OAI211_X1 U16667 ( .C1(n13418), .C2(n14654), .A(n20051), .B(n13342), .ZN(
        P1_U2949) );
  INV_X1 U16668 ( .A(DATAI_9_), .ZN(n13343) );
  MUX2_X1 U16669 ( .A(n13343), .B(n16463), .S(n13565), .Z(n14664) );
  INV_X1 U16670 ( .A(n14664), .ZN(n13344) );
  NAND2_X1 U16671 ( .A1(n13351), .A2(n13344), .ZN(n20047) );
  NAND2_X1 U16672 ( .A1(n13388), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13345) );
  OAI211_X1 U16673 ( .C1(n13418), .C2(n14663), .A(n20047), .B(n13345), .ZN(
        P1_U2946) );
  NOR2_X1 U16674 ( .A1(n13564), .A2(n13346), .ZN(n13347) );
  AOI21_X1 U16675 ( .B1(DATAI_14_), .B2(n13564), .A(n13347), .ZN(n14644) );
  INV_X1 U16676 ( .A(n14644), .ZN(n13348) );
  NAND2_X1 U16677 ( .A1(n13351), .A2(n13348), .ZN(n20055) );
  NAND2_X1 U16678 ( .A1(n13388), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13349) );
  OAI211_X1 U16679 ( .C1(n13418), .C2(n13350), .A(n20055), .B(n13349), .ZN(
        P1_U2951) );
  INV_X1 U16680 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13352) );
  NOR2_X1 U16681 ( .A1(n13564), .A2(n13352), .ZN(n13353) );
  AOI21_X1 U16682 ( .B1(DATAI_15_), .B2(n13564), .A(n13353), .ZN(n14696) );
  INV_X1 U16683 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13354) );
  INV_X1 U16684 ( .A(n13388), .ZN(n13361) );
  OAI222_X1 U16685 ( .A1(n13418), .A2(n20025), .B1(n13387), .B2(n14696), .C1(
        n13354), .C2(n13361), .ZN(P1_U2967) );
  NAND2_X1 U16686 ( .A1(n13564), .A2(DATAI_4_), .ZN(n13356) );
  NAND2_X1 U16687 ( .A1(n13565), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13355) );
  AND2_X1 U16688 ( .A1(n13356), .A2(n13355), .ZN(n16013) );
  NOR2_X1 U16689 ( .A1(n13387), .A2(n16013), .ZN(n13390) );
  AOI21_X1 U16690 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n13388), .A(n13390), 
        .ZN(n13357) );
  OAI21_X1 U16691 ( .B1(n13236), .B2(n13418), .A(n13357), .ZN(P1_U2941) );
  INV_X1 U16692 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20761) );
  NAND2_X1 U16693 ( .A1(n13565), .A2(n20761), .ZN(n13358) );
  OAI21_X1 U16694 ( .B1(n13565), .B2(DATAI_8_), .A(n13358), .ZN(n14668) );
  NOR2_X1 U16695 ( .A1(n13387), .A2(n14668), .ZN(n13407) );
  AOI21_X1 U16696 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n13388), .A(n13407), 
        .ZN(n13359) );
  OAI21_X1 U16697 ( .B1(n13360), .B2(n13418), .A(n13359), .ZN(P1_U2945) );
  NAND2_X1 U16698 ( .A1(n13565), .A2(n16461), .ZN(n13362) );
  OAI21_X1 U16699 ( .B1(n13565), .B2(DATAI_10_), .A(n13362), .ZN(n14659) );
  NOR2_X1 U16700 ( .A1(n13387), .A2(n14659), .ZN(n13404) );
  AOI21_X1 U16701 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n20053), .A(n13404), 
        .ZN(n13363) );
  OAI21_X1 U16702 ( .B1(n13234), .B2(n13418), .A(n13363), .ZN(P1_U2947) );
  NAND2_X1 U16703 ( .A1(n13564), .A2(DATAI_5_), .ZN(n13365) );
  NAND2_X1 U16704 ( .A1(n13565), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13364) );
  AND2_X1 U16705 ( .A1(n13365), .A2(n13364), .ZN(n14684) );
  NOR2_X1 U16706 ( .A1(n13387), .A2(n14684), .ZN(n13414) );
  AOI21_X1 U16707 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n13388), .A(n13414), 
        .ZN(n13366) );
  OAI21_X1 U16708 ( .B1(n20858), .B2(n13418), .A(n13366), .ZN(P1_U2942) );
  NAND2_X1 U16709 ( .A1(n13564), .A2(DATAI_3_), .ZN(n13368) );
  NAND2_X1 U16710 ( .A1(n13565), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13367) );
  AND2_X1 U16711 ( .A1(n13368), .A2(n13367), .ZN(n16017) );
  NOR2_X1 U16712 ( .A1(n13387), .A2(n16017), .ZN(n13409) );
  AOI21_X1 U16713 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n13388), .A(n13409), 
        .ZN(n13369) );
  OAI21_X1 U16714 ( .B1(n13230), .B2(n13418), .A(n13369), .ZN(P1_U2940) );
  NAND2_X1 U16715 ( .A1(n13564), .A2(DATAI_7_), .ZN(n13371) );
  NAND2_X1 U16716 ( .A1(n13565), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13370) );
  AND2_X1 U16717 ( .A1(n13371), .A2(n13370), .ZN(n14674) );
  NOR2_X1 U16718 ( .A1(n13387), .A2(n14674), .ZN(n13416) );
  AOI21_X1 U16719 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n20053), .A(n13416), 
        .ZN(n13372) );
  OAI21_X1 U16720 ( .B1(n14673), .B2(n13418), .A(n13372), .ZN(P1_U2944) );
  INV_X1 U16721 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14649) );
  INV_X1 U16722 ( .A(DATAI_13_), .ZN(n13374) );
  MUX2_X1 U16723 ( .A(n13374), .B(n13373), .S(n13565), .Z(n14698) );
  NOR2_X1 U16724 ( .A1(n13387), .A2(n14698), .ZN(n13401) );
  AOI21_X1 U16725 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n20053), .A(n13401), 
        .ZN(n13375) );
  OAI21_X1 U16726 ( .B1(n14649), .B2(n13418), .A(n13375), .ZN(P1_U2950) );
  NAND2_X1 U16727 ( .A1(n13564), .A2(DATAI_6_), .ZN(n13377) );
  NAND2_X1 U16728 ( .A1(n13565), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13376) );
  AND2_X1 U16729 ( .A1(n13377), .A2(n13376), .ZN(n14680) );
  NOR2_X1 U16730 ( .A1(n13387), .A2(n14680), .ZN(n13412) );
  AOI21_X1 U16731 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n13388), .A(n13412), 
        .ZN(n13378) );
  OAI21_X1 U16732 ( .B1(n14679), .B2(n13418), .A(n13378), .ZN(P1_U2943) );
  NAND2_X1 U16733 ( .A1(n13564), .A2(DATAI_2_), .ZN(n13380) );
  NAND2_X1 U16734 ( .A1(n13565), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13379) );
  AND2_X1 U16735 ( .A1(n13380), .A2(n13379), .ZN(n14689) );
  NOR2_X1 U16736 ( .A1(n13387), .A2(n14689), .ZN(n13398) );
  AOI21_X1 U16737 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n13388), .A(n13398), 
        .ZN(n13381) );
  OAI21_X1 U16738 ( .B1(n13178), .B2(n13418), .A(n13381), .ZN(P1_U2939) );
  NAND2_X1 U16739 ( .A1(n13564), .A2(DATAI_0_), .ZN(n13383) );
  NAND2_X1 U16740 ( .A1(n13565), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13382) );
  AND2_X1 U16741 ( .A1(n13383), .A2(n13382), .ZN(n14212) );
  NOR2_X1 U16742 ( .A1(n13387), .A2(n14212), .ZN(n13392) );
  AOI21_X1 U16743 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n13388), .A(n13392), 
        .ZN(n13384) );
  OAI21_X1 U16744 ( .B1(n13175), .B2(n13418), .A(n13384), .ZN(P1_U2937) );
  NAND2_X1 U16745 ( .A1(n13564), .A2(DATAI_1_), .ZN(n13386) );
  NAND2_X1 U16746 ( .A1(n13565), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13385) );
  AND2_X1 U16747 ( .A1(n13386), .A2(n13385), .ZN(n16021) );
  NOR2_X1 U16748 ( .A1(n13387), .A2(n16021), .ZN(n13395) );
  AOI21_X1 U16749 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n13388), .A(n13395), 
        .ZN(n13389) );
  OAI21_X1 U16750 ( .B1(n13179), .B2(n13418), .A(n13389), .ZN(P1_U2938) );
  INV_X1 U16751 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13738) );
  AOI21_X1 U16752 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n20053), .A(n13390), 
        .ZN(n13391) );
  OAI21_X1 U16753 ( .B1(n13738), .B2(n13418), .A(n13391), .ZN(P1_U2956) );
  INV_X1 U16754 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13394) );
  AOI21_X1 U16755 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n20053), .A(n13392), 
        .ZN(n13393) );
  OAI21_X1 U16756 ( .B1(n13394), .B2(n13418), .A(n13393), .ZN(P1_U2952) );
  AOI21_X1 U16757 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n20053), .A(n13395), 
        .ZN(n13396) );
  OAI21_X1 U16758 ( .B1(n13397), .B2(n13418), .A(n13396), .ZN(P1_U2953) );
  INV_X1 U16759 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13400) );
  AOI21_X1 U16760 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n20053), .A(n13398), 
        .ZN(n13399) );
  OAI21_X1 U16761 ( .B1(n13400), .B2(n13418), .A(n13399), .ZN(P1_U2954) );
  AOI21_X1 U16762 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n20053), .A(n13401), 
        .ZN(n13402) );
  OAI21_X1 U16763 ( .B1(n13403), .B2(n13418), .A(n13402), .ZN(P1_U2965) );
  INV_X1 U16764 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13406) );
  AOI21_X1 U16765 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n20053), .A(n13404), 
        .ZN(n13405) );
  OAI21_X1 U16766 ( .B1(n13406), .B2(n13418), .A(n13405), .ZN(P1_U2962) );
  AOI21_X1 U16767 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n20053), .A(n13407), 
        .ZN(n13408) );
  OAI21_X1 U16768 ( .B1(n13938), .B2(n13418), .A(n13408), .ZN(P1_U2960) );
  AOI21_X1 U16769 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n20053), .A(n13409), 
        .ZN(n13410) );
  OAI21_X1 U16770 ( .B1(n13411), .B2(n13418), .A(n13410), .ZN(P1_U2955) );
  AOI21_X1 U16771 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n20053), .A(n13412), 
        .ZN(n13413) );
  OAI21_X1 U16772 ( .B1(n13846), .B2(n13418), .A(n13413), .ZN(P1_U2958) );
  AOI21_X1 U16773 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n20053), .A(n13414), 
        .ZN(n13415) );
  OAI21_X1 U16774 ( .B1(n13734), .B2(n13418), .A(n13415), .ZN(P1_U2957) );
  INV_X1 U16775 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13419) );
  AOI21_X1 U16776 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n20053), .A(n13416), 
        .ZN(n13417) );
  OAI21_X1 U16777 ( .B1(n13419), .B2(n13418), .A(n13417), .ZN(P1_U2959) );
  OAI21_X1 U16778 ( .B1(n13422), .B2(n13421), .A(n13420), .ZN(n20102) );
  INV_X1 U16779 ( .A(n20001), .ZN(n13424) );
  AOI22_X1 U16780 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U16781 ( .B1(n20066), .B2(n13424), .A(n13423), .ZN(n13425) );
  AOI21_X1 U16782 ( .B1(n13426), .B2(n20062), .A(n13425), .ZN(n13427) );
  OAI21_X1 U16783 ( .B1(n19906), .B2(n20102), .A(n13427), .ZN(P1_U2997) );
  INV_X1 U16784 ( .A(n13448), .ZN(n13464) );
  AND2_X1 U16785 ( .A1(n10266), .A2(n13428), .ZN(n13456) );
  NAND2_X1 U16786 ( .A1(n10120), .A2(n13430), .ZN(n13435) );
  INV_X1 U16787 ( .A(n13431), .ZN(n13474) );
  OR2_X1 U16788 ( .A1(n13474), .A2(n13470), .ZN(n13453) );
  NOR2_X1 U16789 ( .A1(n13432), .A2(n9710), .ZN(n13433) );
  AOI22_X1 U16790 ( .A1(n13453), .A2(n13435), .B1(n13433), .B2(n12374), .ZN(
        n13434) );
  OAI21_X1 U16791 ( .B1(n13456), .B2(n13435), .A(n13434), .ZN(n13436) );
  AOI21_X1 U16792 ( .B1(n13180), .B2(n13464), .A(n13436), .ZN(n13466) );
  INV_X1 U16793 ( .A(n13438), .ZN(n13439) );
  NOR2_X1 U16794 ( .A1(n12165), .A2(n13439), .ZN(n13445) );
  NOR3_X1 U16795 ( .A1(n13445), .A2(n13429), .A3(n13440), .ZN(n13443) );
  NOR2_X1 U16796 ( .A1(n13441), .A2(n13448), .ZN(n13442) );
  AOI211_X1 U16797 ( .C1(n13437), .C2(n12374), .A(n13443), .B(n13442), .ZN(
        n15636) );
  INV_X1 U16798 ( .A(n19547), .ZN(n19296) );
  AOI21_X1 U16799 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n15636), .A(
        n19296), .ZN(n13451) );
  INV_X1 U16800 ( .A(n12374), .ZN(n13446) );
  MUX2_X1 U16801 ( .A(n13446), .B(n13445), .S(n13444), .Z(n13447) );
  OAI21_X1 U16802 ( .B1(n13449), .B2(n13448), .A(n13447), .ZN(n13775) );
  NAND2_X1 U16803 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15636), .ZN(
        n13450) );
  OAI211_X1 U16804 ( .C1(n13451), .C2(n13775), .A(n13485), .B(n13450), .ZN(
        n13452) );
  AOI21_X1 U16805 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13466), .A(
        n13452), .ZN(n13467) );
  AND2_X1 U16806 ( .A1(n13453), .A2(n10120), .ZN(n13458) );
  INV_X1 U16807 ( .A(n13454), .ZN(n13455) );
  NAND2_X1 U16808 ( .A1(n12374), .A2(n13455), .ZN(n13461) );
  OAI211_X1 U16809 ( .C1(n10333), .C2(n13456), .A(n10120), .B(n13461), .ZN(
        n13457) );
  MUX2_X1 U16810 ( .A(n13458), .B(n13457), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13463) );
  INV_X1 U16811 ( .A(n10326), .ZN(n13460) );
  INV_X1 U16812 ( .A(n10354), .ZN(n13459) );
  OAI21_X1 U16813 ( .B1(n13461), .B2(n13460), .A(n13459), .ZN(n13462) );
  NOR2_X1 U16814 ( .A1(n13485), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13465) );
  AOI21_X1 U16815 ( .B1(n15640), .B2(n13485), .A(n13465), .ZN(n13483) );
  OAI21_X1 U16816 ( .B1(n13467), .B2(n19864), .A(n13483), .ZN(n13469) );
  INV_X1 U16817 ( .A(n13466), .ZN(n13841) );
  MUX2_X1 U16818 ( .A(n14352), .B(n13841), .S(n13485), .Z(n13482) );
  NAND2_X1 U16819 ( .A1(n19864), .A2(n19871), .ZN(n19266) );
  INV_X1 U16820 ( .A(n19266), .ZN(n19295) );
  AOI22_X1 U16821 ( .A1(n13482), .A2(n19295), .B1(n13467), .B2(n19864), .ZN(
        n13468) );
  NAND2_X1 U16822 ( .A1(n13469), .A2(n13468), .ZN(n13489) );
  INV_X1 U16823 ( .A(n13470), .ZN(n13472) );
  INV_X1 U16824 ( .A(n13476), .ZN(n13471) );
  OAI22_X1 U16825 ( .A1(n13472), .A2(n13773), .B1(n10238), .B2(n13471), .ZN(
        n13473) );
  AOI21_X1 U16826 ( .B1(n13474), .B2(n13773), .A(n13473), .ZN(n19893) );
  OR2_X1 U16827 ( .A1(n10717), .A2(n13475), .ZN(n19894) );
  OR2_X1 U16828 ( .A1(n14934), .A2(n19787), .ZN(n13477) );
  AOI21_X1 U16829 ( .B1(n13477), .B2(n15862), .A(n13476), .ZN(n13478) );
  NAND2_X1 U16830 ( .A1(n12368), .A2(n13478), .ZN(n18863) );
  NOR2_X1 U16831 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n13479) );
  OR2_X1 U16832 ( .A1(n18863), .A2(n13479), .ZN(n13480) );
  NAND4_X1 U16833 ( .A1(n19893), .A2(n13481), .A3(n19894), .A4(n13480), .ZN(
        n13488) );
  NAND2_X1 U16834 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  OAI21_X1 U16835 ( .B1(n13486), .B2(n13485), .A(n13484), .ZN(n13487) );
  AOI211_X1 U16836 ( .C1(n15870), .C2(n13489), .A(n13488), .B(n13487), .ZN(
        n16371) );
  AOI21_X1 U16837 ( .B1(n16371), .B2(n13837), .A(n16380), .ZN(n13496) );
  NAND2_X1 U16838 ( .A1(n13491), .A2(n13490), .ZN(n13493) );
  NOR2_X1 U16839 ( .A1(n13492), .A2(n19723), .ZN(n14942) );
  OAI21_X1 U16840 ( .B1(n13494), .B2(n13493), .A(n14942), .ZN(n13495) );
  OAI211_X1 U16841 ( .C1(n16367), .C2(n19668), .A(n13497), .B(n15863), .ZN(
        P2_U3593) );
  NOR2_X1 U16842 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16233), .ZN(n13536) );
  INV_X1 U16843 ( .A(n20125), .ZN(n13518) );
  NAND2_X1 U16844 ( .A1(n13498), .A2(n12384), .ZN(n13499) );
  NOR2_X1 U16845 ( .A1(n13499), .A2(n11376), .ZN(n13501) );
  AND3_X1 U16846 ( .A1(n12386), .A2(n13501), .A3(n13500), .ZN(n14907) );
  INV_X1 U16847 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13508) );
  INV_X1 U16848 ( .A(n13503), .ZN(n13504) );
  OAI21_X1 U16849 ( .B1(n13502), .B2(n13508), .A(n13504), .ZN(n13505) );
  NOR2_X1 U16850 ( .A1(n13505), .A2(n11051), .ZN(n14925) );
  INV_X1 U16851 ( .A(n14257), .ZN(n14908) );
  AND2_X1 U16852 ( .A1(n11014), .A2(n13904), .ZN(n13506) );
  NAND2_X1 U16853 ( .A1(n14908), .A2(n13506), .ZN(n13524) );
  MUX2_X1 U16854 ( .A(n13513), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n11113), .Z(n13507) );
  OAI21_X1 U16855 ( .B1(n13503), .B2(n13507), .A(n15802), .ZN(n13515) );
  MUX2_X1 U16856 ( .A(n13503), .B(n13508), .S(n13502), .Z(n13512) );
  INV_X1 U16857 ( .A(n13509), .ZN(n13511) );
  NAND2_X1 U16858 ( .A1(n13511), .A2(n13510), .ZN(n13520) );
  OAI21_X1 U16859 ( .B1(n13513), .B2(n13512), .A(n13520), .ZN(n13514) );
  OAI211_X1 U16860 ( .C1(n14925), .C2(n13524), .A(n13515), .B(n13514), .ZN(
        n13516) );
  INV_X1 U16861 ( .A(n13516), .ZN(n13517) );
  OAI21_X1 U16862 ( .B1(n13518), .B2(n14907), .A(n13517), .ZN(n14924) );
  MUX2_X1 U16863 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14924), .S(
        n15800), .Z(n15814) );
  AOI22_X1 U16864 ( .A1(n13536), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16233), .B2(n15814), .ZN(n13529) );
  OR2_X1 U16865 ( .A1(n13519), .A2(n14907), .ZN(n13527) );
  XNOR2_X1 U16866 ( .A(n13502), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14922) );
  NAND2_X1 U16867 ( .A1(n13520), .A2(n14922), .ZN(n13523) );
  XNOR2_X1 U16868 ( .A(n11113), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13521) );
  NAND2_X1 U16869 ( .A1(n15802), .A2(n13521), .ZN(n13522) );
  OAI211_X1 U16870 ( .C1(n14922), .C2(n13524), .A(n13523), .B(n13522), .ZN(
        n13525) );
  INV_X1 U16871 ( .A(n13525), .ZN(n13526) );
  NAND2_X1 U16872 ( .A1(n13527), .A2(n13526), .ZN(n14918) );
  MUX2_X1 U16873 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14918), .S(
        n15800), .Z(n15809) );
  AOI22_X1 U16874 ( .A1(n15809), .A2(n16233), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13536), .ZN(n13528) );
  OR2_X1 U16875 ( .A1(n13529), .A2(n13528), .ZN(n15822) );
  OR2_X1 U16876 ( .A1(n15822), .A2(n13530), .ZN(n13539) );
  AOI21_X1 U16877 ( .B1(n19981), .B2(n13531), .A(n13533), .ZN(n13532) );
  AOI211_X1 U16878 ( .C1(n13534), .C2(n13533), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13532), .ZN(n13535) );
  AOI21_X1 U16879 ( .B1(n13536), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13535), .ZN(n15824) );
  AND3_X1 U16880 ( .A1(n13539), .A2(n19907), .A3(n15824), .ZN(n13538) );
  NOR2_X1 U16881 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20680) );
  OAI21_X1 U16882 ( .B1(n13538), .B2(n16239), .A(n14046), .ZN(n20113) );
  NAND3_X1 U16883 ( .A1(n13539), .A2(n15824), .A3(n16229), .ZN(n15828) );
  INV_X1 U16884 ( .A(n15828), .ZN(n13542) );
  INV_X1 U16885 ( .A(n11624), .ZN(n13540) );
  INV_X1 U16886 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20439) );
  NAND2_X1 U16887 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20439), .ZN(n13590) );
  INV_X1 U16888 ( .A(n13590), .ZN(n14905) );
  OAI22_X1 U16889 ( .A1(n11622), .A2(n20530), .B1(n13540), .B2(n14905), .ZN(
        n13541) );
  OAI21_X1 U16890 ( .B1(n13542), .B2(n13541), .A(n20113), .ZN(n13543) );
  OAI21_X1 U16891 ( .B1(n20113), .B2(n20317), .A(n13543), .ZN(P1_U3478) );
  AND2_X1 U16892 ( .A1(n13544), .A2(n11008), .ZN(n13547) );
  INV_X1 U16893 ( .A(n13547), .ZN(n13545) );
  AND2_X1 U16894 ( .A1(n13545), .A2(n11010), .ZN(n13546) );
  OAI222_X1 U16895 ( .A1(n16009), .A2(n20075), .B1(n14705), .B2(n16021), .C1(
        n14695), .C2(n13397), .ZN(P1_U2903) );
  OAI222_X1 U16896 ( .A1(n16009), .A2(n13930), .B1(n14705), .B2(n16017), .C1(
        n14695), .C2(n13411), .ZN(P1_U2901) );
  OAI222_X1 U16897 ( .A1(n16009), .A2(n13983), .B1(n14212), .B2(n14705), .C1(
        n14695), .C2(n13394), .ZN(P1_U2904) );
  OAI222_X1 U16898 ( .A1(n16009), .A2(n19999), .B1(n14689), .B2(n14705), .C1(
        n14695), .C2(n13400), .ZN(P1_U2902) );
  NOR2_X1 U16899 ( .A1(n13550), .A2(n13551), .ZN(n13552) );
  OR2_X1 U16900 ( .A1(n13549), .A2(n13552), .ZN(n15555) );
  OAI211_X1 U16901 ( .C1(n13558), .C2(n13557), .A(n13858), .B(n19018), .ZN(
        n13560) );
  NAND2_X1 U16902 ( .A1(n19052), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13559) );
  OAI211_X1 U16903 ( .C1(n15555), .C2(n19052), .A(n13560), .B(n13559), .ZN(
        P2_U2875) );
  NAND2_X1 U16904 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20523) );
  NOR2_X1 U16905 ( .A1(n20523), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13566) );
  OAI21_X1 U16906 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20439), .A(
        n13953), .ZN(n20396) );
  INV_X1 U16907 ( .A(n20396), .ZN(n20536) );
  NAND2_X1 U16908 ( .A1(n20115), .A2(n13587), .ZN(n20529) );
  NOR2_X1 U16909 ( .A1(n13519), .A2(n13561), .ZN(n20522) );
  INV_X1 U16910 ( .A(n13562), .ZN(n20318) );
  NOR3_X1 U16911 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20317), .A3(
        n20523), .ZN(n13570) );
  AOI21_X1 U16912 ( .B1(n20522), .B2(n20318), .A(n13570), .ZN(n13568) );
  OAI211_X1 U16913 ( .C1(n20529), .C2(n20321), .A(n20389), .B(n13568), .ZN(
        n13563) );
  OAI211_X1 U16914 ( .C1(n20538), .C2(n13566), .A(n20536), .B(n13563), .ZN(
        n13718) );
  AOI22_X1 U16915 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13700), .B1(DATAI_27_), 
        .B2(n13699), .ZN(n20461) );
  INV_X1 U16916 ( .A(n11622), .ZN(n13609) );
  OAI22_X1 U16917 ( .A1(n9856), .A2(n20479), .B1(n20491), .B2(n20560), .ZN(
        n13572) );
  NOR2_X2 U16918 ( .A1(n16017), .A2(n14046), .ZN(n20557) );
  INV_X1 U16919 ( .A(n20557), .ZN(n14062) );
  INV_X1 U16920 ( .A(n13566), .ZN(n13567) );
  OAI22_X1 U16921 ( .A1(n13568), .A2(n20530), .B1(n13567), .B2(n20525), .ZN(
        n13569) );
  INV_X1 U16922 ( .A(n13569), .ZN(n13715) );
  INV_X1 U16923 ( .A(n13570), .ZN(n13714) );
  OAI22_X1 U16924 ( .A1(n14062), .A2(n13715), .B1(n20457), .B2(n13714), .ZN(
        n13571) );
  AOI211_X1 U16925 ( .C1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .C2(n13718), .A(
        n13572), .B(n13571), .ZN(n13573) );
  INV_X1 U16926 ( .A(n13573), .ZN(P1_U3140) );
  OAI22_X1 U16927 ( .A1(n20466), .A2(n20479), .B1(n20491), .B2(n20566), .ZN(
        n13576) );
  NOR2_X2 U16928 ( .A1(n16013), .A2(n14046), .ZN(n20562) );
  INV_X1 U16929 ( .A(n20562), .ZN(n14066) );
  AND2_X1 U16930 ( .A1(n13574), .A2(n13701), .ZN(n20561) );
  OAI22_X1 U16931 ( .A1(n14066), .A2(n13715), .B1(n20462), .B2(n13714), .ZN(
        n13575) );
  AOI211_X1 U16932 ( .C1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .C2(n13718), .A(
        n13576), .B(n13575), .ZN(n13577) );
  INV_X1 U16933 ( .A(n13577), .ZN(P1_U3141) );
  AOI22_X1 U16934 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13700), .B1(DATAI_29_), 
        .B2(n13699), .ZN(n20471) );
  OAI22_X1 U16935 ( .A1(n9854), .A2(n20479), .B1(n20491), .B2(n20571), .ZN(
        n13579) );
  NOR2_X2 U16936 ( .A1(n14684), .A2(n14046), .ZN(n20568) );
  INV_X1 U16937 ( .A(n20568), .ZN(n14074) );
  OAI22_X1 U16938 ( .A1(n14074), .A2(n13715), .B1(n20467), .B2(n13714), .ZN(
        n13578) );
  AOI211_X1 U16939 ( .C1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .C2(n13718), .A(
        n13579), .B(n13578), .ZN(n13580) );
  INV_X1 U16940 ( .A(n13580), .ZN(P1_U3142) );
  AOI22_X1 U16941 ( .A1(DATAI_23_), .A2(n13699), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n13700), .ZN(n20588) );
  OAI22_X1 U16942 ( .A1(n20486), .A2(n20479), .B1(n20491), .B2(n9850), .ZN(
        n13582) );
  NOR2_X2 U16943 ( .A1(n14674), .A2(n14046), .ZN(n20581) );
  INV_X1 U16944 ( .A(n20581), .ZN(n14078) );
  OAI22_X1 U16945 ( .A1(n14078), .A2(n13715), .B1(n20477), .B2(n13714), .ZN(
        n13581) );
  AOI211_X1 U16946 ( .C1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .C2(n13718), .A(
        n13582), .B(n13581), .ZN(n13583) );
  INV_X1 U16947 ( .A(n13583), .ZN(P1_U3144) );
  AOI22_X1 U16948 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13700), .B1(DATAI_22_), 
        .B2(n13699), .ZN(n20577) );
  OAI22_X1 U16949 ( .A1(n20476), .A2(n20479), .B1(n20491), .B2(n9852), .ZN(
        n13585) );
  NOR2_X2 U16950 ( .A1(n14680), .A2(n14046), .ZN(n20573) );
  INV_X1 U16951 ( .A(n20573), .ZN(n14093) );
  OAI22_X1 U16952 ( .A1(n14093), .A2(n13715), .B1(n20472), .B2(n13714), .ZN(
        n13584) );
  AOI211_X1 U16953 ( .C1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .C2(n13718), .A(
        n13585), .B(n13584), .ZN(n13586) );
  INV_X1 U16954 ( .A(n13586), .ZN(P1_U3143) );
  INV_X1 U16955 ( .A(n20113), .ZN(n13595) );
  INV_X1 U16956 ( .A(n13587), .ZN(n13588) );
  MUX2_X1 U16957 ( .A(n20529), .B(n20292), .S(n14902), .Z(n13589) );
  NAND3_X1 U16958 ( .A1(n13589), .A2(n20390), .A3(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13592) );
  AOI21_X1 U16959 ( .B1(n20117), .B2(n20321), .A(n20530), .ZN(n13591) );
  AOI22_X1 U16960 ( .A1(n13592), .A2(n13591), .B1(n13590), .B2(n20125), .ZN(
        n13594) );
  NAND2_X1 U16961 ( .A1(n13595), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13593) );
  OAI21_X1 U16962 ( .B1(n13595), .B2(n13594), .A(n13593), .ZN(P1_U3475) );
  OAI21_X1 U16963 ( .B1(n13598), .B2(n13597), .A(n13596), .ZN(n20087) );
  INV_X1 U16964 ( .A(n13930), .ZN(n13601) );
  NAND2_X1 U16965 ( .A1(n20106), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20084) );
  NAND2_X1 U16966 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13599) );
  OAI211_X1 U16967 ( .C1(n20066), .C2(n13923), .A(n20084), .B(n13599), .ZN(
        n13600) );
  AOI21_X1 U16968 ( .B1(n13601), .B2(n20062), .A(n13600), .ZN(n13602) );
  OAI21_X1 U16969 ( .B1(n20087), .B2(n19906), .A(n13602), .ZN(P1_U2996) );
  OR2_X1 U16970 ( .A1(n14902), .A2(n20530), .ZN(n13603) );
  NAND2_X1 U16971 ( .A1(n20389), .A2(n20321), .ZN(n20434) );
  NAND2_X1 U16972 ( .A1(n13603), .A2(n20434), .ZN(n20533) );
  AOI21_X1 U16973 ( .B1(n20292), .B2(n20389), .A(n20533), .ZN(n13608) );
  NOR2_X1 U16974 ( .A1(n13519), .A2(n13604), .ZN(n20289) );
  INV_X1 U16975 ( .A(n20289), .ZN(n13606) );
  NAND2_X1 U16976 ( .A1(n11624), .A2(n13605), .ZN(n20519) );
  OAI21_X1 U16977 ( .B1(n13606), .B2(n20519), .A(n13702), .ZN(n13611) );
  NAND2_X1 U16978 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20288), .ZN(
        n14044) );
  AOI21_X1 U16979 ( .B1(n20530), .B2(n14044), .A(n20396), .ZN(n13607) );
  OAI21_X1 U16980 ( .B1(n13608), .B2(n13611), .A(n13607), .ZN(n13706) );
  NAND2_X1 U16981 ( .A1(n14902), .A2(n13609), .ZN(n20402) );
  NAND2_X1 U16982 ( .A1(n14902), .A2(n11622), .ZN(n20487) );
  OAI22_X1 U16983 ( .A1(n20560), .A2(n13989), .B1(n14089), .B2(n9856), .ZN(
        n13613) );
  INV_X1 U16984 ( .A(n14044), .ZN(n13610) );
  AOI22_X1 U16985 ( .A1(n13611), .A2(n20389), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13610), .ZN(n13703) );
  OAI22_X1 U16986 ( .A1(n14062), .A2(n13703), .B1(n13702), .B2(n20457), .ZN(
        n13612) );
  AOI211_X1 U16987 ( .C1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .C2(n13706), .A(
        n13613), .B(n13612), .ZN(n13614) );
  INV_X1 U16988 ( .A(n13614), .ZN(P1_U3092) );
  OAI22_X1 U16989 ( .A1(n20566), .A2(n13989), .B1(n14089), .B2(n20466), .ZN(
        n13616) );
  OAI22_X1 U16990 ( .A1(n14066), .A2(n13703), .B1(n13702), .B2(n20462), .ZN(
        n13615) );
  AOI211_X1 U16991 ( .C1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .C2(n13706), .A(
        n13616), .B(n13615), .ZN(n13617) );
  INV_X1 U16992 ( .A(n13617), .ZN(P1_U3093) );
  NOR2_X1 U16993 ( .A1(n10032), .A2(n13618), .ZN(n13619) );
  XNOR2_X1 U16994 ( .A(n13619), .B(n15344), .ZN(n13630) );
  XOR2_X1 U16995 ( .A(n13621), .B(n13620), .Z(n19090) );
  INV_X1 U16996 ( .A(n20698), .ZN(n19002) );
  NAND2_X1 U16997 ( .A1(n19090), .A2(n19002), .ZN(n13628) );
  OAI22_X1 U16998 ( .A1(n13623), .A2(n18999), .B1(n19005), .B2(n13622), .ZN(
        n13624) );
  AOI211_X1 U16999 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18986), .A(n13624), .B(
        n18985), .ZN(n13625) );
  INV_X1 U17000 ( .A(n13625), .ZN(n13626) );
  AOI21_X1 U17001 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19012), .A(
        n13626), .ZN(n13627) );
  OAI211_X1 U17002 ( .C1(n15615), .C2(n20705), .A(n13628), .B(n13627), .ZN(
        n13629) );
  AOI21_X1 U17003 ( .B1(n13630), .B2(n19009), .A(n13629), .ZN(n13631) );
  INV_X1 U17004 ( .A(n13631), .ZN(P2_U2848) );
  OAI22_X1 U17005 ( .A1(n20571), .A2(n13989), .B1(n14089), .B2(n9854), .ZN(
        n13633) );
  OAI22_X1 U17006 ( .A1(n14074), .A2(n13703), .B1(n13702), .B2(n20467), .ZN(
        n13632) );
  AOI211_X1 U17007 ( .C1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .C2(n13706), .A(
        n13633), .B(n13632), .ZN(n13634) );
  INV_X1 U17008 ( .A(n13634), .ZN(P1_U3094) );
  OAI22_X1 U17009 ( .A1(n9850), .A2(n13989), .B1(n14089), .B2(n20486), .ZN(
        n13636) );
  OAI22_X1 U17010 ( .A1(n14078), .A2(n13703), .B1(n13702), .B2(n20477), .ZN(
        n13635) );
  AOI211_X1 U17011 ( .C1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .C2(n13706), .A(
        n13636), .B(n13635), .ZN(n13637) );
  INV_X1 U17012 ( .A(n13637), .ZN(P1_U3096) );
  OAI22_X1 U17013 ( .A1(n9852), .A2(n13989), .B1(n14089), .B2(n20476), .ZN(
        n13639) );
  OAI22_X1 U17014 ( .A1(n14093), .A2(n13703), .B1(n13702), .B2(n20472), .ZN(
        n13638) );
  AOI211_X1 U17015 ( .C1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .C2(n13706), .A(
        n13639), .B(n13638), .ZN(n13640) );
  INV_X1 U17016 ( .A(n13640), .ZN(P1_U3095) );
  INV_X1 U17017 ( .A(n20707), .ZN(n13692) );
  NOR2_X1 U17018 ( .A1(n10032), .A2(n13641), .ZN(n13642) );
  XNOR2_X1 U17019 ( .A(n13642), .B(n13803), .ZN(n13643) );
  NAND2_X1 U17020 ( .A1(n13643), .A2(n19009), .ZN(n13655) );
  INV_X1 U17021 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13804) );
  OAI22_X1 U17022 ( .A1(n18999), .A2(n13644), .B1(n13804), .B2(n18981), .ZN(
        n13645) );
  AOI21_X1 U17023 ( .B1(n18986), .B2(P2_REIP_REG_3__SCAN_IN), .A(n13645), .ZN(
        n13646) );
  OAI21_X1 U17024 ( .B1(n13647), .B2(n19005), .A(n13646), .ZN(n13653) );
  OR2_X1 U17025 ( .A1(n13649), .A2(n13648), .ZN(n13651) );
  NAND2_X1 U17026 ( .A1(n13651), .A2(n13650), .ZN(n19861) );
  NOR2_X1 U17027 ( .A1(n19861), .A2(n20698), .ZN(n13652) );
  AOI211_X1 U17028 ( .C1(n19007), .C2(n13207), .A(n13653), .B(n13652), .ZN(
        n13654) );
  OAI211_X1 U17029 ( .C1(n13692), .C2(n19445), .A(n13655), .B(n13654), .ZN(
        P2_U2852) );
  AOI21_X1 U17030 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(n16358) );
  INV_X1 U17031 ( .A(n16358), .ZN(n19046) );
  NAND2_X1 U17032 ( .A1(n10012), .A2(n13660), .ZN(n13661) );
  XNOR2_X1 U17033 ( .A(n16329), .B(n13661), .ZN(n13662) );
  NAND2_X1 U17034 ( .A1(n13662), .A2(n19009), .ZN(n13672) );
  NOR2_X1 U17035 ( .A1(n20697), .A2(n13663), .ZN(n13669) );
  AOI21_X1 U17036 ( .B1(n13666), .B2(n13665), .A(n13664), .ZN(n16353) );
  INV_X1 U17037 ( .A(n16353), .ZN(n19088) );
  AOI22_X1 U17038 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n20694), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19012), .ZN(n13667) );
  OAI211_X1 U17039 ( .C1(n19088), .C2(n20698), .A(n13667), .B(n18933), .ZN(
        n13668) );
  AOI211_X1 U17040 ( .C1(n13670), .C2(n20703), .A(n13669), .B(n13668), .ZN(
        n13671) );
  OAI211_X1 U17041 ( .C1(n19046), .C2(n20705), .A(n13672), .B(n13671), .ZN(
        P2_U2847) );
  OR2_X1 U17042 ( .A1(n9755), .A2(n19037), .ZN(n13673) );
  NAND2_X1 U17043 ( .A1(n13674), .A2(n13673), .ZN(n19105) );
  AND2_X1 U17044 ( .A1(n10012), .A2(n13675), .ZN(n13677) );
  AOI21_X1 U17045 ( .B1(n13932), .B2(n13677), .A(n12836), .ZN(n13676) );
  OAI21_X1 U17046 ( .B1(n13932), .B2(n13677), .A(n13676), .ZN(n13691) );
  NOR2_X1 U17047 ( .A1(n13678), .A2(n13679), .ZN(n13680) );
  OR2_X1 U17048 ( .A1(n13247), .A2(n13680), .ZN(n19051) );
  INV_X1 U17049 ( .A(n19051), .ZN(n13885) );
  INV_X1 U17050 ( .A(n13650), .ZN(n13681) );
  OR2_X1 U17051 ( .A1(n13682), .A2(n13681), .ZN(n13684) );
  INV_X1 U17052 ( .A(n9840), .ZN(n13683) );
  AND2_X1 U17053 ( .A1(n13684), .A2(n13683), .ZN(n19103) );
  AOI22_X1 U17054 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n20694), .B1(n19002), .B2(
        n19103), .ZN(n13685) );
  OAI211_X1 U17055 ( .C1(n20697), .C2(n12251), .A(n13685), .B(n18933), .ZN(
        n13686) );
  AOI21_X1 U17056 ( .B1(n19012), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13686), .ZN(n13687) );
  OAI21_X1 U17057 ( .B1(n13688), .B2(n19005), .A(n13687), .ZN(n13689) );
  AOI21_X1 U17058 ( .B1(n13885), .B2(n19007), .A(n13689), .ZN(n13690) );
  OAI211_X1 U17059 ( .C1(n19105), .C2(n13692), .A(n13691), .B(n13690), .ZN(
        P2_U2851) );
  AOI22_X1 U17060 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n13700), .B1(DATAI_25_), 
        .B2(n13699), .ZN(n20451) );
  OAI22_X1 U17061 ( .A1(n20549), .A2(n13989), .B1(n14089), .B2(n9858), .ZN(
        n13694) );
  NOR2_X2 U17062 ( .A1(n16021), .A2(n14046), .ZN(n20546) );
  INV_X1 U17063 ( .A(n20546), .ZN(n14058) );
  AND2_X1 U17064 ( .A1(n11022), .A2(n13701), .ZN(n20545) );
  OAI22_X1 U17065 ( .A1(n14058), .A2(n13703), .B1(n13702), .B2(n20447), .ZN(
        n13693) );
  AOI211_X1 U17066 ( .C1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .C2(n13706), .A(
        n13694), .B(n13693), .ZN(n13695) );
  INV_X1 U17067 ( .A(n13695), .ZN(P1_U3090) );
  AOI22_X1 U17068 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n13700), .B1(DATAI_18_), 
        .B2(n13699), .ZN(n20555) );
  OAI22_X1 U17069 ( .A1(n20555), .A2(n13989), .B1(n14089), .B2(n20456), .ZN(
        n13697) );
  NOR2_X2 U17070 ( .A1(n14689), .A2(n14046), .ZN(n20551) );
  INV_X1 U17071 ( .A(n20551), .ZN(n14054) );
  AND2_X1 U17072 ( .A1(n11025), .A2(n13701), .ZN(n20550) );
  OAI22_X1 U17073 ( .A1(n14054), .A2(n13703), .B1(n13702), .B2(n20452), .ZN(
        n13696) );
  AOI211_X1 U17074 ( .C1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .C2(n13706), .A(
        n13697), .B(n13696), .ZN(n13698) );
  INV_X1 U17075 ( .A(n13698), .ZN(P1_U3091) );
  AOI22_X1 U17076 ( .A1(DATAI_16_), .A2(n13699), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n13700), .ZN(n20500) );
  OAI22_X1 U17077 ( .A1(n20500), .A2(n13989), .B1(n14089), .B2(n20544), .ZN(
        n13705) );
  NOR2_X2 U17078 ( .A1(n14212), .A2(n14046), .ZN(n20528) );
  INV_X1 U17079 ( .A(n20528), .ZN(n14070) );
  AND2_X1 U17080 ( .A1(n11328), .A2(n13701), .ZN(n20527) );
  OAI22_X1 U17081 ( .A1(n14070), .A2(n13703), .B1(n13702), .B2(n20432), .ZN(
        n13704) );
  AOI211_X1 U17082 ( .C1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .C2(n13706), .A(
        n13705), .B(n13704), .ZN(n13707) );
  INV_X1 U17083 ( .A(n13707), .ZN(P1_U3089) );
  OAI22_X1 U17084 ( .A1(n20456), .A2(n20479), .B1(n20491), .B2(n20555), .ZN(
        n13709) );
  OAI22_X1 U17085 ( .A1(n14054), .A2(n13715), .B1(n20452), .B2(n13714), .ZN(
        n13708) );
  AOI211_X1 U17086 ( .C1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .C2(n13718), .A(
        n13709), .B(n13708), .ZN(n13710) );
  INV_X1 U17087 ( .A(n13710), .ZN(P1_U3139) );
  OAI22_X1 U17088 ( .A1(n9858), .A2(n20479), .B1(n20491), .B2(n20549), .ZN(
        n13712) );
  OAI22_X1 U17089 ( .A1(n14058), .A2(n13715), .B1(n20447), .B2(n13714), .ZN(
        n13711) );
  AOI211_X1 U17090 ( .C1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .C2(n13718), .A(
        n13712), .B(n13711), .ZN(n13713) );
  INV_X1 U17091 ( .A(n13713), .ZN(P1_U3138) );
  OAI22_X1 U17092 ( .A1(n20544), .A2(n20479), .B1(n20491), .B2(n20500), .ZN(
        n13717) );
  OAI22_X1 U17093 ( .A1(n14070), .A2(n13715), .B1(n20432), .B2(n13714), .ZN(
        n13716) );
  AOI211_X1 U17094 ( .C1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .C2(n13718), .A(
        n13717), .B(n13716), .ZN(n13719) );
  INV_X1 U17095 ( .A(n13719), .ZN(P1_U3137) );
  XNOR2_X1 U17096 ( .A(n13720), .B(n13721), .ZN(n13727) );
  AND2_X1 U17097 ( .A1(n13722), .A2(n13723), .ZN(n13724) );
  OR2_X1 U17098 ( .A1(n13724), .A2(n13550), .ZN(n18932) );
  MUX2_X1 U17099 ( .A(n18932), .B(n13725), .S(n19052), .Z(n13726) );
  OAI21_X1 U17100 ( .B1(n13727), .B2(n19041), .A(n13726), .ZN(P2_U2876) );
  NOR2_X1 U17101 ( .A1(n13728), .A2(n13729), .ZN(n13730) );
  OR2_X1 U17102 ( .A1(n9820), .A2(n13730), .ZN(n16101) );
  AND2_X1 U17103 ( .A1(n19977), .A2(n13731), .ZN(n13732) );
  NOR2_X1 U17104 ( .A1(n16218), .A2(n13732), .ZN(n13770) );
  INV_X1 U17105 ( .A(n13770), .ZN(n19966) );
  OAI222_X1 U17106 ( .A1(n16101), .A2(n14635), .B1(n13733), .B2(n20023), .C1(
        n14629), .C2(n19966), .ZN(P1_U2867) );
  OAI222_X1 U17107 ( .A1(n16101), .A2(n16009), .B1(n14684), .B2(n14705), .C1(
        n13734), .C2(n14695), .ZN(P1_U2899) );
  INV_X1 U17108 ( .A(n13735), .ZN(n13736) );
  XNOR2_X1 U17109 ( .A(n13330), .B(n13736), .ZN(n20061) );
  INV_X1 U17110 ( .A(n20061), .ZN(n13737) );
  OAI222_X1 U17111 ( .A1(n13738), .A2(n14695), .B1(n16009), .B2(n13737), .C1(
        n16013), .C2(n14705), .ZN(P1_U2900) );
  NOR2_X1 U17112 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16380), .ZN(n13740) );
  INV_X1 U17113 ( .A(n16367), .ZN(n13743) );
  NAND2_X1 U17114 ( .A1(n13743), .A2(n19793), .ZN(n16375) );
  INV_X1 U17115 ( .A(n16375), .ZN(n13739) );
  AOI21_X1 U17116 ( .B1(n19793), .B2(n13740), .A(n13739), .ZN(n13745) );
  NOR2_X1 U17117 ( .A1(n19793), .A2(n16380), .ZN(n13741) );
  AOI21_X1 U17118 ( .B1(n13840), .B2(n13741), .A(n18862), .ZN(n13742) );
  OR2_X1 U17119 ( .A1(n13743), .A2(n13742), .ZN(n13744) );
  OAI211_X1 U17120 ( .C1(n13745), .C2(n13837), .A(n12836), .B(n13744), .ZN(
        P2_U3177) );
  NAND2_X1 U17121 ( .A1(n13659), .A2(n18941), .ZN(n13746) );
  XNOR2_X1 U17122 ( .A(n15307), .B(n13746), .ZN(n13757) );
  INV_X1 U17123 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13749) );
  AOI22_X1 U17124 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19012), .B1(
        n13747), .B2(n20703), .ZN(n13748) );
  OAI21_X1 U17125 ( .B1(n18999), .B2(n13749), .A(n13748), .ZN(n13750) );
  AOI211_X1 U17126 ( .C1(n18986), .C2(P2_REIP_REG_12__SCAN_IN), .A(n18985), 
        .B(n13750), .ZN(n13755) );
  AOI21_X1 U17127 ( .B1(n13751), .B2(n13753), .A(n13752), .ZN(n19076) );
  NAND2_X1 U17128 ( .A1(n19076), .A2(n19002), .ZN(n13754) );
  OAI211_X1 U17129 ( .C1(n15555), .C2(n20705), .A(n13755), .B(n13754), .ZN(
        n13756) );
  AOI21_X1 U17130 ( .B1(n13757), .B2(n19009), .A(n13756), .ZN(n13758) );
  INV_X1 U17131 ( .A(n13758), .ZN(P2_U2843) );
  INV_X1 U17132 ( .A(n13858), .ZN(n19024) );
  XNOR2_X1 U17133 ( .A(n19024), .B(n19023), .ZN(n13762) );
  OAI21_X1 U17134 ( .B1(n13549), .B2(n13760), .A(n13759), .ZN(n18918) );
  MUX2_X1 U17135 ( .A(n20871), .B(n18918), .S(n19048), .Z(n13761) );
  OAI21_X1 U17136 ( .B1(n13762), .B2(n19041), .A(n13761), .ZN(P2_U2874) );
  OAI21_X1 U17137 ( .B1(n13765), .B2(n13764), .A(n13763), .ZN(n16100) );
  INV_X1 U17138 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n13766) );
  NOR2_X1 U17139 ( .A1(n16209), .A2(n13766), .ZN(n13769) );
  OAI21_X1 U17140 ( .B1(n14158), .B2(n16172), .A(n20100), .ZN(n14884) );
  AOI21_X1 U17141 ( .B1(n16126), .B2(n13767), .A(n14884), .ZN(n16198) );
  AOI21_X1 U17142 ( .B1(n14155), .B2(n20108), .A(n20097), .ZN(n16158) );
  NOR2_X1 U17143 ( .A1(n20093), .A2(n16158), .ZN(n20080) );
  INV_X1 U17144 ( .A(n20080), .ZN(n20092) );
  NAND2_X1 U17145 ( .A1(n14161), .A2(n20890), .ZN(n16199) );
  OAI22_X1 U17146 ( .A1(n16198), .A2(n20890), .B1(n20092), .B2(n16199), .ZN(
        n13768) );
  AOI211_X1 U17147 ( .C1(n20098), .C2(n13770), .A(n13769), .B(n13768), .ZN(
        n13771) );
  OAI21_X1 U17148 ( .B1(n16186), .B2(n16100), .A(n13771), .ZN(P1_U3026) );
  INV_X1 U17149 ( .A(n13772), .ZN(n13774) );
  NAND2_X1 U17150 ( .A1(n13773), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16376) );
  INV_X1 U17151 ( .A(n16376), .ZN(n13839) );
  NOR2_X1 U17152 ( .A1(n10032), .A2(n13786), .ZN(n19010) );
  AOI21_X1 U17153 ( .B1(n10032), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19010), .ZN(n13838) );
  AOI222_X1 U17154 ( .A1(n13775), .A2(n13840), .B1(n13774), .B2(n13839), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n13838), .ZN(n13777) );
  NAND2_X1 U17155 ( .A1(n13843), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13776) );
  OAI21_X1 U17156 ( .B1(n13777), .B2(n13843), .A(n13776), .ZN(P2_U3601) );
  NAND2_X1 U17157 ( .A1(n13780), .A2(n13781), .ZN(n13782) );
  AND2_X1 U17158 ( .A1(n13779), .A2(n13782), .ZN(n19950) );
  INV_X1 U17159 ( .A(n19950), .ZN(n13796) );
  OAI21_X1 U17160 ( .B1(n16220), .B2(n13783), .A(n13895), .ZN(n19945) );
  OAI222_X1 U17161 ( .A1(n13796), .A2(n14635), .B1(n13784), .B2(n20023), .C1(
        n14629), .C2(n19945), .ZN(P1_U2865) );
  OAI211_X1 U17162 ( .C1(n13786), .C2(n13785), .A(n10012), .B(n20691), .ZN(
        n13836) );
  NAND2_X1 U17163 ( .A1(n19879), .A2(n19002), .ZN(n13790) );
  NAND2_X1 U17164 ( .A1(n19009), .A2(n10032), .ZN(n18947) );
  AOI22_X1 U17165 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19012), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n20694), .ZN(n13787) );
  OAI21_X1 U17166 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18947), .A(
        n13787), .ZN(n13788) );
  AOI21_X1 U17167 ( .B1(n18986), .B2(P2_REIP_REG_1__SCAN_IN), .A(n13788), .ZN(
        n13789) );
  OAI211_X1 U17168 ( .C1(n19005), .C2(n13791), .A(n13790), .B(n13789), .ZN(
        n13792) );
  AOI21_X1 U17169 ( .B1(n13793), .B2(n19007), .A(n13792), .ZN(n13795) );
  NAND2_X1 U17170 ( .A1(n19877), .A2(n20707), .ZN(n13794) );
  OAI211_X1 U17171 ( .C1(n13836), .C2(n12836), .A(n13795), .B(n13794), .ZN(
        P2_U2854) );
  OAI222_X1 U17172 ( .A1(n16009), .A2(n13796), .B1(n14674), .B2(n14705), .C1(
        n14695), .C2(n13419), .ZN(P1_U2897) );
  XNOR2_X1 U17173 ( .A(n9716), .B(n13798), .ZN(n13818) );
  NAND2_X1 U17174 ( .A1(n13800), .A2(n13799), .ZN(n13802) );
  XNOR2_X1 U17175 ( .A(n13802), .B(n13801), .ZN(n13815) );
  NAND2_X1 U17176 ( .A1(n13815), .A2(n15335), .ZN(n13808) );
  NOR2_X1 U17177 ( .A1(n19172), .A2(n13803), .ZN(n13806) );
  NAND2_X1 U17178 ( .A1(n18985), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13809) );
  OAI21_X1 U17179 ( .B1(n19184), .B2(n13804), .A(n13809), .ZN(n13805) );
  AOI211_X1 U17180 ( .C1(n13207), .C2(n19176), .A(n13806), .B(n13805), .ZN(
        n13807) );
  OAI211_X1 U17181 ( .C1(n13818), .C2(n19173), .A(n13808), .B(n13807), .ZN(
        P2_U3011) );
  OAI21_X1 U17182 ( .B1(n19861), .B2(n15355), .A(n13809), .ZN(n13814) );
  INV_X1 U17183 ( .A(n13810), .ZN(n13812) );
  INV_X1 U17184 ( .A(n14030), .ZN(n13811) );
  AOI21_X1 U17185 ( .B1(n13812), .B2(n10449), .A(n13811), .ZN(n13813) );
  AOI211_X1 U17186 ( .C1(n12862), .C2(n13207), .A(n13814), .B(n13813), .ZN(
        n13817) );
  NAND2_X1 U17187 ( .A1(n13815), .A2(n16359), .ZN(n13816) );
  OAI211_X1 U17188 ( .C1(n13818), .C2(n15629), .A(n13817), .B(n13816), .ZN(
        P2_U3043) );
  AND2_X1 U17189 ( .A1(n13819), .A2(n13820), .ZN(n13822) );
  OR2_X1 U17190 ( .A1(n13822), .A2(n13821), .ZN(n19073) );
  NAND2_X1 U17191 ( .A1(n13759), .A2(n13824), .ZN(n13825) );
  NAND2_X1 U17192 ( .A1(n13823), .A2(n13825), .ZN(n19030) );
  INV_X1 U17193 ( .A(n19030), .ZN(n13834) );
  AND3_X1 U17194 ( .A1(n19009), .A2(n10012), .A3(n13826), .ZN(n18927) );
  AOI211_X1 U17195 ( .C1(n10012), .C2(n13826), .A(n12836), .B(n13830), .ZN(
        n13829) );
  AOI22_X1 U17196 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19012), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n20694), .ZN(n13827) );
  OAI211_X1 U17197 ( .C1(n19815), .C2(n20697), .A(n13827), .B(n18933), .ZN(
        n13828) );
  AOI211_X1 U17198 ( .C1(n13830), .C2(n18927), .A(n13829), .B(n13828), .ZN(
        n13831) );
  OAI21_X1 U17199 ( .B1(n13832), .B2(n19005), .A(n13831), .ZN(n13833) );
  AOI21_X1 U17200 ( .B1(n13834), .B2(n19007), .A(n13833), .ZN(n13835) );
  OAI21_X1 U17201 ( .B1(n19073), .B2(n20698), .A(n13835), .ZN(P2_U2841) );
  OAI21_X1 U17202 ( .B1(n10012), .B2(n10256), .A(n13836), .ZN(n15637) );
  NOR2_X1 U17203 ( .A1(n13838), .A2(n13837), .ZN(n15635) );
  AOI222_X1 U17204 ( .A1(n13841), .A2(n13840), .B1(n15637), .B2(n15635), .C1(
        n20708), .C2(n13839), .ZN(n13844) );
  NAND2_X1 U17205 ( .A1(n13843), .A2(n14352), .ZN(n13842) );
  OAI21_X1 U17206 ( .B1(n13844), .B2(n13843), .A(n13842), .ZN(P2_U3599) );
  XOR2_X1 U17207 ( .A(n9820), .B(n13845), .Z(n20018) );
  INV_X1 U17208 ( .A(n20018), .ZN(n13847) );
  OAI222_X1 U17209 ( .A1(n16009), .A2(n13847), .B1(n13846), .B2(n14695), .C1(
        n14705), .C2(n14680), .ZN(P1_U2898) );
  AOI22_X1 U17210 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13851) );
  AOI22_X1 U17211 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17212 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13849) );
  AOI22_X1 U17213 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13848) );
  NAND4_X1 U17214 ( .A1(n13851), .A2(n13850), .A3(n13849), .A4(n13848), .ZN(
        n13857) );
  AOI22_X1 U17215 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U17216 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13854) );
  INV_X1 U17217 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n20986) );
  AOI22_X1 U17218 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U17219 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13852) );
  NAND4_X1 U17220 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  NOR2_X1 U17221 ( .A1(n13857), .A2(n13856), .ZN(n13872) );
  NAND2_X1 U17222 ( .A1(n19024), .A2(n10123), .ZN(n13941) );
  AOI22_X1 U17223 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U17224 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13861) );
  AOI22_X1 U17225 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13860) );
  AOI22_X1 U17226 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13859) );
  NAND4_X1 U17227 ( .A1(n13862), .A2(n13861), .A3(n13860), .A4(n13859), .ZN(
        n13868) );
  AOI22_X1 U17228 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U17229 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17230 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17231 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13863) );
  NAND4_X1 U17232 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n13863), .ZN(
        n13867) );
  OR2_X1 U17233 ( .A1(n13868), .A2(n13867), .ZN(n19016) );
  INV_X1 U17234 ( .A(n16292), .ZN(n13871) );
  AOI21_X1 U17235 ( .B1(n13872), .B2(n13869), .A(n13871), .ZN(n14018) );
  NAND2_X1 U17236 ( .A1(n14018), .A2(n19106), .ZN(n13879) );
  INV_X1 U17237 ( .A(n19059), .ZN(n15115) );
  OAI22_X1 U17238 ( .A1(n15115), .A2(n19129), .B1(n13873), .B2(n19095), .ZN(
        n13877) );
  INV_X1 U17239 ( .A(n19060), .ZN(n15119) );
  INV_X1 U17240 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13875) );
  NOR2_X1 U17241 ( .A1(n15119), .A2(n13875), .ZN(n13876) );
  AOI211_X1 U17242 ( .C1(n19061), .C2(BUF1_REG_17__SCAN_IN), .A(n13877), .B(
        n13876), .ZN(n13878) );
  OAI211_X1 U17243 ( .C1(n18905), .C2(n19063), .A(n13879), .B(n13878), .ZN(
        P2_U2902) );
  OAI21_X1 U17244 ( .B1(n9713), .B2(n14006), .A(n9715), .ZN(n13882) );
  INV_X1 U17245 ( .A(n13882), .ZN(n13937) );
  XOR2_X1 U17246 ( .A(n9719), .B(n13884), .Z(n13935) );
  INV_X1 U17247 ( .A(n14028), .ZN(n16362) );
  NAND2_X1 U17248 ( .A1(n16362), .A2(n14006), .ZN(n13889) );
  AOI22_X1 U17249 ( .A1(n16354), .A2(n19103), .B1(n18985), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n13888) );
  NAND3_X1 U17250 ( .A1(n14030), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        n15599), .ZN(n13887) );
  NAND2_X1 U17251 ( .A1(n13885), .A2(n12862), .ZN(n13886) );
  NAND4_X1 U17252 ( .A1(n13889), .A2(n13888), .A3(n13887), .A4(n13886), .ZN(
        n13890) );
  AOI21_X1 U17253 ( .B1(n13935), .B2(n16359), .A(n13890), .ZN(n13891) );
  OAI21_X1 U17254 ( .B1(n13937), .B2(n15629), .A(n13891), .ZN(P2_U3042) );
  AOI21_X1 U17255 ( .B1(n13893), .B2(n13779), .A(n13892), .ZN(n19939) );
  NAND2_X1 U17256 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  NAND2_X1 U17257 ( .A1(n14108), .A2(n13896), .ZN(n19936) );
  OAI22_X1 U17258 ( .A1(n19936), .A2(n14629), .B1(n13897), .B2(n20023), .ZN(
        n13898) );
  AOI21_X1 U17259 ( .B1(n19939), .B2(n12893), .A(n13898), .ZN(n13899) );
  INV_X1 U17260 ( .A(n13899), .ZN(P1_U2864) );
  NAND2_X1 U17261 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16236), .ZN(n13902) );
  OAI221_X1 U17262 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20439), .C1(n16236), 
        .C2(P1_STATE2_REG_3__SCAN_IN), .A(n20680), .ZN(n13900) );
  OAI21_X1 U17263 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13903) );
  INV_X1 U17264 ( .A(n13912), .ZN(n13905) );
  NAND2_X1 U17265 ( .A1(n13905), .A2(n13904), .ZN(n13907) );
  NOR2_X1 U17266 ( .A1(n13916), .A2(n16233), .ZN(n13906) );
  NOR2_X1 U17267 ( .A1(n13912), .A2(n13908), .ZN(n20007) );
  INV_X1 U17268 ( .A(n20086), .ZN(n13927) );
  NAND2_X1 U17269 ( .A1(n20603), .A2(n20321), .ZN(n15793) );
  NAND3_X1 U17270 ( .A1(n13909), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n15793), 
        .ZN(n13910) );
  NOR2_X2 U17271 ( .A1(n13912), .A2(n13910), .ZN(n19993) );
  NOR2_X1 U17272 ( .A1(n13913), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13918) );
  AND2_X1 U17273 ( .A1(n11022), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13914) );
  NOR2_X1 U17274 ( .A1(n13918), .A2(n13914), .ZN(n13915) );
  NAND2_X1 U17275 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13922) );
  OAI221_X1 U17276 ( .B1(n19980), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19980), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20009), .ZN(n13920) );
  NAND2_X1 U17277 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n13920), .ZN(n13921) );
  OAI211_X1 U17278 ( .C1(n19991), .C2(n13923), .A(n13922), .B(n13921), .ZN(
        n13924) );
  AOI21_X1 U17279 ( .B1(n20006), .B2(P1_EBX_REG_3__SCAN_IN), .A(n13924), .ZN(
        n13926) );
  INV_X1 U17280 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20614) );
  NAND4_X1 U17281 ( .A1(n20005), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n20614), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n13925) );
  OAI211_X1 U17282 ( .C1(n13927), .C2(n20010), .A(n13926), .B(n13925), .ZN(
        n13928) );
  AOI21_X1 U17283 ( .B1(n20125), .B2(n20007), .A(n13928), .ZN(n13929) );
  OAI21_X1 U17284 ( .B1(n13930), .B2(n20017), .A(n13929), .ZN(P1_U2837) );
  OAI22_X1 U17285 ( .A1(n19184), .A2(n20984), .B1(n12251), .B2(n18970), .ZN(
        n13931) );
  AOI21_X1 U17286 ( .B1(n16343), .B2(n13932), .A(n13931), .ZN(n13933) );
  OAI21_X1 U17287 ( .B1(n19051), .B2(n15652), .A(n13933), .ZN(n13934) );
  AOI21_X1 U17288 ( .B1(n13935), .B2(n16346), .A(n13934), .ZN(n13936) );
  OAI21_X1 U17289 ( .B1(n13937), .B2(n19173), .A(n13936), .ZN(P2_U3010) );
  INV_X1 U17290 ( .A(n19939), .ZN(n14119) );
  OAI222_X1 U17291 ( .A1(n14119), .A2(n16009), .B1(n13938), .B2(n14695), .C1(
        n14668), .C2(n14705), .ZN(P1_U2896) );
  NAND2_X1 U17292 ( .A1(n13823), .A2(n13939), .ZN(n13940) );
  NAND2_X1 U17293 ( .A1(n14137), .A2(n13940), .ZN(n18912) );
  INV_X1 U17294 ( .A(n18912), .ZN(n13946) );
  NOR2_X1 U17295 ( .A1(n19048), .A2(n18917), .ZN(n13945) );
  AOI211_X1 U17296 ( .C1(n13943), .C2(n19025), .A(n19041), .B(n13942), .ZN(
        n13944) );
  AOI211_X1 U17297 ( .C1(n13946), .C2(n19048), .A(n13945), .B(n13944), .ZN(
        n13947) );
  INV_X1 U17298 ( .A(n13947), .ZN(P2_U2872) );
  AND2_X1 U17299 ( .A1(n20125), .A2(n13519), .ZN(n20352) );
  INV_X1 U17300 ( .A(n20352), .ZN(n20393) );
  INV_X1 U17301 ( .A(n20436), .ZN(n20488) );
  NOR2_X1 U17302 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n11318), .ZN(
        n20392) );
  INV_X1 U17303 ( .A(n20392), .ZN(n13949) );
  NOR2_X1 U17304 ( .A1(n13949), .A2(n20431), .ZN(n13988) );
  INV_X1 U17305 ( .A(n13988), .ZN(n13950) );
  OAI21_X1 U17306 ( .B1(n20393), .B2(n20488), .A(n13950), .ZN(n13954) );
  OR2_X1 U17307 ( .A1(n13952), .A2(n20525), .ZN(n20359) );
  INV_X1 U17308 ( .A(n20359), .ZN(n14045) );
  INV_X1 U17309 ( .A(n20127), .ZN(n13951) );
  INV_X1 U17310 ( .A(n20353), .ZN(n20126) );
  NOR2_X1 U17311 ( .A1(n13951), .A2(n20126), .ZN(n20437) );
  AOI22_X1 U17312 ( .A1(n13954), .A2(n20538), .B1(n14045), .B2(n20437), .ZN(
        n13993) );
  NAND2_X1 U17313 ( .A1(n13952), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20490) );
  NAND2_X1 U17314 ( .A1(n13953), .A2(n20490), .ZN(n20187) );
  AOI21_X1 U17315 ( .B1(n13989), .B2(n20342), .A(n20321), .ZN(n13955) );
  OR2_X1 U17316 ( .A1(n13955), .A2(n13954), .ZN(n13956) );
  AOI22_X1 U17317 ( .A1(n20550), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n13987), .ZN(n13959) );
  INV_X1 U17318 ( .A(n20555), .ZN(n20411) );
  NOR2_X1 U17319 ( .A1(n13989), .A2(n20456), .ZN(n13957) );
  AOI21_X1 U17320 ( .B1(n20345), .B2(n20411), .A(n13957), .ZN(n13958) );
  OAI211_X1 U17321 ( .C1(n14054), .C2(n13993), .A(n13959), .B(n13958), .ZN(
        P1_U3099) );
  AOI22_X1 U17322 ( .A1(n20556), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n13987), .ZN(n13962) );
  INV_X1 U17323 ( .A(n20560), .ZN(n20414) );
  NOR2_X1 U17324 ( .A1(n13989), .A2(n9856), .ZN(n13960) );
  AOI21_X1 U17325 ( .B1(n20345), .B2(n20414), .A(n13960), .ZN(n13961) );
  OAI211_X1 U17326 ( .C1(n14062), .C2(n13993), .A(n13962), .B(n13961), .ZN(
        P1_U3100) );
  AOI22_X1 U17327 ( .A1(n20545), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n13987), .ZN(n13965) );
  INV_X1 U17328 ( .A(n20549), .ZN(n20408) );
  NOR2_X1 U17329 ( .A1(n13989), .A2(n9858), .ZN(n13963) );
  AOI21_X1 U17330 ( .B1(n20345), .B2(n20408), .A(n13963), .ZN(n13964) );
  OAI211_X1 U17331 ( .C1(n14058), .C2(n13993), .A(n13965), .B(n13964), .ZN(
        P1_U3098) );
  AOI22_X1 U17332 ( .A1(n20567), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__5__SCAN_IN), .B2(n13987), .ZN(n13968) );
  INV_X1 U17333 ( .A(n20571), .ZN(n20336) );
  NOR2_X1 U17334 ( .A1(n13989), .A2(n9854), .ZN(n13966) );
  AOI21_X1 U17335 ( .B1(n20345), .B2(n20336), .A(n13966), .ZN(n13967) );
  OAI211_X1 U17336 ( .C1(n14074), .C2(n13993), .A(n13968), .B(n13967), .ZN(
        P1_U3102) );
  AOI22_X1 U17337 ( .A1(n20527), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__0__SCAN_IN), .B2(n13987), .ZN(n13971) );
  INV_X1 U17338 ( .A(n20500), .ZN(n20539) );
  NOR2_X1 U17339 ( .A1(n13989), .A2(n20544), .ZN(n13969) );
  AOI21_X1 U17340 ( .B1(n20345), .B2(n20539), .A(n13969), .ZN(n13970) );
  OAI211_X1 U17341 ( .C1(n14070), .C2(n13993), .A(n13971), .B(n13970), .ZN(
        P1_U3097) );
  AOI22_X1 U17342 ( .A1(n20579), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n13987), .ZN(n13974) );
  NOR2_X1 U17343 ( .A1(n13989), .A2(n20486), .ZN(n13972) );
  AOI21_X1 U17344 ( .B1(n20345), .B2(n9849), .A(n13972), .ZN(n13973) );
  OAI211_X1 U17345 ( .C1(n14078), .C2(n13993), .A(n13974), .B(n13973), .ZN(
        P1_U3104) );
  AOI22_X1 U17346 ( .A1(n20561), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n13987), .ZN(n13977) );
  INV_X1 U17347 ( .A(n20566), .ZN(n20303) );
  NOR2_X1 U17348 ( .A1(n13989), .A2(n20466), .ZN(n13975) );
  AOI21_X1 U17349 ( .B1(n20345), .B2(n20303), .A(n13975), .ZN(n13976) );
  OAI211_X1 U17350 ( .C1(n14066), .C2(n13993), .A(n13977), .B(n13976), .ZN(
        P1_U3101) );
  NAND2_X1 U17351 ( .A1(n19980), .A2(n20009), .ZN(n19949) );
  NAND2_X1 U17352 ( .A1(n19949), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13982) );
  INV_X1 U17353 ( .A(n13978), .ZN(n14894) );
  NAND2_X1 U17354 ( .A1(n19996), .A2(n19991), .ZN(n13979) );
  AOI22_X1 U17355 ( .A1(n19993), .A2(n14894), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13979), .ZN(n13981) );
  NAND2_X1 U17356 ( .A1(n20006), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13980) );
  NAND3_X1 U17357 ( .A1(n13982), .A2(n13981), .A3(n13980), .ZN(n13985) );
  NOR2_X1 U17358 ( .A1(n13983), .A2(n20017), .ZN(n13984) );
  AOI211_X1 U17359 ( .C1(n20007), .C2(n11624), .A(n13985), .B(n13984), .ZN(
        n13986) );
  INV_X1 U17360 ( .A(n13986), .ZN(P1_U2840) );
  AOI22_X1 U17361 ( .A1(n20572), .A2(n13988), .B1(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n13987), .ZN(n13992) );
  NOR2_X1 U17362 ( .A1(n13989), .A2(n20476), .ZN(n13990) );
  AOI21_X1 U17363 ( .B1(n20345), .B2(n9851), .A(n13990), .ZN(n13991) );
  OAI211_X1 U17364 ( .C1(n14093), .C2(n13993), .A(n13992), .B(n13991), .ZN(
        P1_U3103) );
  INV_X1 U17365 ( .A(n13995), .ZN(n13997) );
  NOR2_X1 U17366 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  XOR2_X1 U17367 ( .A(n13994), .B(n13998), .Z(n14017) );
  XOR2_X1 U17368 ( .A(n13999), .B(n14001), .Z(n14015) );
  INV_X1 U17369 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18982) );
  OAI22_X1 U17370 ( .A1(n19184), .A2(n18982), .B1(n19172), .B2(n18990), .ZN(
        n14002) );
  AOI21_X1 U17371 ( .B1(n18985), .B2(P2_REIP_REG_5__SCAN_IN), .A(n14002), .ZN(
        n14003) );
  OAI21_X1 U17372 ( .B1(n15652), .B2(n18991), .A(n14003), .ZN(n14004) );
  AOI21_X1 U17373 ( .B1(n14015), .B2(n16346), .A(n14004), .ZN(n14005) );
  OAI21_X1 U17374 ( .B1(n19173), .B2(n14017), .A(n14005), .ZN(P2_U3009) );
  INV_X1 U17375 ( .A(n14031), .ZN(n15616) );
  AOI211_X1 U17376 ( .C1(n9891), .C2(n14006), .A(n15616), .B(n14028), .ZN(
        n14014) );
  OAI21_X1 U17377 ( .B1(n9840), .B2(n14008), .A(n14007), .ZN(n19101) );
  INV_X1 U17378 ( .A(n18991), .ZN(n14011) );
  NAND3_X1 U17379 ( .A1(n14030), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n15599), .ZN(n14009) );
  OAI21_X1 U17380 ( .B1(n10731), .B2(n18933), .A(n14009), .ZN(n14010) );
  AOI21_X1 U17381 ( .B1(n12862), .B2(n14011), .A(n14010), .ZN(n14012) );
  OAI21_X1 U17382 ( .B1(n19101), .B2(n15355), .A(n14012), .ZN(n14013) );
  AOI211_X1 U17383 ( .C1(n14015), .C2(n16359), .A(n14014), .B(n14013), .ZN(
        n14016) );
  OAI21_X1 U17384 ( .B1(n15629), .B2(n14017), .A(n14016), .ZN(P2_U3041) );
  NAND2_X1 U17385 ( .A1(n14018), .A2(n19018), .ZN(n14020) );
  NAND2_X1 U17386 ( .A1(n19052), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14019) );
  OAI211_X1 U17387 ( .C1(n15253), .C2(n19052), .A(n14020), .B(n14019), .ZN(
        P2_U2870) );
  OAI21_X1 U17388 ( .B1(n14022), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14021), .ZN(n16344) );
  INV_X1 U17389 ( .A(n14023), .ZN(n14025) );
  NAND3_X1 U17390 ( .A1(n14007), .A2(n14025), .A3(n14024), .ZN(n14026) );
  NAND2_X1 U17391 ( .A1(n14027), .A2(n14026), .ZN(n19093) );
  OAI22_X1 U17392 ( .A1(n19093), .A2(n15355), .B1(n10734), .B2(n18933), .ZN(
        n14035) );
  NOR3_X1 U17393 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14028), .A3(
        n14031), .ZN(n14029) );
  INV_X1 U17394 ( .A(n14029), .ZN(n14032) );
  AOI221_X1 U17395 ( .B1(n14031), .B2(n15599), .C1(n14030), .C2(n15599), .A(
        n14029), .ZN(n16352) );
  AOI21_X1 U17396 ( .B1(n14033), .B2(n14032), .A(n16352), .ZN(n14034) );
  AOI211_X1 U17397 ( .C1(n18977), .C2(n12862), .A(n14035), .B(n14034), .ZN(
        n14040) );
  INV_X1 U17398 ( .A(n9722), .ZN(n14037) );
  XNOR2_X1 U17399 ( .A(n14038), .B(n14037), .ZN(n16345) );
  NAND2_X1 U17400 ( .A1(n16345), .A2(n16359), .ZN(n14039) );
  OAI211_X1 U17401 ( .C1(n16344), .C2(n15629), .A(n14040), .B(n14039), .ZN(
        P2_U3040) );
  NAND3_X1 U17402 ( .A1(n14043), .A2(n14089), .A3(n20538), .ZN(n14041) );
  NAND2_X1 U17403 ( .A1(n14041), .A2(n20434), .ZN(n14049) );
  AND2_X1 U17404 ( .A1(n20289), .A2(n20488), .ZN(n14047) );
  INV_X1 U17405 ( .A(n20490), .ZN(n14042) );
  NOR2_X1 U17406 ( .A1(n20353), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20191) );
  INV_X1 U17407 ( .A(n20456), .ZN(n20552) );
  NOR2_X1 U17408 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14044), .ZN(
        n14087) );
  INV_X1 U17409 ( .A(n14047), .ZN(n14048) );
  NOR2_X1 U17410 ( .A1(n20191), .A2(n20525), .ZN(n20188) );
  AOI21_X1 U17411 ( .B1(n14049), .B2(n14048), .A(n20188), .ZN(n14050) );
  OAI211_X1 U17412 ( .C1(n14087), .C2(n20439), .A(n20494), .B(n14050), .ZN(
        n14086) );
  AOI22_X1 U17413 ( .A1(n20550), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n14086), .ZN(n14051) );
  OAI21_X1 U17414 ( .B1(n14089), .B2(n20555), .A(n14051), .ZN(n14052) );
  AOI21_X1 U17415 ( .B1(n20312), .B2(n20552), .A(n14052), .ZN(n14053) );
  OAI21_X1 U17416 ( .B1(n14054), .B2(n14092), .A(n14053), .ZN(P1_U3083) );
  AOI22_X1 U17417 ( .A1(n20545), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n14086), .ZN(n14055) );
  OAI21_X1 U17418 ( .B1(n14089), .B2(n20549), .A(n14055), .ZN(n14056) );
  AOI21_X1 U17419 ( .B1(n20312), .B2(n9857), .A(n14056), .ZN(n14057) );
  OAI21_X1 U17420 ( .B1(n14058), .B2(n14092), .A(n14057), .ZN(P1_U3082) );
  AOI22_X1 U17421 ( .A1(n20556), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n14086), .ZN(n14059) );
  OAI21_X1 U17422 ( .B1(n14089), .B2(n20560), .A(n14059), .ZN(n14060) );
  AOI21_X1 U17423 ( .B1(n20312), .B2(n9855), .A(n14060), .ZN(n14061) );
  OAI21_X1 U17424 ( .B1(n14062), .B2(n14092), .A(n14061), .ZN(P1_U3084) );
  INV_X1 U17425 ( .A(n20466), .ZN(n20563) );
  AOI22_X1 U17426 ( .A1(n20561), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n14086), .ZN(n14063) );
  OAI21_X1 U17427 ( .B1(n14089), .B2(n20566), .A(n14063), .ZN(n14064) );
  AOI21_X1 U17428 ( .B1(n20312), .B2(n20563), .A(n14064), .ZN(n14065) );
  OAI21_X1 U17429 ( .B1(n14066), .B2(n14092), .A(n14065), .ZN(P1_U3085) );
  INV_X1 U17430 ( .A(n20544), .ZN(n20497) );
  AOI22_X1 U17431 ( .A1(n20527), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n14086), .ZN(n14067) );
  OAI21_X1 U17432 ( .B1(n14089), .B2(n20500), .A(n14067), .ZN(n14068) );
  AOI21_X1 U17433 ( .B1(n20312), .B2(n20497), .A(n14068), .ZN(n14069) );
  OAI21_X1 U17434 ( .B1(n14070), .B2(n14092), .A(n14069), .ZN(P1_U3081) );
  AOI22_X1 U17435 ( .A1(n20567), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n14086), .ZN(n14071) );
  OAI21_X1 U17436 ( .B1(n14089), .B2(n20571), .A(n14071), .ZN(n14072) );
  AOI21_X1 U17437 ( .B1(n20312), .B2(n9853), .A(n14072), .ZN(n14073) );
  OAI21_X1 U17438 ( .B1(n14074), .B2(n14092), .A(n14073), .ZN(P1_U3086) );
  INV_X1 U17439 ( .A(n20486), .ZN(n20582) );
  AOI22_X1 U17440 ( .A1(n20579), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n14086), .ZN(n14075) );
  OAI21_X1 U17441 ( .B1(n14089), .B2(n9850), .A(n14075), .ZN(n14076) );
  AOI21_X1 U17442 ( .B1(n20312), .B2(n20582), .A(n14076), .ZN(n14077) );
  OAI21_X1 U17443 ( .B1(n14078), .B2(n14092), .A(n14077), .ZN(P1_U3088) );
  OAI21_X1 U17444 ( .B1(n14079), .B2(n14082), .A(n14081), .ZN(n14817) );
  INV_X1 U17445 ( .A(n14109), .ZN(n14083) );
  AOI21_X1 U17446 ( .B1(n14084), .B2(n14083), .A(n14209), .ZN(n16189) );
  AOI22_X1 U17447 ( .A1(n16189), .A2(n20021), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14642), .ZN(n14085) );
  OAI21_X1 U17448 ( .B1(n14817), .B2(n14635), .A(n14085), .ZN(P1_U2862) );
  INV_X1 U17449 ( .A(n20476), .ZN(n20574) );
  AOI22_X1 U17450 ( .A1(n20572), .A2(n14087), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n14086), .ZN(n14088) );
  OAI21_X1 U17451 ( .B1(n14089), .B2(n9852), .A(n14088), .ZN(n14090) );
  AOI21_X1 U17452 ( .B1(n20312), .B2(n20574), .A(n14090), .ZN(n14091) );
  OAI21_X1 U17453 ( .B1(n14093), .B2(n14092), .A(n14091), .ZN(P1_U3087) );
  INV_X1 U17454 ( .A(n14813), .ZN(n14102) );
  AOI22_X1 U17455 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n20006), .B1(n19993), 
        .B2(n16189), .ZN(n14095) );
  NAND2_X1 U17456 ( .A1(n14094), .A2(n20009), .ZN(n19982) );
  OAI211_X1 U17457 ( .C1(n19996), .C2(n14096), .A(n14095), .B(n19982), .ZN(
        n14101) );
  INV_X1 U17458 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20624) );
  INV_X1 U17459 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20622) );
  NAND3_X1 U17460 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n19933) );
  NOR2_X1 U17461 ( .A1(n20622), .A2(n19933), .ZN(n14097) );
  INV_X1 U17462 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20615) );
  NAND3_X1 U17463 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19979) );
  NOR2_X1 U17464 ( .A1(n20615), .A2(n19979), .ZN(n14098) );
  NAND2_X1 U17465 ( .A1(n20005), .A2(n14098), .ZN(n19932) );
  NAND2_X1 U17466 ( .A1(n14097), .A2(n19964), .ZN(n19924) );
  NOR2_X1 U17467 ( .A1(n20624), .A2(n19924), .ZN(n14099) );
  NAND4_X1 U17468 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n14098), .A4(n14097), .ZN(n14518) );
  INV_X1 U17469 ( .A(n20009), .ZN(n19992) );
  AOI21_X1 U17470 ( .B1(n14518), .B2(n20005), .A(n19992), .ZN(n14173) );
  INV_X1 U17471 ( .A(n14173), .ZN(n15993) );
  MUX2_X1 U17472 ( .A(n14099), .B(n15993), .S(P1_REIP_REG_10__SCAN_IN), .Z(
        n14100) );
  AOI211_X1 U17473 ( .C1(n20013), .C2(n14102), .A(n14101), .B(n14100), .ZN(
        n14103) );
  OAI21_X1 U17474 ( .B1(n15977), .B2(n14817), .A(n14103), .ZN(P1_U2830) );
  INV_X1 U17475 ( .A(n14079), .ZN(n14104) );
  OAI21_X1 U17476 ( .B1(n13892), .B2(n14105), .A(n14104), .ZN(n19927) );
  OAI222_X1 U17477 ( .A1(n19927), .A2(n16009), .B1(n14664), .B2(n14705), .C1(
        n14106), .C2(n14695), .ZN(P1_U2895) );
  AND2_X1 U17478 ( .A1(n14108), .A2(n14107), .ZN(n14110) );
  OR2_X1 U17479 ( .A1(n14110), .A2(n14109), .ZN(n19923) );
  OAI222_X1 U17480 ( .A1(n19927), .A2(n14635), .B1(n14111), .B2(n20023), .C1(
        n14629), .C2(n19923), .ZN(P1_U2863) );
  XNOR2_X1 U17481 ( .A(n14114), .B(n14113), .ZN(n14115) );
  XNOR2_X1 U17482 ( .A(n14112), .B(n14115), .ZN(n16206) );
  NAND2_X1 U17483 ( .A1(n16206), .A2(n20071), .ZN(n14118) );
  NOR2_X1 U17484 ( .A1(n16209), .A2(n20622), .ZN(n16202) );
  NOR2_X1 U17485 ( .A1(n14803), .A2(n20950), .ZN(n14116) );
  AOI211_X1 U17486 ( .C1(n20070), .C2(n19942), .A(n16202), .B(n14116), .ZN(
        n14117) );
  OAI211_X1 U17487 ( .C1(n20076), .C2(n14119), .A(n14118), .B(n14117), .ZN(
        P1_U2991) );
  NAND2_X1 U17488 ( .A1(n9819), .A2(n14120), .ZN(n14121) );
  NAND2_X1 U17489 ( .A1(n15050), .A2(n14121), .ZN(n16296) );
  INV_X1 U17490 ( .A(n15113), .ZN(n14122) );
  AOI21_X1 U17491 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n16311) );
  NAND2_X1 U17492 ( .A1(n16311), .A2(n19002), .ZN(n14131) );
  AOI211_X1 U17493 ( .C1(n15248), .C2(n18900), .A(n14125), .B(n12836), .ZN(
        n14129) );
  AOI22_X1 U17494 ( .A1(n14126), .A2(n20703), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19012), .ZN(n14127) );
  OAI211_X1 U17495 ( .C1(n15245), .C2(n20697), .A(n14127), .B(n18933), .ZN(
        n14128) );
  AOI211_X1 U17496 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n20694), .A(n14129), .B(
        n14128), .ZN(n14130) );
  OAI211_X1 U17497 ( .C1(n16296), .C2(n20705), .A(n14131), .B(n14130), .ZN(
        P2_U2837) );
  NOR2_X1 U17498 ( .A1(n14132), .A2(n14133), .ZN(n14134) );
  OR2_X1 U17499 ( .A1(n14135), .A2(n14134), .ZN(n19064) );
  AND2_X1 U17500 ( .A1(n14137), .A2(n14136), .ZN(n14139) );
  OR2_X1 U17501 ( .A1(n14139), .A2(n14138), .ZN(n19021) );
  INV_X1 U17502 ( .A(n19021), .ZN(n15267) );
  NOR2_X1 U17503 ( .A1(n14140), .A2(n19005), .ZN(n14144) );
  AOI22_X1 U17504 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n20694), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19012), .ZN(n14141) );
  OAI211_X1 U17505 ( .C1(n20697), .C2(n14142), .A(n14141), .B(n18933), .ZN(
        n14143) );
  AOI211_X1 U17506 ( .C1(n15267), .C2(n19007), .A(n14144), .B(n14143), .ZN(
        n14150) );
  NAND2_X1 U17507 ( .A1(n10012), .A2(n14145), .ZN(n14146) );
  XNOR2_X1 U17508 ( .A(n14147), .B(n14146), .ZN(n14148) );
  NAND2_X1 U17509 ( .A1(n14148), .A2(n19009), .ZN(n14149) );
  OAI211_X1 U17510 ( .C1(n19064), .C2(n20698), .A(n14150), .B(n14149), .ZN(
        P2_U2839) );
  OAI222_X1 U17511 ( .A1(n14817), .A2(n16009), .B1(n14695), .B2(n13406), .C1(
        n14659), .C2(n14705), .ZN(P1_U2894) );
  XNOR2_X1 U17512 ( .A(n9750), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14151) );
  XNOR2_X1 U17513 ( .A(n14152), .B(n14151), .ZN(n14167) );
  AOI21_X1 U17514 ( .B1(n20097), .B2(n20093), .A(n14153), .ZN(n14154) );
  OAI21_X1 U17515 ( .B1(n20101), .B2(n14155), .A(n14154), .ZN(n20089) );
  NOR2_X1 U17516 ( .A1(n14156), .A2(n20089), .ZN(n14159) );
  AOI21_X1 U17517 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n16191) );
  OAI22_X1 U17518 ( .A1(n19923), .A2(n16210), .B1(n20624), .B2(n16209), .ZN(
        n14160) );
  AOI21_X1 U17519 ( .B1(n16191), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14160), .ZN(n14163) );
  NAND2_X1 U17520 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16204) );
  NAND3_X1 U17521 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14161), .A3(
        n20080), .ZN(n16225) );
  NOR3_X1 U17522 ( .A1(n16094), .A2(n16204), .A3(n16225), .ZN(n16192) );
  NAND2_X1 U17523 ( .A1(n16192), .A2(n16193), .ZN(n14162) );
  OAI211_X1 U17524 ( .C1(n14167), .C2(n16186), .A(n14163), .B(n14162), .ZN(
        P1_U3022) );
  OAI22_X1 U17525 ( .A1(n14803), .A2(n19922), .B1(n16209), .B2(n20624), .ZN(
        n14165) );
  NOR2_X1 U17526 ( .A1(n19927), .A2(n20076), .ZN(n14164) );
  AOI211_X1 U17527 ( .C1(n20070), .C2(n19928), .A(n14165), .B(n14164), .ZN(
        n14166) );
  OAI21_X1 U17528 ( .B1(n14167), .B2(n19906), .A(n14166), .ZN(P1_U2990) );
  NAND2_X1 U17529 ( .A1(n14168), .A2(n14169), .ZN(n14183) );
  NAND2_X1 U17530 ( .A1(n14168), .A2(n14170), .ZN(n14638) );
  NAND2_X1 U17531 ( .A1(n14638), .A2(n14171), .ZN(n14172) );
  NAND2_X1 U17532 ( .A1(n14183), .A2(n14172), .ZN(n14795) );
  NAND4_X1 U17533 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14198) );
  INV_X1 U17534 ( .A(n14198), .ZN(n14517) );
  OAI21_X1 U17535 ( .B1(n14517), .B2(n19980), .A(n14173), .ZN(n15969) );
  INV_X1 U17536 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20629) );
  NOR2_X1 U17537 ( .A1(n19980), .A2(n14518), .ZN(n15992) );
  NAND3_X1 U17538 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15992), .ZN(n15976) );
  INV_X1 U17539 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20630) );
  OAI21_X1 U17540 ( .B1(n20629), .B2(n15976), .A(n20630), .ZN(n14179) );
  NOR2_X1 U17541 ( .A1(n14791), .A2(n19991), .ZN(n14178) );
  INV_X1 U17542 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14188) );
  INV_X1 U17543 ( .A(n14641), .ZN(n15983) );
  AOI21_X1 U17544 ( .B1(n15983), .B2(n14640), .A(n14174), .ZN(n14175) );
  NOR2_X1 U17545 ( .A1(n14175), .A2(n14186), .ZN(n16157) );
  AOI22_X1 U17546 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20014), .B1(
        n19993), .B2(n16157), .ZN(n14176) );
  OAI211_X1 U17547 ( .C1(n19984), .C2(n14188), .A(n19982), .B(n14176), .ZN(
        n14177) );
  AOI211_X1 U17548 ( .C1(n15969), .C2(n14179), .A(n14178), .B(n14177), .ZN(
        n14180) );
  OAI21_X1 U17549 ( .B1(n14795), .B2(n15977), .A(n14180), .ZN(P1_U2826) );
  INV_X1 U17550 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14181) );
  OAI222_X1 U17551 ( .A1(n14795), .A2(n16009), .B1(n14644), .B2(n14705), .C1(
        n14181), .C2(n14695), .ZN(P1_U2890) );
  AOI21_X1 U17552 ( .B1(n14184), .B2(n14183), .A(n14182), .ZN(n16072) );
  INV_X1 U17553 ( .A(n16072), .ZN(n14697) );
  OAI21_X1 U17554 ( .B1(n14186), .B2(n14185), .A(n14194), .ZN(n16150) );
  INV_X1 U17555 ( .A(n16150), .ZN(n15964) );
  AOI22_X1 U17556 ( .A1(n15964), .A2(n20021), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14642), .ZN(n14187) );
  OAI21_X1 U17557 ( .B1(n14697), .B2(n14635), .A(n14187), .ZN(P1_U2857) );
  INV_X1 U17558 ( .A(n16157), .ZN(n14189) );
  OAI222_X1 U17559 ( .A1(n14189), .A2(n14629), .B1(n14188), .B2(n20023), .C1(
        n14795), .C2(n14635), .ZN(P1_U2858) );
  INV_X1 U17560 ( .A(n14191), .ZN(n15956) );
  OAI21_X1 U17561 ( .B1(n14192), .B2(n14182), .A(n15956), .ZN(n14786) );
  INV_X1 U17562 ( .A(n15959), .ZN(n14193) );
  AOI21_X1 U17563 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n16140) );
  INV_X1 U17564 ( .A(n16140), .ZN(n14197) );
  INV_X1 U17565 ( .A(n14783), .ZN(n14196) );
  OAI22_X1 U17566 ( .A1(n14197), .A2(n20010), .B1(n14196), .B2(n19991), .ZN(
        n14202) );
  INV_X1 U17567 ( .A(n15992), .ZN(n14569) );
  NOR2_X1 U17568 ( .A1(n14198), .A2(n14569), .ZN(n15968) );
  INV_X1 U17569 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20796) );
  INV_X1 U17570 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20633) );
  NOR2_X1 U17571 ( .A1(n20796), .A2(n20633), .ZN(n15953) );
  AOI21_X1 U17572 ( .B1(n20796), .B2(n20633), .A(n15953), .ZN(n14199) );
  AOI22_X1 U17573 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20006), .B1(n15968), 
        .B2(n14199), .ZN(n14200) );
  OAI211_X1 U17574 ( .C1(n19996), .C2(n20907), .A(n14200), .B(n19982), .ZN(
        n14201) );
  AOI211_X1 U17575 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(n15969), .A(n14202), 
        .B(n14201), .ZN(n14203) );
  OAI21_X1 U17576 ( .B1(n14786), .B2(n15977), .A(n14203), .ZN(P1_U2824) );
  AOI22_X1 U17577 ( .A1(n16140), .A2(n20021), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14642), .ZN(n14204) );
  OAI21_X1 U17578 ( .B1(n14786), .B2(n14635), .A(n14204), .ZN(P1_U2856) );
  INV_X1 U17579 ( .A(n14205), .ZN(n14207) );
  OAI21_X1 U17580 ( .B1(n10104), .B2(n14207), .A(n14206), .ZN(n14637) );
  XOR2_X1 U17581 ( .A(n14636), .B(n14637), .Z(n16083) );
  INV_X1 U17582 ( .A(n16083), .ZN(n14218) );
  OR2_X1 U17583 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U17584 ( .A1(n15984), .A2(n14210), .ZN(n15995) );
  OAI222_X1 U17585 ( .A1(n14218), .A2(n14635), .B1(n14211), .B2(n20023), .C1(
        n14629), .C2(n15995), .ZN(P1_U2861) );
  OAI22_X1 U17586 ( .A1(n14690), .A2(n14212), .B1(n14695), .B2(n13175), .ZN(
        n14213) );
  AOI21_X1 U17587 ( .B1(n16025), .B2(DATAI_16_), .A(n14213), .ZN(n14215) );
  NAND2_X1 U17588 ( .A1(n14692), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14214) );
  OAI211_X1 U17589 ( .C1(n14786), .C2(n16009), .A(n14215), .B(n14214), .ZN(
        P1_U2888) );
  OAI222_X1 U17590 ( .A1(n16009), .A2(n14218), .B1(n14705), .B2(n14217), .C1(
        n14216), .C2(n14695), .ZN(P1_U2893) );
  INV_X1 U17591 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16999) );
  INV_X1 U17592 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16790) );
  INV_X1 U17593 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U17594 ( .A1(n18236), .A2(n18218), .ZN(n14219) );
  OAI22_X1 U17595 ( .A1(n15763), .A2(n15764), .B1(n14220), .B2(n14219), .ZN(
        n15871) );
  NAND4_X1 U17596 ( .A1(n18699), .A2(n18835), .A3(n16540), .A4(n15871), .ZN(
        n17228) );
  INV_X1 U17597 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16899) );
  NAND2_X1 U17598 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16911) );
  NOR2_X1 U17599 ( .A1(n16899), .A2(n16911), .ZN(n17209) );
  NAND4_X1 U17600 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(n17207), .ZN(n17194) );
  NAND2_X1 U17601 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17149), .ZN(n17121) );
  NAND3_X1 U17602 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n17048) );
  NAND3_X1 U17603 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .ZN(n14221) );
  NAND2_X1 U17604 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17050), .ZN(n17036) );
  NAND4_X1 U17605 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n15664)
         );
  AND2_X1 U17606 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16960) );
  NAND4_X1 U17607 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n16960), .ZN(n14222) );
  NOR4_X1 U17608 ( .A1(n16999), .A2(n17036), .A3(n15664), .A4(n14222), .ZN(
        n16952) );
  NAND2_X1 U17609 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16952), .ZN(n14223) );
  NOR2_X1 U17610 ( .A1(n17280), .A2(n14223), .ZN(n14225) );
  NAND2_X1 U17611 ( .A1(n17221), .A2(n14223), .ZN(n16953) );
  INV_X1 U17612 ( .A(n16953), .ZN(n14224) );
  MUX2_X1 U17613 ( .A(n14225), .B(n14224), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  INV_X1 U17614 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18640) );
  NAND3_X1 U17615 ( .A1(n15706), .A2(n15766), .A3(n18640), .ZN(n18193) );
  NOR2_X1 U17616 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18193), .ZN(n14226) );
  NAND3_X1 U17617 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18788)
         );
  OAI21_X1 U17618 ( .B1(n14226), .B2(n18788), .A(n18486), .ZN(n18199) );
  INV_X1 U17619 ( .A(n18199), .ZN(n14227) );
  INV_X1 U17620 ( .A(n17773), .ZN(n17829) );
  NOR2_X1 U17621 ( .A1(n17829), .A2(n18842), .ZN(n15755) );
  AOI21_X1 U17622 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15755), .ZN(n15756) );
  NOR2_X1 U17623 ( .A1(n14227), .A2(n15756), .ZN(n14229) );
  NAND2_X1 U17624 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18668), .ZN(n18371) );
  NAND2_X1 U17625 ( .A1(n18371), .A2(n18199), .ZN(n15754) );
  OR2_X1 U17626 ( .A1(n18541), .A2(n15754), .ZN(n14228) );
  MUX2_X1 U17627 ( .A(n14229), .B(n14228), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XNOR2_X1 U17628 ( .A(n14231), .B(n14230), .ZN(n19174) );
  OR2_X1 U17629 ( .A1(n18970), .A2(n20696), .ZN(n19182) );
  OAI21_X1 U17630 ( .B1(n19174), .B2(n15629), .A(n19182), .ZN(n14238) );
  NAND2_X1 U17631 ( .A1(n14233), .A2(n14232), .ZN(n14234) );
  NAND2_X1 U17632 ( .A1(n14235), .A2(n14234), .ZN(n19180) );
  OAI21_X1 U17633 ( .B1(n19180), .B2(n15623), .A(n14236), .ZN(n14237) );
  AOI211_X1 U17634 ( .C1(n14239), .C2(n16354), .A(n14238), .B(n14237), .ZN(
        n14248) );
  OAI21_X1 U17635 ( .B1(n14240), .B2(n14241), .A(n15625), .ZN(n14246) );
  OAI21_X1 U17636 ( .B1(n14242), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14241), .ZN(n14243) );
  AOI21_X1 U17637 ( .B1(n14244), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14243), .ZN(n14245) );
  AOI21_X1 U17638 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14246), .A(
        n14245), .ZN(n14247) );
  OAI211_X1 U17639 ( .C1(n13197), .C2(n15614), .A(n14248), .B(n14247), .ZN(
        P2_U3044) );
  XNOR2_X1 U17640 ( .A(n14250), .B(n14249), .ZN(n15260) );
  NOR2_X1 U17641 ( .A1(n19064), .A2(n15355), .ZN(n14252) );
  NAND2_X1 U17642 ( .A1(n18985), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15264) );
  OAI21_X1 U17643 ( .B1(n19021), .B2(n15614), .A(n15264), .ZN(n14251) );
  AOI211_X1 U17644 ( .C1(n15260), .C2(n16359), .A(n14252), .B(n14251), .ZN(
        n14256) );
  NOR2_X1 U17645 ( .A1(n15286), .A2(n15629), .ZN(n14254) );
  OAI211_X1 U17646 ( .C1(n14254), .C2(n15516), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n15261), .ZN(n14255) );
  INV_X1 U17647 ( .A(n14907), .ZN(n14259) );
  NOR2_X1 U17648 ( .A1(n14257), .A2(n9724), .ZN(n14258) );
  AOI21_X1 U17649 ( .B1(n11624), .B2(n14259), .A(n14258), .ZN(n15804) );
  OAI21_X1 U17650 ( .B1(n15804), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16233), 
        .ZN(n14261) );
  NAND2_X1 U17651 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14920) );
  INV_X1 U17652 ( .A(n15792), .ZN(n14260) );
  AOI22_X1 U17653 ( .A1(n14261), .A2(n14920), .B1(n10881), .B2(n14260), .ZN(
        n14264) );
  AOI21_X1 U17654 ( .B1(n15802), .B2(n14262), .A(n14928), .ZN(n14263) );
  OAI22_X1 U17655 ( .A1(n14264), .A2(n14928), .B1(n14263), .B2(n10881), .ZN(
        P1_U3474) );
  NAND4_X1 U17656 ( .A1(n12904), .A2(n19009), .A3(n13659), .A4(n15132), .ZN(
        n14273) );
  INV_X1 U17657 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14265) );
  OAI22_X1 U17658 ( .A1(n14265), .A2(n18981), .B1(n12842), .B2(n20697), .ZN(
        n14270) );
  NAND2_X1 U17659 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n14266), .ZN(n14268) );
  OAI22_X1 U17660 ( .A1(n19053), .A2(n20698), .B1(n14268), .B2(n14267), .ZN(
        n14269) );
  OAI211_X1 U17661 ( .C1(n16278), .C2(n20705), .A(n14273), .B(n14272), .ZN(
        P2_U2824) );
  NAND2_X1 U17662 ( .A1(n14274), .A2(n15124), .ZN(n14276) );
  XOR2_X1 U17663 ( .A(n14276), .B(n14275), .Z(n14297) );
  NAND2_X1 U17664 ( .A1(n15137), .A2(n14289), .ZN(n14280) );
  INV_X1 U17665 ( .A(n15123), .ZN(n14279) );
  NAND2_X1 U17666 ( .A1(n14287), .A2(n10876), .ZN(n14286) );
  INV_X1 U17667 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U17668 ( .A1(n18985), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14292) );
  OAI21_X1 U17669 ( .B1(n19184), .B2(n14281), .A(n14292), .ZN(n14283) );
  NOR2_X1 U17670 ( .A1(n15001), .A2(n15652), .ZN(n14282) );
  OAI211_X1 U17671 ( .C1(n14297), .C2(n19179), .A(n14286), .B(n14285), .ZN(
        P2_U2985) );
  NAND2_X1 U17672 ( .A1(n14287), .A2(n16357), .ZN(n14296) );
  INV_X1 U17673 ( .A(n15383), .ZN(n15366) );
  OAI21_X1 U17674 ( .B1(n14290), .B2(n15366), .A(n14288), .ZN(n15371) );
  NAND3_X1 U17675 ( .A1(n15383), .A2(n14290), .A3(n14289), .ZN(n14291) );
  OAI211_X1 U17676 ( .C1(n15355), .C2(n15059), .A(n14292), .B(n14291), .ZN(
        n14294) );
  NOR2_X1 U17677 ( .A1(n15001), .A2(n15614), .ZN(n14293) );
  AOI211_X1 U17678 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15371), .A(
        n14294), .B(n14293), .ZN(n14295) );
  OAI211_X1 U17679 ( .C1(n14297), .C2(n15623), .A(n14296), .B(n14295), .ZN(
        P2_U3017) );
  AOI22_X1 U17680 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14301) );
  AOI22_X1 U17681 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14300) );
  AOI22_X1 U17682 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17683 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14298) );
  NAND4_X1 U17684 ( .A1(n14301), .A2(n14300), .A3(n14299), .A4(n14298), .ZN(
        n14307) );
  AOI22_X1 U17685 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14305) );
  AOI22_X1 U17686 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U17687 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17688 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14302) );
  NAND4_X1 U17689 ( .A1(n14305), .A2(n14304), .A3(n14303), .A4(n14302), .ZN(
        n14306) );
  NOR2_X1 U17690 ( .A1(n14307), .A2(n14306), .ZN(n16291) );
  AOI22_X1 U17691 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10452), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U17692 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U17693 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U17694 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14308) );
  NAND4_X1 U17695 ( .A1(n14311), .A2(n14310), .A3(n14309), .A4(n14308), .ZN(
        n14317) );
  AOI22_X1 U17696 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U17697 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U17698 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U17699 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14312) );
  NAND4_X1 U17700 ( .A1(n14315), .A2(n14314), .A3(n14313), .A4(n14312), .ZN(
        n14316) );
  OR2_X1 U17701 ( .A1(n14317), .A2(n14316), .ZN(n15047) );
  AOI22_X1 U17702 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10452), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14321) );
  AOI22_X1 U17703 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U17704 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17705 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14318) );
  NAND4_X1 U17706 ( .A1(n14321), .A2(n14320), .A3(n14319), .A4(n14318), .ZN(
        n14327) );
  AOI22_X1 U17707 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14325) );
  AOI22_X1 U17708 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U17709 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17710 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14322) );
  NAND4_X1 U17711 ( .A1(n14325), .A2(n14324), .A3(n14323), .A4(n14322), .ZN(
        n14326) );
  NOR2_X1 U17712 ( .A1(n14327), .A2(n14326), .ZN(n16279) );
  AOI22_X1 U17713 ( .A1(n10452), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14331) );
  AOI22_X1 U17714 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U17715 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U17716 ( .A1(n10459), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14328) );
  NAND4_X1 U17717 ( .A1(n14331), .A2(n14330), .A3(n14329), .A4(n14328), .ZN(
        n14337) );
  AOI22_X1 U17718 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14335) );
  AOI22_X1 U17719 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U17720 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U17721 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14332) );
  NAND4_X1 U17722 ( .A1(n14335), .A2(n14334), .A3(n14333), .A4(n14332), .ZN(
        n14336) );
  NOR2_X1 U17723 ( .A1(n14337), .A2(n14336), .ZN(n15044) );
  NOR2_X1 U17724 ( .A1(n16279), .A2(n15044), .ZN(n14348) );
  AOI22_X1 U17725 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10452), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17726 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U17727 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U17728 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10459), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14338) );
  NAND4_X1 U17729 ( .A1(n14341), .A2(n14340), .A3(n14339), .A4(n14338), .ZN(
        n14347) );
  AOI22_X1 U17730 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14368), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14345) );
  AOI22_X1 U17731 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10384), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14344) );
  AOI22_X1 U17732 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U17733 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14342) );
  NAND4_X1 U17734 ( .A1(n14345), .A2(n14344), .A3(n14343), .A4(n14342), .ZN(
        n14346) );
  OR2_X1 U17735 ( .A1(n14347), .A2(n14346), .ZN(n16285) );
  AND2_X1 U17736 ( .A1(n14348), .A2(n16285), .ZN(n14349) );
  AOI22_X1 U17737 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U17738 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14350) );
  AND2_X1 U17739 ( .A1(n14351), .A2(n14350), .ZN(n14355) );
  AOI22_X1 U17740 ( .A1(n10147), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14354) );
  INV_X1 U17741 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n20951) );
  AOI22_X1 U17742 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14353) );
  XNOR2_X1 U17743 ( .A(n14352), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14490) );
  NAND4_X1 U17744 ( .A1(n14355), .A2(n14354), .A3(n14353), .A4(n14490), .ZN(
        n14362) );
  AOI22_X1 U17745 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9751), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U17746 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14356) );
  AND2_X1 U17747 ( .A1(n14357), .A2(n14356), .ZN(n14360) );
  INV_X1 U17748 ( .A(n14490), .ZN(n14495) );
  INV_X1 U17749 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19523) );
  AOI22_X1 U17750 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14359) );
  AOI22_X1 U17751 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14358) );
  NAND4_X1 U17752 ( .A1(n14360), .A2(n14495), .A3(n14359), .A4(n14358), .ZN(
        n14361) );
  AND2_X1 U17753 ( .A1(n14362), .A2(n14361), .ZN(n14382) );
  NAND2_X1 U17754 ( .A1(n14382), .A2(n13143), .ZN(n14376) );
  AOI22_X1 U17755 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10452), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17756 ( .A1(n10346), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10379), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U17757 ( .A1(n10453), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10459), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14365) );
  AOI22_X1 U17758 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10354), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14364) );
  NAND4_X1 U17759 ( .A1(n14367), .A2(n14366), .A3(n14365), .A4(n14364), .ZN(
        n14375) );
  AOI22_X1 U17760 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14368), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14373) );
  AOI22_X1 U17761 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12265), .B1(
        n10405), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17762 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14369), .B1(
        n10359), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U17763 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10335), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14370) );
  NAND4_X1 U17764 ( .A1(n14373), .A2(n14372), .A3(n14371), .A4(n14370), .ZN(
        n14374) );
  OR2_X1 U17765 ( .A1(n14375), .A2(n14374), .ZN(n14383) );
  XNOR2_X1 U17766 ( .A(n14376), .B(n14383), .ZN(n14379) );
  INV_X1 U17767 ( .A(n14382), .ZN(n14377) );
  NOR2_X1 U17768 ( .A1(n13143), .A2(n14377), .ZN(n15034) );
  NAND2_X1 U17769 ( .A1(n15035), .A2(n15034), .ZN(n15033) );
  NAND2_X1 U17770 ( .A1(n14380), .A2(n14379), .ZN(n14381) );
  NAND2_X1 U17771 ( .A1(n15033), .A2(n14381), .ZN(n15029) );
  NAND2_X1 U17772 ( .A1(n14383), .A2(n14382), .ZN(n14413) );
  AOI22_X1 U17773 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9751), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U17774 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14384) );
  AND2_X1 U17775 ( .A1(n14385), .A2(n14384), .ZN(n14388) );
  AOI22_X1 U17776 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U17777 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14386) );
  NAND4_X1 U17778 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14490), .ZN(
        n14396) );
  AOI22_X1 U17779 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9693), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U17780 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14390) );
  AND2_X1 U17781 ( .A1(n14391), .A2(n14390), .ZN(n14394) );
  AOI22_X1 U17782 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U17783 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14392) );
  NAND4_X1 U17784 ( .A1(n14394), .A2(n14495), .A3(n14393), .A4(n14392), .ZN(
        n14395) );
  NAND2_X1 U17785 ( .A1(n14396), .A2(n14395), .ZN(n14414) );
  NOR2_X1 U17786 ( .A1(n14413), .A2(n14414), .ZN(n14418) );
  NAND2_X1 U17787 ( .A1(n14418), .A2(n13143), .ZN(n14399) );
  OAI21_X1 U17788 ( .B1(n14397), .B2(n14413), .A(n14414), .ZN(n14398) );
  AND2_X1 U17789 ( .A1(n14399), .A2(n14398), .ZN(n15028) );
  AOI22_X1 U17790 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U17791 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14401) );
  AND2_X1 U17792 ( .A1(n14402), .A2(n14401), .ZN(n14405) );
  AOI22_X1 U17793 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14404) );
  AOI22_X1 U17794 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14403) );
  NAND4_X1 U17795 ( .A1(n14405), .A2(n14404), .A3(n14403), .A4(n14490), .ZN(
        n14412) );
  AOI22_X1 U17796 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9693), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17797 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14406) );
  AND2_X1 U17798 ( .A1(n14407), .A2(n14406), .ZN(n14410) );
  AOI22_X1 U17799 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U17800 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14408) );
  NAND4_X1 U17801 ( .A1(n14410), .A2(n14495), .A3(n14409), .A4(n14408), .ZN(
        n14411) );
  NAND2_X1 U17802 ( .A1(n14412), .A2(n14411), .ZN(n14419) );
  INV_X1 U17803 ( .A(n14419), .ZN(n14417) );
  INV_X1 U17804 ( .A(n14413), .ZN(n14416) );
  NOR2_X1 U17805 ( .A1(n14414), .A2(n14419), .ZN(n14415) );
  NAND2_X1 U17806 ( .A1(n14416), .A2(n14415), .ZN(n14441) );
  OAI211_X1 U17807 ( .C1(n14418), .C2(n14417), .A(n14454), .B(n14441), .ZN(
        n14421) );
  NOR2_X1 U17808 ( .A1(n13143), .A2(n14419), .ZN(n15023) );
  INV_X1 U17809 ( .A(n14420), .ZN(n14423) );
  AOI22_X1 U17810 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U17811 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14425) );
  AND2_X1 U17812 ( .A1(n14426), .A2(n14425), .ZN(n14429) );
  AOI22_X1 U17813 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U17814 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14427) );
  NAND4_X1 U17815 ( .A1(n14429), .A2(n14428), .A3(n14427), .A4(n14490), .ZN(
        n14436) );
  AOI22_X1 U17816 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9751), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U17817 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14430) );
  AND2_X1 U17818 ( .A1(n14431), .A2(n14430), .ZN(n14434) );
  AOI22_X1 U17819 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U17820 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14432) );
  NAND4_X1 U17821 ( .A1(n14434), .A2(n14495), .A3(n14433), .A4(n14432), .ZN(
        n14435) );
  AND2_X1 U17822 ( .A1(n14436), .A2(n14435), .ZN(n14439) );
  XNOR2_X1 U17823 ( .A(n14441), .B(n14439), .ZN(n14437) );
  NAND2_X1 U17824 ( .A1(n9761), .A2(n14439), .ZN(n15014) );
  NOR2_X2 U17825 ( .A1(n15015), .A2(n15014), .ZN(n15013) );
  INV_X1 U17826 ( .A(n14439), .ZN(n14440) );
  NOR2_X1 U17827 ( .A1(n14441), .A2(n14440), .ZN(n14455) );
  AOI22_X1 U17828 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U17829 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14442) );
  AND2_X1 U17830 ( .A1(n14443), .A2(n14442), .ZN(n14446) );
  AOI22_X1 U17831 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14445) );
  AOI22_X1 U17832 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14444) );
  NAND4_X1 U17833 ( .A1(n14446), .A2(n14445), .A3(n14444), .A4(n14490), .ZN(
        n14453) );
  AOI22_X1 U17834 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9693), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U17835 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14447) );
  AND2_X1 U17836 ( .A1(n14448), .A2(n14447), .ZN(n14451) );
  AOI22_X1 U17837 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U17838 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14449) );
  NAND4_X1 U17839 ( .A1(n14451), .A2(n14495), .A3(n14450), .A4(n14449), .ZN(
        n14452) );
  AND2_X1 U17840 ( .A1(n14453), .A2(n14452), .ZN(n14457) );
  NAND2_X1 U17841 ( .A1(n14455), .A2(n14457), .ZN(n15002) );
  OAI211_X1 U17842 ( .C1(n14455), .C2(n14457), .A(n15002), .B(n14454), .ZN(
        n14456) );
  INV_X1 U17843 ( .A(n14457), .ZN(n14458) );
  NOR2_X1 U17844 ( .A1(n13143), .A2(n14458), .ZN(n15009) );
  INV_X1 U17845 ( .A(n14459), .ZN(n15003) );
  AOI22_X1 U17846 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9693), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14461) );
  AOI22_X1 U17847 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14460) );
  AND2_X1 U17848 ( .A1(n14461), .A2(n14460), .ZN(n14464) );
  AOI22_X1 U17849 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14463) );
  AOI22_X1 U17850 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14462) );
  NAND4_X1 U17851 ( .A1(n14464), .A2(n14463), .A3(n14462), .A4(n14490), .ZN(
        n14472) );
  AOI22_X1 U17852 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9751), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U17853 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14465) );
  AND2_X1 U17854 ( .A1(n14466), .A2(n14465), .ZN(n14470) );
  AOI22_X1 U17855 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U17856 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14468) );
  NAND4_X1 U17857 ( .A1(n14470), .A2(n14495), .A3(n14469), .A4(n14468), .ZN(
        n14471) );
  NAND2_X1 U17858 ( .A1(n14472), .A2(n14471), .ZN(n15005) );
  AOI22_X1 U17859 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9751), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14474) );
  AOI22_X1 U17860 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14473) );
  AND2_X1 U17861 ( .A1(n14474), .A2(n14473), .ZN(n14477) );
  AOI22_X1 U17862 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U17863 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14475) );
  NAND4_X1 U17864 ( .A1(n14477), .A2(n14476), .A3(n14475), .A4(n14490), .ZN(
        n14484) );
  AOI22_X1 U17865 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14389), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U17866 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14478) );
  AND2_X1 U17867 ( .A1(n14479), .A2(n14478), .ZN(n14482) );
  AOI22_X1 U17868 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U17869 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14480) );
  NAND4_X1 U17870 ( .A1(n14482), .A2(n14495), .A3(n14481), .A4(n14480), .ZN(
        n14483) );
  NAND2_X1 U17871 ( .A1(n14484), .A2(n14483), .ZN(n14486) );
  OR3_X1 U17872 ( .A1(n15002), .A2(n9761), .A3(n15005), .ZN(n14485) );
  NOR2_X1 U17873 ( .A1(n14485), .A2(n14486), .ZN(n14487) );
  AOI21_X1 U17874 ( .B1(n14486), .B2(n14485), .A(n14487), .ZN(n14996) );
  AOI22_X1 U17875 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U17876 ( .A1(n9698), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14488) );
  NAND2_X1 U17877 ( .A1(n14489), .A2(n14488), .ZN(n14501) );
  AOI22_X1 U17878 ( .A1(n9762), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U17879 ( .A1(n10327), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9693), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14491) );
  NAND3_X1 U17880 ( .A1(n14492), .A2(n14491), .A3(n14490), .ZN(n14500) );
  AOI22_X1 U17881 ( .A1(n9757), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U17882 ( .A1(n14467), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10333), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U17883 ( .A1(n14494), .A2(n14493), .ZN(n14499) );
  AOI22_X1 U17884 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10327), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U17885 ( .A1(n9751), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14400), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14496) );
  NAND3_X1 U17886 ( .A1(n14497), .A2(n14496), .A3(n14495), .ZN(n14498) );
  OAI22_X1 U17887 ( .A1(n14501), .A2(n14500), .B1(n14499), .B2(n14498), .ZN(
        n14502) );
  XNOR2_X1 U17888 ( .A(n14503), .B(n14502), .ZN(n14510) );
  NOR2_X1 U17889 ( .A1(n15361), .A2(n19052), .ZN(n14504) );
  AOI21_X1 U17890 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19052), .A(n14504), .ZN(
        n14505) );
  OAI21_X1 U17891 ( .B1(n14510), .B2(n19041), .A(n14505), .ZN(P2_U2857) );
  AOI22_X1 U17892 ( .A1(n19059), .A2(n19071), .B1(n19119), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14507) );
  AOI22_X1 U17893 ( .A1(n19061), .A2(BUF1_REG_30__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14506) );
  OAI211_X1 U17894 ( .C1(n15356), .C2(n19063), .A(n14507), .B(n14506), .ZN(
        n14508) );
  INV_X1 U17895 ( .A(n14508), .ZN(n14509) );
  OAI21_X1 U17896 ( .B1(n14510), .B2(n19124), .A(n14509), .ZN(P2_U2889) );
  AOI22_X1 U17897 ( .A1(n11401), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14514), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14515) );
  NAND2_X1 U17898 ( .A1(n14516), .A2(n19959), .ZN(n14525) );
  INV_X1 U17899 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20644) );
  INV_X1 U17900 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20837) );
  NAND4_X1 U17901 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14517), .A3(
        P1_REIP_REG_15__SCAN_IN), .A4(P1_REIP_REG_16__SCAN_IN), .ZN(n14570) );
  NOR2_X1 U17902 ( .A1(n14518), .A2(n14570), .ZN(n14571) );
  NAND3_X1 U17903 ( .A1(n14571), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n15914) );
  NAND3_X1 U17904 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n15907) );
  NOR3_X1 U17905 ( .A1(n20837), .A2(n15914), .A3(n15907), .ZN(n14559) );
  NAND3_X1 U17906 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20005), .A3(n14559), 
        .ZN(n15895) );
  NOR2_X1 U17907 ( .A1(n20644), .A2(n15895), .ZN(n15887) );
  NAND2_X1 U17908 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n15887), .ZN(n15878) );
  NAND2_X1 U17909 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14519) );
  NOR2_X1 U17910 ( .A1(n15878), .A2(n14519), .ZN(n14537) );
  AND2_X1 U17911 ( .A1(n14537), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14528) );
  AND2_X1 U17912 ( .A1(n14528), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14520) );
  INV_X1 U17913 ( .A(n19949), .ZN(n19963) );
  NOR2_X1 U17914 ( .A1(n14520), .A2(n19963), .ZN(n14527) );
  INV_X1 U17915 ( .A(n14520), .ZN(n14522) );
  AOI22_X1 U17916 ( .A1(n20006), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20014), .ZN(n14521) );
  OAI21_X1 U17917 ( .B1(n14522), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14521), 
        .ZN(n14523) );
  AOI21_X1 U17918 ( .B1(n14527), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14523), 
        .ZN(n14524) );
  OAI211_X1 U17919 ( .C1(n14818), .C2(n20010), .A(n14525), .B(n14524), .ZN(
        P1_U2809) );
  INV_X1 U17920 ( .A(n14526), .ZN(n14833) );
  OAI21_X1 U17921 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14528), .A(n14527), 
        .ZN(n14530) );
  AOI22_X1 U17922 ( .A1(n14711), .A2(n20013), .B1(n20014), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14529) );
  OAI211_X1 U17923 ( .C1(n19984), .C2(n14531), .A(n14530), .B(n14529), .ZN(
        n14532) );
  AOI21_X1 U17924 ( .B1(n14833), .B2(n19993), .A(n14532), .ZN(n14533) );
  OAI21_X1 U17925 ( .B1(n14648), .B2(n15977), .A(n14533), .ZN(P1_U2810) );
  INV_X1 U17926 ( .A(n14721), .ZN(n14653) );
  INV_X1 U17927 ( .A(n14584), .ZN(n14543) );
  INV_X1 U17928 ( .A(n14537), .ZN(n14553) );
  NAND3_X1 U17929 ( .A1(n14553), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n19949), 
        .ZN(n14541) );
  OAI22_X1 U17930 ( .A1(n14538), .A2(n19996), .B1(n19991), .B2(n14719), .ZN(
        n14539) );
  AOI21_X1 U17931 ( .B1(n20006), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14539), .ZN(
        n14540) );
  OAI211_X1 U17932 ( .C1(n14553), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14541), 
        .B(n14540), .ZN(n14542) );
  AOI21_X1 U17933 ( .B1(n14543), .B2(n19993), .A(n14542), .ZN(n14544) );
  OAI21_X1 U17934 ( .B1(n14653), .B2(n15977), .A(n14544), .ZN(P1_U2811) );
  INV_X1 U17935 ( .A(n14534), .ZN(n14546) );
  INV_X1 U17936 ( .A(n14724), .ZN(n14658) );
  INV_X1 U17937 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20647) );
  OAI22_X1 U17938 ( .A1(n15878), .A2(n20647), .B1(n19963), .B2(n14548), .ZN(
        n14552) );
  AOI22_X1 U17939 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n14728), .ZN(n14550) );
  NAND2_X1 U17940 ( .A1(n20006), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14549) );
  OAI211_X1 U17941 ( .C1(n14586), .C2(n20010), .A(n14550), .B(n14549), .ZN(
        n14551) );
  AOI21_X1 U17942 ( .B1(n14553), .B2(n14552), .A(n14551), .ZN(n14554) );
  OAI21_X1 U17943 ( .B1(n14658), .B2(n15977), .A(n14554), .ZN(P1_U2812) );
  BUF_X1 U17944 ( .A(n14556), .Z(n14557) );
  INV_X1 U17945 ( .A(n14557), .ZN(n14602) );
  AOI21_X1 U17946 ( .B1(n14558), .B2(n14555), .A(n14557), .ZN(n14753) );
  INV_X1 U17947 ( .A(n14753), .ZN(n14672) );
  OAI21_X1 U17948 ( .B1(n19980), .B2(n14559), .A(n20009), .ZN(n15908) );
  NOR2_X1 U17949 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n19980), .ZN(n15901) );
  AOI22_X1 U17950 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(n20006), .B1(n14559), 
        .B2(n15901), .ZN(n14560) );
  OAI21_X1 U17951 ( .B1(n14755), .B2(n19996), .A(n14560), .ZN(n14561) );
  AOI21_X1 U17952 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n15908), .A(n14561), 
        .ZN(n14565) );
  INV_X1 U17953 ( .A(n14757), .ZN(n14562) );
  OAI22_X1 U17954 ( .A1(n14610), .A2(n20010), .B1(n14562), .B2(n19991), .ZN(
        n14563) );
  INV_X1 U17955 ( .A(n14563), .ZN(n14564) );
  OAI211_X1 U17956 ( .C1(n14672), .C2(n15977), .A(n14565), .B(n14564), .ZN(
        P1_U2816) );
  OAI21_X1 U17957 ( .B1(n14566), .B2(n14568), .A(n14567), .ZN(n14773) );
  NOR2_X1 U17958 ( .A1(n14570), .A2(n14569), .ZN(n15942) );
  INV_X1 U17959 ( .A(n14571), .ZN(n14572) );
  AOI21_X1 U17960 ( .B1(n20005), .B2(n14572), .A(n19992), .ZN(n15963) );
  AOI22_X1 U17961 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20014), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(n20006), .ZN(n14573) );
  OAI211_X1 U17962 ( .C1(n15963), .C2(n14771), .A(n14573), .B(n19982), .ZN(
        n14581) );
  INV_X1 U17963 ( .A(n15958), .ZN(n14576) );
  INV_X1 U17964 ( .A(n14574), .ZN(n14575) );
  OAI21_X1 U17965 ( .B1(n15959), .B2(n14576), .A(n14575), .ZN(n14577) );
  AND2_X1 U17966 ( .A1(n14577), .A2(n15950), .ZN(n16122) );
  INV_X1 U17967 ( .A(n16122), .ZN(n14579) );
  INV_X1 U17968 ( .A(n14776), .ZN(n14578) );
  OAI22_X1 U17969 ( .A1(n14579), .A2(n20010), .B1(n14578), .B2(n19991), .ZN(
        n14580) );
  AOI211_X1 U17970 ( .C1(n15942), .C2(n14771), .A(n14581), .B(n14580), .ZN(
        n14582) );
  OAI21_X1 U17971 ( .B1(n14773), .B2(n15977), .A(n14582), .ZN(P1_U2822) );
  INV_X1 U17972 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14583) );
  OAI22_X1 U17973 ( .A1(n14818), .A2(n14629), .B1(n20023), .B2(n14583), .ZN(
        P1_U2841) );
  OAI222_X1 U17974 ( .A1(n14635), .A2(n14653), .B1(n14585), .B2(n20023), .C1(
        n14584), .C2(n14629), .ZN(P1_U2843) );
  INV_X1 U17975 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14587) );
  OAI222_X1 U17976 ( .A1(n14635), .A2(n14658), .B1(n14587), .B2(n20023), .C1(
        n14586), .C2(n14629), .ZN(P1_U2844) );
  OR2_X1 U17977 ( .A1(n14595), .A2(n14588), .ZN(n14589) );
  INV_X1 U17978 ( .A(n16010), .ZN(n14593) );
  NAND2_X1 U17979 ( .A1(n9802), .A2(n14590), .ZN(n14591) );
  NAND2_X1 U17980 ( .A1(n9788), .A2(n14591), .ZN(n15881) );
  OAI222_X1 U17981 ( .A1(n14635), .A2(n14593), .B1(n14592), .B2(n20023), .C1(
        n15881), .C2(n14629), .ZN(P1_U2845) );
  INV_X1 U17982 ( .A(n14595), .ZN(n14596) );
  INV_X1 U17983 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14600) );
  OR2_X1 U17984 ( .A1(n14607), .A2(n14598), .ZN(n14599) );
  NAND2_X1 U17985 ( .A1(n9802), .A2(n14599), .ZN(n15884) );
  AND2_X1 U17986 ( .A1(n14602), .A2(n14601), .ZN(n14603) );
  OR2_X1 U17987 ( .A1(n14603), .A2(n14594), .ZN(n15892) );
  NOR2_X1 U17988 ( .A1(n14605), .A2(n14604), .ZN(n14606) );
  OR2_X1 U17989 ( .A1(n14607), .A2(n14606), .ZN(n15904) );
  OAI22_X1 U17990 ( .A1(n15904), .A2(n14629), .B1(n15893), .B2(n20023), .ZN(
        n14608) );
  INV_X1 U17991 ( .A(n14608), .ZN(n14609) );
  OAI21_X1 U17992 ( .B1(n15892), .B2(n14635), .A(n14609), .ZN(P1_U2847) );
  INV_X1 U17993 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14611) );
  OAI222_X1 U17994 ( .A1(n14635), .A2(n14672), .B1(n14611), .B2(n20023), .C1(
        n14610), .C2(n14629), .ZN(P1_U2848) );
  NAND2_X1 U17996 ( .A1(n14613), .A2(n14614), .ZN(n14615) );
  AND2_X1 U17997 ( .A1(n14555), .A2(n14615), .ZN(n16031) );
  NAND2_X1 U17998 ( .A1(n9792), .A2(n14616), .ZN(n14617) );
  NAND2_X1 U17999 ( .A1(n14618), .A2(n14617), .ZN(n15912) );
  OAI22_X1 U18000 ( .A1(n15912), .A2(n14629), .B1(n15905), .B2(n20023), .ZN(
        n14619) );
  AOI21_X1 U18001 ( .B1(n16031), .B2(n12893), .A(n14619), .ZN(n14620) );
  INV_X1 U18002 ( .A(n14620), .ZN(P1_U2849) );
  OR2_X1 U18003 ( .A1(n9905), .A2(n14621), .ZN(n14622) );
  NAND2_X1 U18004 ( .A1(n9792), .A2(n14622), .ZN(n16107) );
  INV_X1 U18005 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14625) );
  OAI21_X1 U18006 ( .B1(n14623), .B2(n14624), .A(n14613), .ZN(n15916) );
  OAI222_X1 U18007 ( .A1(n16107), .A2(n14629), .B1(n20023), .B2(n14625), .C1(
        n15916), .C2(n14635), .ZN(P1_U2850) );
  AOI21_X1 U18008 ( .B1(n14626), .B2(n9803), .A(n14623), .ZN(n16036) );
  NOR2_X1 U18009 ( .A1(n15856), .A2(n14627), .ZN(n14628) );
  OR2_X1 U18010 ( .A1(n9905), .A2(n14628), .ZN(n15927) );
  OAI22_X1 U18011 ( .A1(n15927), .A2(n14629), .B1(n15924), .B2(n20023), .ZN(
        n14630) );
  AOI21_X1 U18012 ( .B1(n16036), .B2(n12893), .A(n14630), .ZN(n14631) );
  INV_X1 U18013 ( .A(n14631), .ZN(P1_U2851) );
  NOR2_X1 U18014 ( .A1(n20023), .A2(n14632), .ZN(n14633) );
  AOI21_X1 U18015 ( .B1(n16122), .B2(n20021), .A(n14633), .ZN(n14634) );
  OAI21_X1 U18016 ( .B1(n14773), .B2(n14635), .A(n14634), .ZN(P1_U2854) );
  OAI21_X1 U18017 ( .B1(n14637), .B2(n14636), .A(n14206), .ZN(n14699) );
  XNOR2_X1 U18018 ( .A(n14641), .B(n14640), .ZN(n16166) );
  AOI22_X1 U18019 ( .A1(n16166), .A2(n20021), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14642), .ZN(n14643) );
  OAI21_X1 U18020 ( .B1(n15978), .B2(n14635), .A(n14643), .ZN(P1_U2859) );
  OAI22_X1 U18021 ( .A1(n14690), .A2(n14644), .B1(n14695), .B2(n13350), .ZN(
        n14645) );
  AOI21_X1 U18022 ( .B1(n16025), .B2(DATAI_30_), .A(n14645), .ZN(n14647) );
  NAND2_X1 U18023 ( .A1(n14692), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14646) );
  OAI211_X1 U18024 ( .C1(n14648), .C2(n16009), .A(n14647), .B(n14646), .ZN(
        P1_U2874) );
  OAI22_X1 U18025 ( .A1(n14690), .A2(n14698), .B1(n14695), .B2(n14649), .ZN(
        n14650) );
  AOI21_X1 U18026 ( .B1(n16025), .B2(DATAI_29_), .A(n14650), .ZN(n14652) );
  NAND2_X1 U18027 ( .A1(n14692), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14651) );
  OAI211_X1 U18028 ( .C1(n14653), .C2(n16009), .A(n14652), .B(n14651), .ZN(
        P1_U2875) );
  OAI22_X1 U18029 ( .A1(n14690), .A2(n14706), .B1(n14695), .B2(n14654), .ZN(
        n14655) );
  AOI21_X1 U18030 ( .B1(n16025), .B2(DATAI_28_), .A(n14655), .ZN(n14657) );
  NAND2_X1 U18031 ( .A1(n14692), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14656) );
  OAI211_X1 U18032 ( .C1(n14658), .C2(n16009), .A(n14657), .B(n14656), .ZN(
        P1_U2876) );
  OAI22_X1 U18033 ( .A1(n14690), .A2(n14659), .B1(n14695), .B2(n13234), .ZN(
        n14660) );
  AOI21_X1 U18034 ( .B1(n16025), .B2(DATAI_26_), .A(n14660), .ZN(n14662) );
  NAND2_X1 U18035 ( .A1(n14692), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14661) );
  OAI211_X1 U18036 ( .C1(n15885), .C2(n16009), .A(n14662), .B(n14661), .ZN(
        P1_U2878) );
  OAI22_X1 U18037 ( .A1(n14690), .A2(n14664), .B1(n14695), .B2(n14663), .ZN(
        n14665) );
  AOI21_X1 U18038 ( .B1(n16025), .B2(DATAI_25_), .A(n14665), .ZN(n14667) );
  NAND2_X1 U18039 ( .A1(n14692), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14666) );
  OAI211_X1 U18040 ( .C1(n15892), .C2(n16009), .A(n14667), .B(n14666), .ZN(
        P1_U2879) );
  OAI22_X1 U18041 ( .A1(n14690), .A2(n14668), .B1(n14695), .B2(n13360), .ZN(
        n14669) );
  AOI21_X1 U18042 ( .B1(n16025), .B2(DATAI_24_), .A(n14669), .ZN(n14671) );
  NAND2_X1 U18043 ( .A1(n14692), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14670) );
  OAI211_X1 U18044 ( .C1(n14672), .C2(n16009), .A(n14671), .B(n14670), .ZN(
        P1_U2880) );
  INV_X1 U18045 ( .A(n16031), .ZN(n14678) );
  OAI22_X1 U18046 ( .A1(n14690), .A2(n14674), .B1(n14695), .B2(n14673), .ZN(
        n14675) );
  AOI21_X1 U18047 ( .B1(n16025), .B2(DATAI_23_), .A(n14675), .ZN(n14677) );
  NAND2_X1 U18048 ( .A1(n14692), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14676) );
  OAI211_X1 U18049 ( .C1(n14678), .C2(n16009), .A(n14677), .B(n14676), .ZN(
        P1_U2881) );
  OAI22_X1 U18050 ( .A1(n14690), .A2(n14680), .B1(n14695), .B2(n14679), .ZN(
        n14681) );
  AOI21_X1 U18051 ( .B1(n16025), .B2(DATAI_22_), .A(n14681), .ZN(n14683) );
  NAND2_X1 U18052 ( .A1(n14692), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14682) );
  OAI211_X1 U18053 ( .C1(n15916), .C2(n16009), .A(n14683), .B(n14682), .ZN(
        P1_U2882) );
  INV_X1 U18054 ( .A(n16036), .ZN(n14688) );
  OAI22_X1 U18055 ( .A1(n14690), .A2(n14684), .B1(n14695), .B2(n20858), .ZN(
        n14685) );
  AOI21_X1 U18056 ( .B1(n16025), .B2(DATAI_21_), .A(n14685), .ZN(n14687) );
  NAND2_X1 U18057 ( .A1(n14692), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14686) );
  OAI211_X1 U18058 ( .C1(n14688), .C2(n16009), .A(n14687), .B(n14686), .ZN(
        P1_U2883) );
  OAI22_X1 U18059 ( .A1(n14690), .A2(n14689), .B1(n14695), .B2(n13178), .ZN(
        n14691) );
  AOI21_X1 U18060 ( .B1(n16025), .B2(DATAI_18_), .A(n14691), .ZN(n14694) );
  NAND2_X1 U18061 ( .A1(n14692), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14693) );
  OAI211_X1 U18062 ( .C1(n14773), .C2(n16009), .A(n14694), .B(n14693), .ZN(
        P1_U2886) );
  INV_X1 U18063 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20025) );
  OAI222_X1 U18064 ( .A1(n16009), .A2(n14697), .B1(n14705), .B2(n14696), .C1(
        n14695), .C2(n20025), .ZN(P1_U2889) );
  OAI222_X1 U18065 ( .A1(n16009), .A2(n15978), .B1(n14698), .B2(n14705), .C1(
        n14695), .C2(n13403), .ZN(P1_U2891) );
  INV_X1 U18066 ( .A(n14699), .ZN(n14703) );
  INV_X1 U18067 ( .A(n14700), .ZN(n14702) );
  INV_X1 U18068 ( .A(n16079), .ZN(n14707) );
  INV_X1 U18069 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14704) );
  OAI222_X1 U18070 ( .A1(n14707), .A2(n16009), .B1(n14706), .B2(n14705), .C1(
        n14704), .C2(n14695), .ZN(P1_U2892) );
  NAND2_X1 U18071 ( .A1(n14709), .A2(n11604), .ZN(n14710) );
  INV_X1 U18072 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14820) );
  NAND2_X1 U18073 ( .A1(n20070), .A2(n14711), .ZN(n14712) );
  NAND2_X1 U18074 ( .A1(n20106), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14829) );
  OAI211_X1 U18075 ( .C1(n14713), .C2(n14803), .A(n14712), .B(n14829), .ZN(
        n14714) );
  AOI21_X1 U18076 ( .B1(n14715), .B2(n20062), .A(n14714), .ZN(n14716) );
  OAI21_X1 U18077 ( .B1(n19906), .B2(n14835), .A(n14716), .ZN(P1_U2969) );
  AOI21_X1 U18078 ( .B1(n20067), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14717), .ZN(n14718) );
  OAI21_X1 U18079 ( .B1(n20066), .B2(n14719), .A(n14718), .ZN(n14720) );
  AOI21_X1 U18080 ( .B1(n14721), .B2(n20062), .A(n14720), .ZN(n14722) );
  OAI21_X1 U18081 ( .B1(n14723), .B2(n19906), .A(n14722), .ZN(P1_U2970) );
  NAND2_X1 U18082 ( .A1(n14724), .A2(n20062), .ZN(n14730) );
  INV_X1 U18083 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14725) );
  NOR2_X1 U18084 ( .A1(n14803), .A2(n14725), .ZN(n14726) );
  AOI211_X1 U18085 ( .C1(n20070), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        n14729) );
  OAI211_X1 U18086 ( .C1(n14731), .C2(n19906), .A(n14730), .B(n14729), .ZN(
        P1_U2971) );
  MUX2_X1 U18087 ( .A(n14732), .B(n9812), .S(n16056), .Z(n14733) );
  XNOR2_X1 U18088 ( .A(n14733), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14842) );
  NOR2_X1 U18089 ( .A1(n16209), .A2(n20647), .ZN(n14836) );
  AOI21_X1 U18090 ( .B1(n20067), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14836), .ZN(n14734) );
  OAI21_X1 U18091 ( .B1(n20066), .B2(n15875), .A(n14734), .ZN(n14735) );
  AOI21_X1 U18092 ( .B1(n16010), .B2(n20062), .A(n14735), .ZN(n14736) );
  OAI21_X1 U18093 ( .B1(n19906), .B2(n14842), .A(n14736), .ZN(P1_U2972) );
  NOR2_X1 U18094 ( .A1(n14737), .A2(n16056), .ZN(n14739) );
  OAI21_X1 U18095 ( .B1(n14740), .B2(n14739), .A(n14738), .ZN(n14741) );
  XNOR2_X1 U18096 ( .A(n14741), .B(n14844), .ZN(n14852) );
  NAND2_X1 U18097 ( .A1(n20106), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14847) );
  OAI21_X1 U18098 ( .B1(n14803), .B2(n15891), .A(n14847), .ZN(n14743) );
  NOR2_X1 U18099 ( .A1(n15885), .A2(n20076), .ZN(n14742) );
  AOI211_X1 U18100 ( .C1(n20070), .C2(n15882), .A(n14743), .B(n14742), .ZN(
        n14744) );
  OAI21_X1 U18101 ( .B1(n19906), .B2(n14852), .A(n14744), .ZN(P1_U2973) );
  NOR2_X1 U18102 ( .A1(n16209), .A2(n20644), .ZN(n14855) );
  NOR2_X1 U18103 ( .A1(n20066), .A2(n15896), .ZN(n14745) );
  AOI211_X1 U18104 ( .C1(n20067), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14855), .B(n14745), .ZN(n14752) );
  NOR3_X1 U18105 ( .A1(n11536), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14749) );
  INV_X1 U18106 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14746) );
  NOR2_X1 U18107 ( .A1(n14747), .A2(n14746), .ZN(n14748) );
  MUX2_X1 U18108 ( .A(n14749), .B(n14748), .S(n9749), .Z(n14750) );
  XNOR2_X1 U18109 ( .A(n14750), .B(n11534), .ZN(n14853) );
  NAND2_X1 U18110 ( .A1(n14853), .A2(n20071), .ZN(n14751) );
  OAI211_X1 U18111 ( .C1(n15892), .C2(n20076), .A(n14752), .B(n14751), .ZN(
        P1_U2974) );
  NAND2_X1 U18112 ( .A1(n14753), .A2(n20062), .ZN(n14759) );
  INV_X1 U18113 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14754) );
  OAI22_X1 U18114 ( .A1(n14803), .A2(n14755), .B1(n16209), .B2(n14754), .ZN(
        n14756) );
  AOI21_X1 U18115 ( .B1(n20070), .B2(n14757), .A(n14756), .ZN(n14758) );
  OAI211_X1 U18116 ( .C1(n14760), .C2(n19906), .A(n14759), .B(n14758), .ZN(
        P1_U2975) );
  INV_X1 U18117 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14761) );
  OAI22_X1 U18118 ( .A1(n14803), .A2(n15922), .B1(n16209), .B2(n14761), .ZN(
        n14762) );
  AOI21_X1 U18119 ( .B1(n20070), .B2(n15913), .A(n14762), .ZN(n14767) );
  NAND2_X1 U18120 ( .A1(n14763), .A2(n14764), .ZN(n14765) );
  XNOR2_X1 U18121 ( .A(n14765), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16105) );
  NAND2_X1 U18122 ( .A1(n16105), .A2(n20071), .ZN(n14766) );
  OAI211_X1 U18123 ( .C1(n15916), .C2(n20076), .A(n14767), .B(n14766), .ZN(
        P1_U2977) );
  OAI21_X1 U18124 ( .B1(n14768), .B2(n14770), .A(n15845), .ZN(n16121) );
  INV_X1 U18125 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14772) );
  INV_X1 U18126 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14771) );
  OAI22_X1 U18127 ( .A1(n14803), .A2(n14772), .B1(n16209), .B2(n14771), .ZN(
        n14775) );
  NOR2_X1 U18128 ( .A1(n14773), .A2(n20076), .ZN(n14774) );
  AOI211_X1 U18129 ( .C1(n20070), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14777) );
  OAI21_X1 U18130 ( .B1(n19906), .B2(n16121), .A(n14777), .ZN(P1_U2981) );
  OAI21_X1 U18131 ( .B1(n14879), .B2(n14780), .A(n14779), .ZN(n14787) );
  NOR2_X1 U18132 ( .A1(n14787), .A2(n9818), .ZN(n16066) );
  OAI21_X1 U18133 ( .B1(n16066), .B2(n14781), .A(n16067), .ZN(n16055) );
  XNOR2_X1 U18134 ( .A(n16055), .B(n16053), .ZN(n16141) );
  NAND2_X1 U18135 ( .A1(n16141), .A2(n20071), .ZN(n14785) );
  OAI22_X1 U18136 ( .A1(n14803), .A2(n20907), .B1(n16209), .B2(n20633), .ZN(
        n14782) );
  AOI21_X1 U18137 ( .B1(n14783), .B2(n20070), .A(n14782), .ZN(n14784) );
  OAI211_X1 U18138 ( .C1(n20076), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        P1_U2983) );
  OAI21_X1 U18139 ( .B1(n14788), .B2(n9750), .A(n14787), .ZN(n14790) );
  XNOR2_X1 U18140 ( .A(n9750), .B(n16164), .ZN(n14789) );
  XNOR2_X1 U18141 ( .A(n14790), .B(n14789), .ZN(n16159) );
  NAND2_X1 U18142 ( .A1(n16159), .A2(n20071), .ZN(n14794) );
  NOR2_X1 U18143 ( .A1(n16209), .A2(n20630), .ZN(n16156) );
  NOR2_X1 U18144 ( .A1(n20066), .A2(n14791), .ZN(n14792) );
  AOI211_X1 U18145 ( .C1(n20067), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16156), .B(n14792), .ZN(n14793) );
  OAI211_X1 U18146 ( .C1(n20076), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        P1_U2985) );
  INV_X1 U18147 ( .A(n14796), .ZN(n14797) );
  AOI22_X1 U18148 ( .A1(n14879), .A2(n14798), .B1(n16056), .B2(n14797), .ZN(
        n16077) );
  INV_X1 U18149 ( .A(n14800), .ZN(n14799) );
  AOI21_X1 U18150 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16056), .A(
        n14799), .ZN(n16076) );
  NAND2_X1 U18151 ( .A1(n16077), .A2(n16076), .ZN(n16075) );
  NAND2_X1 U18152 ( .A1(n16075), .A2(n14800), .ZN(n14802) );
  XNOR2_X1 U18153 ( .A(n14802), .B(n14801), .ZN(n16174) );
  NAND2_X1 U18154 ( .A1(n16174), .A2(n20071), .ZN(n14806) );
  NOR2_X1 U18155 ( .A1(n16209), .A2(n20629), .ZN(n16165) );
  NOR2_X1 U18156 ( .A1(n14803), .A2(n15975), .ZN(n14804) );
  AOI211_X1 U18157 ( .C1(n20070), .C2(n15981), .A(n16165), .B(n14804), .ZN(
        n14805) );
  OAI211_X1 U18158 ( .C1(n20076), .C2(n15978), .A(n14806), .B(n14805), .ZN(
        P1_U2986) );
  NAND2_X1 U18159 ( .A1(n14809), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14808) );
  XNOR2_X1 U18160 ( .A(n14879), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14807) );
  MUX2_X1 U18161 ( .A(n14808), .B(n14807), .S(n9749), .Z(n14811) );
  INV_X1 U18162 ( .A(n14809), .ZN(n14810) );
  NAND3_X1 U18163 ( .A1(n14810), .A2(n16056), .A3(n16194), .ZN(n14880) );
  NAND2_X1 U18164 ( .A1(n14811), .A2(n14880), .ZN(n16190) );
  NAND2_X1 U18165 ( .A1(n16190), .A2(n20071), .ZN(n14816) );
  INV_X1 U18166 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14812) );
  NOR2_X1 U18167 ( .A1(n16209), .A2(n14812), .ZN(n16188) );
  NOR2_X1 U18168 ( .A1(n20066), .A2(n14813), .ZN(n14814) );
  AOI211_X1 U18169 ( .C1(n20067), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16188), .B(n14814), .ZN(n14815) );
  OAI211_X1 U18170 ( .C1(n20076), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        P1_U2989) );
  NOR4_X1 U18171 ( .A1(n14827), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14820), .A4(n11604), .ZN(n14824) );
  INV_X1 U18172 ( .A(n14856), .ZN(n14843) );
  INV_X1 U18173 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14821) );
  AOI211_X2 U18174 ( .C1(n11604), .C2(n16201), .A(n14820), .B(n14819), .ZN(
        n14830) );
  AOI211_X1 U18175 ( .C1(n16143), .C2(n14843), .A(n14821), .B(n14830), .ZN(
        n14822) );
  OAI21_X1 U18176 ( .B1(n14826), .B2(n16186), .A(n14825), .ZN(P1_U3000) );
  INV_X1 U18177 ( .A(n14827), .ZN(n14828) );
  AOI21_X1 U18178 ( .B1(n14828), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14831) );
  OAI21_X1 U18179 ( .B1(n14831), .B2(n14830), .A(n14829), .ZN(n14832) );
  AOI21_X1 U18180 ( .B1(n14833), .B2(n20098), .A(n14832), .ZN(n14834) );
  OAI21_X1 U18181 ( .B1(n14835), .B2(n16186), .A(n14834), .ZN(P1_U3001) );
  AOI21_X1 U18182 ( .B1(n14837), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14836), .ZN(n14838) );
  OAI21_X1 U18183 ( .B1(n15881), .B2(n16210), .A(n14838), .ZN(n14839) );
  AOI21_X1 U18184 ( .B1(n14840), .B2(n11581), .A(n14839), .ZN(n14841) );
  OAI21_X1 U18185 ( .B1(n14842), .B2(n16186), .A(n14841), .ZN(P1_U3004) );
  INV_X1 U18186 ( .A(n14868), .ZN(n14846) );
  NAND4_X1 U18187 ( .A1(n14846), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n11534), .ZN(n14857) );
  AOI21_X1 U18188 ( .B1(n14857), .B2(n14843), .A(n14844), .ZN(n14850) );
  NAND3_X1 U18189 ( .A1(n14846), .A2(n14845), .A3(n14844), .ZN(n14848) );
  OAI211_X1 U18190 ( .C1(n16210), .C2(n15884), .A(n14848), .B(n14847), .ZN(
        n14849) );
  NOR2_X1 U18191 ( .A1(n14850), .A2(n14849), .ZN(n14851) );
  OAI21_X1 U18192 ( .B1(n14852), .B2(n16186), .A(n14851), .ZN(P1_U3005) );
  INV_X1 U18193 ( .A(n14853), .ZN(n14859) );
  NOR2_X1 U18194 ( .A1(n15904), .A2(n16210), .ZN(n14854) );
  AOI211_X1 U18195 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n14856), .A(
        n14855), .B(n14854), .ZN(n14858) );
  OAI211_X1 U18196 ( .C1(n14859), .C2(n16186), .A(n14858), .B(n14857), .ZN(
        P1_U3006) );
  XNOR2_X1 U18197 ( .A(n9750), .B(n14862), .ZN(n14860) );
  XNOR2_X1 U18198 ( .A(n11536), .B(n14860), .ZN(n16030) );
  NAND2_X1 U18199 ( .A1(n16030), .A2(n20103), .ZN(n14867) );
  INV_X1 U18200 ( .A(n15912), .ZN(n14865) );
  NAND2_X1 U18201 ( .A1(n20106), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14861) );
  OAI21_X1 U18202 ( .B1(n14863), .B2(n14862), .A(n14861), .ZN(n14864) );
  AOI21_X1 U18203 ( .B1(n14865), .B2(n20098), .A(n14864), .ZN(n14866) );
  OAI211_X1 U18204 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14868), .A(
        n14867), .B(n14866), .ZN(P1_U3008) );
  INV_X1 U18205 ( .A(n16106), .ZN(n14877) );
  NOR2_X1 U18206 ( .A1(n9749), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16046) );
  INV_X1 U18207 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16129) );
  OAI21_X1 U18208 ( .B1(n9750), .B2(n16129), .A(n15845), .ZN(n16048) );
  OAI22_X1 U18209 ( .A1(n16048), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16056), .B2(n15845), .ZN(n14869) );
  OAI21_X1 U18210 ( .B1(n11306), .B2(n16046), .A(n14869), .ZN(n14870) );
  XNOR2_X1 U18211 ( .A(n14870), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16035) );
  NAND2_X1 U18212 ( .A1(n16035), .A2(n20103), .ZN(n14876) );
  INV_X1 U18213 ( .A(n14871), .ZN(n14872) );
  NOR2_X1 U18214 ( .A1(n16134), .A2(n14872), .ZN(n16110) );
  INV_X1 U18215 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14873) );
  OAI22_X1 U18216 ( .A1(n15927), .A2(n16210), .B1(n16209), .B2(n14873), .ZN(
        n14874) );
  AOI21_X1 U18217 ( .B1(n16110), .B2(n14878), .A(n14874), .ZN(n14875) );
  OAI211_X1 U18218 ( .C1(n14878), .C2(n14877), .A(n14876), .B(n14875), .ZN(
        P1_U3010) );
  NAND3_X1 U18219 ( .A1(n14879), .A2(n9749), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14881) );
  NAND2_X1 U18220 ( .A1(n14881), .A2(n14880), .ZN(n14882) );
  XOR2_X1 U18221 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n14882), .Z(
        n16084) );
  AOI21_X1 U18222 ( .B1(n14886), .B2(n14883), .A(n20101), .ZN(n14885) );
  AOI211_X1 U18223 ( .C1(n20097), .C2(n16181), .A(n14885), .B(n14884), .ZN(
        n16179) );
  INV_X1 U18224 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14887) );
  NAND2_X1 U18225 ( .A1(n14886), .A2(n14887), .ZN(n16180) );
  OAI22_X1 U18226 ( .A1(n16179), .A2(n14887), .B1(n16225), .B2(n16180), .ZN(
        n14890) );
  INV_X1 U18227 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n14888) );
  OAI22_X1 U18228 ( .A1(n15995), .A2(n16210), .B1(n16209), .B2(n14888), .ZN(
        n14889) );
  AOI211_X1 U18229 ( .C1(n16084), .C2(n20103), .A(n14890), .B(n14889), .ZN(
        n14891) );
  INV_X1 U18230 ( .A(n14891), .ZN(P1_U3020) );
  OR2_X1 U18231 ( .A1(n14892), .A2(n16186), .ZN(n14899) );
  AOI21_X1 U18232 ( .B1(n20098), .B2(n14894), .A(n14893), .ZN(n14898) );
  OAI21_X1 U18233 ( .B1(n16169), .B2(n14895), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14896) );
  NAND4_X1 U18234 ( .A1(n14899), .A2(n14898), .A3(n14897), .A4(n14896), .ZN(
        P1_U3031) );
  OAI21_X1 U18235 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14902), .A(n20533), 
        .ZN(n14900) );
  OAI21_X1 U18236 ( .B1(n14905), .B2(n20436), .A(n14900), .ZN(n14901) );
  MUX2_X1 U18237 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14901), .S(
        n20113), .Z(P1_U3477) );
  NAND3_X1 U18238 ( .A1(n14902), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20538), 
        .ZN(n14903) );
  INV_X1 U18239 ( .A(n20533), .ZN(n20395) );
  MUX2_X1 U18240 ( .A(n14903), .B(n20395), .S(n20115), .Z(n14904) );
  OAI21_X1 U18241 ( .B1(n14905), .B2(n13519), .A(n14904), .ZN(n14906) );
  MUX2_X1 U18242 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14906), .S(
        n20113), .Z(P1_U3476) );
  OR2_X1 U18243 ( .A1(n20436), .A2(n14907), .ZN(n14911) );
  NOR2_X1 U18244 ( .A1(n13530), .A2(n13502), .ZN(n14909) );
  AOI22_X1 U18245 ( .A1(n15802), .A2(n11113), .B1(n14909), .B2(n14908), .ZN(
        n14910) );
  NAND2_X1 U18246 ( .A1(n14911), .A2(n14910), .ZN(n15801) );
  INV_X1 U18247 ( .A(n15801), .ZN(n14915) );
  AOI22_X1 U18248 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n11402), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14821), .ZN(n14919) );
  INV_X1 U18249 ( .A(n14920), .ZN(n14913) );
  NOR3_X1 U18250 ( .A1(n13530), .A2(n13502), .A3(n15792), .ZN(n14912) );
  AOI21_X1 U18251 ( .B1(n14919), .B2(n14913), .A(n14912), .ZN(n14914) );
  OAI21_X1 U18252 ( .B1(n14915), .B2(n14926), .A(n14914), .ZN(n14917) );
  MUX2_X1 U18253 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14917), .S(
        n14916), .Z(P1_U3473) );
  INV_X1 U18254 ( .A(n14918), .ZN(n14921) );
  OAI222_X1 U18255 ( .A1(n14922), .A2(n15792), .B1(n14926), .B2(n14921), .C1(
        n14920), .C2(n14919), .ZN(n14923) );
  MUX2_X1 U18256 ( .A(n14923), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14928), .Z(P1_U3472) );
  INV_X1 U18257 ( .A(n14924), .ZN(n14927) );
  OAI22_X1 U18258 ( .A1(n14927), .A2(n14926), .B1(n14925), .B2(n15792), .ZN(
        n14929) );
  MUX2_X1 U18259 ( .A(n14929), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14928), .Z(P1_U3469) );
  INV_X1 U18260 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n14931) );
  NAND2_X1 U18261 ( .A1(n14931), .A2(n14930), .ZN(n14933) );
  MUX2_X1 U18262 ( .A(n14934), .B(n14933), .S(n14932), .Z(P2_U3612) );
  NAND3_X1 U18263 ( .A1(n14935), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14936), 
        .ZN(n14938) );
  OAI21_X1 U18264 ( .B1(n14936), .B2(n19666), .A(n10231), .ZN(n14937) );
  MUX2_X1 U18265 ( .A(n14938), .B(n14937), .S(n9761), .Z(n14941) );
  OAI21_X1 U18266 ( .B1(n19793), .B2(n19723), .A(n14939), .ZN(n14940) );
  NAND2_X1 U18267 ( .A1(n14941), .A2(n14940), .ZN(n14947) );
  INV_X1 U18268 ( .A(n14942), .ZN(n14945) );
  NOR2_X1 U18269 ( .A1(n19793), .A2(n19156), .ZN(n14944) );
  AOI211_X1 U18270 ( .C1(n19668), .C2(n14945), .A(n14944), .B(n14943), .ZN(
        n14946) );
  MUX2_X1 U18271 ( .A(n14947), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14946), 
        .Z(P2_U3610) );
  AND2_X1 U18272 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  AOI21_X1 U18273 ( .B1(n14951), .B2(n15148), .A(n14952), .ZN(n14953) );
  NAND2_X1 U18274 ( .A1(n14953), .A2(n19009), .ZN(n14961) );
  AOI21_X1 U18275 ( .B1(n14955), .B2(n9777), .A(n9990), .ZN(n15370) );
  NAND2_X1 U18276 ( .A1(n15370), .A2(n19002), .ZN(n14957) );
  AOI22_X1 U18277 ( .A1(n18986), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n20694), .ZN(n14956) );
  OAI211_X1 U18278 ( .C1(n18981), .C2(n10018), .A(n14957), .B(n14956), .ZN(
        n14958) );
  AOI21_X1 U18279 ( .B1(n14959), .B2(n20703), .A(n14958), .ZN(n14960) );
  OAI211_X1 U18280 ( .C1(n20705), .C2(n15374), .A(n14961), .B(n14960), .ZN(
        P2_U2827) );
  NOR2_X1 U18281 ( .A1(n15037), .A2(n14963), .ZN(n14964) );
  OR2_X1 U18282 ( .A1(n14962), .A2(n14964), .ZN(n15187) );
  OR2_X1 U18283 ( .A1(n14966), .A2(n14967), .ZN(n14968) );
  NAND2_X1 U18284 ( .A1(n14965), .A2(n14968), .ZN(n15091) );
  OR2_X1 U18285 ( .A1(n20697), .A2(n15183), .ZN(n14970) );
  NAND2_X1 U18286 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n20694), .ZN(n14969) );
  OAI211_X1 U18287 ( .C1(n15091), .C2(n20698), .A(n14970), .B(n14969), .ZN(
        n14971) );
  AOI21_X1 U18288 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19012), .A(
        n14971), .ZN(n14972) );
  OAI21_X1 U18289 ( .B1(n14973), .B2(n19005), .A(n14972), .ZN(n14977) );
  AOI211_X1 U18290 ( .C1(n15184), .C2(n14974), .A(n12836), .B(n14975), .ZN(
        n14976) );
  AOI211_X1 U18291 ( .C1(n15416), .C2(n19007), .A(n14977), .B(n14976), .ZN(
        n14978) );
  INV_X1 U18292 ( .A(n14978), .ZN(P2_U2831) );
  NOR2_X1 U18293 ( .A1(n14980), .A2(n14979), .ZN(n14981) );
  OR2_X1 U18294 ( .A1(n12953), .A2(n14981), .ZN(n16305) );
  AOI211_X1 U18295 ( .C1(n14984), .C2(n14982), .A(n14983), .B(n12836), .ZN(
        n14985) );
  INV_X1 U18296 ( .A(n14985), .ZN(n14994) );
  NOR2_X1 U18297 ( .A1(n15049), .A2(n14986), .ZN(n14987) );
  OR2_X1 U18298 ( .A1(n12956), .A2(n14987), .ZN(n16290) );
  INV_X1 U18299 ( .A(n16290), .ZN(n15484) );
  NAND2_X1 U18300 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n20694), .ZN(n14988) );
  OAI21_X1 U18301 ( .B1(n20697), .B2(n19824), .A(n14988), .ZN(n14989) );
  AOI21_X1 U18302 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19012), .A(
        n14989), .ZN(n14990) );
  OAI21_X1 U18303 ( .B1(n14991), .B2(n19005), .A(n14990), .ZN(n14992) );
  AOI21_X1 U18304 ( .B1(n15484), .B2(n19007), .A(n14992), .ZN(n14993) );
  OAI211_X1 U18305 ( .C1(n16305), .C2(n20698), .A(n14994), .B(n14993), .ZN(
        P2_U2835) );
  NOR2_X1 U18306 ( .A1(n14995), .A2(n14996), .ZN(n15055) );
  INV_X1 U18307 ( .A(n15055), .ZN(n14998) );
  INV_X1 U18308 ( .A(n15054), .ZN(n14997) );
  NAND3_X1 U18309 ( .A1(n14998), .A2(n14997), .A3(n19018), .ZN(n15000) );
  NAND2_X1 U18310 ( .A1(n19052), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14999) );
  OAI211_X1 U18311 ( .C1(n19052), .C2(n15001), .A(n15000), .B(n14999), .ZN(
        P2_U2858) );
  NAND2_X1 U18312 ( .A1(n15003), .A2(n15002), .ZN(n15004) );
  XOR2_X1 U18313 ( .A(n15005), .B(n15004), .Z(n15066) );
  NOR2_X1 U18314 ( .A1(n15374), .A2(n19052), .ZN(n15006) );
  AOI21_X1 U18315 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19052), .A(n15006), .ZN(
        n15007) );
  OAI21_X1 U18316 ( .B1(n15066), .B2(n19041), .A(n15007), .ZN(P2_U2859) );
  OAI21_X1 U18317 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15072) );
  NOR2_X1 U18318 ( .A1(n15386), .A2(n19052), .ZN(n15011) );
  AOI21_X1 U18319 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19052), .A(n15011), .ZN(
        n15012) );
  OAI21_X1 U18320 ( .B1(n15072), .B2(n19041), .A(n15012), .ZN(P2_U2860) );
  AOI21_X1 U18321 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15073) );
  NAND2_X1 U18322 ( .A1(n15073), .A2(n19018), .ZN(n15020) );
  AOI21_X1 U18323 ( .B1(n15018), .B2(n15016), .A(n11591), .ZN(n16243) );
  NAND2_X1 U18324 ( .A1(n16243), .A2(n19048), .ZN(n15019) );
  OAI211_X1 U18325 ( .C1(n19048), .C2(n20956), .A(n15020), .B(n15019), .ZN(
        P2_U2861) );
  OAI21_X1 U18326 ( .B1(n15021), .B2(n15023), .A(n15022), .ZN(n15081) );
  OR2_X1 U18327 ( .A1(n14962), .A2(n15024), .ZN(n15025) );
  NAND2_X1 U18328 ( .A1(n15016), .A2(n15025), .ZN(n16254) );
  MUX2_X1 U18329 ( .A(n16254), .B(n15026), .S(n19052), .Z(n15027) );
  OAI21_X1 U18330 ( .B1(n15081), .B2(n19041), .A(n15027), .ZN(P2_U2862) );
  INV_X1 U18331 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15032) );
  OR2_X1 U18332 ( .A1(n15029), .A2(n15028), .ZN(n15089) );
  NAND3_X1 U18333 ( .A1(n15089), .A2(n19018), .A3(n14420), .ZN(n15031) );
  NAND2_X1 U18334 ( .A1(n15416), .A2(n19048), .ZN(n15030) );
  OAI211_X1 U18335 ( .C1(n19048), .C2(n15032), .A(n15031), .B(n15030), .ZN(
        P2_U2863) );
  OAI21_X1 U18336 ( .B1(n15035), .B2(n15034), .A(n15033), .ZN(n15103) );
  AND2_X1 U18337 ( .A1(n15451), .A2(n15036), .ZN(n15038) );
  OR2_X1 U18338 ( .A1(n15038), .A2(n15037), .ZN(n16267) );
  NOR2_X1 U18339 ( .A1(n16267), .A2(n19052), .ZN(n15039) );
  AOI21_X1 U18340 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n19052), .A(n15039), .ZN(
        n15040) );
  OAI21_X1 U18341 ( .B1(n15103), .B2(n19041), .A(n15040), .ZN(P2_U2864) );
  NAND2_X1 U18342 ( .A1(n15042), .A2(n16285), .ZN(n16287) );
  INV_X1 U18343 ( .A(n16280), .ZN(n15043) );
  AOI21_X1 U18344 ( .B1(n15044), .B2(n16287), .A(n15043), .ZN(n15104) );
  NAND2_X1 U18345 ( .A1(n15104), .A2(n19018), .ZN(n15046) );
  NAND2_X1 U18346 ( .A1(n19052), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15045) );
  OAI211_X1 U18347 ( .C1(n15462), .C2(n19052), .A(n15046), .B(n15045), .ZN(
        P2_U2866) );
  NOR2_X1 U18348 ( .A1(n16294), .A2(n15047), .ZN(n15048) );
  OR2_X1 U18349 ( .A1(n15042), .A2(n15048), .ZN(n15122) );
  NAND2_X1 U18350 ( .A1(n19052), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15053) );
  AOI21_X1 U18351 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n18883) );
  NAND2_X1 U18352 ( .A1(n18883), .A2(n19048), .ZN(n15052) );
  OAI211_X1 U18353 ( .C1(n15122), .C2(n19041), .A(n15053), .B(n15052), .ZN(
        P2_U2868) );
  NOR3_X1 U18354 ( .A1(n15055), .A2(n15054), .A3(n19124), .ZN(n15061) );
  AOI22_X1 U18355 ( .A1(n19061), .A2(BUF1_REG_29__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U18356 ( .A1(n19059), .A2(n15056), .B1(n19119), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15057) );
  OAI211_X1 U18357 ( .C1(n19063), .C2(n15059), .A(n15058), .B(n15057), .ZN(
        n15060) );
  OR2_X1 U18358 ( .A1(n15061), .A2(n15060), .ZN(P2_U2890) );
  INV_X1 U18359 ( .A(n19077), .ZN(n15062) );
  OAI22_X1 U18360 ( .A1(n15115), .A2(n15062), .B1(n19095), .B2(n13059), .ZN(
        n15063) );
  AOI21_X1 U18361 ( .B1(n15370), .B2(n19120), .A(n15063), .ZN(n15065) );
  AOI22_X1 U18362 ( .A1(n19061), .A2(BUF1_REG_28__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15064) );
  OAI211_X1 U18363 ( .C1(n15066), .C2(n19124), .A(n15065), .B(n15064), .ZN(
        P2_U2891) );
  AOI22_X1 U18364 ( .A1(n19061), .A2(BUF1_REG_27__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U18365 ( .A1(n19059), .A2(n15067), .B1(n19119), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15068) );
  OAI211_X1 U18366 ( .C1(n19063), .C2(n15385), .A(n15069), .B(n15068), .ZN(
        n15070) );
  INV_X1 U18367 ( .A(n15070), .ZN(n15071) );
  OAI21_X1 U18368 ( .B1(n15072), .B2(n19124), .A(n15071), .ZN(P2_U2892) );
  NAND2_X1 U18369 ( .A1(n15073), .A2(n19106), .ZN(n15080) );
  AOI22_X1 U18370 ( .A1(n19059), .A2(n19082), .B1(n19119), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U18371 ( .A1(n19061), .A2(BUF1_REG_26__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15078) );
  OR2_X1 U18372 ( .A1(n15075), .A2(n15074), .ZN(n15076) );
  AND2_X1 U18373 ( .A1(n12943), .A2(n15076), .ZN(n16251) );
  NAND2_X1 U18374 ( .A1(n19120), .A2(n16251), .ZN(n15077) );
  NAND4_X1 U18375 ( .A1(n15080), .A2(n15079), .A3(n15078), .A4(n15077), .ZN(
        P2_U2893) );
  OR2_X1 U18376 ( .A1(n15081), .A2(n19124), .ZN(n15088) );
  AOI22_X1 U18377 ( .A1(n19059), .A2(n19085), .B1(n19119), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U18378 ( .A1(n19061), .A2(BUF1_REG_25__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15086) );
  INV_X1 U18379 ( .A(n15082), .ZN(n15083) );
  XNOR2_X1 U18380 ( .A(n14965), .B(n15083), .ZN(n16255) );
  INV_X1 U18381 ( .A(n16255), .ZN(n15084) );
  OR2_X1 U18382 ( .A1(n19063), .A2(n15084), .ZN(n15085) );
  NAND4_X1 U18383 ( .A1(n15088), .A2(n15087), .A3(n15086), .A4(n15085), .ZN(
        P2_U2894) );
  NAND3_X1 U18384 ( .A1(n15089), .A2(n19106), .A3(n14420), .ZN(n15095) );
  AOI22_X1 U18385 ( .A1(n19059), .A2(n15090), .B1(n19119), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U18386 ( .A1(n19061), .A2(BUF1_REG_24__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15093) );
  INV_X1 U18387 ( .A(n15091), .ZN(n15419) );
  NAND2_X1 U18388 ( .A1(n19120), .A2(n15419), .ZN(n15092) );
  NAND4_X1 U18389 ( .A1(n15095), .A2(n15094), .A3(n15093), .A4(n15092), .ZN(
        P2_U2895) );
  NOR2_X1 U18390 ( .A1(n15097), .A2(n15096), .ZN(n15098) );
  OR2_X1 U18391 ( .A1(n14966), .A2(n15098), .ZN(n16266) );
  AOI22_X1 U18392 ( .A1(n19061), .A2(BUF1_REG_23__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U18393 ( .A1(n19059), .A2(n19220), .B1(n19119), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15099) );
  OAI211_X1 U18394 ( .C1(n19063), .C2(n16266), .A(n15100), .B(n15099), .ZN(
        n15101) );
  INV_X1 U18395 ( .A(n15101), .ZN(n15102) );
  OAI21_X1 U18396 ( .B1(n15103), .B2(n19124), .A(n15102), .ZN(P2_U2896) );
  NAND2_X1 U18397 ( .A1(n15104), .A2(n19106), .ZN(n15111) );
  OAI22_X1 U18398 ( .A1(n15115), .A2(n15106), .B1(n15105), .B2(n19095), .ZN(
        n15109) );
  INV_X1 U18399 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15107) );
  NOR2_X1 U18400 ( .A1(n15119), .A2(n15107), .ZN(n15108) );
  AOI211_X1 U18401 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n19061), .A(n15109), .B(
        n15108), .ZN(n15110) );
  OAI211_X1 U18402 ( .C1(n15467), .C2(n19063), .A(n15111), .B(n15110), .ZN(
        P2_U2898) );
  XNOR2_X1 U18403 ( .A(n15113), .B(n15112), .ZN(n15494) );
  INV_X1 U18404 ( .A(n15494), .ZN(n18884) );
  INV_X1 U18405 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15118) );
  OAI22_X1 U18406 ( .A1(n15115), .A2(n19118), .B1(n15114), .B2(n19095), .ZN(
        n15116) );
  AOI21_X1 U18407 ( .B1(n19061), .B2(BUF1_REG_19__SCAN_IN), .A(n15116), .ZN(
        n15117) );
  OAI21_X1 U18408 ( .B1(n15119), .B2(n15118), .A(n15117), .ZN(n15120) );
  AOI21_X1 U18409 ( .B1(n18884), .B2(n19120), .A(n15120), .ZN(n15121) );
  OAI21_X1 U18410 ( .B1(n19124), .B2(n15122), .A(n15121), .ZN(P2_U2900) );
  XNOR2_X1 U18411 ( .A(n15123), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15365) );
  NAND2_X1 U18412 ( .A1(n15125), .A2(n15124), .ZN(n15130) );
  INV_X1 U18413 ( .A(n15126), .ZN(n15128) );
  NAND2_X1 U18414 ( .A1(n15128), .A2(n15127), .ZN(n15129) );
  XNOR2_X1 U18415 ( .A(n15130), .B(n15129), .ZN(n15363) );
  NOR2_X1 U18416 ( .A1(n18970), .A2(n15131), .ZN(n15352) );
  NOR2_X1 U18417 ( .A1(n19172), .A2(n15132), .ZN(n15133) );
  AOI211_X1 U18418 ( .C1(n16322), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15352), .B(n15133), .ZN(n15134) );
  OAI21_X1 U18419 ( .B1(n15361), .B2(n15652), .A(n15134), .ZN(n15135) );
  AOI21_X1 U18420 ( .B1(n15363), .B2(n16346), .A(n15135), .ZN(n15136) );
  OAI21_X1 U18421 ( .B1(n15365), .B2(n19173), .A(n15136), .ZN(P2_U2984) );
  OAI21_X1 U18422 ( .B1(n15138), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15137), .ZN(n15378) );
  INV_X1 U18423 ( .A(n15139), .ZN(n15141) );
  AOI22_X1 U18424 ( .A1(n15142), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n15141), .B2(n15140), .ZN(n15145) );
  XOR2_X1 U18425 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15143), .Z(
        n15144) );
  XNOR2_X1 U18426 ( .A(n15145), .B(n15144), .ZN(n15376) );
  NOR2_X1 U18427 ( .A1(n18970), .A2(n15146), .ZN(n15369) );
  NOR2_X1 U18428 ( .A1(n19184), .A2(n10018), .ZN(n15147) );
  AOI211_X1 U18429 ( .C1(n15148), .C2(n16343), .A(n15369), .B(n15147), .ZN(
        n15149) );
  OAI21_X1 U18430 ( .B1(n15374), .B2(n15652), .A(n15149), .ZN(n15150) );
  AOI21_X1 U18431 ( .B1(n15376), .B2(n16346), .A(n15150), .ZN(n15151) );
  OAI21_X1 U18432 ( .B1(n15378), .B2(n19173), .A(n15151), .ZN(P2_U2986) );
  BUF_X1 U18433 ( .A(n15152), .Z(n15153) );
  OAI21_X1 U18434 ( .B1(n15153), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14278), .ZN(n15403) );
  OAI21_X1 U18435 ( .B1(n15154), .B2(n15164), .A(n15165), .ZN(n15155) );
  XNOR2_X1 U18436 ( .A(n15156), .B(n15155), .ZN(n15401) );
  NAND2_X1 U18437 ( .A1(n16243), .A2(n19176), .ZN(n15158) );
  NOR2_X1 U18438 ( .A1(n18933), .A2(n19833), .ZN(n15396) );
  AOI21_X1 U18439 ( .B1(n16322), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15396), .ZN(n15157) );
  OAI211_X1 U18440 ( .C1(n19172), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15160) );
  AOI21_X1 U18441 ( .B1(n15401), .B2(n16346), .A(n15160), .ZN(n15161) );
  OAI21_X1 U18442 ( .B1(n15403), .B2(n19173), .A(n15161), .ZN(P2_U2988) );
  INV_X1 U18443 ( .A(n15153), .ZN(n15163) );
  OAI21_X1 U18444 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15162), .A(
        n15163), .ZN(n15414) );
  INV_X1 U18445 ( .A(n15164), .ZN(n15166) );
  NAND2_X1 U18446 ( .A1(n15166), .A2(n15165), .ZN(n15167) );
  XOR2_X1 U18447 ( .A(n15167), .B(n15154), .Z(n15412) );
  NAND2_X1 U18448 ( .A1(n18985), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15404) );
  OAI21_X1 U18449 ( .B1(n19184), .B2(n15168), .A(n15404), .ZN(n15169) );
  AOI21_X1 U18450 ( .B1(n16343), .B2(n16259), .A(n15169), .ZN(n15170) );
  OAI21_X1 U18451 ( .B1(n16254), .B2(n15652), .A(n15170), .ZN(n15171) );
  AOI21_X1 U18452 ( .B1(n15412), .B2(n16346), .A(n15171), .ZN(n15172) );
  OAI21_X1 U18453 ( .B1(n15414), .B2(n19173), .A(n15172), .ZN(P2_U2989) );
  INV_X1 U18454 ( .A(n15162), .ZN(n15174) );
  OAI21_X1 U18455 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15173), .A(
        n15174), .ZN(n15427) );
  NAND2_X1 U18456 ( .A1(n15175), .A2(n15447), .ZN(n15193) );
  XNOR2_X1 U18457 ( .A(n15177), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15192) );
  NAND2_X1 U18458 ( .A1(n15193), .A2(n15192), .ZN(n15435) );
  OAI21_X1 U18459 ( .B1(n15177), .B2(n15176), .A(n15435), .ZN(n15182) );
  INV_X1 U18460 ( .A(n15178), .ZN(n15180) );
  NAND2_X1 U18461 ( .A1(n15180), .A2(n15179), .ZN(n15181) );
  XNOR2_X1 U18462 ( .A(n15182), .B(n15181), .ZN(n15425) );
  NOR2_X1 U18463 ( .A1(n18933), .A2(n15183), .ZN(n15418) );
  AOI21_X1 U18464 ( .B1(n16322), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15418), .ZN(n15186) );
  NAND2_X1 U18465 ( .A1(n16343), .A2(n15184), .ZN(n15185) );
  OAI211_X1 U18466 ( .C1(n15187), .C2(n15652), .A(n15186), .B(n15185), .ZN(
        n15188) );
  AOI21_X1 U18467 ( .B1(n15425), .B2(n16346), .A(n15188), .ZN(n15189) );
  OAI21_X1 U18468 ( .B1(n15427), .B2(n19173), .A(n15189), .ZN(P2_U2990) );
  INV_X1 U18469 ( .A(n15173), .ZN(n15191) );
  OAI21_X1 U18470 ( .B1(n15443), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15191), .ZN(n15442) );
  NOR2_X1 U18471 ( .A1(n15193), .A2(n15192), .ZN(n15437) );
  NOR2_X1 U18472 ( .A1(n15437), .A2(n19179), .ZN(n15197) );
  OAI22_X1 U18473 ( .A1(n19184), .A2(n10833), .B1(n10792), .B2(n18970), .ZN(
        n15194) );
  AOI21_X1 U18474 ( .B1(n16343), .B2(n16271), .A(n15194), .ZN(n15195) );
  OAI21_X1 U18475 ( .B1(n16267), .B2(n15652), .A(n15195), .ZN(n15196) );
  AOI21_X1 U18476 ( .B1(n15197), .B2(n15435), .A(n15196), .ZN(n15198) );
  OAI21_X1 U18477 ( .B1(n15442), .B2(n19173), .A(n15198), .ZN(P2_U2991) );
  OAI21_X1 U18478 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15243) );
  NAND2_X1 U18479 ( .A1(n15243), .A2(n15202), .ZN(n15220) );
  NAND3_X1 U18480 ( .A1(n15220), .A2(n15219), .A3(n15218), .ZN(n15203) );
  NAND2_X1 U18481 ( .A1(n15203), .A2(n15217), .ZN(n15207) );
  NOR2_X1 U18482 ( .A1(n15204), .A2(n10861), .ZN(n15205) );
  XNOR2_X1 U18483 ( .A(n15205), .B(n15465), .ZN(n15206) );
  XNOR2_X1 U18484 ( .A(n15207), .B(n15206), .ZN(n15474) );
  NAND2_X1 U18485 ( .A1(n18985), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15463) );
  OAI21_X1 U18486 ( .B1(n19184), .B2(n15208), .A(n15463), .ZN(n15210) );
  NOR2_X1 U18487 ( .A1(n15462), .A2(n15652), .ZN(n15209) );
  AOI211_X1 U18488 ( .C1(n16343), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15215) );
  OR2_X1 U18489 ( .A1(n15212), .A2(n15475), .ZN(n15216) );
  INV_X1 U18490 ( .A(n15190), .ZN(n15213) );
  AOI21_X1 U18491 ( .B1(n15465), .B2(n15216), .A(n15213), .ZN(n15471) );
  NAND2_X1 U18492 ( .A1(n15471), .A2(n10876), .ZN(n15214) );
  OAI211_X1 U18493 ( .C1(n15474), .C2(n19179), .A(n15215), .B(n15214), .ZN(
        P2_U2993) );
  OAI21_X1 U18494 ( .B1(n10113), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15216), .ZN(n15489) );
  NAND2_X1 U18495 ( .A1(n15218), .A2(n15217), .ZN(n15222) );
  NAND2_X1 U18496 ( .A1(n15220), .A2(n15219), .ZN(n15221) );
  XOR2_X1 U18497 ( .A(n15222), .B(n15221), .Z(n15487) );
  NOR2_X1 U18498 ( .A1(n18933), .A2(n19824), .ZN(n15479) );
  NOR2_X1 U18499 ( .A1(n19172), .A2(n15223), .ZN(n15224) );
  AOI211_X1 U18500 ( .C1(n16322), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15479), .B(n15224), .ZN(n15225) );
  OAI21_X1 U18501 ( .B1(n16290), .B2(n15652), .A(n15225), .ZN(n15226) );
  AOI21_X1 U18502 ( .B1(n15487), .B2(n16346), .A(n15226), .ZN(n15227) );
  OAI21_X1 U18503 ( .B1(n19173), .B2(n15489), .A(n15227), .ZN(P2_U2994) );
  NAND2_X1 U18504 ( .A1(n15229), .A2(n15228), .ZN(n15232) );
  INV_X1 U18505 ( .A(n15242), .ZN(n15230) );
  AOI21_X1 U18506 ( .B1(n15243), .B2(n15241), .A(n15230), .ZN(n15231) );
  XOR2_X1 U18507 ( .A(n15232), .B(n15231), .Z(n15500) );
  NAND2_X1 U18508 ( .A1(n18886), .A2(n16343), .ZN(n15233) );
  NAND2_X1 U18509 ( .A1(n18985), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15491) );
  OAI211_X1 U18510 ( .C1(n19184), .C2(n15234), .A(n15233), .B(n15491), .ZN(
        n15235) );
  AOI21_X1 U18511 ( .B1(n18883), .B2(n19176), .A(n15235), .ZN(n15238) );
  AOI21_X1 U18512 ( .B1(n15236), .B2(n15212), .A(n10113), .ZN(n15497) );
  NAND2_X1 U18513 ( .A1(n15497), .A2(n10876), .ZN(n15237) );
  OAI211_X1 U18514 ( .C1(n15500), .C2(n19179), .A(n15238), .B(n15237), .ZN(
        P2_U2995) );
  INV_X1 U18515 ( .A(n15239), .ZN(n15240) );
  OAI21_X1 U18516 ( .B1(n15240), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15212), .ZN(n15510) );
  NAND2_X1 U18517 ( .A1(n15242), .A2(n15241), .ZN(n15244) );
  XOR2_X1 U18518 ( .A(n15244), .B(n15243), .Z(n15501) );
  OR2_X1 U18519 ( .A1(n18970), .A2(n15245), .ZN(n15502) );
  OAI21_X1 U18520 ( .B1(n19184), .B2(n15246), .A(n15502), .ZN(n15247) );
  AOI21_X1 U18521 ( .B1(n15248), .B2(n16343), .A(n15247), .ZN(n15249) );
  OAI21_X1 U18522 ( .B1(n16296), .B2(n15652), .A(n15249), .ZN(n15250) );
  AOI21_X1 U18523 ( .B1(n15501), .B2(n16346), .A(n15250), .ZN(n15251) );
  OAI21_X1 U18524 ( .B1(n19173), .B2(n15510), .A(n15251), .ZN(P2_U2996) );
  INV_X1 U18525 ( .A(n15252), .ZN(n15259) );
  OAI211_X1 U18526 ( .C1(n10119), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10876), .B(n15239), .ZN(n15258) );
  INV_X1 U18527 ( .A(n15253), .ZN(n18899) );
  NAND2_X1 U18528 ( .A1(n16322), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15254) );
  OAI211_X1 U18529 ( .C1(n18901), .C2(n19172), .A(n15255), .B(n15254), .ZN(
        n15256) );
  AOI21_X1 U18530 ( .B1(n18899), .B2(n19176), .A(n15256), .ZN(n15257) );
  OAI211_X1 U18531 ( .C1(n15259), .C2(n19179), .A(n15258), .B(n15257), .ZN(
        P2_U2997) );
  INV_X1 U18532 ( .A(n15260), .ZN(n15270) );
  OAI21_X1 U18533 ( .B1(n15286), .B2(n15515), .A(n15261), .ZN(n15262) );
  NAND3_X1 U18534 ( .A1(n9868), .A2(n10876), .A3(n15262), .ZN(n15269) );
  NAND2_X1 U18535 ( .A1(n16322), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15263) );
  OAI211_X1 U18536 ( .C1(n15265), .C2(n19172), .A(n15264), .B(n15263), .ZN(
        n15266) );
  AOI21_X1 U18537 ( .B1(n15267), .B2(n19176), .A(n15266), .ZN(n15268) );
  OAI211_X1 U18538 ( .C1(n15270), .C2(n19179), .A(n15269), .B(n15268), .ZN(
        P2_U2998) );
  XNOR2_X1 U18539 ( .A(n15286), .B(n15515), .ZN(n15523) );
  NAND2_X1 U18540 ( .A1(n15272), .A2(n15271), .ZN(n15276) );
  INV_X1 U18541 ( .A(n15283), .ZN(n15273) );
  NOR2_X1 U18542 ( .A1(n15274), .A2(n15273), .ZN(n15275) );
  XOR2_X1 U18543 ( .A(n15276), .B(n15275), .Z(n15521) );
  NOR2_X1 U18544 ( .A1(n18933), .A2(n19817), .ZN(n15513) );
  AOI21_X1 U18545 ( .B1(n16322), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15513), .ZN(n15279) );
  NAND2_X1 U18546 ( .A1(n15277), .A2(n16343), .ZN(n15278) );
  OAI211_X1 U18547 ( .C1(n18912), .C2(n15652), .A(n15279), .B(n15278), .ZN(
        n15280) );
  AOI21_X1 U18548 ( .B1(n15521), .B2(n16346), .A(n15280), .ZN(n15281) );
  OAI21_X1 U18549 ( .B1(n15523), .B2(n19173), .A(n15281), .ZN(P2_U2999) );
  NAND2_X1 U18550 ( .A1(n15283), .A2(n15282), .ZN(n15284) );
  XNOR2_X1 U18551 ( .A(n15285), .B(n15284), .ZN(n15535) );
  AOI21_X1 U18552 ( .B1(n15529), .B2(n9780), .A(n14253), .ZN(n15524) );
  NAND2_X1 U18553 ( .A1(n15524), .A2(n10876), .ZN(n15292) );
  NAND2_X1 U18554 ( .A1(n18985), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n15527) );
  OAI21_X1 U18555 ( .B1(n19184), .B2(n15287), .A(n15527), .ZN(n15289) );
  NOR2_X1 U18556 ( .A1(n19030), .A2(n15652), .ZN(n15288) );
  AOI211_X1 U18557 ( .C1(n16343), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        n15291) );
  OAI211_X1 U18558 ( .C1(n19179), .C2(n15535), .A(n15292), .B(n15291), .ZN(
        P2_U3000) );
  NAND2_X1 U18559 ( .A1(n15293), .A2(n9780), .ZN(n15548) );
  NAND2_X1 U18560 ( .A1(n15296), .A2(n15295), .ZN(n15297) );
  XNOR2_X1 U18561 ( .A(n15294), .B(n15297), .ZN(n15546) );
  NOR2_X1 U18562 ( .A1(n18933), .A2(n15298), .ZN(n15540) );
  NOR2_X1 U18563 ( .A1(n19172), .A2(n18928), .ZN(n15299) );
  AOI211_X1 U18564 ( .C1(n16322), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15540), .B(n15299), .ZN(n15300) );
  OAI21_X1 U18565 ( .B1(n18918), .B2(n15652), .A(n15300), .ZN(n15301) );
  AOI21_X1 U18566 ( .B1(n15546), .B2(n16346), .A(n15301), .ZN(n15302) );
  OAI21_X1 U18567 ( .B1(n15548), .B2(n19173), .A(n15302), .ZN(P2_U3001) );
  NAND2_X1 U18568 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  XNOR2_X1 U18569 ( .A(n9732), .B(n15306), .ZN(n15557) );
  AOI22_X1 U18570 ( .A1(n16322), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18985), .ZN(n15309) );
  NAND2_X1 U18571 ( .A1(n16343), .A2(n15307), .ZN(n15308) );
  OAI211_X1 U18572 ( .C1(n15555), .C2(n15652), .A(n15309), .B(n15308), .ZN(
        n15310) );
  AOI21_X1 U18573 ( .B1(n15557), .B2(n16346), .A(n15310), .ZN(n15311) );
  OAI21_X1 U18574 ( .B1(n15559), .B2(n19173), .A(n15311), .ZN(P2_U3002) );
  NOR2_X1 U18575 ( .A1(n15312), .A2(n15594), .ZN(n15584) );
  NAND2_X1 U18576 ( .A1(n15314), .A2(n15313), .ZN(n15334) );
  INV_X1 U18577 ( .A(n15315), .ZN(n15332) );
  NOR2_X1 U18578 ( .A1(n15334), .A2(n15332), .ZN(n15581) );
  INV_X1 U18579 ( .A(n15581), .ZN(n15318) );
  INV_X1 U18580 ( .A(n15316), .ZN(n15579) );
  OAI21_X1 U18581 ( .B1(n15318), .B2(n15579), .A(n15317), .ZN(n15322) );
  NAND2_X1 U18582 ( .A1(n15320), .A2(n15319), .ZN(n15321) );
  XNOR2_X1 U18583 ( .A(n15322), .B(n15321), .ZN(n15575) );
  NOR2_X1 U18584 ( .A1(n18933), .A2(n19811), .ZN(n15570) );
  NOR2_X1 U18585 ( .A1(n19184), .A2(n15323), .ZN(n15324) );
  AOI211_X1 U18586 ( .C1(n15325), .C2(n16343), .A(n15570), .B(n15324), .ZN(
        n15326) );
  OAI21_X1 U18587 ( .B1(n18932), .B2(n15652), .A(n15326), .ZN(n15327) );
  AOI21_X1 U18588 ( .B1(n15575), .B2(n16346), .A(n15327), .ZN(n15328) );
  OAI21_X1 U18589 ( .B1(n15577), .B2(n19173), .A(n15328), .ZN(P2_U3003) );
  NOR2_X1 U18590 ( .A1(n18933), .A2(n15329), .ZN(n15602) );
  INV_X1 U18591 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15330) );
  OAI22_X1 U18592 ( .A1(n19184), .A2(n15330), .B1(n19172), .B2(n18961), .ZN(
        n15331) );
  AOI211_X1 U18593 ( .C1(n18964), .C2(n19176), .A(n15602), .B(n15331), .ZN(
        n15337) );
  NOR2_X1 U18594 ( .A1(n15580), .A2(n15332), .ZN(n15333) );
  XNOR2_X1 U18595 ( .A(n15334), .B(n15333), .ZN(n15609) );
  NAND2_X1 U18596 ( .A1(n15609), .A2(n15335), .ZN(n15336) );
  OAI211_X1 U18597 ( .C1(n15612), .C2(n19173), .A(n15337), .B(n15336), .ZN(
        P2_U3005) );
  OR2_X1 U18598 ( .A1(n9717), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15613) );
  NAND3_X1 U18599 ( .A1(n15613), .A2(n15339), .A3(n10876), .ZN(n15351) );
  NAND2_X1 U18600 ( .A1(n15340), .A2(n15341), .ZN(n16331) );
  INV_X1 U18601 ( .A(n16330), .ZN(n15343) );
  AND2_X1 U18602 ( .A1(n16330), .A2(n15341), .ZN(n15342) );
  OAI22_X1 U18603 ( .A1(n16331), .A2(n15343), .B1(n15342), .B2(n15340), .ZN(
        n15624) );
  NOR2_X1 U18604 ( .A1(n15624), .A2(n19179), .ZN(n15349) );
  NOR2_X1 U18605 ( .A1(n15615), .A2(n15652), .ZN(n15348) );
  INV_X1 U18606 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15345) );
  OAI22_X1 U18607 ( .A1(n19184), .A2(n15345), .B1(n19172), .B2(n15344), .ZN(
        n15347) );
  NAND2_X1 U18608 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n18985), .ZN(n15617) );
  INV_X1 U18609 ( .A(n15617), .ZN(n15346) );
  NOR4_X1 U18610 ( .A1(n15349), .A2(n15348), .A3(n15347), .A4(n15346), .ZN(
        n15350) );
  NAND2_X1 U18611 ( .A1(n15351), .A2(n15350), .ZN(P2_U3007) );
  INV_X1 U18612 ( .A(n16354), .ZN(n15355) );
  INV_X1 U18613 ( .A(n15352), .ZN(n15354) );
  INV_X1 U18614 ( .A(n15357), .ZN(n15360) );
  NAND2_X1 U18615 ( .A1(n15358), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15359) );
  OAI211_X1 U18616 ( .C1(n15361), .C2(n15614), .A(n15360), .B(n15359), .ZN(
        n15362) );
  AOI21_X1 U18617 ( .B1(n15363), .B2(n16359), .A(n15362), .ZN(n15364) );
  OAI21_X1 U18618 ( .B1(n15365), .B2(n15629), .A(n15364), .ZN(P2_U3016) );
  NOR3_X1 U18619 ( .A1(n15367), .A2(n15382), .A3(n15366), .ZN(n15368) );
  AOI211_X1 U18620 ( .C1(n15370), .C2(n16354), .A(n15369), .B(n15368), .ZN(
        n15373) );
  NAND2_X1 U18621 ( .A1(n15371), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15372) );
  OAI211_X1 U18622 ( .C1(n15374), .C2(n15614), .A(n15373), .B(n15372), .ZN(
        n15375) );
  AOI21_X1 U18623 ( .B1(n15376), .B2(n16359), .A(n15375), .ZN(n15377) );
  OAI21_X1 U18624 ( .B1(n15378), .B2(n15629), .A(n15377), .ZN(P2_U3018) );
  NAND3_X1 U18625 ( .A1(n15380), .A2(n16357), .A3(n15379), .ZN(n15391) );
  AOI21_X1 U18626 ( .B1(n15383), .B2(n15382), .A(n15381), .ZN(n15384) );
  OAI21_X1 U18627 ( .B1(n15355), .B2(n15385), .A(n15384), .ZN(n15388) );
  NOR2_X1 U18628 ( .A1(n15386), .A2(n15614), .ZN(n15387) );
  AOI211_X1 U18629 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15389), .A(
        n15388), .B(n15387), .ZN(n15390) );
  OAI211_X1 U18630 ( .C1(n15392), .C2(n15623), .A(n15391), .B(n15390), .ZN(
        P2_U3019) );
  NAND2_X1 U18631 ( .A1(n16243), .A2(n12862), .ZN(n15398) );
  INV_X1 U18632 ( .A(n15393), .ZN(n15405) );
  AOI211_X1 U18633 ( .C1(n15399), .C2(n15406), .A(n15394), .B(n15405), .ZN(
        n15395) );
  AOI211_X1 U18634 ( .C1(n16354), .C2(n16251), .A(n15396), .B(n15395), .ZN(
        n15397) );
  OAI211_X1 U18635 ( .C1(n15407), .C2(n15399), .A(n15398), .B(n15397), .ZN(
        n15400) );
  AOI21_X1 U18636 ( .B1(n15401), .B2(n16359), .A(n15400), .ZN(n15402) );
  OAI21_X1 U18637 ( .B1(n15403), .B2(n15629), .A(n15402), .ZN(P2_U3020) );
  OAI21_X1 U18638 ( .B1(n15405), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15404), .ZN(n15409) );
  NOR2_X1 U18639 ( .A1(n15407), .A2(n15406), .ZN(n15408) );
  AOI211_X1 U18640 ( .C1(n16354), .C2(n16255), .A(n15409), .B(n15408), .ZN(
        n15410) );
  OAI21_X1 U18641 ( .B1(n16254), .B2(n15614), .A(n15410), .ZN(n15411) );
  AOI21_X1 U18642 ( .B1(n15412), .B2(n16359), .A(n15411), .ZN(n15413) );
  OAI21_X1 U18643 ( .B1(n15414), .B2(n15629), .A(n15413), .ZN(P2_U3021) );
  AOI21_X1 U18644 ( .B1(n15430), .B2(n15415), .A(n15457), .ZN(n15423) );
  NAND2_X1 U18645 ( .A1(n15416), .A2(n12862), .ZN(n15421) );
  NOR3_X1 U18646 ( .A1(n15430), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15455), .ZN(n15417) );
  AOI211_X1 U18647 ( .C1(n16354), .C2(n15419), .A(n15418), .B(n15417), .ZN(
        n15420) );
  OAI211_X1 U18648 ( .C1(n15423), .C2(n15422), .A(n15421), .B(n15420), .ZN(
        n15424) );
  AOI21_X1 U18649 ( .B1(n15425), .B2(n16359), .A(n15424), .ZN(n15426) );
  OAI21_X1 U18650 ( .B1(n15427), .B2(n15629), .A(n15426), .ZN(P2_U3022) );
  INV_X1 U18651 ( .A(n16267), .ZN(n15440) );
  NAND2_X1 U18652 ( .A1(n15457), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15434) );
  INV_X1 U18653 ( .A(n16266), .ZN(n15428) );
  NAND2_X1 U18654 ( .A1(n16354), .A2(n15428), .ZN(n15433) );
  OR2_X1 U18655 ( .A1(n10792), .A2(n18970), .ZN(n15432) );
  OAI211_X1 U18656 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15430), .B(n15429), .ZN(
        n15431) );
  NAND4_X1 U18657 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15439) );
  INV_X1 U18658 ( .A(n15435), .ZN(n15436) );
  NOR3_X1 U18659 ( .A1(n15437), .A2(n15436), .A3(n15623), .ZN(n15438) );
  AOI211_X1 U18660 ( .C1(n15440), .C2(n12862), .A(n15439), .B(n15438), .ZN(
        n15441) );
  OAI21_X1 U18661 ( .B1(n15629), .B2(n15442), .A(n15441), .ZN(P2_U3023) );
  AOI21_X1 U18662 ( .B1(n20823), .B2(n15190), .A(n15443), .ZN(n16316) );
  INV_X1 U18663 ( .A(n16316), .ZN(n15461) );
  NAND2_X1 U18664 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  XNOR2_X1 U18665 ( .A(n15445), .B(n15448), .ZN(n16318) );
  NAND2_X1 U18666 ( .A1(n12955), .A2(n15449), .ZN(n15450) );
  NAND2_X1 U18667 ( .A1(n15451), .A2(n15450), .ZN(n16315) );
  AOI21_X1 U18668 ( .B1(n15452), .B2(n9776), .A(n15096), .ZN(n15782) );
  NAND2_X1 U18669 ( .A1(n16354), .A2(n15782), .ZN(n15454) );
  NAND2_X1 U18670 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18985), .ZN(n15453) );
  OAI211_X1 U18671 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15455), .A(
        n15454), .B(n15453), .ZN(n15456) );
  AOI21_X1 U18672 ( .B1(n15457), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15456), .ZN(n15458) );
  OAI21_X1 U18673 ( .B1(n16315), .B2(n15614), .A(n15458), .ZN(n15459) );
  AOI21_X1 U18674 ( .B1(n16318), .B2(n16359), .A(n15459), .ZN(n15460) );
  OAI21_X1 U18675 ( .B1(n15461), .B2(n15629), .A(n15460), .ZN(P2_U3024) );
  INV_X1 U18676 ( .A(n15462), .ZN(n15470) );
  OAI211_X1 U18677 ( .C1(n15466), .C2(n15465), .A(n15464), .B(n15463), .ZN(
        n15469) );
  NOR2_X1 U18678 ( .A1(n15467), .A2(n15355), .ZN(n15468) );
  AOI211_X1 U18679 ( .C1(n15470), .C2(n12862), .A(n15469), .B(n15468), .ZN(
        n15473) );
  NAND2_X1 U18680 ( .A1(n15471), .A2(n16357), .ZN(n15472) );
  OAI211_X1 U18681 ( .C1(n15474), .C2(n15623), .A(n15473), .B(n15472), .ZN(
        P2_U3025) );
  OAI21_X1 U18682 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15475), .ZN(n15482) );
  OR2_X1 U18683 ( .A1(n15476), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15503) );
  NOR2_X1 U18684 ( .A1(n15626), .A2(n15477), .ZN(n15478) );
  NOR2_X1 U18685 ( .A1(n15514), .A2(n15478), .ZN(n15505) );
  NAND2_X1 U18686 ( .A1(n15503), .A2(n15505), .ZN(n15490) );
  NAND2_X1 U18687 ( .A1(n15490), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15481) );
  INV_X1 U18688 ( .A(n15479), .ZN(n15480) );
  OAI211_X1 U18689 ( .C1(n15482), .C2(n15493), .A(n15481), .B(n15480), .ZN(
        n15483) );
  AOI21_X1 U18690 ( .B1(n15484), .B2(n12862), .A(n15483), .ZN(n15485) );
  OAI21_X1 U18691 ( .B1(n16305), .B2(n15355), .A(n15485), .ZN(n15486) );
  AOI21_X1 U18692 ( .B1(n15487), .B2(n16359), .A(n15486), .ZN(n15488) );
  OAI21_X1 U18693 ( .B1(n15629), .B2(n15489), .A(n15488), .ZN(P2_U3026) );
  NAND2_X1 U18694 ( .A1(n15490), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15492) );
  OAI211_X1 U18695 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15493), .A(
        n15492), .B(n15491), .ZN(n15496) );
  NOR2_X1 U18696 ( .A1(n15494), .A2(n15355), .ZN(n15495) );
  AOI211_X1 U18697 ( .C1(n18883), .C2(n12862), .A(n15496), .B(n15495), .ZN(
        n15499) );
  NAND2_X1 U18698 ( .A1(n15497), .A2(n16357), .ZN(n15498) );
  OAI211_X1 U18699 ( .C1(n15500), .C2(n15623), .A(n15499), .B(n15498), .ZN(
        P2_U3027) );
  NAND2_X1 U18700 ( .A1(n15501), .A2(n16359), .ZN(n15509) );
  NOR2_X1 U18701 ( .A1(n16296), .A2(n15614), .ZN(n15507) );
  OAI211_X1 U18702 ( .C1(n15505), .C2(n15504), .A(n15503), .B(n15502), .ZN(
        n15506) );
  AOI211_X1 U18703 ( .C1(n16311), .C2(n16354), .A(n15507), .B(n15506), .ZN(
        n15508) );
  OAI211_X1 U18704 ( .C1(n15510), .C2(n15629), .A(n15509), .B(n15508), .ZN(
        P2_U3028) );
  INV_X1 U18705 ( .A(n14132), .ZN(n15511) );
  OAI21_X1 U18706 ( .B1(n13821), .B2(n15512), .A(n15511), .ZN(n19069) );
  NOR2_X1 U18707 ( .A1(n19069), .A2(n15355), .ZN(n15520) );
  AOI21_X1 U18708 ( .B1(n15514), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15513), .ZN(n15518) );
  NAND2_X1 U18709 ( .A1(n15516), .A2(n15515), .ZN(n15517) );
  OAI211_X1 U18710 ( .C1(n18912), .C2(n15614), .A(n15518), .B(n15517), .ZN(
        n15519) );
  AOI211_X1 U18711 ( .C1(n15521), .C2(n16359), .A(n15520), .B(n15519), .ZN(
        n15522) );
  OAI21_X1 U18712 ( .B1(n15523), .B2(n15629), .A(n15522), .ZN(P2_U3031) );
  NAND2_X1 U18713 ( .A1(n15524), .A2(n16357), .ZN(n15534) );
  INV_X1 U18714 ( .A(n19073), .ZN(n15532) );
  NOR2_X1 U18715 ( .A1(n19030), .A2(n15614), .ZN(n15531) );
  INV_X1 U18716 ( .A(n15607), .ZN(n15563) );
  NAND2_X1 U18717 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15568), .ZN(
        n15525) );
  OAI21_X1 U18718 ( .B1(n15563), .B2(n15525), .A(n15599), .ZN(n15552) );
  INV_X1 U18719 ( .A(n15567), .ZN(n15592) );
  XNOR2_X1 U18720 ( .A(n15539), .B(n15529), .ZN(n15526) );
  NAND3_X1 U18721 ( .A1(n15592), .A2(n15568), .A3(n15526), .ZN(n15528) );
  OAI211_X1 U18722 ( .C1(n15529), .C2(n15552), .A(n15528), .B(n15527), .ZN(
        n15530) );
  AOI211_X1 U18723 ( .C1(n15532), .C2(n16354), .A(n15531), .B(n15530), .ZN(
        n15533) );
  OAI211_X1 U18724 ( .C1(n15535), .C2(n15623), .A(n15534), .B(n15533), .ZN(
        P2_U3032) );
  OAI21_X1 U18725 ( .B1(n13752), .B2(n15536), .A(n13819), .ZN(n19074) );
  NAND3_X1 U18726 ( .A1(n15592), .A2(n15568), .A3(n15551), .ZN(n15550) );
  AOI21_X1 U18727 ( .B1(n15550), .B2(n15552), .A(n15537), .ZN(n15543) );
  NOR2_X1 U18728 ( .A1(n18918), .A2(n15614), .ZN(n15542) );
  NOR4_X1 U18729 ( .A1(n15567), .A2(n15539), .A3(n15538), .A4(n15551), .ZN(
        n15541) );
  NOR4_X1 U18730 ( .A1(n15543), .A2(n15542), .A3(n15541), .A4(n15540), .ZN(
        n15544) );
  OAI21_X1 U18731 ( .B1(n19074), .B2(n15355), .A(n15544), .ZN(n15545) );
  AOI21_X1 U18732 ( .B1(n15546), .B2(n16359), .A(n15545), .ZN(n15547) );
  OAI21_X1 U18733 ( .B1(n15548), .B2(n15629), .A(n15547), .ZN(P2_U3033) );
  NAND2_X1 U18734 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18985), .ZN(n15549) );
  OAI211_X1 U18735 ( .C1(n15552), .C2(n15551), .A(n15550), .B(n15549), .ZN(
        n15553) );
  AOI21_X1 U18736 ( .B1(n16354), .B2(n19076), .A(n15553), .ZN(n15554) );
  OAI21_X1 U18737 ( .B1(n15614), .B2(n15555), .A(n15554), .ZN(n15556) );
  AOI21_X1 U18738 ( .B1(n15557), .B2(n16359), .A(n15556), .ZN(n15558) );
  OAI21_X1 U18739 ( .B1(n15559), .B2(n15629), .A(n15558), .ZN(P2_U3034) );
  NOR2_X1 U18740 ( .A1(n18932), .A2(n15614), .ZN(n15574) );
  NAND2_X1 U18741 ( .A1(n15561), .A2(n15560), .ZN(n15605) );
  INV_X1 U18742 ( .A(n15605), .ZN(n15562) );
  AOI21_X1 U18743 ( .B1(n15599), .B2(n15563), .A(n15562), .ZN(n15595) );
  OR2_X1 U18744 ( .A1(n15564), .A2(n15565), .ZN(n15566) );
  NAND2_X1 U18745 ( .A1(n13751), .A2(n15566), .ZN(n19080) );
  INV_X1 U18746 ( .A(n19080), .ZN(n18936) );
  AOI211_X1 U18747 ( .C1(n15572), .C2(n15594), .A(n15568), .B(n15567), .ZN(
        n15569) );
  AOI211_X1 U18748 ( .C1(n16354), .C2(n18936), .A(n15570), .B(n15569), .ZN(
        n15571) );
  OAI21_X1 U18749 ( .B1(n15595), .B2(n15572), .A(n15571), .ZN(n15573) );
  AOI211_X1 U18750 ( .C1(n15575), .C2(n16359), .A(n15574), .B(n15573), .ZN(
        n15576) );
  OAI21_X1 U18751 ( .B1(n15577), .B2(n15629), .A(n15576), .ZN(P2_U3035) );
  NOR2_X1 U18752 ( .A1(n15579), .A2(n15578), .ZN(n15583) );
  NOR2_X1 U18753 ( .A1(n15581), .A2(n15580), .ZN(n15582) );
  XOR2_X1 U18754 ( .A(n15583), .B(n15582), .Z(n16323) );
  AOI21_X1 U18755 ( .B1(n15594), .B2(n15312), .A(n15584), .ZN(n16324) );
  NAND2_X1 U18756 ( .A1(n16324), .A2(n16357), .ZN(n15598) );
  INV_X1 U18757 ( .A(n13722), .ZN(n15585) );
  AOI21_X1 U18758 ( .B1(n15586), .B2(n13306), .A(n15585), .ZN(n19033) );
  NOR2_X1 U18759 ( .A1(n15587), .A2(n15588), .ZN(n15589) );
  OR2_X1 U18760 ( .A1(n15564), .A2(n15589), .ZN(n19084) );
  NOR2_X1 U18761 ( .A1(n15355), .A2(n19084), .ZN(n15591) );
  NOR2_X1 U18762 ( .A1(n12298), .A2(n18970), .ZN(n15590) );
  AOI211_X1 U18763 ( .C1(n15592), .C2(n15594), .A(n15591), .B(n15590), .ZN(
        n15593) );
  OAI21_X1 U18764 ( .B1(n15595), .B2(n15594), .A(n15593), .ZN(n15596) );
  AOI21_X1 U18765 ( .B1(n12862), .B2(n19033), .A(n15596), .ZN(n15597) );
  OAI211_X1 U18766 ( .C1(n16323), .C2(n15623), .A(n15598), .B(n15597), .ZN(
        P2_U3036) );
  NAND2_X1 U18767 ( .A1(n15599), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15606) );
  NOR2_X1 U18768 ( .A1(n15600), .A2(n13664), .ZN(n15601) );
  OR2_X1 U18769 ( .A1(n15587), .A2(n15601), .ZN(n19087) );
  INV_X1 U18770 ( .A(n19087), .ZN(n15603) );
  AOI21_X1 U18771 ( .B1(n16354), .B2(n15603), .A(n15602), .ZN(n15604) );
  OAI211_X1 U18772 ( .C1(n15607), .C2(n15606), .A(n15605), .B(n15604), .ZN(
        n15608) );
  AOI21_X1 U18773 ( .B1(n12862), .B2(n18964), .A(n15608), .ZN(n15611) );
  NAND2_X1 U18774 ( .A1(n15609), .A2(n16359), .ZN(n15610) );
  OAI211_X1 U18775 ( .C1(n15612), .C2(n15629), .A(n15611), .B(n15610), .ZN(
        P2_U3037) );
  NAND3_X1 U18776 ( .A1(n15613), .A2(n15339), .A3(n16357), .ZN(n15622) );
  NOR2_X1 U18777 ( .A1(n15615), .A2(n15614), .ZN(n15620) );
  NAND4_X1 U18778 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16362), .A3(
        n15616), .A4(n15618), .ZN(n16351) );
  OAI211_X1 U18779 ( .C1(n16352), .C2(n15618), .A(n16351), .B(n15617), .ZN(
        n15619) );
  AOI211_X1 U18780 ( .C1(n16354), .C2(n19090), .A(n15620), .B(n15619), .ZN(
        n15621) );
  OAI211_X1 U18781 ( .C1(n15624), .C2(n15623), .A(n15622), .B(n15621), .ZN(
        P2_U3039) );
  MUX2_X1 U18782 ( .A(n15626), .B(n15625), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n15634) );
  AOI22_X1 U18783 ( .A1(n12862), .A2(n19008), .B1(n16359), .B2(n15627), .ZN(
        n15633) );
  NOR2_X1 U18784 ( .A1(n15629), .A2(n15628), .ZN(n15630) );
  AOI211_X1 U18785 ( .C1(n19001), .C2(n16354), .A(n15631), .B(n15630), .ZN(
        n15632) );
  NAND3_X1 U18786 ( .A1(n15634), .A2(n15633), .A3(n15632), .ZN(P2_U3046) );
  INV_X1 U18787 ( .A(n15635), .ZN(n15638) );
  OAI222_X1 U18788 ( .A1(n16376), .A2(n19874), .B1(n15638), .B2(n15637), .C1(
        n19854), .C2(n15636), .ZN(n15639) );
  MUX2_X1 U18789 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15639), .S(
        n15641), .Z(P2_U3600) );
  OAI22_X1 U18790 ( .A1(n19445), .A2(n16376), .B1(n15640), .B2(n19854), .ZN(
        n15642) );
  MUX2_X1 U18791 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15642), .S(
        n15641), .Z(P2_U3596) );
  OAI21_X1 U18792 ( .B1(n19777), .B2(n19262), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15643) );
  NAND2_X1 U18793 ( .A1(n15643), .A2(n19852), .ZN(n15646) );
  NOR2_X1 U18794 ( .A1(n19447), .A2(n19266), .ZN(n19190) );
  INV_X1 U18795 ( .A(n19190), .ZN(n19217) );
  AND2_X1 U18796 ( .A1(n19721), .A2(n19217), .ZN(n15649) );
  OAI21_X1 U18797 ( .B1(n15647), .B2(n19190), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15644) );
  INV_X1 U18798 ( .A(n19224), .ZN(n15663) );
  AND2_X1 U18799 ( .A1(n15645), .A2(n19621), .ZN(n19749) );
  INV_X1 U18800 ( .A(n19749), .ZN(n19635) );
  INV_X1 U18801 ( .A(n15646), .ZN(n15650) );
  INV_X1 U18802 ( .A(n19621), .ZN(n19730) );
  AOI211_X1 U18803 ( .C1(n15647), .C2(n19668), .A(n19190), .B(n19852), .ZN(
        n15648) );
  AOI211_X2 U18804 ( .C1(n15650), .C2(n15649), .A(n19730), .B(n15648), .ZN(
        n19228) );
  INV_X1 U18805 ( .A(n19228), .ZN(n15661) );
  INV_X1 U18806 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16453) );
  AND2_X1 U18807 ( .A1(n19216), .A2(n15654), .ZN(n19748) );
  AOI22_X1 U18808 ( .A1(n19750), .A2(n19262), .B1(n19190), .B2(n19748), .ZN(
        n15655) );
  OAI21_X1 U18809 ( .B1(n19218), .B2(n19753), .A(n15655), .ZN(n15656) );
  AOI21_X1 U18810 ( .B1(n15661), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n15656), .ZN(n15657) );
  OAI21_X1 U18811 ( .B1(n15663), .B2(n19635), .A(n15657), .ZN(P2_U3051) );
  AND2_X1 U18812 ( .A1(n16303), .A2(n19621), .ZN(n19755) );
  INV_X1 U18813 ( .A(n19755), .ZN(n19639) );
  AOI22_X1 U18814 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19213), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19214), .ZN(n19759) );
  INV_X1 U18815 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16451) );
  INV_X1 U18816 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18219) );
  OAI22_X1 U18817 ( .A1(n16451), .A2(n19223), .B1(n18219), .B2(n19221), .ZN(
        n19756) );
  AND2_X1 U18818 ( .A1(n19216), .A2(n15658), .ZN(n19754) );
  AOI22_X1 U18819 ( .A1(n19756), .A2(n19262), .B1(n19190), .B2(n19754), .ZN(
        n15659) );
  OAI21_X1 U18820 ( .B1(n19218), .B2(n19759), .A(n15659), .ZN(n15660) );
  AOI21_X1 U18821 ( .B1(n15661), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n15660), .ZN(n15662) );
  OAI21_X1 U18822 ( .B1(n15663), .B2(n19639), .A(n15662), .ZN(P2_U3052) );
  INV_X1 U18823 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17011) );
  NAND2_X1 U18824 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17023), .ZN(n17012) );
  NAND2_X1 U18825 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16969), .ZN(n15739) );
  NAND2_X1 U18826 ( .A1(n18236), .A2(n17227), .ZN(n17231) );
  INV_X1 U18827 ( .A(n16969), .ZN(n16964) );
  NAND2_X1 U18828 ( .A1(n17221), .A2(n16964), .ZN(n16967) );
  OAI21_X1 U18829 ( .B1(n16960), .B2(n17231), .A(n16967), .ZN(n16958) );
  AOI22_X1 U18830 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15668) );
  AOI22_X1 U18831 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U18832 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18833 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15665) );
  NAND4_X1 U18834 ( .A1(n15668), .A2(n15667), .A3(n15666), .A4(n15665), .ZN(
        n15674) );
  AOI22_X1 U18835 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15672) );
  AOI22_X1 U18836 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U18837 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U18838 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15669) );
  NAND4_X1 U18839 ( .A1(n15672), .A2(n15671), .A3(n15670), .A4(n15669), .ZN(
        n15673) );
  NOR2_X1 U18840 ( .A1(n15674), .A2(n15673), .ZN(n15737) );
  AOI22_X1 U18841 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U18842 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18843 ( .A1(n15746), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U18844 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15675) );
  NAND4_X1 U18845 ( .A1(n15678), .A2(n15677), .A3(n15676), .A4(n15675), .ZN(
        n15684) );
  AOI22_X1 U18846 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18847 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15681) );
  AOI22_X1 U18848 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18849 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15679) );
  NAND4_X1 U18850 ( .A1(n15682), .A2(n15681), .A3(n15680), .A4(n15679), .ZN(
        n15683) );
  NOR2_X1 U18851 ( .A1(n15684), .A2(n15683), .ZN(n16965) );
  AOI22_X1 U18852 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17173), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15688) );
  AOI22_X1 U18853 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9697), .ZN(n15687) );
  AOI22_X1 U18854 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18855 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17175), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15685) );
  NAND4_X1 U18856 ( .A1(n15688), .A2(n15687), .A3(n15686), .A4(n15685), .ZN(
        n15694) );
  AOI22_X1 U18857 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15692) );
  AOI22_X1 U18858 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17176), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15691) );
  AOI22_X1 U18859 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17162), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U18860 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17159), .ZN(n15689) );
  NAND4_X1 U18861 ( .A1(n15692), .A2(n15691), .A3(n15690), .A4(n15689), .ZN(
        n15693) );
  NOR2_X1 U18862 ( .A1(n15694), .A2(n15693), .ZN(n16976) );
  AOI22_X1 U18863 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U18864 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18865 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15695) );
  OAI21_X1 U18866 ( .B1(n16878), .B2(n20872), .A(n15695), .ZN(n15701) );
  AOI22_X1 U18867 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U18868 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15698) );
  AOI22_X1 U18869 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15697) );
  AOI22_X1 U18870 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15696) );
  NAND4_X1 U18871 ( .A1(n15699), .A2(n15698), .A3(n15697), .A4(n15696), .ZN(
        n15700) );
  AOI211_X1 U18872 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n15701), .B(n15700), .ZN(n15702) );
  NAND3_X1 U18873 ( .A1(n15704), .A2(n15703), .A3(n15702), .ZN(n16981) );
  AOI22_X1 U18874 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15715) );
  AOI22_X1 U18875 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U18876 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15705) );
  OAI21_X1 U18877 ( .B1(n15706), .B2(n17198), .A(n15705), .ZN(n15712) );
  AOI22_X1 U18878 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U18879 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U18880 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15708) );
  AOI22_X1 U18881 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15707) );
  NAND4_X1 U18882 ( .A1(n15710), .A2(n15709), .A3(n15708), .A4(n15707), .ZN(
        n15711) );
  AOI211_X1 U18883 ( .C1(n17151), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15712), .B(n15711), .ZN(n15713) );
  NAND3_X1 U18884 ( .A1(n15715), .A2(n15714), .A3(n15713), .ZN(n16982) );
  NAND2_X1 U18885 ( .A1(n16981), .A2(n16982), .ZN(n16980) );
  NOR2_X1 U18886 ( .A1(n16976), .A2(n16980), .ZN(n16973) );
  AOI22_X1 U18887 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U18888 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15724) );
  INV_X1 U18889 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20869) );
  AOI22_X1 U18890 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15716) );
  OAI21_X1 U18891 ( .B1(n9793), .B2(n20869), .A(n15716), .ZN(n15722) );
  AOI22_X1 U18892 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18893 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18894 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15718) );
  AOI22_X1 U18895 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15717) );
  NAND4_X1 U18896 ( .A1(n15720), .A2(n15719), .A3(n15718), .A4(n15717), .ZN(
        n15721) );
  AOI211_X1 U18897 ( .C1(n17172), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n15722), .B(n15721), .ZN(n15723) );
  NAND3_X1 U18898 ( .A1(n15725), .A2(n15724), .A3(n15723), .ZN(n16972) );
  NAND2_X1 U18899 ( .A1(n16973), .A2(n16972), .ZN(n16971) );
  NOR2_X1 U18900 ( .A1(n16965), .A2(n16971), .ZN(n17254) );
  AOI22_X1 U18901 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15736) );
  AOI22_X1 U18902 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15735) );
  INV_X1 U18903 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20921) );
  AOI22_X1 U18904 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15726) );
  OAI21_X1 U18905 ( .B1(n15727), .B2(n20921), .A(n15726), .ZN(n15733) );
  AOI22_X1 U18906 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15731) );
  AOI22_X1 U18907 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U18908 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15729) );
  AOI22_X1 U18909 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15728) );
  NAND4_X1 U18910 ( .A1(n15731), .A2(n15730), .A3(n15729), .A4(n15728), .ZN(
        n15732) );
  AOI211_X1 U18911 ( .C1(n12484), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n15733), .B(n15732), .ZN(n15734) );
  NAND3_X1 U18912 ( .A1(n15736), .A2(n15735), .A3(n15734), .ZN(n17253) );
  NAND2_X1 U18913 ( .A1(n17254), .A2(n17253), .ZN(n17252) );
  NOR2_X1 U18914 ( .A1(n15737), .A2(n17252), .ZN(n16957) );
  AOI21_X1 U18915 ( .B1(n15737), .B2(n17252), .A(n16957), .ZN(n17248) );
  AOI22_X1 U18916 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16958), .B1(n17229), 
        .B2(n17248), .ZN(n15738) );
  OAI21_X1 U18917 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15739), .A(n15738), .ZN(
        P3_U2675) );
  AOI22_X1 U18918 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U18919 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15743) );
  AOI22_X1 U18920 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15742) );
  AOI22_X1 U18921 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15741) );
  NAND4_X1 U18922 ( .A1(n15744), .A2(n15743), .A3(n15742), .A4(n15741), .ZN(
        n15752) );
  AOI22_X1 U18923 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18924 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15745), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U18925 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U18926 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15747) );
  NAND4_X1 U18927 ( .A1(n15750), .A2(n15749), .A3(n15748), .A4(n15747), .ZN(
        n15751) );
  NOR2_X1 U18928 ( .A1(n15752), .A2(n15751), .ZN(n17327) );
  INV_X2 U18929 ( .A(n17229), .ZN(n17221) );
  INV_X1 U18930 ( .A(n17119), .ZN(n17105) );
  INV_X1 U18931 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20779) );
  OAI221_X1 U18932 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17105), .C1(n20779), 
        .C2(n17119), .A(n17221), .ZN(n15753) );
  OAI21_X1 U18933 ( .B1(n17327), .B2(n17221), .A(n15753), .ZN(P3_U2690) );
  NAND2_X1 U18934 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18348) );
  AOI221_X1 U18935 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18348), .C1(n15755), 
        .C2(n18348), .A(n15754), .ZN(n18198) );
  NOR2_X1 U18936 ( .A1(n15756), .A2(n20932), .ZN(n15757) );
  OAI21_X1 U18937 ( .B1(n15757), .B2(n18541), .A(n18199), .ZN(n18196) );
  AOI22_X1 U18938 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18198), .B1(
        n18196), .B2(n18674), .ZN(P3_U2865) );
  INV_X1 U18939 ( .A(n18632), .ZN(n16520) );
  NOR2_X1 U18940 ( .A1(n16520), .A2(n18837), .ZN(n15760) );
  NOR2_X1 U18941 ( .A1(n18835), .A2(n17441), .ZN(n17442) );
  NOR2_X1 U18942 ( .A1(n16537), .A2(n17442), .ZN(n15758) );
  AOI21_X1 U18943 ( .B1(n15760), .B2(n17380), .A(n15759), .ZN(n15762) );
  OAI21_X1 U18944 ( .B1(n18206), .B2(n17441), .A(n10050), .ZN(n15761) );
  NAND3_X1 U18945 ( .A1(n18632), .A2(n18844), .A3(n15761), .ZN(n15873) );
  OAI211_X1 U18946 ( .C1(n15764), .C2(n15763), .A(n15762), .B(n15873), .ZN(
        n18662) );
  INV_X1 U18947 ( .A(n18662), .ZN(n18672) );
  NAND2_X1 U18948 ( .A1(n18840), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18202) );
  INV_X1 U18949 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18194) );
  OR2_X1 U18950 ( .A1(n18194), .A2(n18788), .ZN(n15765) );
  OAI211_X1 U18951 ( .C1(n18692), .C2(n18672), .A(n18202), .B(n15765), .ZN(
        n18819) );
  INV_X1 U18952 ( .A(n18803), .ZN(n18817) );
  AOI21_X1 U18953 ( .B1(n15766), .B2(n18640), .A(n10050), .ZN(n18684) );
  NAND3_X1 U18954 ( .A1(n18819), .A2(n18817), .A3(n18684), .ZN(n15767) );
  OAI21_X1 U18955 ( .B1(n18819), .B2(n18640), .A(n15767), .ZN(P3_U3284) );
  INV_X1 U18956 ( .A(n18107), .ZN(n17913) );
  OAI22_X1 U18957 ( .A1(n16421), .A2(n18190), .B1(n16420), .B2(n17913), .ZN(
        n15768) );
  NOR2_X1 U18958 ( .A1(n15769), .A2(n15768), .ZN(n15837) );
  INV_X1 U18959 ( .A(n18076), .ZN(n17999) );
  AOI21_X1 U18960 ( .B1(n17999), .B2(n17887), .A(n15770), .ZN(n16423) );
  INV_X1 U18961 ( .A(n15771), .ZN(n16383) );
  INV_X1 U18962 ( .A(n15772), .ZN(n16382) );
  AOI22_X1 U18963 ( .A1(n18107), .A2(n16383), .B1(n18150), .B2(n16382), .ZN(
        n15840) );
  OAI21_X1 U18964 ( .B1(n18186), .B2(n16423), .A(n15840), .ZN(n15773) );
  AOI21_X1 U18965 ( .B1(n15774), .B2(n17500), .A(n15773), .ZN(n15779) );
  INV_X2 U18966 ( .A(n18184), .ZN(n18186) );
  NOR2_X1 U18967 ( .A1(n15776), .A2(n15775), .ZN(n15777) );
  XNOR2_X1 U18968 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15777), .ZN(
        n16403) );
  AOI22_X1 U18969 ( .A1(n18186), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18089), 
        .B2(n16403), .ZN(n15778) );
  OAI221_X1 U18970 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15837), 
        .C1(n16400), .C2(n15779), .A(n15778), .ZN(P3_U2833) );
  AOI22_X1 U18971 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19012), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18986), .ZN(n15791) );
  INV_X1 U18972 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16282) );
  OAI22_X1 U18973 ( .A1(n15780), .A2(n19005), .B1(n18999), .B2(n16282), .ZN(
        n15781) );
  INV_X1 U18974 ( .A(n15781), .ZN(n15790) );
  INV_X1 U18975 ( .A(n15782), .ZN(n16297) );
  OAI22_X1 U18976 ( .A1(n16315), .A2(n20705), .B1(n20698), .B2(n16297), .ZN(
        n15783) );
  INV_X1 U18977 ( .A(n15783), .ZN(n15789) );
  AOI21_X1 U18978 ( .B1(n15786), .B2(n15784), .A(n15785), .ZN(n15787) );
  NAND2_X1 U18979 ( .A1(n19009), .A2(n15787), .ZN(n15788) );
  NAND4_X1 U18980 ( .A1(n15791), .A2(n15790), .A3(n15789), .A4(n15788), .ZN(
        P2_U2833) );
  NOR2_X1 U18981 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15792), .ZN(n15833) );
  INV_X1 U18982 ( .A(n15793), .ZN(n15794) );
  NAND2_X1 U18983 ( .A1(n15795), .A2(n15794), .ZN(n15796) );
  OR2_X1 U18984 ( .A1(n15797), .A2(n15796), .ZN(n15798) );
  NAND2_X1 U18985 ( .A1(n20603), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15799) );
  AND2_X1 U18986 ( .A1(n15798), .A2(n15799), .ZN(n15826) );
  INV_X1 U18987 ( .A(n15826), .ZN(n15831) );
  INV_X1 U18988 ( .A(n15799), .ZN(n20683) );
  OAI21_X1 U18989 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20593), .A(n20525), 
        .ZN(n16226) );
  NAND2_X1 U18990 ( .A1(n15801), .A2(n15800), .ZN(n15808) );
  AOI21_X1 U18991 ( .B1(n15802), .B2(n9724), .A(n20317), .ZN(n15803) );
  AND2_X1 U18992 ( .A1(n15804), .A2(n15803), .ZN(n15806) );
  INV_X1 U18993 ( .A(n15806), .ZN(n15805) );
  NAND2_X1 U18994 ( .A1(n15805), .A2(n20524), .ZN(n15807) );
  AOI22_X1 U18995 ( .A1(n15808), .A2(n15807), .B1(n15806), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15811) );
  OAI21_X1 U18996 ( .B1(n15811), .B2(n15810), .A(n15809), .ZN(n15813) );
  NAND2_X1 U18997 ( .A1(n15811), .A2(n15810), .ZN(n15812) );
  NAND2_X1 U18998 ( .A1(n15813), .A2(n15812), .ZN(n15815) );
  AOI222_X1 U18999 ( .A1(n15815), .A2(n11318), .B1(n15815), .B2(n15814), .C1(
        n11318), .C2(n15814), .ZN(n15825) );
  NAND2_X1 U19000 ( .A1(n19907), .A2(n15816), .ZN(n15817) );
  NAND2_X1 U19001 ( .A1(n15818), .A2(n15817), .ZN(n15820) );
  AND4_X1 U19002 ( .A1(n15822), .A2(n15821), .A3(n15820), .A4(n15819), .ZN(
        n15823) );
  OAI211_X1 U19003 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15825), .A(
        n15824), .B(n15823), .ZN(n16234) );
  OAI21_X1 U19004 ( .B1(n20589), .B2(n20684), .A(n15826), .ZN(n16235) );
  NAND2_X1 U19005 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16235), .ZN(n15827) );
  AOI21_X1 U19006 ( .B1(n20589), .B2(n16234), .A(n15827), .ZN(n15829) );
  OAI211_X1 U19007 ( .C1(n20683), .C2(n16226), .A(n15829), .B(n15828), .ZN(
        n15830) );
  OAI21_X1 U19008 ( .B1(n15831), .B2(n20046), .A(n15830), .ZN(n15832) );
  AOI21_X1 U19009 ( .B1(n20680), .B2(n15833), .A(n15832), .ZN(P1_U3161) );
  NAND2_X1 U19010 ( .A1(n15835), .A2(n15834), .ZN(n15836) );
  XNOR2_X1 U19011 ( .A(n15836), .B(n16394), .ZN(n16392) );
  INV_X1 U19012 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18775) );
  NOR2_X1 U19013 ( .A1(n18184), .A2(n18775), .ZN(n16386) );
  NOR3_X1 U19014 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15837), .A3(
        n16400), .ZN(n15838) );
  AOI211_X1 U19015 ( .C1(n18089), .C2(n16392), .A(n16386), .B(n15838), .ZN(
        n15839) );
  OAI221_X1 U19016 ( .B1(n16394), .B2(n15841), .C1(n16394), .C2(n15840), .A(
        n15839), .ZN(P3_U2832) );
  INV_X1 U19017 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20609) );
  OAI221_X1 U19018 ( .B1(n20593), .B2(HOLD), .C1(n20593), .C2(n20609), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n15844) );
  INV_X1 U19019 ( .A(HOLD), .ZN(n20594) );
  OAI211_X1 U19020 ( .C1(n20609), .C2(n20594), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15842) );
  NAND3_X1 U19021 ( .A1(n15844), .A2(n15843), .A3(n15842), .ZN(P1_U3195) );
  INV_X1 U19022 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16510) );
  NOR2_X1 U19023 ( .A1(n20044), .A2(n16510), .ZN(P1_U2905) );
  AND2_X1 U19024 ( .A1(n9750), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16045) );
  INV_X1 U19025 ( .A(n15845), .ZN(n15848) );
  INV_X1 U19026 ( .A(n16046), .ZN(n15846) );
  NOR3_X1 U19027 ( .A1(n14768), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15846), .ZN(n15847) );
  AOI21_X1 U19028 ( .B1(n16045), .B2(n15848), .A(n15847), .ZN(n15849) );
  XNOR2_X1 U19029 ( .A(n15849), .B(n11308), .ZN(n16044) );
  INV_X1 U19030 ( .A(n15850), .ZN(n15852) );
  OAI21_X1 U19031 ( .B1(n15852), .B2(n16172), .A(n9692), .ZN(n16115) );
  AOI22_X1 U19032 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16115), .B1(
        n20106), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15861) );
  NAND2_X1 U19033 ( .A1(n15854), .A2(n15853), .ZN(n15858) );
  AOI21_X1 U19034 ( .B1(n9907), .B2(n15949), .A(n15855), .ZN(n15857) );
  OR2_X1 U19035 ( .A1(n15857), .A2(n15856), .ZN(n15938) );
  OAI22_X1 U19036 ( .A1(n16120), .A2(n15858), .B1(n16210), .B2(n15938), .ZN(
        n15859) );
  INV_X1 U19037 ( .A(n15859), .ZN(n15860) );
  OAI211_X1 U19038 ( .C1(n16044), .C2(n16186), .A(n15861), .B(n15860), .ZN(
        P1_U3011) );
  NOR3_X1 U19039 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15865) );
  INV_X1 U19040 ( .A(n16377), .ZN(n15864) );
  NOR3_X1 U19041 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16380), .A3(n15862), 
        .ZN(n16372) );
  INV_X1 U19042 ( .A(n15863), .ZN(n15869) );
  NOR4_X1 U19043 ( .A1(n15865), .A2(n15864), .A3(n16372), .A4(n15869), .ZN(
        P2_U3178) );
  INV_X1 U19044 ( .A(n15866), .ZN(n15868) );
  AOI211_X1 U19045 ( .C1(n15869), .C2(n15868), .A(n15867), .B(n19621), .ZN(
        n19891) );
  INV_X1 U19046 ( .A(n19891), .ZN(n19888) );
  NOR2_X1 U19047 ( .A1(n15870), .A2(n19888), .ZN(P2_U3047) );
  NAND3_X1 U19048 ( .A1(n18203), .A2(n18206), .A3(n15871), .ZN(n15872) );
  NAND2_X1 U19049 ( .A1(n18236), .A2(n17379), .ZN(n17348) );
  INV_X1 U19050 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20811) );
  NAND2_X2 U19051 ( .A1(n18664), .A2(n17379), .ZN(n17368) );
  AOI22_X1 U19052 ( .A1(n17373), .A2(BUF2_REG_0__SCAN_IN), .B1(n17372), .B2(
        n17869), .ZN(n15874) );
  OAI221_X1 U19053 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17348), .C1(n20811), 
        .C2(n17379), .A(n15874), .ZN(P3_U2735) );
  NAND2_X1 U19054 ( .A1(n19949), .A2(n15878), .ZN(n15883) );
  OAI22_X1 U19055 ( .A1(n12028), .A2(n19996), .B1(n15875), .B2(n19991), .ZN(
        n15876) );
  AOI21_X1 U19056 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n20006), .A(n15876), .ZN(
        n15877) );
  OAI221_X1 U19057 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n15878), .C1(n20647), 
        .C2(n15883), .A(n15877), .ZN(n15879) );
  AOI21_X1 U19058 ( .B1(n16010), .B2(n19959), .A(n15879), .ZN(n15880) );
  OAI21_X1 U19059 ( .B1(n15881), .B2(n20010), .A(n15880), .ZN(P1_U2813) );
  AOI22_X1 U19060 ( .A1(n15882), .A2(n20013), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n20006), .ZN(n15890) );
  INV_X1 U19061 ( .A(n15883), .ZN(n15888) );
  OAI22_X1 U19062 ( .A1(n15885), .A2(n15977), .B1(n15884), .B2(n20010), .ZN(
        n15886) );
  OAI211_X1 U19063 ( .C1(n15891), .C2(n19996), .A(n15890), .B(n15889), .ZN(
        P1_U2814) );
  NOR2_X1 U19064 ( .A1(n15892), .A2(n15977), .ZN(n15900) );
  NOR2_X1 U19065 ( .A1(n19984), .A2(n15893), .ZN(n15899) );
  INV_X1 U19066 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15894) );
  NOR2_X1 U19067 ( .A1(n19996), .A2(n15894), .ZN(n15898) );
  OAI22_X1 U19068 ( .A1(n19991), .A2(n15896), .B1(P1_REIP_REG_25__SCAN_IN), 
        .B2(n15895), .ZN(n15897) );
  NOR4_X1 U19069 ( .A1(n15900), .A2(n15899), .A3(n15898), .A4(n15897), .ZN(
        n15903) );
  OAI21_X1 U19070 ( .B1(n15901), .B2(n15908), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15902) );
  OAI211_X1 U19071 ( .C1(n20010), .C2(n15904), .A(n15903), .B(n15902), .ZN(
        P1_U2815) );
  OAI22_X1 U19072 ( .A1(n16034), .A2(n19991), .B1(n15905), .B2(n19984), .ZN(
        n15906) );
  AOI21_X1 U19073 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20014), .A(
        n15906), .ZN(n15911) );
  NAND3_X1 U19074 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(n15942), .ZN(n15932) );
  OAI21_X1 U19075 ( .B1(n15907), .B2(n15932), .A(n20837), .ZN(n15909) );
  AOI22_X1 U19076 ( .A1(n16031), .A2(n19959), .B1(n15909), .B2(n15908), .ZN(
        n15910) );
  OAI211_X1 U19077 ( .C1(n20010), .C2(n15912), .A(n15911), .B(n15910), .ZN(
        P1_U2817) );
  AOI22_X1 U19078 ( .A1(n15913), .A2(n20013), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n20006), .ZN(n15921) );
  INV_X1 U19079 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20639) );
  OR2_X1 U19080 ( .A1(n15914), .A2(n20639), .ZN(n15923) );
  AOI21_X1 U19081 ( .B1(n20005), .B2(n15923), .A(n19992), .ZN(n15931) );
  OAI21_X1 U19082 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19980), .A(n15931), 
        .ZN(n15919) );
  NAND2_X1 U19083 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15915) );
  NOR3_X1 U19084 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15915), .A3(n15932), 
        .ZN(n15918) );
  OAI22_X1 U19085 ( .A1(n15916), .A2(n15977), .B1(n20010), .B2(n16107), .ZN(
        n15917) );
  AOI211_X1 U19086 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n15919), .A(n15918), 
        .B(n15917), .ZN(n15920) );
  OAI211_X1 U19087 ( .C1(n15922), .C2(n19996), .A(n15921), .B(n15920), .ZN(
        P1_U2818) );
  NOR3_X1 U19088 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19980), .A3(n15923), 
        .ZN(n15926) );
  OAI22_X1 U19089 ( .A1(n15931), .A2(n14873), .B1(n15924), .B2(n19984), .ZN(
        n15925) );
  AOI211_X1 U19090 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15926), .B(n15925), .ZN(n15930) );
  INV_X1 U19091 ( .A(n15927), .ZN(n15928) );
  AOI22_X1 U19092 ( .A1(n16036), .A2(n19959), .B1(n19993), .B2(n15928), .ZN(
        n15929) );
  OAI211_X1 U19093 ( .C1(n16039), .C2(n19991), .A(n15930), .B(n15929), .ZN(
        P1_U2819) );
  AOI21_X1 U19094 ( .B1(n20639), .B2(n15932), .A(n15931), .ZN(n15935) );
  OAI22_X1 U19095 ( .A1(n15933), .A2(n19996), .B1(n16001), .B2(n19984), .ZN(
        n15934) );
  AOI211_X1 U19096 ( .C1(n20013), .C2(n16040), .A(n15935), .B(n15934), .ZN(
        n15940) );
  INV_X1 U19097 ( .A(n15936), .ZN(n15948) );
  XOR2_X1 U19098 ( .A(n15937), .B(n15948), .Z(n16041) );
  INV_X1 U19099 ( .A(n15938), .ZN(n15999) );
  AOI22_X1 U19100 ( .A1(n16041), .A2(n19959), .B1(n19993), .B2(n15999), .ZN(
        n15939) );
  NAND2_X1 U19101 ( .A1(n15940), .A2(n15939), .ZN(P1_U2820) );
  INV_X1 U19102 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20636) );
  OAI22_X1 U19103 ( .A1(n15963), .A2(n20636), .B1(n16052), .B2(n19991), .ZN(
        n15945) );
  NAND2_X1 U19104 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15941) );
  OAI211_X1 U19105 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n15942), .B(n15941), .ZN(n15943) );
  OAI211_X1 U19106 ( .C1(n19984), .C2(n16003), .A(n19982), .B(n15943), .ZN(
        n15944) );
  AOI211_X1 U19107 ( .C1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n20014), .A(
        n15945), .B(n15944), .ZN(n15952) );
  NAND2_X1 U19108 ( .A1(n14567), .A2(n15946), .ZN(n15947) );
  AND2_X1 U19109 ( .A1(n15948), .A2(n15947), .ZN(n16049) );
  XNOR2_X1 U19110 ( .A(n15950), .B(n15949), .ZN(n16116) );
  AOI22_X1 U19111 ( .A1(n16049), .A2(n19959), .B1(n19993), .B2(n16116), .ZN(
        n15951) );
  NAND2_X1 U19112 ( .A1(n15952), .A2(n15951), .ZN(P1_U2821) );
  AOI21_X1 U19113 ( .B1(n15953), .B2(n15968), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n15962) );
  INV_X1 U19114 ( .A(n19982), .ZN(n19957) );
  OAI22_X1 U19115 ( .A1(n11830), .A2(n19996), .B1(n16005), .B2(n19984), .ZN(
        n15954) );
  AOI211_X1 U19116 ( .C1(n20013), .C2(n16060), .A(n19957), .B(n15954), .ZN(
        n15961) );
  INV_X1 U19117 ( .A(n15955), .ZN(n15957) );
  AOI21_X1 U19118 ( .B1(n15957), .B2(n15956), .A(n14566), .ZN(n16061) );
  XNOR2_X1 U19119 ( .A(n15959), .B(n15958), .ZN(n16133) );
  AOI22_X1 U19120 ( .A1(n16061), .A2(n19959), .B1(n19993), .B2(n16133), .ZN(
        n15960) );
  OAI211_X1 U19121 ( .C1(n15963), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        P1_U2823) );
  AOI22_X1 U19122 ( .A1(n16071), .A2(n20013), .B1(n19993), .B2(n15964), .ZN(
        n15972) );
  OAI22_X1 U19123 ( .A1(n15966), .A2(n19996), .B1(n15965), .B2(n19984), .ZN(
        n15967) );
  AOI211_X1 U19124 ( .C1(n15968), .C2(n20796), .A(n19957), .B(n15967), .ZN(
        n15971) );
  AOI22_X1 U19125 ( .A1(n16072), .A2(n19959), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15969), .ZN(n15970) );
  NAND3_X1 U19126 ( .A1(n15972), .A2(n15971), .A3(n15970), .ZN(P1_U2825) );
  NAND2_X1 U19127 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15973) );
  AOI21_X1 U19128 ( .B1(n20005), .B2(n15973), .A(n15993), .ZN(n15991) );
  AOI22_X1 U19129 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20006), .B1(n19993), 
        .B2(n16166), .ZN(n15974) );
  OAI211_X1 U19130 ( .C1(n19996), .C2(n15975), .A(n15974), .B(n19982), .ZN(
        n15980) );
  OAI22_X1 U19131 ( .A1(n15978), .A2(n15977), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15976), .ZN(n15979) );
  AOI211_X1 U19132 ( .C1(n15981), .C2(n20013), .A(n15980), .B(n15979), .ZN(
        n15982) );
  OAI21_X1 U19133 ( .B1(n15991), .B2(n20629), .A(n15982), .ZN(P1_U2827) );
  AOI21_X1 U19134 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15992), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15990) );
  AOI21_X1 U19135 ( .B1(n15985), .B2(n15984), .A(n15983), .ZN(n16178) );
  OAI22_X1 U19136 ( .A1(n15986), .A2(n19996), .B1(n16007), .B2(n19984), .ZN(
        n15987) );
  AOI211_X1 U19137 ( .C1(n16178), .C2(n19993), .A(n19957), .B(n15987), .ZN(
        n15989) );
  AOI22_X1 U19138 ( .A1(n16080), .A2(n20013), .B1(n19959), .B2(n16079), .ZN(
        n15988) );
  OAI211_X1 U19139 ( .C1(n15991), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        P1_U2828) );
  AOI22_X1 U19140 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n20006), .B1(n15992), 
        .B2(n14888), .ZN(n15998) );
  AOI22_X1 U19141 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n20014), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n15993), .ZN(n15994) );
  OAI211_X1 U19142 ( .C1(n15995), .C2(n20010), .A(n15994), .B(n19982), .ZN(
        n15996) );
  AOI21_X1 U19143 ( .B1(n19959), .B2(n16083), .A(n15996), .ZN(n15997) );
  OAI211_X1 U19144 ( .C1(n16087), .C2(n19991), .A(n15998), .B(n15997), .ZN(
        P1_U2829) );
  AOI22_X1 U19145 ( .A1(n16041), .A2(n12893), .B1(n20021), .B2(n15999), .ZN(
        n16000) );
  OAI21_X1 U19146 ( .B1(n20023), .B2(n16001), .A(n16000), .ZN(P1_U2852) );
  AOI22_X1 U19147 ( .A1(n16049), .A2(n12893), .B1(n20021), .B2(n16116), .ZN(
        n16002) );
  OAI21_X1 U19148 ( .B1(n20023), .B2(n16003), .A(n16002), .ZN(P1_U2853) );
  AOI22_X1 U19149 ( .A1(n16061), .A2(n12893), .B1(n20021), .B2(n16133), .ZN(
        n16004) );
  OAI21_X1 U19150 ( .B1(n20023), .B2(n16005), .A(n16004), .ZN(P1_U2855) );
  AOI22_X1 U19151 ( .A1(n16079), .A2(n12893), .B1(n20021), .B2(n16178), .ZN(
        n16006) );
  OAI21_X1 U19152 ( .B1(n20023), .B2(n16007), .A(n16006), .ZN(P1_U2860) );
  INV_X1 U19153 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16438) );
  AOI22_X1 U19154 ( .A1(n16024), .A2(n16008), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16022), .ZN(n16012) );
  INV_X1 U19155 ( .A(n16009), .ZN(n16026) );
  AOI22_X1 U19156 ( .A1(n16010), .A2(n16026), .B1(n16025), .B2(DATAI_27_), 
        .ZN(n16011) );
  OAI211_X1 U19157 ( .C1(n16438), .C2(n16029), .A(n16012), .B(n16011), .ZN(
        P1_U2877) );
  INV_X1 U19158 ( .A(n16013), .ZN(n16014) );
  AOI22_X1 U19159 ( .A1(n16024), .A2(n16014), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16022), .ZN(n16016) );
  AOI22_X1 U19160 ( .A1(n16041), .A2(n16026), .B1(n16025), .B2(DATAI_20_), 
        .ZN(n16015) );
  OAI211_X1 U19161 ( .C1(n16029), .C2(n16451), .A(n16016), .B(n16015), .ZN(
        P1_U2884) );
  INV_X1 U19162 ( .A(n16017), .ZN(n16018) );
  AOI22_X1 U19163 ( .A1(n16024), .A2(n16018), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16022), .ZN(n16020) );
  AOI22_X1 U19164 ( .A1(n16049), .A2(n16026), .B1(n16025), .B2(DATAI_19_), 
        .ZN(n16019) );
  OAI211_X1 U19165 ( .C1(n16029), .C2(n16453), .A(n16020), .B(n16019), .ZN(
        P1_U2885) );
  INV_X1 U19166 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19192) );
  INV_X1 U19167 ( .A(n16021), .ZN(n16023) );
  AOI22_X1 U19168 ( .A1(n16024), .A2(n16023), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16022), .ZN(n16028) );
  AOI22_X1 U19169 ( .A1(n16061), .A2(n16026), .B1(n16025), .B2(DATAI_17_), 
        .ZN(n16027) );
  OAI211_X1 U19170 ( .C1(n16029), .C2(n19192), .A(n16028), .B(n16027), .ZN(
        P1_U2887) );
  AOI22_X1 U19171 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16033) );
  AOI22_X1 U19172 ( .A1(n16031), .A2(n20062), .B1(n20071), .B2(n16030), .ZN(
        n16032) );
  OAI211_X1 U19173 ( .C1(n20066), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        P1_U2976) );
  AOI22_X1 U19174 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16038) );
  AOI22_X1 U19175 ( .A1(n16036), .A2(n20062), .B1(n20071), .B2(n16035), .ZN(
        n16037) );
  OAI211_X1 U19176 ( .C1(n20066), .C2(n16039), .A(n16038), .B(n16037), .ZN(
        P1_U2978) );
  AOI22_X1 U19177 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16043) );
  AOI22_X1 U19178 ( .A1(n16041), .A2(n20062), .B1(n20070), .B2(n16040), .ZN(
        n16042) );
  OAI211_X1 U19179 ( .C1(n16044), .C2(n19906), .A(n16043), .B(n16042), .ZN(
        P1_U2979) );
  AOI22_X1 U19180 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16051) );
  NOR2_X1 U19181 ( .A1(n16046), .A2(n16045), .ZN(n16047) );
  XNOR2_X1 U19182 ( .A(n16048), .B(n16047), .ZN(n16117) );
  AOI22_X1 U19183 ( .A1(n20071), .A2(n16117), .B1(n16049), .B2(n20062), .ZN(
        n16050) );
  OAI211_X1 U19184 ( .C1(n20066), .C2(n16052), .A(n16051), .B(n16050), .ZN(
        P1_U2980) );
  INV_X1 U19185 ( .A(n16053), .ZN(n16054) );
  NOR2_X1 U19186 ( .A1(n16055), .A2(n16054), .ZN(n16058) );
  NOR2_X1 U19187 ( .A1(n16058), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16057) );
  MUX2_X1 U19188 ( .A(n16058), .B(n16057), .S(n16056), .Z(n16059) );
  XNOR2_X1 U19189 ( .A(n16059), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16139) );
  AOI22_X1 U19190 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16063) );
  AOI22_X1 U19191 ( .A1(n16061), .A2(n20062), .B1(n16060), .B2(n20070), .ZN(
        n16062) );
  OAI211_X1 U19192 ( .C1(n19906), .C2(n16139), .A(n16063), .B(n16062), .ZN(
        P1_U2982) );
  INV_X1 U19193 ( .A(n16064), .ZN(n16065) );
  NOR2_X1 U19194 ( .A1(n16066), .A2(n16065), .ZN(n16070) );
  NAND2_X1 U19195 ( .A1(n16068), .A2(n16067), .ZN(n16069) );
  XNOR2_X1 U19196 ( .A(n16070), .B(n16069), .ZN(n16155) );
  AOI22_X1 U19197 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U19198 ( .A1(n16072), .A2(n20062), .B1(n16071), .B2(n20070), .ZN(
        n16073) );
  OAI211_X1 U19199 ( .C1(n16155), .C2(n19906), .A(n16074), .B(n16073), .ZN(
        P1_U2984) );
  OAI21_X1 U19200 ( .B1(n16077), .B2(n16076), .A(n16075), .ZN(n16078) );
  INV_X1 U19201 ( .A(n16078), .ZN(n16187) );
  AOI22_X1 U19202 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16082) );
  AOI22_X1 U19203 ( .A1(n20070), .A2(n16080), .B1(n20062), .B2(n16079), .ZN(
        n16081) );
  OAI211_X1 U19204 ( .C1(n16187), .C2(n19906), .A(n16082), .B(n16081), .ZN(
        P1_U2987) );
  AOI22_X1 U19205 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16086) );
  AOI22_X1 U19206 ( .A1(n20071), .A2(n16084), .B1(n20062), .B2(n16083), .ZN(
        n16085) );
  OAI211_X1 U19207 ( .C1(n20066), .C2(n16087), .A(n16086), .B(n16085), .ZN(
        P1_U2988) );
  AOI22_X1 U19208 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16093) );
  NAND2_X1 U19209 ( .A1(n16090), .A2(n16089), .ZN(n16091) );
  XNOR2_X1 U19210 ( .A(n16088), .B(n16091), .ZN(n16212) );
  AOI22_X1 U19211 ( .A1(n16212), .A2(n20071), .B1(n20062), .B2(n19950), .ZN(
        n16092) );
  OAI211_X1 U19212 ( .C1(n20066), .C2(n19953), .A(n16093), .B(n16092), .ZN(
        P1_U2992) );
  AOI22_X1 U19213 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16099) );
  XNOR2_X1 U19214 ( .A(n16095), .B(n16094), .ZN(n16096) );
  XNOR2_X1 U19215 ( .A(n16097), .B(n16096), .ZN(n16222) );
  AOI22_X1 U19216 ( .A1(n16222), .A2(n20071), .B1(n20062), .B2(n20018), .ZN(
        n16098) );
  OAI211_X1 U19217 ( .C1(n20066), .C2(n19962), .A(n16099), .B(n16098), .ZN(
        P1_U2993) );
  AOI22_X1 U19218 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16104) );
  INV_X1 U19219 ( .A(n16100), .ZN(n16102) );
  INV_X1 U19220 ( .A(n16101), .ZN(n19968) );
  AOI22_X1 U19221 ( .A1(n16102), .A2(n20071), .B1(n20062), .B2(n19968), .ZN(
        n16103) );
  OAI211_X1 U19222 ( .C1(n20066), .C2(n19971), .A(n16104), .B(n16103), .ZN(
        P1_U2994) );
  AOI22_X1 U19223 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16106), .B1(
        n20103), .B2(n16105), .ZN(n16114) );
  NAND2_X1 U19224 ( .A1(n20106), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16113) );
  INV_X1 U19225 ( .A(n16107), .ZN(n16108) );
  NAND2_X1 U19226 ( .A1(n16108), .A2(n20098), .ZN(n16112) );
  OAI211_X1 U19227 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16110), .B(n16109), .ZN(
        n16111) );
  NAND4_X1 U19228 ( .A1(n16114), .A2(n16113), .A3(n16112), .A4(n16111), .ZN(
        P1_U3009) );
  AOI22_X1 U19229 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16115), .B1(
        n20106), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16119) );
  AOI22_X1 U19230 ( .A1(n16117), .A2(n20103), .B1(n20098), .B2(n16116), .ZN(
        n16118) );
  OAI211_X1 U19231 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16120), .A(
        n16119), .B(n16118), .ZN(P1_U3012) );
  INV_X1 U19232 ( .A(n16121), .ZN(n16123) );
  AOI22_X1 U19233 ( .A1(n16123), .A2(n20103), .B1(n20098), .B2(n16122), .ZN(
        n16132) );
  AOI21_X1 U19234 ( .B1(n16126), .B2(n16125), .A(n16124), .ZN(n16177) );
  OAI21_X1 U19235 ( .B1(n16143), .B2(n16127), .A(n16177), .ZN(n16135) );
  NOR2_X1 U19236 ( .A1(n16209), .A2(n14771), .ZN(n16128) );
  AOI221_X1 U19237 ( .B1(n16130), .B2(n16129), .C1(n16135), .C2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(n16128), .ZN(n16131) );
  NAND2_X1 U19238 ( .A1(n16132), .A2(n16131), .ZN(P1_U3013) );
  AOI22_X1 U19239 ( .A1(n16133), .A2(n20098), .B1(n20106), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16138) );
  INV_X1 U19240 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16144) );
  NOR2_X1 U19241 ( .A1(n16142), .A2(n16144), .ZN(n16136) );
  NOR2_X1 U19242 ( .A1(n16134), .A2(n16164), .ZN(n16145) );
  OAI221_X1 U19243 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16136), 
        .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n16145), .A(n16135), .ZN(
        n16137) );
  OAI211_X1 U19244 ( .C1(n16139), .C2(n16186), .A(n16138), .B(n16137), .ZN(
        P1_U3014) );
  AOI22_X1 U19245 ( .A1(n16141), .A2(n20103), .B1(n20098), .B2(n16140), .ZN(
        n16149) );
  NAND2_X1 U19246 ( .A1(n20106), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16148) );
  AND2_X1 U19247 ( .A1(n16142), .A2(n16145), .ZN(n16152) );
  OAI21_X1 U19248 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16143), .A(
        n16177), .ZN(n16153) );
  OAI21_X1 U19249 ( .B1(n16152), .B2(n16153), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16147) );
  NAND3_X1 U19250 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16145), .A3(
        n16144), .ZN(n16146) );
  NAND4_X1 U19251 ( .A1(n16149), .A2(n16148), .A3(n16147), .A4(n16146), .ZN(
        P1_U3015) );
  OAI22_X1 U19252 ( .A1(n16150), .A2(n16210), .B1(n20796), .B2(n16209), .ZN(
        n16151) );
  AOI211_X1 U19253 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16153), .A(
        n16152), .B(n16151), .ZN(n16154) );
  OAI21_X1 U19254 ( .B1(n16155), .B2(n16186), .A(n16154), .ZN(P1_U3016) );
  AOI21_X1 U19255 ( .B1(n16157), .B2(n20098), .A(n16156), .ZN(n16163) );
  NOR2_X1 U19256 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16158), .ZN(
        n16160) );
  AOI22_X1 U19257 ( .A1(n16161), .A2(n16160), .B1(n20103), .B2(n16159), .ZN(
        n16162) );
  OAI211_X1 U19258 ( .C1(n16177), .C2(n16164), .A(n16163), .B(n16162), .ZN(
        P1_U3017) );
  AOI21_X1 U19259 ( .B1(n16166), .B2(n20098), .A(n16165), .ZN(n16176) );
  OAI221_X1 U19260 ( .B1(n16169), .B2(n16168), .C1(n16169), .C2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16167), .ZN(n16170) );
  OAI21_X1 U19261 ( .B1(n16172), .B2(n16171), .A(n16170), .ZN(n16173) );
  AOI22_X1 U19262 ( .A1(n16174), .A2(n20103), .B1(n14788), .B2(n16173), .ZN(
        n16175) );
  OAI211_X1 U19263 ( .C1(n16177), .C2(n14788), .A(n16176), .B(n16175), .ZN(
        P1_U3018) );
  AOI22_X1 U19264 ( .A1(n16178), .A2(n20098), .B1(n20106), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16185) );
  INV_X1 U19265 ( .A(n20108), .ZN(n16200) );
  OAI21_X1 U19266 ( .B1(n16200), .B2(n16180), .A(n16179), .ZN(n16183) );
  OAI21_X1 U19267 ( .B1(n16181), .B2(n16225), .A(n11303), .ZN(n16182) );
  OAI21_X1 U19268 ( .B1(n11303), .B2(n16183), .A(n16182), .ZN(n16184) );
  OAI211_X1 U19269 ( .C1(n16187), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        P1_U3019) );
  AOI21_X1 U19270 ( .B1(n16189), .B2(n20098), .A(n16188), .ZN(n16197) );
  AOI22_X1 U19271 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16191), .B1(
        n20103), .B2(n16190), .ZN(n16196) );
  OAI221_X1 U19272 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16194), .C2(n16193), .A(
        n16192), .ZN(n16195) );
  NAND3_X1 U19273 ( .A1(n16197), .A2(n16196), .A3(n16195), .ZN(P1_U3021) );
  OAI21_X1 U19274 ( .B1(n16200), .B2(n16199), .A(n16198), .ZN(n16221) );
  AOI21_X1 U19275 ( .B1(n16094), .B2(n16201), .A(n16221), .ZN(n16214) );
  INV_X1 U19276 ( .A(n19936), .ZN(n16203) );
  AOI21_X1 U19277 ( .B1(n16203), .B2(n20098), .A(n16202), .ZN(n16208) );
  AOI211_X1 U19278 ( .C1(n14113), .C2(n16215), .A(n16094), .B(n16225), .ZN(
        n16205) );
  AOI22_X1 U19279 ( .A1(n16206), .A2(n20103), .B1(n16205), .B2(n16204), .ZN(
        n16207) );
  OAI211_X1 U19280 ( .C1(n16214), .C2(n14113), .A(n16208), .B(n16207), .ZN(
        P1_U3023) );
  OR2_X1 U19281 ( .A1(n16094), .A2(n16225), .ZN(n16216) );
  INV_X1 U19282 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20620) );
  OAI22_X1 U19283 ( .A1(n19945), .A2(n16210), .B1(n20620), .B2(n16209), .ZN(
        n16211) );
  AOI21_X1 U19284 ( .B1(n16212), .B2(n20103), .A(n16211), .ZN(n16213) );
  OAI221_X1 U19285 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16216), .C1(
        n16215), .C2(n16214), .A(n16213), .ZN(P1_U3024) );
  NOR2_X1 U19286 ( .A1(n16218), .A2(n16217), .ZN(n16219) );
  AOI22_X1 U19287 ( .A1(n9831), .A2(n20098), .B1(n20106), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16224) );
  AOI22_X1 U19288 ( .A1(n16222), .A2(n20103), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16221), .ZN(n16223) );
  OAI211_X1 U19289 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16225), .A(
        n16224), .B(n16223), .ZN(P1_U3025) );
  OAI211_X1 U19290 ( .C1(n16234), .C2(n16235), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n16226), .ZN(n16232) );
  AOI21_X1 U19291 ( .B1(n20683), .B2(n16228), .A(n16227), .ZN(n20590) );
  INV_X1 U19292 ( .A(n16229), .ZN(n16230) );
  NAND2_X1 U19293 ( .A1(n20590), .A2(n16230), .ZN(n16231) );
  AOI22_X1 U19294 ( .A1(n16233), .A2(n16232), .B1(n16235), .B2(n16231), .ZN(
        P1_U3162) );
  NOR2_X1 U19295 ( .A1(n16235), .A2(n16234), .ZN(n16237) );
  OAI21_X1 U19296 ( .B1(n16237), .B2(n16236), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n16238) );
  NAND2_X1 U19297 ( .A1(n16239), .A2(n16238), .ZN(P1_U3466) );
  AOI211_X1 U19298 ( .C1(n16242), .C2(n16240), .A(n12836), .B(n16241), .ZN(
        n16250) );
  INV_X1 U19299 ( .A(n16243), .ZN(n16248) );
  AOI22_X1 U19300 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19012), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n20694), .ZN(n16244) );
  OAI21_X1 U19301 ( .B1(n20697), .B2(n19833), .A(n16244), .ZN(n16245) );
  AOI21_X1 U19302 ( .B1(n16246), .B2(n20703), .A(n16245), .ZN(n16247) );
  OAI21_X1 U19303 ( .B1(n16248), .B2(n20705), .A(n16247), .ZN(n16249) );
  AOI211_X1 U19304 ( .C1(n19002), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        n16252) );
  INV_X1 U19305 ( .A(n16252), .ZN(P2_U2829) );
  AOI22_X1 U19306 ( .A1(n16253), .A2(n20703), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n18986), .ZN(n16264) );
  AOI22_X1 U19307 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n20694), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19012), .ZN(n16263) );
  INV_X1 U19308 ( .A(n16254), .ZN(n16256) );
  AOI22_X1 U19309 ( .A1(n16256), .A2(n19007), .B1(n19002), .B2(n16255), .ZN(
        n16262) );
  AOI21_X1 U19310 ( .B1(n16259), .B2(n16257), .A(n16258), .ZN(n16260) );
  NAND2_X1 U19311 ( .A1(n19009), .A2(n16260), .ZN(n16261) );
  NAND4_X1 U19312 ( .A1(n16264), .A2(n16263), .A3(n16262), .A4(n16261), .ZN(
        P2_U2830) );
  AOI22_X1 U19313 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19012), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18986), .ZN(n16276) );
  AOI22_X1 U19314 ( .A1(n16265), .A2(n20703), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n20694), .ZN(n16275) );
  OAI22_X1 U19315 ( .A1(n16267), .A2(n20705), .B1(n20698), .B2(n16266), .ZN(
        n16268) );
  INV_X1 U19316 ( .A(n16268), .ZN(n16274) );
  AOI21_X1 U19317 ( .B1(n16271), .B2(n16269), .A(n16270), .ZN(n16272) );
  NAND2_X1 U19318 ( .A1(n19009), .A2(n16272), .ZN(n16273) );
  NAND4_X1 U19319 ( .A1(n16276), .A2(n16275), .A3(n16274), .A4(n16273), .ZN(
        P2_U2832) );
  INV_X1 U19320 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16277) );
  AOI22_X1 U19321 ( .A1(n19048), .A2(n16278), .B1(n16277), .B2(n19052), .ZN(
        P2_U2856) );
  NAND2_X1 U19322 ( .A1(n16280), .A2(n16279), .ZN(n16281) );
  NAND2_X1 U19323 ( .A1(n14378), .A2(n16281), .ZN(n16298) );
  OAI22_X1 U19324 ( .A1(n16298), .A2(n19041), .B1(n19048), .B2(n16282), .ZN(
        n16283) );
  INV_X1 U19325 ( .A(n16283), .ZN(n16284) );
  OAI21_X1 U19326 ( .B1(n19052), .B2(n16315), .A(n16284), .ZN(P2_U2865) );
  OR2_X1 U19327 ( .A1(n15042), .A2(n16285), .ZN(n16286) );
  NAND2_X1 U19328 ( .A1(n16287), .A2(n16286), .ZN(n16304) );
  INV_X1 U19329 ( .A(n16304), .ZN(n16288) );
  AOI22_X1 U19330 ( .A1(n16288), .A2(n19018), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19052), .ZN(n16289) );
  OAI21_X1 U19331 ( .B1(n19052), .B2(n16290), .A(n16289), .ZN(P2_U2867) );
  AND2_X1 U19332 ( .A1(n16292), .A2(n16291), .ZN(n16293) );
  NOR2_X1 U19333 ( .A1(n16294), .A2(n16293), .ZN(n16310) );
  AOI22_X1 U19334 ( .A1(n16310), .A2(n19018), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19052), .ZN(n16295) );
  OAI21_X1 U19335 ( .B1(n19052), .B2(n16296), .A(n16295), .ZN(P2_U2869) );
  AOI22_X1 U19336 ( .A1(n19059), .A2(n19207), .B1(n19119), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16302) );
  AOI22_X1 U19337 ( .A1(n19061), .A2(BUF1_REG_22__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16301) );
  OAI22_X1 U19338 ( .A1(n16298), .A2(n19124), .B1(n19063), .B2(n16297), .ZN(
        n16299) );
  INV_X1 U19339 ( .A(n16299), .ZN(n16300) );
  NAND3_X1 U19340 ( .A1(n16302), .A2(n16301), .A3(n16300), .ZN(P2_U2897) );
  AOI22_X1 U19341 ( .A1(n19059), .A2(n16303), .B1(n19119), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16309) );
  AOI22_X1 U19342 ( .A1(n19061), .A2(BUF1_REG_20__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16308) );
  OAI22_X1 U19343 ( .A1(n16305), .A2(n19063), .B1(n19124), .B2(n16304), .ZN(
        n16306) );
  INV_X1 U19344 ( .A(n16306), .ZN(n16307) );
  NAND3_X1 U19345 ( .A1(n16309), .A2(n16308), .A3(n16307), .ZN(P2_U2899) );
  AOI22_X1 U19346 ( .A1(n19059), .A2(n19197), .B1(n19119), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16314) );
  AOI22_X1 U19347 ( .A1(n19061), .A2(BUF1_REG_18__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16313) );
  AOI22_X1 U19348 ( .A1(n16311), .A2(n19120), .B1(n19106), .B2(n16310), .ZN(
        n16312) );
  NAND3_X1 U19349 ( .A1(n16314), .A2(n16313), .A3(n16312), .ZN(P2_U2901) );
  AOI22_X1 U19350 ( .A1(n16322), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18985), .ZN(n16320) );
  INV_X1 U19351 ( .A(n16315), .ZN(n16317) );
  AOI222_X1 U19352 ( .A1(n16318), .A2(n16346), .B1(n19176), .B2(n16317), .C1(
        n10876), .C2(n16316), .ZN(n16319) );
  AOI22_X1 U19353 ( .A1(n16322), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18985), .ZN(n16327) );
  INV_X1 U19354 ( .A(n16323), .ZN(n16325) );
  AOI222_X1 U19355 ( .A1(n16325), .A2(n16346), .B1(n19176), .B2(n19033), .C1(
        n10876), .C2(n16324), .ZN(n16326) );
  OAI211_X1 U19356 ( .C1(n19172), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        P2_U3004) );
  AOI22_X1 U19357 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18985), .B1(n16343), 
        .B2(n16329), .ZN(n16341) );
  NAND2_X1 U19358 ( .A1(n16331), .A2(n16330), .ZN(n16335) );
  NAND2_X1 U19359 ( .A1(n16333), .A2(n16332), .ZN(n16334) );
  XNOR2_X1 U19360 ( .A(n16335), .B(n16334), .ZN(n16360) );
  OAI21_X1 U19361 ( .B1(n16336), .B2(n16338), .A(n16337), .ZN(n16339) );
  INV_X1 U19362 ( .A(n16339), .ZN(n16356) );
  AOI222_X1 U19363 ( .A1(n16360), .A2(n16346), .B1(n19176), .B2(n16358), .C1(
        n10876), .C2(n16356), .ZN(n16340) );
  OAI211_X1 U19364 ( .C1(n19184), .C2(n16342), .A(n16341), .B(n16340), .ZN(
        P2_U3006) );
  AOI22_X1 U19365 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18985), .B1(n16343), 
        .B2(n18976), .ZN(n16349) );
  INV_X1 U19366 ( .A(n16344), .ZN(n16347) );
  AOI222_X1 U19367 ( .A1(n16347), .A2(n10876), .B1(n16346), .B2(n16345), .C1(
        n19176), .C2(n18977), .ZN(n16348) );
  OAI211_X1 U19368 ( .C1(n19184), .C2(n16350), .A(n16349), .B(n16348), .ZN(
        P2_U3008) );
  NAND2_X1 U19369 ( .A1(n16352), .A2(n16351), .ZN(n16355) );
  AOI22_X1 U19370 ( .A1(n16355), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16354), .B2(n16353), .ZN(n16366) );
  AOI222_X1 U19371 ( .A1(n16360), .A2(n16359), .B1(n12862), .B2(n16358), .C1(
        n16357), .C2(n16356), .ZN(n16365) );
  NAND2_X1 U19372 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18985), .ZN(n16364) );
  NAND3_X1 U19373 ( .A1(n16362), .A2(n16361), .A3(n20760), .ZN(n16363) );
  NAND4_X1 U19374 ( .A1(n16366), .A2(n16365), .A3(n16364), .A4(n16363), .ZN(
        P2_U3038) );
  INV_X1 U19375 ( .A(n19886), .ZN(n16369) );
  OAI21_X1 U19376 ( .B1(n16369), .B2(n16368), .A(n16367), .ZN(n16370) );
  INV_X1 U19377 ( .A(n16370), .ZN(n16381) );
  INV_X1 U19378 ( .A(n16371), .ZN(n16374) );
  AOI211_X1 U19379 ( .C1(n18862), .C2(n16374), .A(n16373), .B(n16372), .ZN(
        n16379) );
  OAI211_X1 U19380 ( .C1(n16377), .C2(n16376), .A(n16380), .B(n16375), .ZN(
        n16378) );
  OAI211_X1 U19381 ( .C1(n16381), .C2(n16380), .A(n16379), .B(n16378), .ZN(
        P2_U3176) );
  NAND2_X1 U19382 ( .A1(n17839), .A2(n16382), .ZN(n16398) );
  NAND2_X1 U19383 ( .A1(n17781), .A2(n16383), .ZN(n16399) );
  NAND2_X1 U19384 ( .A1(n17980), .A2(n17582), .ZN(n17580) );
  INV_X1 U19385 ( .A(n17580), .ZN(n17938) );
  INV_X1 U19386 ( .A(n17739), .ZN(n18061) );
  INV_X1 U19387 ( .A(n17662), .ZN(n17986) );
  NOR3_X1 U19388 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16385), .A3(
        n17519), .ZN(n16391) );
  INV_X1 U19389 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16574) );
  XOR2_X1 U19390 ( .A(n16404), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16571) );
  AOI21_X1 U19391 ( .B1(n17687), .B2(n16571), .A(n16386), .ZN(n16387) );
  OAI221_X1 U19392 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16389), .C1(
        n16574), .C2(n16388), .A(n16387), .ZN(n16390) );
  AOI211_X1 U19393 ( .C1(n17765), .C2(n16392), .A(n16391), .B(n16390), .ZN(
        n16393) );
  OAI221_X1 U19394 ( .B1(n16394), .B2(n16398), .C1(n16394), .C2(n16399), .A(
        n16393), .ZN(P3_U2800) );
  OAI21_X1 U19395 ( .B1(n18488), .B2(n16395), .A(n16584), .ZN(n16396) );
  AOI22_X1 U19396 ( .A1(n18186), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16397), 
        .B2(n16396), .ZN(n16409) );
  AOI21_X1 U19397 ( .B1(n16421), .B2(n16400), .A(n16398), .ZN(n16402) );
  AOI21_X1 U19398 ( .B1(n16400), .B2(n16420), .A(n16399), .ZN(n16401) );
  AOI211_X1 U19399 ( .C1(n17765), .C2(n16403), .A(n16402), .B(n16401), .ZN(
        n16408) );
  AOI21_X1 U19400 ( .B1(n16405), .B2(n16584), .A(n16404), .ZN(n16583) );
  OAI21_X1 U19401 ( .B1(n17687), .B2(n16406), .A(n16583), .ZN(n16407) );
  NAND3_X1 U19402 ( .A1(n16409), .A2(n16408), .A3(n16407), .ZN(P3_U2801) );
  AOI21_X1 U19403 ( .B1(n17603), .B2(n17512), .A(n16426), .ZN(n17499) );
  AOI22_X1 U19404 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17770), .B1(
        n17603), .B2(n17500), .ZN(n17498) );
  NOR2_X1 U19405 ( .A1(n17499), .A2(n17498), .ZN(n17497) );
  INV_X1 U19406 ( .A(n18188), .ZN(n18174) );
  NAND2_X1 U19407 ( .A1(n17603), .A2(n18174), .ZN(n16414) );
  NOR2_X1 U19408 ( .A1(n18636), .A2(n16417), .ZN(n18041) );
  AOI22_X1 U19409 ( .A1(n18630), .A2(n18061), .B1(n16384), .B2(n18041), .ZN(
        n17985) );
  INV_X1 U19410 ( .A(n16410), .ZN(n16411) );
  OAI21_X1 U19411 ( .B1(n17985), .B2(n17986), .A(n16411), .ZN(n17915) );
  NAND2_X1 U19412 ( .A1(n16412), .A2(n17915), .ZN(n17892) );
  OAI22_X1 U19413 ( .A1(n17497), .A2(n16414), .B1(n16413), .B2(n17892), .ZN(
        n16415) );
  AOI22_X1 U19414 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18186), .B1(n17500), 
        .B2(n16415), .ZN(n16429) );
  INV_X1 U19415 ( .A(n16416), .ZN(n16419) );
  OAI211_X1 U19416 ( .C1(n16419), .C2(n17512), .A(n16418), .B(n16417), .ZN(
        n16424) );
  AOI22_X1 U19417 ( .A1(n18630), .A2(n16421), .B1(n18041), .B2(n16420), .ZN(
        n16422) );
  OAI211_X1 U19418 ( .C1(n17497), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        n16425) );
  NAND3_X1 U19419 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18184), .A3(
        n16425), .ZN(n16428) );
  NAND3_X1 U19420 ( .A1(n18089), .A2(n16426), .A3(n17498), .ZN(n16427) );
  NAND3_X1 U19421 ( .A1(n16429), .A2(n16428), .A3(n16427), .ZN(P3_U2834) );
  NOR3_X1 U19422 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16431) );
  NOR4_X1 U19423 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16430) );
  NAND4_X1 U19424 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16431), .A3(n16430), .A4(
        U215), .ZN(U213) );
  INV_X1 U19425 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19130) );
  INV_X1 U19426 ( .A(U214), .ZN(n16473) );
  NOR2_X1 U19427 ( .A1(n16473), .A2(n16432), .ZN(n16476) );
  CLKBUF_X1 U19428 ( .A(n16475), .Z(n16479) );
  OAI222_X1 U19429 ( .A1(U212), .A2(n19130), .B1(n16479), .B2(n19054), .C1(
        U214), .C2(n16510), .ZN(U216) );
  INV_X1 U19430 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19431 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16472), .ZN(n16433) );
  OAI21_X1 U19432 ( .B1(n16434), .B2(n16479), .A(n16433), .ZN(U217) );
  INV_X1 U19433 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19201) );
  AOI22_X1 U19434 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16472), .ZN(n16435) );
  OAI21_X1 U19435 ( .B1(n19201), .B2(n16479), .A(n16435), .ZN(U218) );
  INV_X1 U19436 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16437) );
  AOI22_X1 U19437 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16472), .ZN(n16436) );
  OAI21_X1 U19438 ( .B1(n16437), .B2(n16479), .A(n16436), .ZN(U219) );
  INV_X1 U19439 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n16439) );
  INV_X1 U19440 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n20936) );
  OAI222_X1 U19441 ( .A1(U214), .A2(n16439), .B1(n16479), .B2(n16438), .C1(
        U212), .C2(n20936), .ZN(U220) );
  INV_X1 U19442 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16441) );
  AOI22_X1 U19443 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16472), .ZN(n16440) );
  OAI21_X1 U19444 ( .B1(n16441), .B2(n16479), .A(n16440), .ZN(U221) );
  INV_X1 U19445 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16443) );
  AOI22_X1 U19446 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16472), .ZN(n16442) );
  OAI21_X1 U19447 ( .B1(n16443), .B2(n16479), .A(n16442), .ZN(U222) );
  INV_X1 U19448 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U19449 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16472), .ZN(n16444) );
  OAI21_X1 U19450 ( .B1(n16445), .B2(n16479), .A(n16444), .ZN(U223) );
  INV_X1 U19451 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20807) );
  INV_X1 U19452 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n16446) );
  OAI222_X1 U19453 ( .A1(U212), .A2(n16502), .B1(n16479), .B2(n20807), .C1(
        U214), .C2(n16446), .ZN(U224) );
  INV_X1 U19454 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19209) );
  AOI22_X1 U19455 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16472), .ZN(n16447) );
  OAI21_X1 U19456 ( .B1(n19209), .B2(n16479), .A(n16447), .ZN(U225) );
  INV_X1 U19457 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16449) );
  AOI22_X1 U19458 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16472), .ZN(n16448) );
  OAI21_X1 U19459 ( .B1(n16449), .B2(n16479), .A(n16448), .ZN(U226) );
  AOI22_X1 U19460 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16472), .ZN(n16450) );
  OAI21_X1 U19461 ( .B1(n16451), .B2(n16475), .A(n16450), .ZN(U227) );
  AOI22_X1 U19462 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16472), .ZN(n16452) );
  OAI21_X1 U19463 ( .B1(n16453), .B2(n16479), .A(n16452), .ZN(U228) );
  AOI222_X1 U19464 ( .A1(n16473), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n16476), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n16472), .C2(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n16454) );
  INV_X1 U19465 ( .A(n16454), .ZN(U229) );
  INV_X1 U19466 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16497) );
  OAI222_X1 U19467 ( .A1(U212), .A2(n16497), .B1(n16479), .B2(n19192), .C1(
        U214), .C2(n20804), .ZN(U230) );
  INV_X1 U19468 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n19187) );
  AOI22_X1 U19469 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16472), .ZN(n16455) );
  OAI21_X1 U19470 ( .B1(n19187), .B2(n16475), .A(n16455), .ZN(U231) );
  AOI22_X1 U19471 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16472), .ZN(n16456) );
  OAI21_X1 U19472 ( .B1(n13352), .B2(n16479), .A(n16456), .ZN(U232) );
  INV_X1 U19473 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16493) );
  INV_X1 U19474 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n20731) );
  OAI222_X1 U19475 ( .A1(U212), .A2(n16493), .B1(n16479), .B2(n13346), .C1(
        U214), .C2(n20731), .ZN(U233) );
  AOI22_X1 U19476 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16472), .ZN(n16457) );
  OAI21_X1 U19477 ( .B1(n13373), .B2(n16475), .A(n16457), .ZN(U234) );
  INV_X1 U19478 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16491) );
  INV_X1 U19479 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n20824) );
  OAI222_X1 U19480 ( .A1(U212), .A2(n16491), .B1(n16479), .B2(n16458), .C1(
        U214), .C2(n20824), .ZN(U235) );
  AOI22_X1 U19481 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16472), .ZN(n16459) );
  OAI21_X1 U19482 ( .B1(n13337), .B2(n16479), .A(n16459), .ZN(U236) );
  AOI22_X1 U19483 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16472), .ZN(n16460) );
  OAI21_X1 U19484 ( .B1(n16461), .B2(n16475), .A(n16460), .ZN(U237) );
  AOI22_X1 U19485 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16472), .ZN(n16462) );
  OAI21_X1 U19486 ( .B1(n16463), .B2(n16479), .A(n16462), .ZN(U238) );
  AOI22_X1 U19487 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16472), .ZN(n16464) );
  OAI21_X1 U19488 ( .B1(n20761), .B2(n16479), .A(n16464), .ZN(U239) );
  INV_X1 U19489 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16466) );
  AOI22_X1 U19490 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16472), .ZN(n16465) );
  OAI21_X1 U19491 ( .B1(n16466), .B2(n16475), .A(n16465), .ZN(U240) );
  AOI222_X1 U19492 ( .A1(n16473), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n16476), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n16472), .C2(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n16467) );
  INV_X1 U19493 ( .A(n16467), .ZN(U241) );
  INV_X1 U19494 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19495 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16476), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16472), .ZN(n16468) );
  OAI21_X1 U19496 ( .B1(n16469), .B2(U214), .A(n16468), .ZN(U242) );
  INV_X1 U19497 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20748) );
  AOI22_X1 U19498 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16472), .ZN(n16470) );
  OAI21_X1 U19499 ( .B1(n20748), .B2(n16479), .A(n16470), .ZN(U243) );
  INV_X1 U19500 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n20040) );
  AOI22_X1 U19501 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16476), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16472), .ZN(n16471) );
  OAI21_X1 U19502 ( .B1(n20040), .B2(U214), .A(n16471), .ZN(U244) );
  AOI22_X1 U19503 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16473), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16472), .ZN(n16474) );
  OAI21_X1 U19504 ( .B1(n20904), .B2(n16475), .A(n16474), .ZN(U245) );
  INV_X1 U19505 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n20867) );
  AOI22_X1 U19506 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16476), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16472), .ZN(n16477) );
  OAI21_X1 U19507 ( .B1(n20867), .B2(U214), .A(n16477), .ZN(U246) );
  INV_X1 U19508 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16480) );
  INV_X1 U19509 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n20043) );
  OAI222_X1 U19510 ( .A1(U212), .A2(n16480), .B1(n16479), .B2(n16478), .C1(
        U214), .C2(n20043), .ZN(U247) );
  AOI22_X1 U19511 ( .A1(n16509), .A2(n16480), .B1(n18200), .B2(U215), .ZN(U251) );
  OAI22_X1 U19512 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16509), .ZN(n16481) );
  INV_X1 U19513 ( .A(n16481), .ZN(U252) );
  INV_X1 U19514 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19515 ( .A1(n16494), .A2(n16482), .B1(n18210), .B2(U215), .ZN(U253) );
  OAI22_X1 U19516 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16509), .ZN(n16483) );
  INV_X1 U19517 ( .A(n16483), .ZN(U254) );
  INV_X1 U19518 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16484) );
  INV_X1 U19519 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18220) );
  AOI22_X1 U19520 ( .A1(n16494), .A2(n16484), .B1(n18220), .B2(U215), .ZN(U255) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16485) );
  INV_X1 U19522 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18224) );
  AOI22_X1 U19523 ( .A1(n16509), .A2(n16485), .B1(n18224), .B2(U215), .ZN(U256) );
  INV_X1 U19524 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n20749) );
  INV_X1 U19525 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18229) );
  AOI22_X1 U19526 ( .A1(n16494), .A2(n20749), .B1(n18229), .B2(U215), .ZN(U257) );
  INV_X1 U19527 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16486) );
  INV_X1 U19528 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U19529 ( .A1(n16494), .A2(n16486), .B1(n18233), .B2(U215), .ZN(U258) );
  INV_X1 U19530 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16487) );
  INV_X1 U19531 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19532 ( .A1(n16494), .A2(n16487), .B1(n17471), .B2(U215), .ZN(U259) );
  INV_X1 U19533 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16488) );
  INV_X1 U19534 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U19535 ( .A1(n16494), .A2(n16488), .B1(n17473), .B2(U215), .ZN(U260) );
  INV_X1 U19536 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16489) );
  INV_X1 U19537 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U19538 ( .A1(n16494), .A2(n16489), .B1(n17475), .B2(U215), .ZN(U261) );
  INV_X1 U19539 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16490) );
  INV_X1 U19540 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U19541 ( .A1(n16494), .A2(n16490), .B1(n17477), .B2(U215), .ZN(U262) );
  INV_X1 U19542 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U19543 ( .A1(n16509), .A2(n16491), .B1(n17479), .B2(U215), .ZN(U263) );
  INV_X1 U19544 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16492) );
  INV_X1 U19545 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U19546 ( .A1(n16494), .A2(n16492), .B1(n17482), .B2(U215), .ZN(U264) );
  INV_X1 U19547 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U19548 ( .A1(n16494), .A2(n16493), .B1(n17487), .B2(U215), .ZN(U265) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16509), .ZN(n16495) );
  INV_X1 U19550 ( .A(n16495), .ZN(U266) );
  INV_X1 U19551 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16496) );
  INV_X1 U19552 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19186) );
  AOI22_X1 U19553 ( .A1(n16509), .A2(n16496), .B1(n19186), .B2(U215), .ZN(U267) );
  AOI22_X1 U19554 ( .A1(n16509), .A2(n16497), .B1(n13875), .B2(U215), .ZN(U268) );
  INV_X1 U19555 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n20783) );
  INV_X1 U19556 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U19557 ( .A1(n16509), .A2(n20783), .B1(n18211), .B2(U215), .ZN(U269) );
  INV_X1 U19558 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16498) );
  AOI22_X1 U19559 ( .A1(n16509), .A2(n16498), .B1(n15118), .B2(U215), .ZN(U270) );
  INV_X1 U19560 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16499) );
  AOI22_X1 U19561 ( .A1(n16509), .A2(n16499), .B1(n18219), .B2(U215), .ZN(U271) );
  INV_X1 U19562 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16500) );
  AOI22_X1 U19563 ( .A1(n16509), .A2(n16500), .B1(n15107), .B2(U215), .ZN(U272) );
  INV_X1 U19564 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16501) );
  INV_X1 U19565 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19208) );
  AOI22_X1 U19566 ( .A1(n16509), .A2(n16501), .B1(n19208), .B2(U215), .ZN(U273) );
  INV_X1 U19567 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U19568 ( .A1(n16509), .A2(n16502), .B1(n19222), .B2(U215), .ZN(U274) );
  OAI22_X1 U19569 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16509), .ZN(n16503) );
  INV_X1 U19570 ( .A(n16503), .ZN(U275) );
  OAI22_X1 U19571 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16509), .ZN(n16504) );
  INV_X1 U19572 ( .A(n16504), .ZN(U276) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16509), .ZN(n16505) );
  INV_X1 U19574 ( .A(n16505), .ZN(U277) );
  INV_X1 U19575 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U19576 ( .A1(n16509), .A2(n20936), .B1(n18215), .B2(U215), .ZN(U278) );
  OAI22_X1 U19577 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16509), .ZN(n16506) );
  INV_X1 U19578 ( .A(n16506), .ZN(U279) );
  INV_X1 U19579 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16507) );
  INV_X1 U19580 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19200) );
  AOI22_X1 U19581 ( .A1(n16509), .A2(n16507), .B1(n19200), .B2(U215), .ZN(U280) );
  INV_X1 U19582 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16508) );
  INV_X1 U19583 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n20757) );
  AOI22_X1 U19584 ( .A1(n16509), .A2(n16508), .B1(n20757), .B2(U215), .ZN(U281) );
  INV_X1 U19585 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U19586 ( .A1(n16509), .A2(n19130), .B1(n18232), .B2(U215), .ZN(U282) );
  INV_X1 U19587 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17382) );
  AOI222_X1 U19588 ( .A1(n17382), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n16510), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n19130), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n16511) );
  INV_X2 U19589 ( .A(n16513), .ZN(n16512) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20803) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U19592 ( .A1(n16512), .A2(n20803), .B1(n19810), .B2(n16513), .ZN(
        U347) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20920) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19595 ( .A1(n16512), .A2(n20920), .B1(n19809), .B2(n16513), .ZN(
        U348) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18733) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19808) );
  AOI22_X1 U19598 ( .A1(n16512), .A2(n18733), .B1(n19808), .B2(n16513), .ZN(
        U349) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18732) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U19601 ( .A1(n16512), .A2(n18732), .B1(n19807), .B2(n16513), .ZN(
        U350) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18730) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U19604 ( .A1(n16512), .A2(n18730), .B1(n19806), .B2(n16513), .ZN(
        U351) );
  INV_X1 U19605 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U19606 ( .A1(n16512), .A2(n20793), .B1(n19805), .B2(n16513), .ZN(
        U352) );
  INV_X1 U19607 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18728) );
  INV_X1 U19608 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U19609 ( .A1(n16512), .A2(n18728), .B1(n19804), .B2(n16513), .ZN(
        U353) );
  INV_X1 U19610 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18726) );
  INV_X1 U19611 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19803) );
  AOI22_X1 U19612 ( .A1(n16512), .A2(n18726), .B1(n19803), .B2(n16513), .ZN(
        U354) );
  INV_X1 U19613 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18774) );
  INV_X1 U19614 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19841) );
  AOI22_X1 U19615 ( .A1(n16512), .A2(n18774), .B1(n19841), .B2(n16513), .ZN(
        U355) );
  INV_X1 U19616 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18771) );
  INV_X1 U19617 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19839) );
  AOI22_X1 U19618 ( .A1(n16512), .A2(n18771), .B1(n19839), .B2(n16513), .ZN(
        U356) );
  INV_X1 U19619 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18768) );
  INV_X1 U19620 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19837) );
  AOI22_X1 U19621 ( .A1(n16512), .A2(n18768), .B1(n19837), .B2(n16513), .ZN(
        U357) );
  INV_X1 U19622 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20891) );
  INV_X1 U19623 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19835) );
  AOI22_X1 U19624 ( .A1(n16512), .A2(n20891), .B1(n19835), .B2(n16513), .ZN(
        U358) );
  INV_X1 U19625 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18766) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19834) );
  AOI22_X1 U19627 ( .A1(n16512), .A2(n18766), .B1(n19834), .B2(n16513), .ZN(
        U359) );
  INV_X1 U19628 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18764) );
  INV_X1 U19629 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19832) );
  AOI22_X1 U19630 ( .A1(n16512), .A2(n18764), .B1(n19832), .B2(n16513), .ZN(
        U360) );
  INV_X1 U19631 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18763) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U19633 ( .A1(n16512), .A2(n18763), .B1(n19830), .B2(n16513), .ZN(
        U361) );
  INV_X1 U19634 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18761) );
  INV_X1 U19635 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U19636 ( .A1(n16512), .A2(n18761), .B1(n19829), .B2(n16513), .ZN(
        U362) );
  INV_X1 U19637 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18759) );
  INV_X1 U19638 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19828) );
  AOI22_X1 U19639 ( .A1(n16512), .A2(n18759), .B1(n19828), .B2(n16513), .ZN(
        U363) );
  INV_X1 U19640 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18757) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19827) );
  AOI22_X1 U19642 ( .A1(n16512), .A2(n18757), .B1(n19827), .B2(n16513), .ZN(
        U364) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18724) );
  INV_X1 U19644 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20821) );
  AOI22_X1 U19645 ( .A1(n16512), .A2(n18724), .B1(n20821), .B2(n16513), .ZN(
        U365) );
  INV_X1 U19646 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18755) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U19648 ( .A1(n16512), .A2(n18755), .B1(n19825), .B2(n16513), .ZN(
        U366) );
  INV_X1 U19649 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18753) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U19651 ( .A1(n16512), .A2(n18753), .B1(n19823), .B2(n16513), .ZN(
        U367) );
  INV_X1 U19652 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18751) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U19654 ( .A1(n16512), .A2(n18751), .B1(n19821), .B2(n16513), .ZN(
        U368) );
  INV_X1 U19655 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18749) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19820) );
  AOI22_X1 U19657 ( .A1(n16512), .A2(n18749), .B1(n19820), .B2(n16513), .ZN(
        U369) );
  INV_X1 U19658 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18748) );
  INV_X1 U19659 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U19660 ( .A1(n16512), .A2(n18748), .B1(n19818), .B2(n16513), .ZN(
        U370) );
  INV_X1 U19661 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18746) );
  INV_X1 U19662 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20728) );
  AOI22_X1 U19663 ( .A1(n16512), .A2(n18746), .B1(n20728), .B2(n16513), .ZN(
        U371) );
  INV_X1 U19664 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18743) );
  INV_X1 U19665 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19816) );
  AOI22_X1 U19666 ( .A1(n16512), .A2(n18743), .B1(n19816), .B2(n16513), .ZN(
        U372) );
  INV_X1 U19667 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18742) );
  INV_X1 U19668 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U19669 ( .A1(n16512), .A2(n18742), .B1(n19814), .B2(n16513), .ZN(
        U373) );
  INV_X1 U19670 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18739) );
  INV_X1 U19671 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19813) );
  AOI22_X1 U19672 ( .A1(n16512), .A2(n18739), .B1(n19813), .B2(n16513), .ZN(
        U374) );
  INV_X1 U19673 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18738) );
  INV_X1 U19674 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19812) );
  AOI22_X1 U19675 ( .A1(n16512), .A2(n18738), .B1(n19812), .B2(n16513), .ZN(
        U375) );
  INV_X1 U19676 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18722) );
  INV_X1 U19677 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20721) );
  AOI22_X1 U19678 ( .A1(n16512), .A2(n18722), .B1(n20721), .B2(n16513), .ZN(
        U376) );
  INV_X1 U19679 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16514) );
  NOR2_X1 U19680 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18719), .ZN(n18708) );
  OAI22_X1 U19681 ( .A1(n18705), .A2(n18708), .B1(n18719), .B2(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18703) );
  INV_X1 U19682 ( .A(n18703), .ZN(n18786) );
  OAI21_X1 U19683 ( .B1(n18719), .B2(n16514), .A(n18783), .ZN(P3_U2633) );
  INV_X1 U19684 ( .A(n18851), .ZN(n16515) );
  NOR2_X1 U19685 ( .A1(n18840), .A2(n16515), .ZN(n18698) );
  AOI221_X1 U19686 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n17443), .C1(
        P3_CODEFETCH_REG_SCAN_IN), .C2(n16521), .A(n18698), .ZN(n16516) );
  INV_X1 U19687 ( .A(n16516), .ZN(P3_U2634) );
  INV_X1 U19688 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18721) );
  AOI21_X1 U19689 ( .B1(n18719), .B2(n18721), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16517) );
  AOI22_X1 U19690 ( .A1(n18848), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16517), 
        .B2(n18849), .ZN(P3_U2635) );
  NOR2_X1 U19691 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16518) );
  OAI21_X1 U19692 ( .B1(n16518), .B2(BS16), .A(n18786), .ZN(n18784) );
  OAI21_X1 U19693 ( .B1(n18786), .B2(n16545), .A(n18784), .ZN(P3_U2636) );
  NOR3_X1 U19694 ( .A1(n16521), .A2(n16520), .A3(n16519), .ZN(n18637) );
  NOR2_X1 U19695 ( .A1(n18637), .A2(n18692), .ZN(n18831) );
  OAI21_X1 U19696 ( .B1(n18831), .B2(n18194), .A(n16522), .ZN(P3_U2637) );
  NOR4_X1 U19697 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_18__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16526) );
  NOR4_X1 U19698 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n16525) );
  NOR4_X1 U19699 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16524) );
  NOR4_X1 U19700 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16523) );
  NAND4_X1 U19701 ( .A1(n16526), .A2(n16525), .A3(n16524), .A4(n16523), .ZN(
        n16532) );
  NOR4_X1 U19702 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16530) );
  AOI211_X1 U19703 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_14__SCAN_IN), .B(
        P3_DATAWIDTH_REG_28__SCAN_IN), .ZN(n16529) );
  NOR4_X1 U19704 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16528) );
  NOR4_X1 U19705 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16527) );
  NAND4_X1 U19706 ( .A1(n16530), .A2(n16529), .A3(n16528), .A4(n16527), .ZN(
        n16531) );
  NOR2_X1 U19707 ( .A1(n16532), .A2(n16531), .ZN(n18829) );
  INV_X1 U19708 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18779) );
  NOR3_X1 U19709 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16534) );
  OAI21_X1 U19710 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16534), .A(n18829), .ZN(
        n16533) );
  OAI21_X1 U19711 ( .B1(n18829), .B2(n18779), .A(n16533), .ZN(P3_U2638) );
  INV_X1 U19712 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20926) );
  INV_X1 U19713 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18785) );
  AOI21_X1 U19714 ( .B1(n20926), .B2(n18785), .A(n16534), .ZN(n16535) );
  INV_X1 U19715 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20791) );
  INV_X1 U19716 ( .A(n18829), .ZN(n18824) );
  AOI22_X1 U19717 ( .A1(n18829), .A2(n16535), .B1(n20791), .B2(n18824), .ZN(
        P3_U2639) );
  NOR2_X2 U19718 ( .A1(n18789), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18569) );
  NAND2_X1 U19719 ( .A1(n18800), .A2(n18569), .ZN(n18685) );
  INV_X1 U19720 ( .A(n18685), .ZN(n18689) );
  NOR3_X1 U19721 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18694) );
  NAND2_X1 U19722 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18694), .ZN(n16889) );
  AOI211_X1 U19723 ( .C1(P3_STATE2_REG_0__SCAN_IN), .C2(n18689), .A(n16905), 
        .B(n18853), .ZN(n16539) );
  AOI211_X1 U19724 ( .C1(n18206), .C2(n18833), .A(n18837), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16541) );
  AOI211_X4 U19725 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18835), .A(n16541), .B(
        n16544), .ZN(n16928) );
  INV_X1 U19726 ( .A(n16541), .ZN(n18686) );
  INV_X1 U19727 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20745) );
  INV_X1 U19728 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18760) );
  INV_X1 U19729 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18756) );
  INV_X1 U19730 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18750) );
  INV_X1 U19731 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18740) );
  INV_X1 U19732 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18734) );
  INV_X1 U19733 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18723) );
  NOR2_X1 U19734 ( .A1(n20926), .A2(n18723), .ZN(n16895) );
  AND2_X1 U19735 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n16895), .ZN(n16870) );
  NAND3_X1 U19736 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n16870), .ZN(n16827) );
  NAND2_X1 U19737 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16835) );
  NOR3_X1 U19738 ( .A1(n18734), .A2(n16827), .A3(n16835), .ZN(n16793) );
  NAND4_X1 U19739 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16793), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16771) );
  NOR2_X1 U19740 ( .A1(n18740), .A2(n16771), .ZN(n16710) );
  NAND3_X1 U19741 ( .A1(n16710), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .ZN(n16744) );
  NAND2_X1 U19742 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16728) );
  NOR3_X1 U19743 ( .A1(n18750), .A2(n16744), .A3(n16728), .ZN(n16688) );
  NAND4_X1 U19744 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16688), .A3(
        P3_REIP_REG_18__SCAN_IN), .A4(P3_REIP_REG_19__SCAN_IN), .ZN(n16673) );
  NOR2_X1 U19745 ( .A1(n18756), .A2(n16673), .ZN(n16662) );
  NAND2_X1 U19746 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16662), .ZN(n16645) );
  NOR2_X1 U19747 ( .A1(n18760), .A2(n16645), .ZN(n16636) );
  NAND2_X1 U19748 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16636), .ZN(n16625) );
  NOR2_X1 U19749 ( .A1(n20745), .A2(n16625), .ZN(n16613) );
  NAND2_X1 U19750 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16613), .ZN(n16560) );
  NOR2_X1 U19751 ( .A1(n16921), .A2(n16560), .ZN(n16607) );
  NAND4_X1 U19752 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16607), .ZN(n16562) );
  NOR3_X1 U19753 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18775), .A3(n16562), 
        .ZN(n16542) );
  AOI21_X1 U19754 ( .B1(n16928), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16542), .ZN(
        n16568) );
  NAND2_X1 U19755 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18835), .ZN(n16543) );
  AOI211_X4 U19756 ( .C1(n16545), .C2(n18844), .A(n16544), .B(n16543), .ZN(
        n16927) );
  NOR3_X1 U19757 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16897) );
  INV_X1 U19758 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17210) );
  NAND2_X1 U19759 ( .A1(n16897), .A2(n17210), .ZN(n16880) );
  NAND2_X1 U19760 ( .A1(n16869), .A2(n17203), .ZN(n16855) );
  INV_X1 U19761 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17193) );
  NAND2_X1 U19762 ( .A1(n16846), .A2(n17193), .ZN(n16831) );
  NAND2_X1 U19763 ( .A1(n16821), .A2(n16811), .ZN(n16809) );
  NAND2_X1 U19764 ( .A1(n16801), .A2(n16790), .ZN(n16789) );
  NAND2_X1 U19765 ( .A1(n16769), .A2(n20779), .ZN(n16765) );
  INV_X1 U19766 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16739) );
  NAND2_X1 U19767 ( .A1(n16750), .A2(n16739), .ZN(n16737) );
  INV_X1 U19768 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17049) );
  NAND2_X1 U19769 ( .A1(n16724), .A2(n17049), .ZN(n16718) );
  INV_X1 U19770 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16694) );
  NAND2_X1 U19771 ( .A1(n16709), .A2(n16694), .ZN(n16693) );
  NAND2_X1 U19772 ( .A1(n16678), .A2(n17011), .ZN(n16668) );
  INV_X1 U19773 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U19774 ( .A1(n16656), .A2(n16966), .ZN(n16653) );
  INV_X1 U19775 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16631) );
  NAND2_X1 U19776 ( .A1(n16637), .A2(n16631), .ZN(n16630) );
  NOR2_X1 U19777 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16630), .ZN(n16614) );
  INV_X1 U19778 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16963) );
  NAND2_X1 U19779 ( .A1(n16614), .A2(n16963), .ZN(n16608) );
  NOR2_X1 U19780 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16608), .ZN(n16593) );
  INV_X1 U19781 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16959) );
  NAND2_X1 U19782 ( .A1(n16593), .A2(n16959), .ZN(n16570) );
  NOR2_X1 U19783 ( .A1(n16868), .A2(n16570), .ZN(n16578) );
  INV_X1 U19784 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16566) );
  INV_X1 U19785 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16548) );
  NAND2_X1 U19786 ( .A1(n16559), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16558) );
  AOI21_X1 U19787 ( .B1(n16548), .B2(n16558), .A(n16547), .ZN(n17496) );
  INV_X1 U19788 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16622) );
  NAND2_X1 U19789 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17525), .ZN(
        n17495) );
  AOI21_X1 U19790 ( .B1(n16622), .B2(n17495), .A(n16559), .ZN(n17526) );
  NOR2_X1 U19791 ( .A1(n17866), .A2(n17612), .ZN(n16686) );
  INV_X1 U19792 ( .A(n16686), .ZN(n17587) );
  NAND2_X1 U19793 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16552), .ZN(
        n16551) );
  NAND2_X1 U19794 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17535), .ZN(
        n16555) );
  XOR2_X1 U19795 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n16555), .Z(
        n17561) );
  INV_X1 U19796 ( .A(n17561), .ZN(n16640) );
  AOI21_X1 U19797 ( .B1(n16549), .B2(n16551), .A(n17535), .ZN(n17586) );
  INV_X1 U19798 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16923) );
  AND2_X1 U19799 ( .A1(n16686), .A2(n16923), .ZN(n16550) );
  AOI21_X1 U19800 ( .B1(n17611), .B2(n17587), .A(n16552), .ZN(n17615) );
  NOR2_X1 U19801 ( .A1(n16676), .A2(n9696), .ZN(n16667) );
  OAI21_X1 U19802 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16552), .A(
        n16551), .ZN(n16553) );
  INV_X1 U19803 ( .A(n16553), .ZN(n17601) );
  NOR2_X1 U19804 ( .A1(n16666), .A2(n9696), .ZN(n16658) );
  NOR2_X1 U19805 ( .A1(n17586), .A2(n16658), .ZN(n16657) );
  NOR2_X1 U19806 ( .A1(n16657), .A2(n9696), .ZN(n16647) );
  OAI21_X1 U19807 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17535), .A(
        n16555), .ZN(n16554) );
  INV_X1 U19808 ( .A(n16554), .ZN(n17568) );
  NOR2_X1 U19809 ( .A1(n16646), .A2(n9696), .ZN(n16639) );
  NOR2_X1 U19810 ( .A1(n16640), .A2(n16639), .ZN(n16638) );
  NOR2_X1 U19811 ( .A1(n16638), .A2(n9696), .ZN(n16624) );
  INV_X1 U19812 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16626) );
  INV_X1 U19813 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20938) );
  OR2_X1 U19814 ( .A1(n20938), .A2(n16555), .ZN(n16557) );
  INV_X1 U19815 ( .A(n17495), .ZN(n16556) );
  AOI21_X1 U19816 ( .B1(n16626), .B2(n16557), .A(n16556), .ZN(n17537) );
  NOR2_X1 U19817 ( .A1(n16623), .A2(n9696), .ZN(n16616) );
  NOR2_X1 U19818 ( .A1(n16615), .A2(n9696), .ZN(n16603) );
  OAI21_X1 U19819 ( .B1(n16559), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16558), .ZN(n17514) );
  INV_X1 U19820 ( .A(n17514), .ZN(n16604) );
  NOR2_X1 U19821 ( .A1(n16602), .A2(n9696), .ZN(n16595) );
  NOR2_X1 U19822 ( .A1(n17496), .A2(n16595), .ZN(n16594) );
  NOR2_X1 U19823 ( .A1(n16594), .A2(n9696), .ZN(n16582) );
  NOR2_X1 U19824 ( .A1(n16581), .A2(n9696), .ZN(n16573) );
  NAND2_X1 U19825 ( .A1(n16887), .A2(n16905), .ZN(n16914) );
  NOR3_X1 U19826 ( .A1(n16571), .A2(n16573), .A3(n16914), .ZN(n16565) );
  NAND3_X1 U19827 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16561) );
  AND2_X1 U19828 ( .A1(n16871), .A2(n16560), .ZN(n16612) );
  NOR2_X1 U19829 ( .A1(n16924), .A2(n16612), .ZN(n16611) );
  INV_X1 U19830 ( .A(n16611), .ZN(n16619) );
  AOI21_X1 U19831 ( .B1(n16871), .B2(n16561), .A(n16619), .ZN(n16592) );
  NOR2_X1 U19832 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16562), .ZN(n16576) );
  INV_X1 U19833 ( .A(n16576), .ZN(n16563) );
  AOI21_X1 U19834 ( .B1(n16592), .B2(n16563), .A(n18773), .ZN(n16564) );
  AOI211_X1 U19835 ( .C1(n16578), .C2(n16566), .A(n16565), .B(n16564), .ZN(
        n16567) );
  OAI211_X1 U19836 ( .C1(n16569), .C2(n16913), .A(n16568), .B(n16567), .ZN(
        P3_U2640) );
  NAND2_X1 U19837 ( .A1(n16927), .A2(n16570), .ZN(n16588) );
  OAI22_X1 U19838 ( .A1(n16592), .A2(n18775), .B1(n16574), .B2(n16913), .ZN(
        n16575) );
  OAI21_X1 U19839 ( .B1(n16928), .B2(n16578), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16579) );
  OAI211_X1 U19840 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16588), .A(n16580), .B(
        n16579), .ZN(P3_U2641) );
  INV_X1 U19841 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18770) );
  AOI211_X1 U19842 ( .C1(n16583), .C2(n16582), .A(n16581), .B(n16889), .ZN(
        n16587) );
  NAND3_X1 U19843 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16607), .ZN(n16585) );
  OAI22_X1 U19844 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16585), .B1(n16584), 
        .B2(n16913), .ZN(n16586) );
  AOI211_X1 U19845 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16928), .A(n16587), .B(
        n16586), .ZN(n16591) );
  INV_X1 U19846 ( .A(n16588), .ZN(n16589) );
  OAI21_X1 U19847 ( .B1(n16593), .B2(n16959), .A(n16589), .ZN(n16590) );
  OAI211_X1 U19848 ( .C1(n16592), .C2(n18770), .A(n16591), .B(n16590), .ZN(
        P3_U2642) );
  AOI22_X1 U19849 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16896), .B1(
        n16928), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16601) );
  AOI211_X1 U19850 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16608), .A(n16593), .B(
        n16868), .ZN(n16597) );
  AOI211_X1 U19851 ( .C1(n17496), .C2(n16595), .A(n16594), .B(n16889), .ZN(
        n16596) );
  AOI211_X1 U19852 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16619), .A(n16597), 
        .B(n16596), .ZN(n16600) );
  NAND2_X1 U19853 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16598) );
  OAI211_X1 U19854 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16607), .B(n16598), .ZN(n16599) );
  NAND3_X1 U19855 ( .A1(n16601), .A2(n16600), .A3(n16599), .ZN(P3_U2643) );
  INV_X1 U19856 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18767) );
  AOI211_X1 U19857 ( .C1(n16604), .C2(n16603), .A(n16602), .B(n16889), .ZN(
        n16606) );
  INV_X1 U19858 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17517) );
  OAI22_X1 U19859 ( .A1(n17517), .A2(n16913), .B1(n16915), .B2(n16963), .ZN(
        n16605) );
  AOI211_X1 U19860 ( .C1(n16607), .C2(n18767), .A(n16606), .B(n16605), .ZN(
        n16610) );
  OAI211_X1 U19861 ( .C1(n16614), .C2(n16963), .A(n16927), .B(n16608), .ZN(
        n16609) );
  OAI211_X1 U19862 ( .C1(n16611), .C2(n18767), .A(n16610), .B(n16609), .ZN(
        P3_U2644) );
  AOI22_X1 U19863 ( .A1(n16928), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16613), 
        .B2(n16612), .ZN(n16621) );
  AOI211_X1 U19864 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16630), .A(n16614), .B(
        n16868), .ZN(n16618) );
  AOI211_X1 U19865 ( .C1(n17526), .C2(n16616), .A(n16615), .B(n16889), .ZN(
        n16617) );
  AOI211_X1 U19866 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16619), .A(n16618), 
        .B(n16617), .ZN(n16620) );
  OAI211_X1 U19867 ( .C1(n16622), .C2(n16913), .A(n16621), .B(n16620), .ZN(
        P3_U2645) );
  INV_X1 U19868 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18762) );
  OAI21_X1 U19869 ( .B1(n16636), .B2(n16921), .A(n16922), .ZN(n16652) );
  AOI21_X1 U19870 ( .B1(n16871), .B2(n18762), .A(n16652), .ZN(n16634) );
  AOI211_X1 U19871 ( .C1(n17537), .C2(n16624), .A(n16623), .B(n16889), .ZN(
        n16629) );
  NOR3_X1 U19872 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16921), .A3(n16625), 
        .ZN(n16628) );
  OAI22_X1 U19873 ( .A1(n16626), .A2(n16913), .B1(n16915), .B2(n16631), .ZN(
        n16627) );
  NOR3_X1 U19874 ( .A1(n16629), .A2(n16628), .A3(n16627), .ZN(n16633) );
  OAI211_X1 U19875 ( .C1(n16637), .C2(n16631), .A(n16927), .B(n16630), .ZN(
        n16632) );
  OAI211_X1 U19876 ( .C1(n16634), .C2(n20745), .A(n16633), .B(n16632), .ZN(
        P3_U2646) );
  NOR2_X1 U19877 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16921), .ZN(n16635) );
  AOI22_X1 U19878 ( .A1(n16928), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16636), 
        .B2(n16635), .ZN(n16644) );
  AOI211_X1 U19879 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16653), .A(n16637), .B(
        n16868), .ZN(n16642) );
  AOI211_X1 U19880 ( .C1(n16640), .C2(n16639), .A(n16638), .B(n16889), .ZN(
        n16641) );
  AOI211_X1 U19881 ( .C1(n16652), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16642), 
        .B(n16641), .ZN(n16643) );
  OAI211_X1 U19882 ( .C1(n20938), .C2(n16913), .A(n16644), .B(n16643), .ZN(
        P3_U2647) );
  OAI21_X1 U19883 ( .B1(n16921), .B2(n16645), .A(n18760), .ZN(n16651) );
  AOI211_X1 U19884 ( .C1(n17568), .C2(n16647), .A(n16646), .B(n16889), .ZN(
        n16650) );
  INV_X1 U19885 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16648) );
  OAI22_X1 U19886 ( .A1(n16648), .A2(n16913), .B1(n16915), .B2(n16966), .ZN(
        n16649) );
  AOI211_X1 U19887 ( .C1(n16652), .C2(n16651), .A(n16650), .B(n16649), .ZN(
        n16655) );
  OAI211_X1 U19888 ( .C1(n16656), .C2(n16966), .A(n16927), .B(n16653), .ZN(
        n16654) );
  NAND2_X1 U19889 ( .A1(n16655), .A2(n16654), .ZN(P3_U2648) );
  AOI221_X1 U19890 ( .B1(n18756), .B2(n16871), .C1(n16673), .C2(n16871), .A(
        n16924), .ZN(n16665) );
  INV_X1 U19891 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18758) );
  AOI22_X1 U19892 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16896), .B1(
        n16928), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16664) );
  NOR2_X1 U19893 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16921), .ZN(n16661) );
  AOI211_X1 U19894 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16668), .A(n16656), .B(
        n16868), .ZN(n16660) );
  AOI211_X1 U19895 ( .C1(n17586), .C2(n16658), .A(n16657), .B(n16889), .ZN(
        n16659) );
  AOI211_X1 U19896 ( .C1(n16662), .C2(n16661), .A(n16660), .B(n16659), .ZN(
        n16663) );
  OAI211_X1 U19897 ( .C1(n16665), .C2(n18758), .A(n16664), .B(n16663), .ZN(
        P3_U2649) );
  AOI21_X1 U19898 ( .B1(n16673), .B2(n16871), .A(n16924), .ZN(n16685) );
  INV_X1 U19899 ( .A(n16685), .ZN(n16672) );
  AOI211_X1 U19900 ( .C1(n17601), .C2(n16667), .A(n16666), .B(n16889), .ZN(
        n16671) );
  INV_X1 U19901 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17597) );
  OAI211_X1 U19902 ( .C1(n16678), .C2(n17011), .A(n16927), .B(n16668), .ZN(
        n16669) );
  OAI21_X1 U19903 ( .B1(n16913), .B2(n17597), .A(n16669), .ZN(n16670) );
  AOI211_X1 U19904 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16672), .A(n16671), 
        .B(n16670), .ZN(n16675) );
  OR3_X1 U19905 ( .A1(n16921), .A2(n16673), .A3(P3_REIP_REG_21__SCAN_IN), .ZN(
        n16674) );
  OAI211_X1 U19906 ( .C1(n17011), .C2(n16915), .A(n16675), .B(n16674), .ZN(
        P3_U2650) );
  INV_X1 U19907 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18754) );
  AOI211_X1 U19908 ( .C1(n17615), .C2(n16677), .A(n16676), .B(n16889), .ZN(
        n16683) );
  AOI211_X1 U19909 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16693), .A(n16678), .B(
        n16868), .ZN(n16682) );
  INV_X1 U19910 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20902) );
  INV_X1 U19911 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18752) );
  NAND2_X1 U19912 ( .A1(n16871), .A2(n16688), .ZN(n16679) );
  NOR4_X1 U19913 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20902), .A3(n18752), 
        .A4(n16679), .ZN(n16681) );
  OAI22_X1 U19914 ( .A1(n17611), .A2(n16913), .B1(n16915), .B2(n16999), .ZN(
        n16680) );
  NOR4_X1 U19915 ( .A1(n16683), .A2(n16682), .A3(n16681), .A4(n16680), .ZN(
        n16684) );
  OAI21_X1 U19916 ( .B1(n16685), .B2(n18754), .A(n16684), .ZN(P3_U2651) );
  INV_X1 U19917 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16697) );
  INV_X1 U19918 ( .A(n16700), .ZN(n17629) );
  NOR2_X1 U19919 ( .A1(n17866), .A2(n17629), .ZN(n17621) );
  NAND2_X1 U19920 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17621), .ZN(
        n16699) );
  AOI21_X1 U19921 ( .B1(n16697), .B2(n16699), .A(n16686), .ZN(n17622) );
  CLKBUF_X1 U19922 ( .A(n16687), .Z(n17678) );
  NAND2_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17678), .ZN(
        n17664) );
  NOR2_X1 U19924 ( .A1(n17680), .A2(n17664), .ZN(n16732) );
  AOI21_X1 U19925 ( .B1(n16732), .B2(n16923), .A(n9696), .ZN(n16722) );
  AOI21_X1 U19926 ( .B1(n16887), .B2(n16699), .A(n16722), .ZN(n16702) );
  XNOR2_X1 U19927 ( .A(n17622), .B(n16702), .ZN(n16692) );
  OAI21_X1 U19928 ( .B1(n16921), .B2(n16688), .A(n16922), .ZN(n16706) );
  INV_X1 U19929 ( .A(n16706), .ZN(n16715) );
  NAND3_X1 U19930 ( .A1(n16688), .A2(n16871), .A3(n20902), .ZN(n16703) );
  AOI21_X1 U19931 ( .B1(n16715), .B2(n16703), .A(n18752), .ZN(n16691) );
  NAND4_X1 U19932 ( .A1(n16688), .A2(n16871), .A3(P3_REIP_REG_18__SCAN_IN), 
        .A4(n18752), .ZN(n16689) );
  OAI211_X1 U19933 ( .C1(n16915), .C2(n16694), .A(n18184), .B(n16689), .ZN(
        n16690) );
  AOI211_X1 U19934 ( .C1(n16905), .C2(n16692), .A(n16691), .B(n16690), .ZN(
        n16696) );
  OAI211_X1 U19935 ( .C1(n16709), .C2(n16694), .A(n16927), .B(n16693), .ZN(
        n16695) );
  OAI211_X1 U19936 ( .C1(n16913), .C2(n16697), .A(n16696), .B(n16695), .ZN(
        P3_U2652) );
  AOI21_X1 U19937 ( .B1(n16718), .B2(P3_EBX_REG_18__SCAN_IN), .A(n16868), .ZN(
        n16698) );
  AOI21_X1 U19938 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16928), .A(n16698), .ZN(
        n16708) );
  OAI21_X1 U19939 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17621), .A(
        n16699), .ZN(n17639) );
  NAND2_X1 U19940 ( .A1(n16905), .A2(n9696), .ZN(n16909) );
  NOR2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17866), .ZN(
        n16906) );
  OAI221_X1 U19942 ( .B1(n17639), .B2(n16700), .C1(n17639), .C2(n16906), .A(
        n16905), .ZN(n16701) );
  AOI22_X1 U19943 ( .A1(n16702), .A2(n17639), .B1(n16909), .B2(n16701), .ZN(
        n16705) );
  INV_X1 U19944 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17642) );
  OAI211_X1 U19945 ( .C1(n17642), .C2(n16913), .A(n18184), .B(n16703), .ZN(
        n16704) );
  AOI211_X1 U19946 ( .C1(n16706), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16705), 
        .B(n16704), .ZN(n16707) );
  OAI21_X1 U19947 ( .B1(n16709), .B2(n16708), .A(n16707), .ZN(P3_U2653) );
  INV_X1 U19948 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18744) );
  INV_X1 U19949 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18741) );
  NAND2_X1 U19950 ( .A1(n16871), .A2(n16710), .ZN(n16761) );
  NOR3_X1 U19951 ( .A1(n18744), .A2(n18741), .A3(n16761), .ZN(n16729) );
  INV_X1 U19952 ( .A(n16729), .ZN(n16743) );
  OAI21_X1 U19953 ( .B1(n16728), .B2(n16743), .A(n18750), .ZN(n16711) );
  INV_X1 U19954 ( .A(n16711), .ZN(n16716) );
  INV_X1 U19955 ( .A(n17664), .ZN(n16712) );
  NAND2_X1 U19956 ( .A1(n17667), .A2(n16712), .ZN(n16721) );
  AOI21_X1 U19957 ( .B1(n17651), .B2(n16721), .A(n17621), .ZN(n17655) );
  NOR2_X1 U19958 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17664), .ZN(
        n16733) );
  AOI21_X1 U19959 ( .B1(n17667), .B2(n16733), .A(n9696), .ZN(n16713) );
  XNOR2_X1 U19960 ( .A(n17655), .B(n16713), .ZN(n16714) );
  OAI22_X1 U19961 ( .A1(n16716), .A2(n16715), .B1(n16889), .B2(n16714), .ZN(
        n16717) );
  AOI211_X1 U19962 ( .C1(n16928), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18186), .B(
        n16717), .ZN(n16720) );
  OAI211_X1 U19963 ( .C1(n16724), .C2(n17049), .A(n16927), .B(n16718), .ZN(
        n16719) );
  OAI211_X1 U19964 ( .C1(n16913), .C2(n17651), .A(n16720), .B(n16719), .ZN(
        P3_U2654) );
  AOI21_X1 U19965 ( .B1(n16871), .B2(n16744), .A(n16924), .ZN(n16755) );
  INV_X1 U19966 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18747) );
  OAI21_X1 U19967 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16732), .A(
        n16721), .ZN(n17668) );
  INV_X1 U19968 ( .A(n17668), .ZN(n16723) );
  INV_X1 U19969 ( .A(n16722), .ZN(n16735) );
  AOI221_X1 U19970 ( .B1(n16723), .B2(n16722), .C1(n17668), .C2(n16735), .A(
        n16889), .ZN(n16727) );
  AOI211_X1 U19971 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16737), .A(n16724), .B(
        n16868), .ZN(n16726) );
  INV_X1 U19972 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17076) );
  OAI22_X1 U19973 ( .A1(n17665), .A2(n16913), .B1(n16915), .B2(n17076), .ZN(
        n16725) );
  NOR4_X1 U19974 ( .A1(n18186), .A2(n16727), .A3(n16726), .A4(n16725), .ZN(
        n16731) );
  OAI211_X1 U19975 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16729), .B(n16728), .ZN(n16730) );
  OAI211_X1 U19976 ( .C1(n16755), .C2(n18747), .A(n16731), .B(n16730), .ZN(
        P3_U2655) );
  INV_X1 U19977 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18745) );
  AOI21_X1 U19978 ( .B1(n17680), .B2(n17664), .A(n16732), .ZN(n17686) );
  INV_X1 U19979 ( .A(n17686), .ZN(n16736) );
  OAI21_X1 U19980 ( .B1(n16733), .B2(n16736), .A(n16905), .ZN(n16734) );
  AOI22_X1 U19981 ( .A1(n16736), .A2(n16735), .B1(n16909), .B2(n16734), .ZN(
        n16741) );
  OAI211_X1 U19982 ( .C1(n16750), .C2(n16739), .A(n16927), .B(n16737), .ZN(
        n16738) );
  OAI211_X1 U19983 ( .C1(n16915), .C2(n16739), .A(n18184), .B(n16738), .ZN(
        n16740) );
  AOI211_X1 U19984 ( .C1(n16896), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16741), .B(n16740), .ZN(n16742) );
  OAI221_X1 U19985 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16743), .C1(n18745), 
        .C2(n16755), .A(n16742), .ZN(P3_U2656) );
  INV_X1 U19986 ( .A(n16744), .ZN(n16745) );
  NOR3_X1 U19987 ( .A1(n16745), .A2(n16761), .A3(n18741), .ZN(n16746) );
  AOI211_X1 U19988 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n16896), .A(
        n18186), .B(n16746), .ZN(n16754) );
  NAND2_X1 U19989 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17708), .ZN(
        n17704) );
  NOR2_X1 U19990 ( .A1(n17709), .A2(n17704), .ZN(n16756) );
  OAI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16756), .A(
        n17664), .ZN(n17702) );
  INV_X1 U19992 ( .A(n16906), .ZN(n16865) );
  OAI21_X1 U19993 ( .B1(n17691), .B2(n16865), .A(n16887), .ZN(n16749) );
  OAI21_X1 U19994 ( .B1(n17702), .B2(n16749), .A(n16905), .ZN(n16748) );
  AOI21_X1 U19995 ( .B1(n17702), .B2(n16749), .A(n16748), .ZN(n16752) );
  AOI211_X1 U19996 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16765), .A(n16750), .B(
        n16868), .ZN(n16751) );
  AOI211_X1 U19997 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16928), .A(n16752), .B(
        n16751), .ZN(n16753) );
  OAI211_X1 U19998 ( .C1(n18744), .C2(n16755), .A(n16754), .B(n16753), .ZN(
        P3_U2657) );
  INV_X1 U19999 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16768) );
  AOI21_X1 U20000 ( .B1(n16871), .B2(n16771), .A(n16924), .ZN(n16787) );
  NAND2_X1 U20001 ( .A1(n16871), .A2(n18740), .ZN(n16770) );
  AOI21_X1 U20002 ( .B1(n16787), .B2(n16770), .A(n18741), .ZN(n16764) );
  INV_X1 U20003 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20733) );
  NOR2_X1 U20004 ( .A1(n20733), .A2(n17704), .ZN(n16758) );
  INV_X1 U20005 ( .A(n16756), .ZN(n16757) );
  OAI21_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16758), .A(
        n16757), .ZN(n17711) );
  INV_X1 U20007 ( .A(n16758), .ZN(n16773) );
  OAI21_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16773), .A(
        n16887), .ZN(n16760) );
  OAI21_X1 U20009 ( .B1(n17711), .B2(n16760), .A(n16905), .ZN(n16759) );
  AOI21_X1 U20010 ( .B1(n17711), .B2(n16760), .A(n16759), .ZN(n16763) );
  OAI22_X1 U20011 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16761), .B1(n16915), 
        .B2(n20779), .ZN(n16762) );
  NOR4_X1 U20012 ( .A1(n18186), .A2(n16764), .A3(n16763), .A4(n16762), .ZN(
        n16767) );
  OAI211_X1 U20013 ( .C1(n16769), .C2(n20779), .A(n16927), .B(n16765), .ZN(
        n16766) );
  OAI211_X1 U20014 ( .C1(n16913), .C2(n16768), .A(n16767), .B(n16766), .ZN(
        P3_U2658) );
  AOI211_X1 U20015 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16789), .A(n16769), .B(
        n16868), .ZN(n16777) );
  INV_X1 U20016 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16772) );
  OAI22_X1 U20017 ( .A1(n16915), .A2(n16772), .B1(n16771), .B2(n16770), .ZN(
        n16776) );
  INV_X1 U20018 ( .A(n17704), .ZN(n16779) );
  OAI21_X1 U20019 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16779), .A(
        n16773), .ZN(n17721) );
  OAI21_X1 U20020 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16773), .A(
        n17721), .ZN(n16774) );
  OAI22_X1 U20021 ( .A1(n20733), .A2(n16913), .B1(n16914), .B2(n16774), .ZN(
        n16775) );
  NOR4_X1 U20022 ( .A1(n18186), .A2(n16777), .A3(n16776), .A4(n16775), .ZN(
        n16781) );
  INV_X1 U20023 ( .A(n17721), .ZN(n16778) );
  AOI21_X1 U20024 ( .B1(n16887), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16889), .ZN(n16918) );
  OAI211_X1 U20025 ( .C1(n16779), .C2(n9696), .A(n16778), .B(n16918), .ZN(
        n16780) );
  OAI211_X1 U20026 ( .C1(n16787), .C2(n18740), .A(n16781), .B(n16780), .ZN(
        P3_U2659) );
  INV_X1 U20027 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18736) );
  INV_X1 U20028 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18735) );
  NOR2_X1 U20029 ( .A1(n18736), .A2(n18735), .ZN(n16795) );
  NAND2_X1 U20030 ( .A1(n16871), .A2(n16793), .ZN(n16812) );
  INV_X1 U20031 ( .A(n16812), .ZN(n16782) );
  AOI21_X1 U20032 ( .B1(n16795), .B2(n16782), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16786) );
  INV_X1 U20033 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16798) );
  CLKBUF_X1 U20034 ( .A(n16783), .Z(n17785) );
  NAND3_X1 U20035 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17785), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16828) );
  NOR2_X1 U20036 ( .A1(n17774), .A2(n16828), .ZN(n16817) );
  NAND2_X1 U20037 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16817), .ZN(
        n16806) );
  NOR2_X1 U20038 ( .A1(n16798), .A2(n16806), .ZN(n16797) );
  AOI21_X1 U20039 ( .B1(n16797), .B2(n16923), .A(n9696), .ZN(n16784) );
  OAI21_X1 U20040 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16797), .A(
        n17704), .ZN(n17735) );
  XOR2_X1 U20041 ( .A(n16784), .B(n17735), .Z(n16785) );
  OAI22_X1 U20042 ( .A1(n16787), .A2(n16786), .B1(n16889), .B2(n16785), .ZN(
        n16788) );
  AOI211_X1 U20043 ( .C1(n16928), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18186), .B(
        n16788), .ZN(n16792) );
  OAI211_X1 U20044 ( .C1(n16801), .C2(n16790), .A(n16927), .B(n16789), .ZN(
        n16791) );
  OAI211_X1 U20045 ( .C1(n16913), .C2(n17737), .A(n16792), .B(n16791), .ZN(
        P3_U2660) );
  OAI21_X1 U20046 ( .B1(n16921), .B2(n16793), .A(n16922), .ZN(n16794) );
  INV_X1 U20047 ( .A(n16794), .ZN(n16820) );
  AOI211_X1 U20048 ( .C1(n18736), .C2(n18735), .A(n16795), .B(n16812), .ZN(
        n16796) );
  AOI211_X1 U20049 ( .C1(n16928), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18186), .B(
        n16796), .ZN(n16805) );
  AOI21_X1 U20050 ( .B1(n16798), .B2(n16806), .A(n16797), .ZN(n17752) );
  OAI21_X1 U20051 ( .B1(n16806), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16887), .ZN(n16808) );
  INV_X1 U20052 ( .A(n16808), .ZN(n16800) );
  OAI21_X1 U20053 ( .B1(n17752), .B2(n16800), .A(n16905), .ZN(n16799) );
  AOI21_X1 U20054 ( .B1(n17752), .B2(n16800), .A(n16799), .ZN(n16803) );
  AOI211_X1 U20055 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16809), .A(n16801), .B(
        n16868), .ZN(n16802) );
  AOI211_X1 U20056 ( .C1(n16896), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16803), .B(n16802), .ZN(n16804) );
  OAI211_X1 U20057 ( .C1(n16820), .C2(n18736), .A(n16805), .B(n16804), .ZN(
        P3_U2661) );
  OAI21_X1 U20058 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16817), .A(
        n16806), .ZN(n17762) );
  NAND2_X1 U20059 ( .A1(n17785), .A2(n16906), .ZN(n16842) );
  NOR2_X1 U20060 ( .A1(n17787), .A2(n16842), .ZN(n16818) );
  OAI221_X1 U20061 ( .B1(n17762), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(
        n17762), .C2(n16818), .A(n16905), .ZN(n16807) );
  AOI22_X1 U20062 ( .A1(n17762), .A2(n16808), .B1(n16909), .B2(n16807), .ZN(
        n16815) );
  OAI211_X1 U20063 ( .C1(n16821), .C2(n16811), .A(n16927), .B(n16809), .ZN(
        n16810) );
  OAI21_X1 U20064 ( .B1(n16811), .B2(n16915), .A(n16810), .ZN(n16814) );
  INV_X1 U20065 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17760) );
  OAI22_X1 U20066 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16812), .B1(n17760), 
        .B2(n16913), .ZN(n16813) );
  NOR4_X1 U20067 ( .A1(n18186), .A2(n16815), .A3(n16814), .A4(n16813), .ZN(
        n16816) );
  OAI21_X1 U20068 ( .B1(n16820), .B2(n18735), .A(n16816), .ZN(P3_U2662) );
  AOI21_X1 U20069 ( .B1(n17774), .B2(n16828), .A(n16817), .ZN(n17778) );
  NOR2_X1 U20070 ( .A1(n16818), .A2(n9696), .ZN(n16819) );
  XNOR2_X1 U20071 ( .A(n17778), .B(n16819), .ZN(n16826) );
  AOI21_X1 U20072 ( .B1(n16928), .B2(P3_EBX_REG_8__SCAN_IN), .A(n18186), .ZN(
        n16825) );
  NAND4_X1 U20073 ( .A1(n16871), .A2(P3_REIP_REG_5__SCAN_IN), .A3(
        P3_REIP_REG_4__SCAN_IN), .A4(n16870), .ZN(n16851) );
  AOI221_X1 U20074 ( .B1(n16835), .B2(n18734), .C1(n16851), .C2(n18734), .A(
        n16820), .ZN(n16823) );
  AOI211_X1 U20075 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16831), .A(n16821), .B(
        n16868), .ZN(n16822) );
  AOI211_X1 U20076 ( .C1(n16896), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16823), .B(n16822), .ZN(n16824) );
  OAI211_X1 U20077 ( .C1(n16889), .C2(n16826), .A(n16825), .B(n16824), .ZN(
        P3_U2663) );
  AOI21_X1 U20078 ( .B1(n16871), .B2(n16827), .A(n16924), .ZN(n16853) );
  INV_X1 U20079 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18731) );
  NOR2_X1 U20080 ( .A1(n17866), .A2(n17801), .ZN(n16852) );
  INV_X1 U20081 ( .A(n16852), .ZN(n16840) );
  NOR2_X1 U20082 ( .A1(n17808), .A2(n16840), .ZN(n16839) );
  OAI21_X1 U20083 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16839), .A(
        n16828), .ZN(n17797) );
  NAND2_X1 U20084 ( .A1(n16887), .A2(n16842), .ZN(n16830) );
  OAI21_X1 U20085 ( .B1(n17797), .B2(n16830), .A(n16905), .ZN(n16829) );
  AOI21_X1 U20086 ( .B1(n17797), .B2(n16830), .A(n16829), .ZN(n16834) );
  OAI211_X1 U20087 ( .C1(n16846), .C2(n17193), .A(n16927), .B(n16831), .ZN(
        n16832) );
  OAI211_X1 U20088 ( .C1(n16915), .C2(n17193), .A(n18184), .B(n16832), .ZN(
        n16833) );
  AOI211_X1 U20089 ( .C1(n16896), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16834), .B(n16833), .ZN(n16838) );
  INV_X1 U20090 ( .A(n16851), .ZN(n16836) );
  OAI211_X1 U20091 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16836), .B(n16835), .ZN(n16837) );
  OAI211_X1 U20092 ( .C1(n16853), .C2(n18731), .A(n16838), .B(n16837), .ZN(
        P3_U2664) );
  INV_X1 U20093 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18729) );
  AOI21_X1 U20094 ( .B1(n17808), .B2(n16840), .A(n16839), .ZN(n17805) );
  OAI21_X1 U20095 ( .B1(n16852), .B2(n9696), .A(n16918), .ZN(n16845) );
  INV_X1 U20096 ( .A(n17805), .ZN(n16844) );
  INV_X1 U20097 ( .A(n16842), .ZN(n16843) );
  AOI221_X1 U20098 ( .B1(n17805), .B2(n16845), .C1(n16844), .C2(n16914), .A(
        n16843), .ZN(n16849) );
  AOI211_X1 U20099 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16855), .A(n16846), .B(
        n16868), .ZN(n16848) );
  INV_X1 U20100 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17192) );
  OAI22_X1 U20101 ( .A1(n17808), .A2(n16913), .B1(n16915), .B2(n17192), .ZN(
        n16847) );
  NOR4_X1 U20102 ( .A1(n18186), .A2(n16849), .A3(n16848), .A4(n16847), .ZN(
        n16850) );
  OAI221_X1 U20103 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16851), .C1(n18729), 
        .C2(n16853), .A(n16850), .ZN(P3_U2665) );
  INV_X1 U20104 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U20105 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17809), .ZN(
        n16862) );
  AOI21_X1 U20106 ( .B1(n16857), .B2(n16862), .A(n16852), .ZN(n17816) );
  OAI21_X1 U20107 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16862), .A(
        n16887), .ZN(n16866) );
  XNOR2_X1 U20108 ( .A(n17816), .B(n16866), .ZN(n16860) );
  INV_X1 U20109 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20797) );
  NAND3_X1 U20110 ( .A1(n16871), .A2(P3_REIP_REG_4__SCAN_IN), .A3(n16870), 
        .ZN(n16854) );
  AOI21_X1 U20111 ( .B1(n20797), .B2(n16854), .A(n16853), .ZN(n16859) );
  OAI211_X1 U20112 ( .C1(n16869), .C2(n17203), .A(n16927), .B(n16855), .ZN(
        n16856) );
  OAI21_X1 U20113 ( .B1(n16913), .B2(n16857), .A(n16856), .ZN(n16858) );
  AOI211_X1 U20114 ( .C1(n16905), .C2(n16860), .A(n16859), .B(n16858), .ZN(
        n16861) );
  OAI211_X1 U20115 ( .C1(n16915), .C2(n17203), .A(n16861), .B(n18184), .ZN(
        P3_U2666) );
  NOR2_X1 U20116 ( .A1(n16870), .A2(n16921), .ZN(n16884) );
  NOR2_X1 U20117 ( .A1(n16924), .A2(n16884), .ZN(n16893) );
  INV_X1 U20118 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18727) );
  NAND2_X1 U20119 ( .A1(n18203), .A2(n18853), .ZN(n18856) );
  AOI21_X1 U20120 ( .B1(n16878), .B2(n18640), .A(n18856), .ZN(n16864) );
  NOR2_X1 U20121 ( .A1(n17866), .A2(n17828), .ZN(n16885) );
  OAI21_X1 U20122 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16885), .A(
        n16862), .ZN(n17831) );
  OAI22_X1 U20123 ( .A1(n17830), .A2(n16913), .B1(n17831), .B2(n16909), .ZN(
        n16863) );
  NOR3_X1 U20124 ( .A1(n18186), .A2(n16864), .A3(n16863), .ZN(n16877) );
  INV_X1 U20125 ( .A(n17831), .ZN(n16867) );
  OR2_X1 U20126 ( .A1(n17828), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17835) );
  OAI22_X1 U20127 ( .A1(n16867), .A2(n16866), .B1(n16865), .B2(n17835), .ZN(
        n16875) );
  AOI211_X1 U20128 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16880), .A(n16869), .B(
        n16868), .ZN(n16874) );
  NAND2_X1 U20129 ( .A1(n16871), .A2(n16870), .ZN(n16872) );
  INV_X1 U20130 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20716) );
  OAI22_X1 U20131 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16872), .B1(n16915), 
        .B2(n20716), .ZN(n16873) );
  AOI211_X1 U20132 ( .C1(n16905), .C2(n16875), .A(n16874), .B(n16873), .ZN(
        n16876) );
  OAI211_X1 U20133 ( .C1(n16893), .C2(n18727), .A(n16877), .B(n16876), .ZN(
        P3_U2667) );
  INV_X1 U20134 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18725) );
  INV_X1 U20135 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16886) );
  OAI22_X1 U20136 ( .A1(n16886), .A2(n16913), .B1(n16915), .B2(n17210), .ZN(
        n16883) );
  NOR2_X1 U20137 ( .A1(n12634), .A2(n18807), .ZN(n18658) );
  INV_X1 U20138 ( .A(n18658), .ZN(n18643) );
  NOR2_X1 U20139 ( .A1(n18821), .A2(n18643), .ZN(n16879) );
  OAI21_X1 U20140 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16879), .A(
        n16878), .ZN(n18793) );
  OAI211_X1 U20141 ( .C1(n16897), .C2(n17210), .A(n16927), .B(n16880), .ZN(
        n16881) );
  OAI21_X1 U20142 ( .B1(n18856), .B2(n18793), .A(n16881), .ZN(n16882) );
  AOI211_X1 U20143 ( .C1(n16895), .C2(n16884), .A(n16883), .B(n16882), .ZN(
        n16892) );
  NAND2_X1 U20144 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16894) );
  AOI21_X1 U20145 ( .B1(n16886), .B2(n16894), .A(n16885), .ZN(n17845) );
  OAI21_X1 U20146 ( .B1(n16894), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16887), .ZN(n16888) );
  INV_X1 U20147 ( .A(n16888), .ZN(n16904) );
  AOI21_X1 U20148 ( .B1(n17845), .B2(n16904), .A(n16889), .ZN(n16890) );
  OAI21_X1 U20149 ( .B1(n17845), .B2(n16904), .A(n16890), .ZN(n16891) );
  OAI211_X1 U20150 ( .C1(n16893), .C2(n18725), .A(n16892), .B(n16891), .ZN(
        P3_U2668) );
  OAI21_X1 U20151 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16894), .ZN(n17854) );
  AOI211_X1 U20152 ( .C1(n20926), .C2(n18723), .A(n16895), .B(n16921), .ZN(
        n16903) );
  NAND2_X1 U20153 ( .A1(n18807), .A2(n18657), .ZN(n18641) );
  OAI21_X1 U20154 ( .B1(n18821), .B2(n18643), .A(n18641), .ZN(n18801) );
  AOI22_X1 U20155 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16896), .B1(
        n16924), .B2(P3_REIP_REG_2__SCAN_IN), .ZN(n16901) );
  NOR2_X1 U20156 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16912) );
  INV_X1 U20157 ( .A(n16897), .ZN(n16898) );
  OAI211_X1 U20158 ( .C1(n16912), .C2(n16899), .A(n16927), .B(n16898), .ZN(
        n16900) );
  OAI211_X1 U20159 ( .C1(n18856), .C2(n18801), .A(n16901), .B(n16900), .ZN(
        n16902) );
  AOI211_X1 U20160 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16928), .A(n16903), .B(
        n16902), .ZN(n16908) );
  OAI211_X1 U20161 ( .C1(n16906), .C2(n17854), .A(n16905), .B(n16904), .ZN(
        n16907) );
  OAI211_X1 U20162 ( .C1(n16909), .C2(n17854), .A(n16908), .B(n16907), .ZN(
        P3_U2669) );
  NAND2_X1 U20163 ( .A1(n18657), .A2(n16910), .ZN(n18808) );
  INV_X1 U20164 ( .A(n16911), .ZN(n17218) );
  NOR2_X1 U20165 ( .A1(n16912), .A2(n17218), .ZN(n17223) );
  AOI22_X1 U20166 ( .A1(n16927), .A2(n17223), .B1(n16924), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n16920) );
  OAI21_X1 U20167 ( .B1(n16923), .B2(n16914), .A(n16913), .ZN(n16917) );
  INV_X1 U20168 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17226) );
  OAI22_X1 U20169 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16921), .B1(n16915), 
        .B2(n17226), .ZN(n16916) );
  AOI221_X1 U20170 ( .B1(n16918), .B2(n17866), .C1(n16917), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16916), .ZN(n16919) );
  OAI211_X1 U20171 ( .C1(n18808), .C2(n18856), .A(n16920), .B(n16919), .ZN(
        P3_U2670) );
  NAND2_X1 U20172 ( .A1(n16922), .A2(n16921), .ZN(n16926) );
  NOR2_X1 U20173 ( .A1(n16924), .A2(n16923), .ZN(n16925) );
  AOI22_X1 U20174 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16926), .B1(n16925), 
        .B2(n18803), .ZN(n16930) );
  OAI21_X1 U20175 ( .B1(n16928), .B2(n16927), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16929) );
  OAI211_X1 U20176 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18856), .A(
        n16930), .B(n16929), .ZN(P3_U2671) );
  AOI22_X1 U20177 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20178 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20179 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20180 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16931) );
  NAND4_X1 U20181 ( .A1(n16934), .A2(n16933), .A3(n16932), .A4(n16931), .ZN(
        n16940) );
  AOI22_X1 U20182 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20183 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20184 ( .A1(n15746), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20185 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16935) );
  NAND4_X1 U20186 ( .A1(n16938), .A2(n16937), .A3(n16936), .A4(n16935), .ZN(
        n16939) );
  NOR2_X1 U20187 ( .A1(n16940), .A2(n16939), .ZN(n16951) );
  AOI22_X1 U20188 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16950) );
  AOI22_X1 U20189 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20190 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16941) );
  OAI21_X1 U20191 ( .B1(n9791), .B2(n20874), .A(n16941), .ZN(n16947) );
  AOI22_X1 U20192 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20193 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20194 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20195 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16942) );
  NAND4_X1 U20196 ( .A1(n16945), .A2(n16944), .A3(n16943), .A4(n16942), .ZN(
        n16946) );
  AOI211_X1 U20197 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16947), .B(n16946), .ZN(n16948) );
  NAND3_X1 U20198 ( .A1(n16950), .A2(n16949), .A3(n16948), .ZN(n16956) );
  NAND2_X1 U20199 ( .A1(n16957), .A2(n16956), .ZN(n16955) );
  XNOR2_X1 U20200 ( .A(n16951), .B(n16955), .ZN(n17242) );
  NOR2_X1 U20201 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16952), .ZN(n16954) );
  OAI22_X1 U20202 ( .A1(n17242), .A2(n17221), .B1(n16954), .B2(n16953), .ZN(
        P3_U2673) );
  OAI21_X1 U20203 ( .B1(n16957), .B2(n16956), .A(n16955), .ZN(n17247) );
  OAI222_X1 U20204 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16969), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n16960), .C1(n16959), .C2(n16958), .ZN(
        n16961) );
  OAI21_X1 U20205 ( .B1(n17247), .B2(n17221), .A(n16961), .ZN(P3_U2674) );
  OAI211_X1 U20206 ( .C1(n17254), .C2(n17253), .A(n17229), .B(n17252), .ZN(
        n16962) );
  OAI221_X1 U20207 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16964), .C1(n16963), 
        .C2(n16967), .A(n16962), .ZN(P3_U2676) );
  XNOR2_X1 U20208 ( .A(n16965), .B(n16971), .ZN(n17262) );
  NAND3_X1 U20209 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n16984), .ZN(n16970) );
  INV_X1 U20210 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16968) );
  OAI222_X1 U20211 ( .A1(n17262), .A2(n17221), .B1(n16970), .B2(n16969), .C1(
        n16968), .C2(n16967), .ZN(P3_U2677) );
  INV_X1 U20212 ( .A(n16970), .ZN(n16975) );
  AOI22_X1 U20213 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17221), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n16984), .ZN(n16974) );
  OAI21_X1 U20214 ( .B1(n16973), .B2(n16972), .A(n16971), .ZN(n17267) );
  OAI22_X1 U20215 ( .A1(n16975), .A2(n16974), .B1(n17221), .B2(n17267), .ZN(
        P3_U2678) );
  INV_X1 U20216 ( .A(n16984), .ZN(n16978) );
  XNOR2_X1 U20217 ( .A(n16976), .B(n16980), .ZN(n17272) );
  NAND3_X1 U20218 ( .A1(n16978), .A2(P3_EBX_REG_24__SCAN_IN), .A3(n17221), 
        .ZN(n16977) );
  OAI221_X1 U20219 ( .B1(n16978), .B2(P3_EBX_REG_24__SCAN_IN), .C1(n17221), 
        .C2(n17272), .A(n16977), .ZN(P3_U2679) );
  INV_X1 U20220 ( .A(n16979), .ZN(n16998) );
  AOI21_X1 U20221 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17221), .A(n16998), .ZN(
        n16983) );
  OAI21_X1 U20222 ( .B1(n16982), .B2(n16981), .A(n16980), .ZN(n17277) );
  OAI22_X1 U20223 ( .A1(n16984), .A2(n16983), .B1(n17221), .B2(n17277), .ZN(
        P3_U2680) );
  AOI21_X1 U20224 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17221), .A(n16985), .ZN(
        n16997) );
  AOI22_X1 U20225 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20226 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20227 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16986) );
  OAI21_X1 U20228 ( .B1(n12410), .B2(n20874), .A(n16986), .ZN(n16992) );
  AOI22_X1 U20229 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20230 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20231 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20232 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16987) );
  NAND4_X1 U20233 ( .A1(n16990), .A2(n16989), .A3(n16988), .A4(n16987), .ZN(
        n16991) );
  AOI211_X1 U20234 ( .C1(n17181), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n16992), .B(n16991), .ZN(n16993) );
  NAND3_X1 U20235 ( .A1(n16995), .A2(n16994), .A3(n16993), .ZN(n17278) );
  INV_X1 U20236 ( .A(n17278), .ZN(n16996) );
  OAI22_X1 U20237 ( .A1(n16998), .A2(n16997), .B1(n16996), .B2(n17221), .ZN(
        P3_U2681) );
  OAI21_X1 U20238 ( .B1(n16999), .B2(n17036), .A(n17221), .ZN(n17024) );
  AOI22_X1 U20239 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20240 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20241 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20242 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17000) );
  NAND4_X1 U20243 ( .A1(n17003), .A2(n17002), .A3(n17001), .A4(n17000), .ZN(
        n17009) );
  AOI22_X1 U20244 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20245 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20246 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20247 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17004) );
  NAND4_X1 U20248 ( .A1(n17007), .A2(n17006), .A3(n17005), .A4(n17004), .ZN(
        n17008) );
  NOR2_X1 U20249 ( .A1(n17009), .A2(n17008), .ZN(n17287) );
  OR2_X1 U20250 ( .A1(n17287), .A2(n17221), .ZN(n17010) );
  OAI221_X1 U20251 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17012), .C1(n17011), 
        .C2(n17024), .A(n17010), .ZN(P3_U2682) );
  AOI22_X1 U20252 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20253 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20254 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20255 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17013) );
  NAND4_X1 U20256 ( .A1(n17016), .A2(n17015), .A3(n17014), .A4(n17013), .ZN(
        n17022) );
  AOI22_X1 U20257 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20258 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20259 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20260 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17017) );
  NAND4_X1 U20261 ( .A1(n17020), .A2(n17019), .A3(n17018), .A4(n17017), .ZN(
        n17021) );
  NOR2_X1 U20262 ( .A1(n17022), .A2(n17021), .ZN(n17294) );
  NOR2_X1 U20263 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17023), .ZN(n17025) );
  OAI22_X1 U20264 ( .A1(n17294), .A2(n17221), .B1(n17025), .B2(n17024), .ZN(
        P3_U2683) );
  AOI22_X1 U20265 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20266 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20267 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20268 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17026) );
  NAND4_X1 U20269 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17035) );
  AOI22_X1 U20270 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20271 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20272 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20273 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17030) );
  NAND4_X1 U20274 ( .A1(n17033), .A2(n17032), .A3(n17031), .A4(n17030), .ZN(
        n17034) );
  NOR2_X1 U20275 ( .A1(n17035), .A2(n17034), .ZN(n17300) );
  OAI21_X1 U20276 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17050), .A(n17036), .ZN(
        n17037) );
  AOI22_X1 U20277 ( .A1(n17229), .A2(n17300), .B1(n17037), .B2(n17221), .ZN(
        P3_U2684) );
  AOI22_X1 U20278 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20279 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20280 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20281 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17038) );
  NAND4_X1 U20282 ( .A1(n17041), .A2(n17040), .A3(n17039), .A4(n17038), .ZN(
        n17047) );
  AOI22_X1 U20283 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20284 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20285 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20286 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U20287 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17046) );
  NOR2_X1 U20288 ( .A1(n17047), .A2(n17046), .ZN(n17304) );
  NOR3_X1 U20289 ( .A1(n17280), .A2(n17119), .A3(n17048), .ZN(n17077) );
  NAND2_X1 U20290 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17077), .ZN(n17065) );
  NOR2_X1 U20291 ( .A1(n17049), .A2(n17065), .ZN(n17052) );
  NOR2_X1 U20292 ( .A1(n17229), .A2(n17050), .ZN(n17051) );
  OAI21_X1 U20293 ( .B1(n17052), .B2(P3_EBX_REG_18__SCAN_IN), .A(n17051), .ZN(
        n17053) );
  OAI21_X1 U20294 ( .B1(n17304), .B2(n17221), .A(n17053), .ZN(P3_U2685) );
  AOI22_X1 U20295 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20296 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17154), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n15746), .ZN(n17056) );
  AOI22_X1 U20297 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17183), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20298 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17152), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17175), .ZN(n17054) );
  NAND4_X1 U20299 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17063) );
  AOI22_X1 U20300 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20301 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17173), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17176), .ZN(n17060) );
  AOI22_X1 U20302 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9697), .ZN(n17059) );
  AOI22_X1 U20303 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17174), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17162), .ZN(n17058) );
  NAND4_X1 U20304 ( .A1(n17061), .A2(n17060), .A3(n17059), .A4(n17058), .ZN(
        n17062) );
  NOR2_X1 U20305 ( .A1(n17063), .A2(n17062), .ZN(n17310) );
  NAND3_X1 U20306 ( .A1(n17065), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17221), 
        .ZN(n17064) );
  OAI221_X1 U20307 ( .B1(n17065), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17221), 
        .C2(n17310), .A(n17064), .ZN(P3_U2686) );
  AOI22_X1 U20308 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20309 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20310 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20311 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17066) );
  NAND4_X1 U20312 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n17075) );
  AOI22_X1 U20313 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20314 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20315 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20316 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20317 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  NOR2_X1 U20318 ( .A1(n17075), .A2(n17074), .ZN(n17316) );
  NOR2_X1 U20319 ( .A1(n17229), .A2(n17077), .ZN(n17089) );
  AOI22_X1 U20320 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17089), .B1(n17077), 
        .B2(n17076), .ZN(n17078) );
  OAI21_X1 U20321 ( .B1(n17316), .B2(n17221), .A(n17078), .ZN(P3_U2687) );
  AOI22_X1 U20322 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20323 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20324 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20325 ( .A1(n15746), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17079) );
  NAND4_X1 U20326 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        n17088) );
  AOI22_X1 U20327 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20328 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20329 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20330 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17083) );
  NAND4_X1 U20331 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17087) );
  NOR2_X1 U20332 ( .A1(n17088), .A2(n17087), .ZN(n17320) );
  INV_X1 U20333 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17104) );
  NOR2_X1 U20334 ( .A1(n17104), .A2(n20779), .ZN(n17090) );
  OAI221_X1 U20335 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17105), .C1(
        P3_EBX_REG_15__SCAN_IN), .C2(n17090), .A(n17089), .ZN(n17091) );
  OAI21_X1 U20336 ( .B1(n17320), .B2(n17221), .A(n17091), .ZN(P3_U2688) );
  AOI21_X1 U20337 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17105), .A(n17229), .ZN(
        n17103) );
  AOI22_X1 U20338 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20339 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20340 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17092) );
  OAI21_X1 U20341 ( .B1(n17093), .B2(n20874), .A(n17092), .ZN(n17099) );
  AOI22_X1 U20342 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20343 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20344 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20345 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17094) );
  NAND4_X1 U20346 ( .A1(n17097), .A2(n17096), .A3(n17095), .A4(n17094), .ZN(
        n17098) );
  AOI211_X1 U20347 ( .C1(n9704), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17099), .B(n17098), .ZN(n17100) );
  NAND3_X1 U20348 ( .A1(n17102), .A2(n17101), .A3(n17100), .ZN(n17322) );
  AOI22_X1 U20349 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17103), .B1(n17229), 
        .B2(n17322), .ZN(n17107) );
  NAND4_X1 U20350 ( .A1(n18236), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17105), 
        .A4(n17104), .ZN(n17106) );
  NAND2_X1 U20351 ( .A1(n17107), .A2(n17106), .ZN(P3_U2689) );
  AOI22_X1 U20352 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20353 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20354 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20355 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17109) );
  NAND4_X1 U20356 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17118) );
  AOI22_X1 U20357 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20358 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20359 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20360 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17113) );
  NAND4_X1 U20361 ( .A1(n17116), .A2(n17115), .A3(n17114), .A4(n17113), .ZN(
        n17117) );
  NOR2_X1 U20362 ( .A1(n17118), .A2(n17117), .ZN(n17331) );
  OAI21_X1 U20363 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17135), .A(n17119), .ZN(
        n17120) );
  AOI22_X1 U20364 ( .A1(n17229), .A2(n17331), .B1(n17120), .B2(n17221), .ZN(
        P3_U2691) );
  INV_X1 U20365 ( .A(n17121), .ZN(n17122) );
  OAI21_X1 U20366 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17122), .A(n17221), .ZN(
        n17134) );
  AOI22_X1 U20367 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20368 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20369 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15746), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20370 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17124) );
  NAND4_X1 U20371 ( .A1(n17127), .A2(n17126), .A3(n17125), .A4(n17124), .ZN(
        n17133) );
  AOI22_X1 U20372 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20373 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20374 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17129) );
  AOI22_X1 U20375 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17128) );
  NAND4_X1 U20376 ( .A1(n17131), .A2(n17130), .A3(n17129), .A4(n17128), .ZN(
        n17132) );
  NOR2_X1 U20377 ( .A1(n17133), .A2(n17132), .ZN(n17334) );
  OAI22_X1 U20378 ( .A1(n17135), .A2(n17134), .B1(n17334), .B2(n17221), .ZN(
        P3_U2692) );
  AOI22_X1 U20379 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20380 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20381 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20382 ( .A1(n15746), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17136) );
  NAND4_X1 U20383 ( .A1(n17139), .A2(n17138), .A3(n17137), .A4(n17136), .ZN(
        n17147) );
  AOI22_X1 U20384 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20385 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20386 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20387 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9697), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17142) );
  NAND4_X1 U20388 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17146) );
  NOR2_X1 U20389 ( .A1(n17147), .A2(n17146), .ZN(n17340) );
  NOR2_X1 U20390 ( .A1(n17229), .A2(n17149), .ZN(n17169) );
  NOR2_X1 U20391 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17280), .ZN(n17148) );
  AOI22_X1 U20392 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17169), .B1(n17149), 
        .B2(n17148), .ZN(n17150) );
  OAI21_X1 U20393 ( .B1(n17340), .B2(n17221), .A(n17150), .ZN(P3_U2693) );
  AOI22_X1 U20394 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17152), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20395 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17173), .ZN(n17157) );
  AOI22_X1 U20396 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20397 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17175), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17154), .ZN(n17155) );
  NAND4_X1 U20398 ( .A1(n17158), .A2(n17157), .A3(n17156), .A4(n17155), .ZN(
        n17168) );
  AOI22_X1 U20399 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17159), .ZN(n17166) );
  AOI22_X1 U20400 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n15746), .ZN(n17165) );
  AOI22_X1 U20401 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20402 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9697), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17163) );
  NAND4_X1 U20403 ( .A1(n17166), .A2(n17165), .A3(n17164), .A4(n17163), .ZN(
        n17167) );
  NOR2_X1 U20404 ( .A1(n17168), .A2(n17167), .ZN(n17342) );
  INV_X1 U20405 ( .A(n17194), .ZN(n17170) );
  OAI21_X1 U20406 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17170), .A(n17169), .ZN(
        n17171) );
  OAI21_X1 U20407 ( .B1(n17342), .B2(n17221), .A(n17171), .ZN(P3_U2694) );
  AOI22_X1 U20408 ( .A1(n17172), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12485), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20409 ( .A1(n12462), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20410 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20411 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17177) );
  NAND4_X1 U20412 ( .A1(n17180), .A2(n17179), .A3(n17178), .A4(n17177), .ZN(
        n17191) );
  AOI22_X1 U20413 ( .A1(n12464), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20414 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20415 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20416 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17186) );
  NAND4_X1 U20417 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17190) );
  NOR2_X1 U20418 ( .A1(n17191), .A2(n17190), .ZN(n17345) );
  NOR2_X1 U20419 ( .A1(n17193), .A2(n17192), .ZN(n17195) );
  NOR3_X1 U20420 ( .A1(n17280), .A2(n17203), .A3(n17208), .ZN(n17200) );
  OAI221_X1 U20421 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17195), .C1(
        P3_EBX_REG_8__SCAN_IN), .C2(n17200), .A(n17194), .ZN(n17196) );
  AOI22_X1 U20422 ( .A1(n17229), .A2(n17345), .B1(n17196), .B2(n17221), .ZN(
        P3_U2695) );
  NAND2_X1 U20423 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17200), .ZN(n17199) );
  NAND3_X1 U20424 ( .A1(n17199), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n17221), .ZN(
        n17197) );
  OAI221_X1 U20425 ( .B1(n17199), .B2(P3_EBX_REG_7__SCAN_IN), .C1(n17221), 
        .C2(n17198), .A(n17197), .ZN(P3_U2696) );
  INV_X1 U20426 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17202) );
  OAI211_X1 U20427 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17200), .A(n17199), .B(
        n17221), .ZN(n17201) );
  OAI21_X1 U20428 ( .B1(n17221), .B2(n17202), .A(n17201), .ZN(P3_U2697) );
  AOI21_X1 U20429 ( .B1(n17203), .B2(n17208), .A(n17229), .ZN(n17204) );
  INV_X1 U20430 ( .A(n17204), .ZN(n17206) );
  INV_X1 U20431 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17205) );
  OAI22_X1 U20432 ( .A1(n17207), .A2(n17206), .B1(n17205), .B2(n17221), .ZN(
        P3_U2698) );
  INV_X1 U20433 ( .A(n17208), .ZN(n17213) );
  INV_X1 U20434 ( .A(n17231), .ZN(n17224) );
  NAND2_X1 U20435 ( .A1(n17209), .A2(n17224), .ZN(n17214) );
  NOR2_X1 U20436 ( .A1(n17210), .A2(n17214), .ZN(n17217) );
  AOI21_X1 U20437 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17221), .A(n17217), .ZN(
        n17212) );
  INV_X1 U20438 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17211) );
  OAI22_X1 U20439 ( .A1(n17213), .A2(n17212), .B1(n17211), .B2(n17221), .ZN(
        P3_U2699) );
  INV_X1 U20440 ( .A(n17214), .ZN(n17219) );
  AOI21_X1 U20441 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17221), .A(n17219), .ZN(
        n17216) );
  INV_X1 U20442 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17215) );
  OAI22_X1 U20443 ( .A1(n17217), .A2(n17216), .B1(n17215), .B2(n17221), .ZN(
        P3_U2700) );
  AOI21_X1 U20444 ( .B1(n17227), .B2(n17218), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17222) );
  INV_X1 U20445 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17220) );
  AOI221_X1 U20446 ( .B1(n17222), .B2(n17221), .C1(n17220), .C2(n17229), .A(
        n17219), .ZN(P3_U2701) );
  AOI22_X1 U20447 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17229), .B1(
        n17224), .B2(n17223), .ZN(n17225) );
  OAI21_X1 U20448 ( .B1(n17227), .B2(n17226), .A(n17225), .ZN(P3_U2702) );
  AOI22_X1 U20449 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17229), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17228), .ZN(n17230) );
  OAI21_X1 U20450 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17231), .A(n17230), .ZN(
        P3_U2703) );
  INV_X1 U20451 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17387) );
  INV_X1 U20452 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17391) );
  INV_X1 U20453 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17397) );
  INV_X1 U20454 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17492) );
  INV_X1 U20455 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20941) );
  NOR2_X1 U20456 ( .A1(n20811), .A2(n20941), .ZN(n17374) );
  INV_X1 U20457 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17424) );
  INV_X1 U20458 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17426) );
  INV_X1 U20459 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17428) );
  INV_X1 U20460 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17434) );
  NOR4_X1 U20461 ( .A1(n17424), .A2(n17426), .A3(n17428), .A4(n17434), .ZN(
        n17232) );
  NAND4_X1 U20462 ( .A1(n17374), .A2(P3_EAX_REG_4__SCAN_IN), .A3(
        P3_EAX_REG_3__SCAN_IN), .A4(n17232), .ZN(n17321) );
  NAND4_X1 U20463 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17233)
         );
  INV_X1 U20464 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17399) );
  INV_X1 U20465 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17401) );
  NOR2_X1 U20466 ( .A1(n17399), .A2(n17401), .ZN(n17234) );
  NAND4_X1 U20467 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17234), .ZN(n17279) );
  NAND2_X1 U20468 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17244), .ZN(n17243) );
  NAND2_X1 U20469 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17239), .ZN(n17238) );
  NAND3_X1 U20470 ( .A1(n17366), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17238), 
        .ZN(n17237) );
  NOR2_X2 U20471 ( .A1(n17235), .A2(n17366), .ZN(n17311) );
  NAND2_X1 U20472 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17311), .ZN(n17236) );
  OAI211_X1 U20473 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17238), .A(n17237), .B(
        n17236), .ZN(P3_U2704) );
  NOR2_X2 U20474 ( .A1(n18223), .A2(n17366), .ZN(n17312) );
  AOI22_X1 U20475 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17311), .ZN(n17241) );
  OAI211_X1 U20476 ( .C1(n17239), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17366), .B(
        n17238), .ZN(n17240) );
  OAI211_X1 U20477 ( .C1(n17242), .C2(n17368), .A(n17241), .B(n17240), .ZN(
        P3_U2705) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17311), .ZN(n17246) );
  OAI211_X1 U20479 ( .C1(n17244), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17366), .B(
        n17243), .ZN(n17245) );
  OAI211_X1 U20480 ( .C1(n17247), .C2(n17368), .A(n17246), .B(n17245), .ZN(
        P3_U2706) );
  INV_X1 U20481 ( .A(n17312), .ZN(n17285) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17311), .B1(n17372), .B2(
        n17248), .ZN(n17251) );
  OAI211_X1 U20483 ( .C1(n9796), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17366), .B(
        n17249), .ZN(n17250) );
  OAI211_X1 U20484 ( .C1(n17285), .C2(n17479), .A(n17251), .B(n17250), .ZN(
        P3_U2707) );
  OAI21_X1 U20485 ( .B1(n17254), .B2(n17253), .A(n17252), .ZN(n17258) );
  AOI22_X1 U20486 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17311), .ZN(n17257) );
  AOI211_X1 U20487 ( .C1(n17387), .C2(n17259), .A(n9796), .B(n17295), .ZN(
        n17255) );
  INV_X1 U20488 ( .A(n17255), .ZN(n17256) );
  OAI211_X1 U20489 ( .C1(n17258), .C2(n17368), .A(n17257), .B(n17256), .ZN(
        P3_U2708) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17311), .ZN(n17261) );
  OAI211_X1 U20491 ( .C1(n17263), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17366), .B(
        n17259), .ZN(n17260) );
  OAI211_X1 U20492 ( .C1(n17262), .C2(n17368), .A(n17261), .B(n17260), .ZN(
        P3_U2709) );
  AOI22_X1 U20493 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17311), .ZN(n17266) );
  AOI211_X1 U20494 ( .C1(n17391), .C2(n17268), .A(n17263), .B(n17295), .ZN(
        n17264) );
  INV_X1 U20495 ( .A(n17264), .ZN(n17265) );
  OAI211_X1 U20496 ( .C1(n17267), .C2(n17368), .A(n17266), .B(n17265), .ZN(
        P3_U2710) );
  AOI22_X1 U20497 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17311), .ZN(n17271) );
  OAI211_X1 U20498 ( .C1(n17269), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17366), .B(
        n17268), .ZN(n17270) );
  OAI211_X1 U20499 ( .C1(n17272), .C2(n17368), .A(n17271), .B(n17270), .ZN(
        P3_U2711) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17311), .ZN(n17276) );
  OAI211_X1 U20501 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17274), .A(n17366), .B(
        n17273), .ZN(n17275) );
  OAI211_X1 U20502 ( .C1(n17277), .C2(n17368), .A(n17276), .B(n17275), .ZN(
        P3_U2712) );
  AOI22_X1 U20503 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17311), .B1(n17372), .B2(
        n17278), .ZN(n17284) );
  INV_X1 U20504 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17449) );
  INV_X1 U20505 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17446) );
  NAND2_X1 U20506 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17305), .ZN(n17301) );
  NAND2_X1 U20507 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17296), .ZN(n17291) );
  NAND2_X1 U20508 ( .A1(n17366), .A2(n17291), .ZN(n17290) );
  OAI21_X1 U20509 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17348), .A(n17290), .ZN(
        n17282) );
  NOR3_X1 U20510 ( .A1(n17280), .A2(n17313), .A3(n17279), .ZN(n17281) );
  AOI22_X1 U20511 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17282), .B1(n17281), 
        .B2(n17397), .ZN(n17283) );
  OAI211_X1 U20512 ( .C1(n18229), .C2(n17285), .A(n17284), .B(n17283), .ZN(
        P3_U2713) );
  INV_X1 U20513 ( .A(n17311), .ZN(n17286) );
  OAI22_X1 U20514 ( .A1(n17287), .A2(n17368), .B1(n15107), .B2(n17286), .ZN(
        n17288) );
  AOI21_X1 U20515 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17312), .A(n17288), .ZN(
        n17289) );
  OAI221_X1 U20516 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17291), .C1(n17399), 
        .C2(n17290), .A(n17289), .ZN(P3_U2714) );
  AOI22_X1 U20517 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17311), .ZN(n17293) );
  OAI211_X1 U20518 ( .C1(n17296), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17366), .B(
        n17291), .ZN(n17292) );
  OAI211_X1 U20519 ( .C1(n17294), .C2(n17368), .A(n17293), .B(n17292), .ZN(
        P3_U2715) );
  AOI22_X1 U20520 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17311), .ZN(n17299) );
  AOI211_X1 U20521 ( .C1(n17449), .C2(n17301), .A(n17296), .B(n17295), .ZN(
        n17297) );
  INV_X1 U20522 ( .A(n17297), .ZN(n17298) );
  OAI211_X1 U20523 ( .C1(n17300), .C2(n17368), .A(n17299), .B(n17298), .ZN(
        P3_U2716) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17311), .ZN(n17303) );
  OAI211_X1 U20525 ( .C1(n17305), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17366), .B(
        n17301), .ZN(n17302) );
  OAI211_X1 U20526 ( .C1(n17304), .C2(n17368), .A(n17303), .B(n17302), .ZN(
        P3_U2717) );
  AOI22_X1 U20527 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17311), .ZN(n17309) );
  INV_X1 U20528 ( .A(n17313), .ZN(n17307) );
  INV_X1 U20529 ( .A(n17305), .ZN(n17306) );
  OAI211_X1 U20530 ( .C1(n17307), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17366), .B(
        n17306), .ZN(n17308) );
  OAI211_X1 U20531 ( .C1(n17310), .C2(n17368), .A(n17309), .B(n17308), .ZN(
        P3_U2718) );
  AOI22_X1 U20532 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17312), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17311), .ZN(n17315) );
  OAI211_X1 U20533 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17317), .A(n17366), .B(
        n17313), .ZN(n17314) );
  OAI211_X1 U20534 ( .C1(n17316), .C2(n17368), .A(n17315), .B(n17314), .ZN(
        P3_U2719) );
  AOI21_X1 U20535 ( .B1(n17492), .B2(n17323), .A(n17317), .ZN(n17318) );
  AOI22_X1 U20536 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17373), .B1(n17318), .B2(
        n17366), .ZN(n17319) );
  OAI21_X1 U20537 ( .B1(n17320), .B2(n17368), .A(n17319), .ZN(P3_U2720) );
  INV_X1 U20538 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17415) );
  INV_X1 U20539 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17420) );
  NOR2_X1 U20540 ( .A1(n17321), .A2(n17348), .ZN(n17351) );
  NAND2_X1 U20541 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17351), .ZN(n17341) );
  NAND3_X1 U20542 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(n17344), .ZN(n17330) );
  NOR2_X1 U20543 ( .A1(n17415), .A2(n17330), .ZN(n17333) );
  NAND2_X1 U20544 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17333), .ZN(n17326) );
  AOI22_X1 U20545 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17373), .B1(n17372), .B2(
        n17322), .ZN(n17325) );
  NAND3_X1 U20546 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17366), .A3(n17323), 
        .ZN(n17324) );
  OAI211_X1 U20547 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17326), .A(n17325), .B(
        n17324), .ZN(P3_U2721) );
  INV_X1 U20548 ( .A(n17326), .ZN(n17329) );
  AOI21_X1 U20549 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17366), .A(n17333), .ZN(
        n17328) );
  OAI222_X1 U20550 ( .A1(n17371), .A2(n17482), .B1(n17329), .B2(n17328), .C1(
        n17368), .C2(n17327), .ZN(P3_U2722) );
  INV_X1 U20551 ( .A(n17330), .ZN(n17336) );
  AOI21_X1 U20552 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17366), .A(n17336), .ZN(
        n17332) );
  OAI222_X1 U20553 ( .A1(n17371), .A2(n17479), .B1(n17333), .B2(n17332), .C1(
        n17368), .C2(n17331), .ZN(P3_U2723) );
  AOI22_X1 U20554 ( .A1(n17344), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17366), .ZN(n17335) );
  OAI222_X1 U20555 ( .A1(n17371), .A2(n17477), .B1(n17336), .B2(n17335), .C1(
        n17368), .C2(n17334), .ZN(P3_U2724) );
  NAND2_X1 U20556 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17344), .ZN(n17337) );
  OAI211_X1 U20557 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17344), .A(n17366), .B(
        n17337), .ZN(n17339) );
  NAND2_X1 U20558 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17373), .ZN(n17338) );
  OAI211_X1 U20559 ( .C1(n17340), .C2(n17368), .A(n17339), .B(n17338), .ZN(
        P3_U2725) );
  INV_X1 U20560 ( .A(n17341), .ZN(n17347) );
  AOI21_X1 U20561 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17366), .A(n17347), .ZN(
        n17343) );
  OAI222_X1 U20562 ( .A1(n17371), .A2(n17473), .B1(n17344), .B2(n17343), .C1(
        n17368), .C2(n17342), .ZN(P3_U2726) );
  AOI21_X1 U20563 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17366), .A(n17351), .ZN(
        n17346) );
  OAI222_X1 U20564 ( .A1(n17371), .A2(n17471), .B1(n17347), .B2(n17346), .C1(
        n17368), .C2(n17345), .ZN(P3_U2727) );
  NAND2_X1 U20565 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n17349) );
  INV_X1 U20566 ( .A(n17348), .ZN(n17376) );
  NAND3_X1 U20567 ( .A1(n17374), .A2(P3_EAX_REG_2__SCAN_IN), .A3(n17376), .ZN(
        n17365) );
  NOR2_X1 U20568 ( .A1(n17349), .A2(n17365), .ZN(n17361) );
  NAND2_X1 U20569 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17361), .ZN(n17352) );
  NOR2_X1 U20570 ( .A1(n17426), .A2(n17352), .ZN(n17354) );
  AOI21_X1 U20571 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17366), .A(n17354), .ZN(
        n17350) );
  OAI222_X1 U20572 ( .A1(n17371), .A2(n18233), .B1(n17351), .B2(n17350), .C1(
        n17368), .C2(n10049), .ZN(P3_U2728) );
  INV_X1 U20573 ( .A(n17352), .ZN(n17358) );
  AOI21_X1 U20574 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17366), .A(n17358), .ZN(
        n17355) );
  OAI222_X1 U20575 ( .A1(n17371), .A2(n18229), .B1(n17355), .B2(n17354), .C1(
        n17368), .C2(n17353), .ZN(P3_U2729) );
  AOI21_X1 U20576 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17366), .A(n17361), .ZN(
        n17357) );
  OAI222_X1 U20577 ( .A1(n18224), .A2(n17371), .B1(n17358), .B2(n17357), .C1(
        n17368), .C2(n17356), .ZN(P3_U2730) );
  INV_X1 U20578 ( .A(n17365), .ZN(n17370) );
  AOI22_X1 U20579 ( .A1(n17370), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17366), .ZN(n17360) );
  OAI222_X1 U20580 ( .A1(n18220), .A2(n17371), .B1(n17361), .B2(n17360), .C1(
        n17368), .C2(n17359), .ZN(P3_U2731) );
  NAND3_X1 U20581 ( .A1(n17366), .A2(P3_EAX_REG_3__SCAN_IN), .A3(n17365), .ZN(
        n17364) );
  AOI22_X1 U20582 ( .A1(n17373), .A2(BUF2_REG_3__SCAN_IN), .B1(n17372), .B2(
        n17362), .ZN(n17363) );
  OAI211_X1 U20583 ( .C1(P3_EAX_REG_3__SCAN_IN), .C2(n17365), .A(n17364), .B(
        n17363), .ZN(P3_U2732) );
  AOI22_X1 U20584 ( .A1(n17376), .A2(n17374), .B1(P3_EAX_REG_2__SCAN_IN), .B2(
        n17366), .ZN(n17369) );
  OAI222_X1 U20585 ( .A1(n18210), .A2(n17371), .B1(n17370), .B2(n17369), .C1(
        n17368), .C2(n17367), .ZN(P3_U2733) );
  AOI22_X1 U20586 ( .A1(n17373), .A2(BUF2_REG_1__SCAN_IN), .B1(n17372), .B2(
        n12511), .ZN(n17378) );
  INV_X1 U20587 ( .A(n17374), .ZN(n17375) );
  OAI211_X1 U20588 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(P3_EAX_REG_1__SCAN_IN), 
        .A(n17376), .B(n17375), .ZN(n17377) );
  OAI211_X1 U20589 ( .C1(n17379), .C2(n20941), .A(n17378), .B(n17377), .ZN(
        P3_U2734) );
  OR2_X1 U20590 ( .A1(n18800), .A2(n17870), .ZN(n17438) );
  INV_X1 U20591 ( .A(n17443), .ZN(n17381) );
  NOR2_X1 U20592 ( .A1(n17439), .A2(n17382), .ZN(P3_U2736) );
  INV_X1 U20593 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n20925) );
  NOR2_X1 U20594 ( .A1(n18203), .A2(n17440), .ZN(n17407) );
  INV_X1 U20595 ( .A(n17438), .ZN(n18845) );
  AOI22_X1 U20596 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17407), .B1(n18845), 
        .B2(P3_UWORD_REG_14__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20597 ( .B1(n20925), .B2(n17439), .A(n17383), .ZN(P3_U2737) );
  INV_X1 U20598 ( .A(P3_UWORD_REG_13__SCAN_IN), .ZN(n20743) );
  INV_X2 U20599 ( .A(n17439), .ZN(n17435) );
  AOI22_X1 U20600 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17407), .B1(n17435), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20601 ( .B1(n20743), .B2(n17438), .A(n17384), .ZN(P3_U2738) );
  INV_X1 U20602 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20855) );
  AOI22_X1 U20603 ( .A1(n18845), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20604 ( .B1(n20855), .B2(n17406), .A(n17385), .ZN(P3_U2739) );
  AOI22_X1 U20605 ( .A1(n17436), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17386) );
  OAI21_X1 U20606 ( .B1(n17387), .B2(n17406), .A(n17386), .ZN(P3_U2740) );
  INV_X1 U20607 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20608 ( .A1(n17436), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20609 ( .B1(n17389), .B2(n17406), .A(n17388), .ZN(P3_U2741) );
  AOI22_X1 U20610 ( .A1(n17436), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20611 ( .B1(n17391), .B2(n17406), .A(n17390), .ZN(P3_U2742) );
  INV_X1 U20612 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U20613 ( .A1(n17436), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20614 ( .B1(n17393), .B2(n17406), .A(n17392), .ZN(P3_U2743) );
  INV_X1 U20615 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20616 ( .A1(n17436), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17394) );
  OAI21_X1 U20617 ( .B1(n17395), .B2(n17406), .A(n17394), .ZN(P3_U2744) );
  AOI22_X1 U20618 ( .A1(n17436), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20619 ( .B1(n17397), .B2(n17406), .A(n17396), .ZN(P3_U2745) );
  AOI22_X1 U20620 ( .A1(n17436), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20621 ( .B1(n17399), .B2(n17406), .A(n17398), .ZN(P3_U2746) );
  AOI22_X1 U20622 ( .A1(n17436), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20623 ( .B1(n17401), .B2(n17406), .A(n17400), .ZN(P3_U2747) );
  AOI22_X1 U20624 ( .A1(n17436), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20625 ( .B1(n17449), .B2(n17406), .A(n17402), .ZN(P3_U2748) );
  INV_X1 U20626 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20627 ( .A1(n17436), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20628 ( .B1(n17404), .B2(n17406), .A(n17403), .ZN(P3_U2749) );
  AOI22_X1 U20629 ( .A1(n17436), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20630 ( .B1(n17446), .B2(n17406), .A(n17405), .ZN(P3_U2750) );
  INV_X1 U20631 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n20765) );
  AOI22_X1 U20632 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17407), .B1(n18845), 
        .B2(P3_UWORD_REG_0__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20633 ( .B1(n20765), .B2(n17439), .A(n17408), .ZN(P3_U2751) );
  AOI22_X1 U20634 ( .A1(n17436), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20635 ( .B1(n17492), .B2(n17440), .A(n17409), .ZN(P3_U2752) );
  INV_X1 U20636 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20637 ( .A1(n17436), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20638 ( .B1(n17411), .B2(n17440), .A(n17410), .ZN(P3_U2753) );
  INV_X1 U20639 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20640 ( .A1(n17436), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20641 ( .B1(n17413), .B2(n17440), .A(n17412), .ZN(P3_U2754) );
  AOI22_X1 U20642 ( .A1(n17436), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20643 ( .B1(n17415), .B2(n17440), .A(n17414), .ZN(P3_U2755) );
  INV_X1 U20644 ( .A(P3_LWORD_REG_11__SCAN_IN), .ZN(n20843) );
  INV_X1 U20645 ( .A(n17440), .ZN(n17431) );
  AOI22_X1 U20646 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17431), .B1(n17435), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17416) );
  OAI21_X1 U20647 ( .B1(n20843), .B2(n17438), .A(n17416), .ZN(P3_U2756) );
  INV_X1 U20648 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20649 ( .A1(n17436), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17417) );
  OAI21_X1 U20650 ( .B1(n17418), .B2(n17440), .A(n17417), .ZN(P3_U2757) );
  AOI22_X1 U20651 ( .A1(n17436), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17419) );
  OAI21_X1 U20652 ( .B1(n17420), .B2(n17440), .A(n17419), .ZN(P3_U2758) );
  INV_X1 U20653 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20654 ( .A1(n17436), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20655 ( .B1(n17422), .B2(n17440), .A(n17421), .ZN(P3_U2759) );
  AOI22_X1 U20656 ( .A1(n17436), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17423) );
  OAI21_X1 U20657 ( .B1(n17424), .B2(n17440), .A(n17423), .ZN(P3_U2760) );
  AOI22_X1 U20658 ( .A1(n17436), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20659 ( .B1(n17426), .B2(n17440), .A(n17425), .ZN(P3_U2761) );
  AOI22_X1 U20660 ( .A1(n17436), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17427) );
  OAI21_X1 U20661 ( .B1(n17428), .B2(n17440), .A(n17427), .ZN(P3_U2762) );
  INV_X1 U20662 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20663 ( .A1(n17436), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20664 ( .B1(n17430), .B2(n17440), .A(n17429), .ZN(P3_U2763) );
  INV_X1 U20665 ( .A(P3_LWORD_REG_3__SCAN_IN), .ZN(n20953) );
  AOI22_X1 U20666 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17431), .B1(n17435), .B2(
        P3_DATAO_REG_3__SCAN_IN), .ZN(n17432) );
  OAI21_X1 U20667 ( .B1(n20953), .B2(n17438), .A(n17432), .ZN(P3_U2764) );
  AOI22_X1 U20668 ( .A1(n18845), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20669 ( .B1(n17434), .B2(n17440), .A(n17433), .ZN(P3_U2765) );
  AOI22_X1 U20670 ( .A1(n17436), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17435), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20671 ( .B1(n20941), .B2(n17440), .A(n17437), .ZN(P3_U2766) );
  INV_X1 U20672 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n20939) );
  INV_X1 U20673 ( .A(P3_LWORD_REG_0__SCAN_IN), .ZN(n20806) );
  OAI222_X1 U20674 ( .A1(n17440), .A2(n20811), .B1(n17439), .B2(n20939), .C1(
        n17438), .C2(n20806), .ZN(P3_U2767) );
  AOI211_X1 U20675 ( .C1(n18837), .C2(n18835), .A(n17441), .B(n17443), .ZN(
        n17465) );
  NAND2_X1 U20676 ( .A1(n17465), .A2(n18835), .ZN(n17486) );
  INV_X1 U20677 ( .A(n17442), .ZN(n18687) );
  INV_X2 U20678 ( .A(n17491), .ZN(n17484) );
  INV_X1 U20679 ( .A(n17465), .ZN(n17488) );
  AOI22_X1 U20680 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17483), .ZN(n17444) );
  OAI21_X1 U20681 ( .B1(n18200), .B2(n17486), .A(n17444), .ZN(P3_U2768) );
  INV_X1 U20682 ( .A(n17486), .ZN(n17489) );
  AOI22_X1 U20683 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17489), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17488), .ZN(n17445) );
  OAI21_X1 U20684 ( .B1(n17446), .B2(n17491), .A(n17445), .ZN(P3_U2769) );
  AOI22_X1 U20685 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17483), .ZN(n17447) );
  OAI21_X1 U20686 ( .B1(n18210), .B2(n17486), .A(n17447), .ZN(P3_U2770) );
  AOI22_X1 U20687 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17489), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17488), .ZN(n17448) );
  OAI21_X1 U20688 ( .B1(n17449), .B2(n17491), .A(n17448), .ZN(P3_U2771) );
  AOI22_X1 U20689 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17483), .ZN(n17450) );
  OAI21_X1 U20690 ( .B1(n18220), .B2(n17486), .A(n17450), .ZN(P3_U2772) );
  AOI22_X1 U20691 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17483), .ZN(n17451) );
  OAI21_X1 U20692 ( .B1(n18224), .B2(n17486), .A(n17451), .ZN(P3_U2773) );
  AOI22_X1 U20693 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17483), .ZN(n17452) );
  OAI21_X1 U20694 ( .B1(n18229), .B2(n17486), .A(n17452), .ZN(P3_U2774) );
  AOI22_X1 U20695 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17488), .ZN(n17453) );
  OAI21_X1 U20696 ( .B1(n18233), .B2(n17486), .A(n17453), .ZN(P3_U2775) );
  AOI22_X1 U20697 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17488), .ZN(n17454) );
  OAI21_X1 U20698 ( .B1(n17471), .B2(n17486), .A(n17454), .ZN(P3_U2776) );
  AOI22_X1 U20699 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17488), .ZN(n17455) );
  OAI21_X1 U20700 ( .B1(n17473), .B2(n17486), .A(n17455), .ZN(P3_U2777) );
  AOI22_X1 U20701 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17488), .ZN(n17456) );
  OAI21_X1 U20702 ( .B1(n17475), .B2(n17486), .A(n17456), .ZN(P3_U2778) );
  AOI22_X1 U20703 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17488), .ZN(n17457) );
  OAI21_X1 U20704 ( .B1(n17477), .B2(n17486), .A(n17457), .ZN(P3_U2779) );
  AOI22_X1 U20705 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17488), .ZN(n17458) );
  OAI21_X1 U20706 ( .B1(n17479), .B2(n17486), .A(n17458), .ZN(P3_U2780) );
  AOI22_X1 U20707 ( .A1(P3_UWORD_REG_13__SCAN_IN), .A2(n17483), .B1(
        P3_EAX_REG_29__SCAN_IN), .B2(n17484), .ZN(n17459) );
  OAI21_X1 U20708 ( .B1(n17482), .B2(n17481), .A(n17459), .ZN(P3_U2781) );
  AOI22_X1 U20709 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17484), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17483), .ZN(n17460) );
  OAI21_X1 U20710 ( .B1(n17487), .B2(n17481), .A(n17460), .ZN(P3_U2782) );
  AOI22_X1 U20711 ( .A1(P3_LWORD_REG_0__SCAN_IN), .A2(n17483), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n17484), .ZN(n17461) );
  OAI21_X1 U20712 ( .B1(n18200), .B2(n17481), .A(n17461), .ZN(P3_U2783) );
  AOI22_X1 U20713 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17489), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17488), .ZN(n17462) );
  OAI21_X1 U20714 ( .B1(n20941), .B2(n17491), .A(n17462), .ZN(P3_U2784) );
  AOI22_X1 U20715 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17488), .ZN(n17463) );
  OAI21_X1 U20716 ( .B1(n18210), .B2(n17481), .A(n17463), .ZN(P3_U2785) );
  AOI22_X1 U20717 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17489), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n17484), .ZN(n17464) );
  OAI21_X1 U20718 ( .B1(n17465), .B2(n20953), .A(n17464), .ZN(P3_U2786) );
  AOI22_X1 U20719 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17483), .ZN(n17466) );
  OAI21_X1 U20720 ( .B1(n18220), .B2(n17481), .A(n17466), .ZN(P3_U2787) );
  AOI22_X1 U20721 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17483), .ZN(n17467) );
  OAI21_X1 U20722 ( .B1(n18224), .B2(n17481), .A(n17467), .ZN(P3_U2788) );
  AOI22_X1 U20723 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17488), .ZN(n17468) );
  OAI21_X1 U20724 ( .B1(n18229), .B2(n17481), .A(n17468), .ZN(P3_U2789) );
  AOI22_X1 U20725 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17483), .ZN(n17469) );
  OAI21_X1 U20726 ( .B1(n18233), .B2(n17481), .A(n17469), .ZN(P3_U2790) );
  AOI22_X1 U20727 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17483), .ZN(n17470) );
  OAI21_X1 U20728 ( .B1(n17471), .B2(n17481), .A(n17470), .ZN(P3_U2791) );
  AOI22_X1 U20729 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17483), .ZN(n17472) );
  OAI21_X1 U20730 ( .B1(n17473), .B2(n17481), .A(n17472), .ZN(P3_U2792) );
  AOI22_X1 U20731 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17483), .ZN(n17474) );
  OAI21_X1 U20732 ( .B1(n17475), .B2(n17481), .A(n17474), .ZN(P3_U2793) );
  AOI22_X1 U20733 ( .A1(P3_LWORD_REG_11__SCAN_IN), .A2(n17483), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17484), .ZN(n17476) );
  OAI21_X1 U20734 ( .B1(n17477), .B2(n17481), .A(n17476), .ZN(P3_U2794) );
  AOI22_X1 U20735 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17483), .ZN(n17478) );
  OAI21_X1 U20736 ( .B1(n17479), .B2(n17481), .A(n17478), .ZN(P3_U2795) );
  AOI22_X1 U20737 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17483), .ZN(n17480) );
  OAI21_X1 U20738 ( .B1(n17482), .B2(n17481), .A(n17480), .ZN(P3_U2796) );
  AOI22_X1 U20739 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17484), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17483), .ZN(n17485) );
  OAI21_X1 U20740 ( .B1(n17487), .B2(n17486), .A(n17485), .ZN(P3_U2797) );
  AOI22_X1 U20741 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17489), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17488), .ZN(n17490) );
  OAI21_X1 U20742 ( .B1(n17492), .B2(n17491), .A(n17490), .ZN(P3_U2798) );
  OAI21_X1 U20743 ( .B1(n17493), .B2(n17773), .A(n17871), .ZN(n17494) );
  AOI21_X1 U20744 ( .B1(n17705), .B2(n17495), .A(n17494), .ZN(n17530) );
  OAI21_X1 U20745 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17610), .A(
        n17530), .ZN(n17516) );
  AOI22_X1 U20746 ( .A1(n17687), .A2(n17496), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17516), .ZN(n17510) );
  AOI21_X1 U20747 ( .B1(n17499), .B2(n17498), .A(n17497), .ZN(n17504) );
  NOR3_X1 U20748 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17887), .A3(
        n17519), .ZN(n17503) );
  NOR2_X1 U20749 ( .A1(n17839), .A2(n17781), .ZN(n17578) );
  INV_X1 U20750 ( .A(n17781), .ZN(n17714) );
  OAI22_X1 U20751 ( .A1(n17877), .A2(n17875), .B1(n17883), .B2(n17714), .ZN(
        n17532) );
  NOR2_X1 U20752 ( .A1(n17887), .A2(n17532), .ZN(n17501) );
  NOR3_X1 U20753 ( .A1(n17578), .A2(n17501), .A3(n17500), .ZN(n17502) );
  AOI211_X1 U20754 ( .C1(n17765), .C2(n17504), .A(n17503), .B(n17502), .ZN(
        n17509) );
  NAND2_X1 U20755 ( .A1(n18186), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17508) );
  NOR2_X1 U20756 ( .A1(n17630), .A2(n17505), .ZN(n17518) );
  OAI211_X1 U20757 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17518), .B(n17506), .ZN(n17507) );
  NAND4_X1 U20758 ( .A1(n17510), .A2(n17509), .A3(n17508), .A4(n17507), .ZN(
        P3_U2802) );
  NAND2_X1 U20759 ( .A1(n17512), .A2(n17511), .ZN(n17513) );
  XNOR2_X1 U20760 ( .A(n17603), .B(n17513), .ZN(n17891) );
  OAI22_X1 U20761 ( .A1(n18184), .A2(n18767), .B1(n17722), .B2(n17514), .ZN(
        n17515) );
  AOI221_X1 U20762 ( .B1(n17518), .B2(n17517), .C1(n17516), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17515), .ZN(n17522) );
  INV_X1 U20763 ( .A(n17519), .ZN(n17520) );
  AOI22_X1 U20764 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17532), .B1(
        n17520), .B2(n17887), .ZN(n17521) );
  OAI211_X1 U20765 ( .C1(n17891), .C2(n17784), .A(n17522), .B(n17521), .ZN(
        P3_U2803) );
  AOI21_X1 U20766 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17524), .A(
        n17523), .ZN(n17900) );
  INV_X1 U20767 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17894) );
  AOI21_X1 U20768 ( .B1(n17525), .B2(n18575), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17529) );
  INV_X1 U20769 ( .A(n17610), .ZN(n17527) );
  OAI21_X1 U20770 ( .B1(n17687), .B2(n17527), .A(n17526), .ZN(n17528) );
  NAND2_X1 U20771 ( .A1(n18186), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17898) );
  OAI211_X1 U20772 ( .C1(n17530), .C2(n17529), .A(n17528), .B(n17898), .ZN(
        n17531) );
  AOI221_X1 U20773 ( .B1(n17533), .B2(n17894), .C1(n17532), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17531), .ZN(n17534) );
  OAI21_X1 U20774 ( .B1(n17900), .B2(n17784), .A(n17534), .ZN(P3_U2804) );
  OAI21_X1 U20775 ( .B1(n17535), .B2(n17870), .A(n17871), .ZN(n17536) );
  AOI21_X1 U20776 ( .B1(n18575), .B2(n17545), .A(n17536), .ZN(n17571) );
  OAI21_X1 U20777 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17610), .A(
        n17571), .ZN(n17551) );
  AOI22_X1 U20778 ( .A1(n17687), .A2(n17537), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17551), .ZN(n17549) );
  XNOR2_X1 U20779 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17538), .ZN(
        n17911) );
  NOR2_X1 U20780 ( .A1(n17566), .A2(n12724), .ZN(n17575) );
  NAND2_X1 U20781 ( .A1(n20775), .A2(n17879), .ZN(n17905) );
  INV_X1 U20782 ( .A(n17905), .ZN(n17539) );
  AOI22_X1 U20783 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17540), .B1(
        n17575), .B2(n17539), .ZN(n17914) );
  OAI21_X1 U20784 ( .B1(n17770), .B2(n17542), .A(n17541), .ZN(n17543) );
  XNOR2_X1 U20785 ( .A(n17543), .B(n20775), .ZN(n17909) );
  OAI22_X1 U20786 ( .A1(n17914), .A2(n17714), .B1(n17784), .B2(n17909), .ZN(
        n17544) );
  AOI21_X1 U20787 ( .B1(n17839), .B2(n17911), .A(n17544), .ZN(n17548) );
  NAND2_X1 U20788 ( .A1(n18186), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17907) );
  NOR2_X1 U20789 ( .A1(n17630), .A2(n17545), .ZN(n17552) );
  OAI211_X1 U20790 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17552), .B(n17546), .ZN(n17547) );
  NAND4_X1 U20791 ( .A1(n17549), .A2(n17548), .A3(n17907), .A4(n17547), .ZN(
        P3_U2805) );
  NOR2_X1 U20792 ( .A1(n18184), .A2(n18762), .ZN(n17550) );
  AOI221_X1 U20793 ( .B1(n17552), .B2(n20938), .C1(n17551), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17550), .ZN(n17560) );
  OAI21_X1 U20794 ( .B1(n17554), .B2(n17556), .A(n17553), .ZN(n17916) );
  NOR2_X1 U20795 ( .A1(n17920), .A2(n17875), .ZN(n17574) );
  AOI21_X1 U20796 ( .B1(n17781), .B2(n17917), .A(n17574), .ZN(n17557) );
  INV_X1 U20797 ( .A(n17657), .ZN(n17673) );
  NAND2_X1 U20798 ( .A1(n17555), .A2(n17556), .ZN(n17928) );
  OAI22_X1 U20799 ( .A1(n17557), .A2(n17556), .B1(n17673), .B2(n17928), .ZN(
        n17558) );
  AOI21_X1 U20800 ( .B1(n17765), .B2(n17916), .A(n17558), .ZN(n17559) );
  OAI211_X1 U20801 ( .C1(n17722), .C2(n17561), .A(n17560), .B(n17559), .ZN(
        P3_U2806) );
  OAI22_X1 U20802 ( .A1(n17603), .A2(n17942), .B1(n17583), .B2(n17562), .ZN(
        n17564) );
  NOR2_X1 U20803 ( .A1(n17564), .A2(n17563), .ZN(n17565) );
  XNOR2_X1 U20804 ( .A(n17565), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17933) );
  OAI21_X1 U20805 ( .B1(n17566), .B2(n17940), .A(n17922), .ZN(n17573) );
  AOI21_X1 U20806 ( .B1(n17567), .B2(n18575), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17570) );
  OAI21_X1 U20807 ( .B1(n17687), .B2(n17527), .A(n17568), .ZN(n17569) );
  NAND2_X1 U20808 ( .A1(n18186), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17932) );
  OAI211_X1 U20809 ( .C1(n17571), .C2(n17570), .A(n17569), .B(n17932), .ZN(
        n17572) );
  AOI21_X1 U20810 ( .B1(n17574), .B2(n17573), .A(n17572), .ZN(n17577) );
  OAI211_X1 U20811 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17575), .A(
        n17781), .B(n17917), .ZN(n17576) );
  OAI211_X1 U20812 ( .C1(n17933), .C2(n17784), .A(n17577), .B(n17576), .ZN(
        P3_U2807) );
  INV_X1 U20813 ( .A(n17578), .ZN(n17617) );
  INV_X1 U20814 ( .A(n17940), .ZN(n18009) );
  OAI22_X1 U20815 ( .A1(n18009), .A2(n17875), .B1(n17579), .B2(n17714), .ZN(
        n17644) );
  AOI21_X1 U20816 ( .B1(n17617), .B2(n17580), .A(n17644), .ZN(n17609) );
  INV_X1 U20817 ( .A(n17563), .ZN(n17581) );
  OAI221_X1 U20818 ( .B1(n17583), .B2(n17582), .C1(n17583), .C2(n17602), .A(
        n17581), .ZN(n17584) );
  XNOR2_X1 U20819 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17584), .ZN(
        n17946) );
  NOR3_X1 U20820 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17630), .A3(
        n17585), .ZN(n17594) );
  INV_X1 U20821 ( .A(n17586), .ZN(n17592) );
  NAND2_X1 U20822 ( .A1(n18186), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17947) );
  AND3_X1 U20823 ( .A1(n17597), .A2(n17707), .A3(n17589), .ZN(n17600) );
  NAND2_X1 U20824 ( .A1(n17705), .A2(n17587), .ZN(n17588) );
  OAI211_X1 U20825 ( .C1(n17589), .C2(n17773), .A(n17871), .B(n17588), .ZN(
        n17614) );
  AOI21_X1 U20826 ( .B1(n17527), .B2(n17611), .A(n17614), .ZN(n17598) );
  INV_X1 U20827 ( .A(n17598), .ZN(n17590) );
  OAI21_X1 U20828 ( .B1(n17600), .B2(n17590), .A(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17591) );
  OAI211_X1 U20829 ( .C1(n17592), .C2(n17722), .A(n17947), .B(n17591), .ZN(
        n17593) );
  AOI211_X1 U20830 ( .C1(n17946), .C2(n17765), .A(n17594), .B(n17593), .ZN(
        n17595) );
  OAI221_X1 U20831 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17596), 
        .C1(n17942), .C2(n17609), .A(n17595), .ZN(P3_U2808) );
  OAI22_X1 U20832 ( .A1(n17598), .A2(n17597), .B1(n18184), .B2(n18756), .ZN(
        n17599) );
  AOI211_X1 U20833 ( .C1(n17601), .C2(n17687), .A(n17600), .B(n17599), .ZN(
        n17608) );
  NAND3_X1 U20834 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17603), .A3(
        n17602), .ZN(n17624) );
  INV_X1 U20835 ( .A(n17604), .ZN(n17637) );
  OAI22_X1 U20836 ( .A1(n17939), .A2(n17624), .B1(n17605), .B2(n17637), .ZN(
        n17606) );
  XNOR2_X1 U20837 ( .A(n17945), .B(n17606), .ZN(n17958) );
  NAND2_X1 U20838 ( .A1(n17980), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17623) );
  NOR3_X1 U20839 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17939), .A3(
        n17623), .ZN(n17957) );
  AOI22_X1 U20840 ( .A1(n17765), .A2(n17958), .B1(n17657), .B2(n17957), .ZN(
        n17607) );
  OAI211_X1 U20841 ( .C1(n17609), .C2(n17945), .A(n17608), .B(n17607), .ZN(
        P3_U2809) );
  NAND2_X1 U20842 ( .A1(n17722), .A2(n17610), .ZN(n17844) );
  OAI21_X1 U20843 ( .B1(n17612), .B2(n18488), .A(n17611), .ZN(n17613) );
  AOI22_X1 U20844 ( .A1(n17615), .A2(n17844), .B1(n17614), .B2(n17613), .ZN(
        n17620) );
  INV_X1 U20845 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17626) );
  XNOR2_X1 U20846 ( .A(n17616), .B(n17936), .ZN(n17961) );
  INV_X1 U20847 ( .A(n17623), .ZN(n17951) );
  NAND2_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17951), .ZN(
        n17963) );
  AOI21_X1 U20849 ( .B1(n17617), .B2(n17963), .A(n17644), .ZN(n17627) );
  OR2_X1 U20850 ( .A1(n17963), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17970) );
  OAI22_X1 U20851 ( .A1(n17627), .A2(n17936), .B1(n17673), .B2(n17970), .ZN(
        n17618) );
  AOI21_X1 U20852 ( .B1(n17765), .B2(n17961), .A(n17618), .ZN(n17619) );
  OAI211_X1 U20853 ( .C1(n18184), .C2(n18754), .A(n17620), .B(n17619), .ZN(
        P3_U2810) );
  INV_X1 U20854 ( .A(n17871), .ZN(n17827) );
  OAI21_X1 U20855 ( .B1(n17827), .B2(n17629), .A(n17798), .ZN(n17650) );
  OAI21_X1 U20856 ( .B1(n17621), .B2(n17870), .A(n17650), .ZN(n17641) );
  AOI22_X1 U20857 ( .A1(n17687), .A2(n17622), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17641), .ZN(n17634) );
  NOR2_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17623), .ZN(
        n17971) );
  OAI21_X1 U20859 ( .B1(n17637), .B2(n17635), .A(n17624), .ZN(n17625) );
  XNOR2_X1 U20860 ( .A(n17625), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17976) );
  OAI22_X1 U20861 ( .A1(n17976), .A2(n17784), .B1(n17627), .B2(n17626), .ZN(
        n17628) );
  AOI21_X1 U20862 ( .B1(n17657), .B2(n17971), .A(n17628), .ZN(n17633) );
  NAND2_X1 U20863 ( .A1(n18186), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17974) );
  NOR2_X1 U20864 ( .A1(n17630), .A2(n17629), .ZN(n17643) );
  NAND2_X1 U20865 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17631) );
  OAI211_X1 U20866 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17643), .B(n17631), .ZN(n17632) );
  NAND4_X1 U20867 ( .A1(n17634), .A2(n17633), .A3(n17974), .A4(n17632), .ZN(
        P3_U2811) );
  OAI21_X1 U20868 ( .B1(n17770), .B2(n17636), .A(n17635), .ZN(n17638) );
  XNOR2_X1 U20869 ( .A(n17638), .B(n17637), .ZN(n17991) );
  NAND2_X1 U20870 ( .A1(n18186), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17989) );
  OAI21_X1 U20871 ( .B1(n17722), .B2(n17639), .A(n17989), .ZN(n17640) );
  AOI221_X1 U20872 ( .B1(n17643), .B2(n17642), .C1(n17641), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17640), .ZN(n17647) );
  INV_X1 U20873 ( .A(n17644), .ZN(n17672) );
  OAI21_X1 U20874 ( .B1(n17980), .B2(n17673), .A(n17672), .ZN(n17656) );
  NOR2_X1 U20875 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17645), .ZN(
        n17987) );
  AOI22_X1 U20876 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17656), .B1(
        n17657), .B2(n17987), .ZN(n17646) );
  OAI211_X1 U20877 ( .C1(n17784), .C2(n17991), .A(n17647), .B(n17646), .ZN(
        P3_U2812) );
  AOI21_X1 U20878 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17649), .A(
        n17648), .ZN(n17996) );
  NOR2_X1 U20879 ( .A1(n18184), .A2(n18750), .ZN(n17654) );
  AOI221_X1 U20880 ( .B1(n17652), .B2(n17651), .C1(n18488), .C2(n17651), .A(
        n17650), .ZN(n17653) );
  AOI211_X1 U20881 ( .C1(n17655), .C2(n17844), .A(n17654), .B(n17653), .ZN(
        n17659) );
  OAI221_X1 U20882 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17657), .A(n17656), .ZN(
        n17658) );
  OAI211_X1 U20883 ( .C1(n17996), .C2(n17784), .A(n17659), .B(n17658), .ZN(
        P3_U2813) );
  NOR2_X1 U20884 ( .A1(n17770), .A2(n17660), .ZN(n17716) );
  AOI22_X1 U20885 ( .A1(n17716), .A2(n17662), .B1(n17661), .B2(n17770), .ZN(
        n17663) );
  XNOR2_X1 U20886 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17663), .ZN(
        n18005) );
  OAI211_X1 U20887 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17678), .B(n17707), .ZN(n17666) );
  OAI21_X1 U20888 ( .B1(n17678), .B2(n17773), .A(n17871), .ZN(n17693) );
  AOI21_X1 U20889 ( .B1(n17705), .B2(n17664), .A(n17693), .ZN(n17679) );
  OAI22_X1 U20890 ( .A1(n17667), .A2(n17666), .B1(n17679), .B2(n17665), .ZN(
        n17670) );
  OAI22_X1 U20891 ( .A1(n18184), .A2(n18747), .B1(n17722), .B2(n17668), .ZN(
        n17669) );
  AOI211_X1 U20892 ( .C1(n17765), .C2(n18005), .A(n17670), .B(n17669), .ZN(
        n17671) );
  OAI221_X1 U20893 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17673), 
        .C1(n18003), .C2(n17672), .A(n17671), .ZN(P3_U2814) );
  NAND3_X1 U20894 ( .A1(n17769), .A2(n17755), .A3(n17770), .ZN(n17741) );
  NOR2_X1 U20895 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17741), .ZN(
        n17726) );
  INV_X1 U20896 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17703) );
  NOR3_X1 U20897 ( .A1(n18039), .A2(n17674), .A3(n17660), .ZN(n17675) );
  AOI21_X1 U20898 ( .B1(n17726), .B2(n17703), .A(n17675), .ZN(n17676) );
  AOI221_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18059), 
        .C1(n17770), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17676), .ZN(
        n17677) );
  XOR2_X1 U20900 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17677), .Z(
        n18017) );
  INV_X1 U20901 ( .A(n18017), .ZN(n17689) );
  NAND2_X1 U20902 ( .A1(n17678), .A2(n17707), .ZN(n17681) );
  NAND2_X1 U20903 ( .A1(n18186), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18018) );
  OAI221_X1 U20904 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17681), .C1(
        n17680), .C2(n17679), .A(n18018), .ZN(n17685) );
  NOR2_X1 U20905 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17695), .ZN(
        n18014) );
  NAND2_X1 U20906 ( .A1(n17781), .A2(n12724), .ZN(n17683) );
  NOR2_X1 U20907 ( .A1(n17697), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18008) );
  NAND2_X1 U20908 ( .A1(n17839), .A2(n17940), .ZN(n17682) );
  OAI22_X1 U20909 ( .A1(n18014), .A2(n17683), .B1(n18008), .B2(n17682), .ZN(
        n17684) );
  AOI211_X1 U20910 ( .C1(n17687), .C2(n17686), .A(n17685), .B(n17684), .ZN(
        n17688) );
  OAI21_X1 U20911 ( .B1(n17784), .B2(n17689), .A(n17688), .ZN(P3_U2815) );
  OAI21_X1 U20912 ( .B1(n17691), .B2(n18488), .A(n17690), .ZN(n17692) );
  AOI22_X1 U20913 ( .A1(n18186), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17693), 
        .B2(n17692), .ZN(n17701) );
  INV_X1 U20914 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18029) );
  AOI221_X1 U20915 ( .B1(n17703), .B2(n18029), .C1(n17694), .C2(n18029), .A(
        n17695), .ZN(n18035) );
  NAND2_X1 U20916 ( .A1(n17726), .A2(n18059), .ZN(n17717) );
  NAND2_X1 U20917 ( .A1(n18022), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18026) );
  INV_X1 U20918 ( .A(n17716), .ZN(n17756) );
  OAI22_X1 U20919 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17717), .B1(
        n18026), .B2(n17756), .ZN(n17696) );
  XNOR2_X1 U20920 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17696), .ZN(
        n18033) );
  INV_X1 U20921 ( .A(n18022), .ZN(n18023) );
  NOR2_X1 U20922 ( .A1(n17739), .A2(n18023), .ZN(n18043) );
  INV_X1 U20923 ( .A(n17697), .ZN(n17698) );
  OAI221_X1 U20924 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18043), .A(n17698), .ZN(
        n18032) );
  OAI22_X1 U20925 ( .A1(n18033), .A2(n17784), .B1(n17875), .B2(n18032), .ZN(
        n17699) );
  AOI21_X1 U20926 ( .B1(n17781), .B2(n18035), .A(n17699), .ZN(n17700) );
  OAI211_X1 U20927 ( .C1(n17867), .C2(n17702), .A(n17701), .B(n17700), .ZN(
        P3_U2816) );
  NAND2_X1 U20928 ( .A1(n18022), .A2(n17703), .ZN(n18048) );
  AOI21_X1 U20929 ( .B1(n17705), .B2(n17704), .A(n17827), .ZN(n17706) );
  OAI21_X1 U20930 ( .B1(n17708), .B2(n17773), .A(n17706), .ZN(n17725) );
  NOR2_X1 U20931 ( .A1(n18184), .A2(n18741), .ZN(n17713) );
  NAND2_X1 U20932 ( .A1(n17708), .A2(n17707), .ZN(n17723) );
  OAI21_X1 U20933 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17709), .ZN(n17710) );
  OAI22_X1 U20934 ( .A1(n17722), .A2(n17711), .B1(n17723), .B2(n17710), .ZN(
        n17712) );
  AOI211_X1 U20935 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17725), .A(
        n17713), .B(n17712), .ZN(n17720) );
  INV_X1 U20936 ( .A(n17694), .ZN(n17715) );
  OAI22_X1 U20937 ( .A1(n17715), .A2(n17714), .B1(n18043), .B2(n17875), .ZN(
        n17730) );
  INV_X1 U20938 ( .A(n18039), .ZN(n18051) );
  NAND2_X1 U20939 ( .A1(n18051), .A2(n17716), .ZN(n17728) );
  OAI21_X1 U20940 ( .B1(n18059), .B2(n17728), .A(n17717), .ZN(n17718) );
  XOR2_X1 U20941 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17718), .Z(
        n18038) );
  AOI22_X1 U20942 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17730), .B1(
        n17765), .B2(n18038), .ZN(n17719) );
  OAI211_X1 U20943 ( .C1(n17768), .C2(n18048), .A(n17720), .B(n17719), .ZN(
        P3_U2817) );
  NAND2_X1 U20944 ( .A1(n18051), .A2(n18059), .ZN(n17733) );
  NOR2_X1 U20945 ( .A1(n18184), .A2(n18740), .ZN(n18056) );
  OAI22_X1 U20946 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17723), .B1(
        n17722), .B2(n17721), .ZN(n17724) );
  AOI211_X1 U20947 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17725), .A(
        n18056), .B(n17724), .ZN(n17732) );
  INV_X1 U20948 ( .A(n17726), .ZN(n17727) );
  NAND2_X1 U20949 ( .A1(n17728), .A2(n17727), .ZN(n17729) );
  XNOR2_X1 U20950 ( .A(n17729), .B(n18059), .ZN(n18057) );
  AOI22_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17730), .B1(
        n17765), .B2(n18057), .ZN(n17731) );
  OAI211_X1 U20952 ( .C1(n17768), .C2(n17733), .A(n17732), .B(n17731), .ZN(
        P3_U2818) );
  INV_X1 U20953 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18044) );
  NAND2_X1 U20954 ( .A1(n17740), .A2(n18044), .ZN(n18073) );
  NOR2_X1 U20955 ( .A1(n17734), .A2(n18488), .ZN(n17748) );
  NOR2_X1 U20956 ( .A1(n17737), .A2(n17748), .ZN(n17738) );
  INV_X1 U20957 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18737) );
  OAI22_X1 U20958 ( .A1(n17867), .A2(n17735), .B1(n18184), .B2(n18737), .ZN(
        n17736) );
  AOI221_X1 U20959 ( .B1(n17798), .B2(n17738), .C1(n17737), .C2(n17748), .A(
        n17736), .ZN(n17745) );
  AOI22_X1 U20960 ( .A1(n17839), .A2(n17739), .B1(n17781), .B2(n17660), .ZN(
        n17767) );
  OAI21_X1 U20961 ( .B1(n17740), .B2(n17768), .A(n17767), .ZN(n17743) );
  INV_X1 U20962 ( .A(n17740), .ZN(n18068) );
  OAI21_X1 U20963 ( .B1(n17756), .B2(n18068), .A(n17741), .ZN(n17742) );
  XNOR2_X1 U20964 ( .A(n17742), .B(n18044), .ZN(n18060) );
  AOI22_X1 U20965 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17743), .B1(
        n17765), .B2(n18060), .ZN(n17744) );
  OAI211_X1 U20966 ( .C1(n17768), .C2(n18073), .A(n17745), .B(n17744), .ZN(
        P3_U2819) );
  INV_X1 U20967 ( .A(n17768), .ZN(n17746) );
  NAND2_X1 U20968 ( .A1(n18068), .A2(n17746), .ZN(n17754) );
  NAND3_X1 U20969 ( .A1(n17785), .A2(n17771), .A3(n18575), .ZN(n17761) );
  NOR2_X1 U20970 ( .A1(n17760), .A2(n17761), .ZN(n17759) );
  AOI21_X1 U20971 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17798), .A(
        n17759), .ZN(n17747) );
  OAI22_X1 U20972 ( .A1(n17748), .A2(n17747), .B1(n18184), .B2(n18736), .ZN(
        n17751) );
  NAND2_X1 U20973 ( .A1(n17769), .A2(n17770), .ZN(n17757) );
  AOI22_X1 U20974 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17756), .B1(
        n17757), .B2(n18092), .ZN(n17749) );
  XNOR2_X1 U20975 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17749), .ZN(
        n18080) );
  OAI22_X1 U20976 ( .A1(n18080), .A2(n17784), .B1(n17767), .B2(n18074), .ZN(
        n17750) );
  AOI211_X1 U20977 ( .C1(n17752), .C2(n17844), .A(n17751), .B(n17750), .ZN(
        n17753) );
  OAI21_X1 U20978 ( .B1(n17755), .B2(n17754), .A(n17753), .ZN(P3_U2820) );
  NAND2_X1 U20979 ( .A1(n17757), .A2(n17756), .ZN(n17758) );
  XNOR2_X1 U20980 ( .A(n17758), .B(n18092), .ZN(n18088) );
  INV_X1 U20981 ( .A(n17798), .ZN(n17865) );
  AOI211_X1 U20982 ( .C1(n17761), .C2(n17760), .A(n17865), .B(n17759), .ZN(
        n17764) );
  OAI22_X1 U20983 ( .A1(n17867), .A2(n17762), .B1(n18184), .B2(n18735), .ZN(
        n17763) );
  AOI211_X1 U20984 ( .C1(n17765), .C2(n18088), .A(n17764), .B(n17763), .ZN(
        n17766) );
  OAI221_X1 U20985 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17768), .C1(
        n18092), .C2(n17767), .A(n17766), .ZN(P3_U2821) );
  NOR2_X1 U20986 ( .A1(n16384), .A2(n17769), .ZN(n18106) );
  XNOR2_X1 U20987 ( .A(n18106), .B(n17770), .ZN(n18111) );
  NAND2_X1 U20988 ( .A1(n17785), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17772) );
  AOI211_X1 U20989 ( .C1(n17774), .C2(n17772), .A(n17771), .B(n18488), .ZN(
        n17777) );
  OAI21_X1 U20990 ( .B1(n17773), .B2(n17785), .A(n17871), .ZN(n17786) );
  INV_X1 U20991 ( .A(n17786), .ZN(n17775) );
  OAI22_X1 U20992 ( .A1(n17775), .A2(n17774), .B1(n18184), .B2(n18734), .ZN(
        n17776) );
  AOI211_X1 U20993 ( .C1(n17778), .C2(n17844), .A(n17777), .B(n17776), .ZN(
        n17783) );
  AOI21_X1 U20994 ( .B1(n17780), .B2(n18103), .A(n17779), .ZN(n18105) );
  AOI22_X1 U20995 ( .A1(n17839), .A2(n18105), .B1(n17781), .B2(n18106), .ZN(
        n17782) );
  OAI211_X1 U20996 ( .C1(n18111), .C2(n17784), .A(n17783), .B(n17782), .ZN(
        P3_U2822) );
  AND2_X1 U20997 ( .A1(n17785), .A2(n18575), .ZN(n17788) );
  NOR2_X1 U20998 ( .A1(n18184), .A2(n18731), .ZN(n18113) );
  AOI221_X1 U20999 ( .B1(n17788), .B2(n17787), .C1(n17786), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18113), .ZN(n17796) );
  NAND2_X1 U21000 ( .A1(n17790), .A2(n17789), .ZN(n17791) );
  XNOR2_X1 U21001 ( .A(n17791), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18114) );
  AOI21_X1 U21002 ( .B1(n17794), .B2(n17793), .A(n17792), .ZN(n18115) );
  AOI22_X1 U21003 ( .A1(n17839), .A2(n18114), .B1(n17863), .B2(n18115), .ZN(
        n17795) );
  OAI211_X1 U21004 ( .C1(n17867), .C2(n17797), .A(n17796), .B(n17795), .ZN(
        P3_U2823) );
  OAI21_X1 U21005 ( .B1(n17801), .B2(n18488), .A(n17798), .ZN(n17819) );
  AOI21_X1 U21006 ( .B1(n9839), .B2(n17800), .A(n17799), .ZN(n18127) );
  NOR2_X1 U21007 ( .A1(n18184), .A2(n18729), .ZN(n18123) );
  NOR3_X1 U21008 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17801), .A3(
        n18488), .ZN(n17802) );
  AOI211_X1 U21009 ( .C1(n17863), .C2(n18127), .A(n18123), .B(n17802), .ZN(
        n17807) );
  AOI21_X1 U21010 ( .B1(n18124), .B2(n17804), .A(n17803), .ZN(n18126) );
  AOI22_X1 U21011 ( .A1(n17839), .A2(n18126), .B1(n17805), .B2(n17844), .ZN(
        n17806) );
  OAI211_X1 U21012 ( .C1(n17808), .C2(n17819), .A(n17807), .B(n17806), .ZN(
        P3_U2824) );
  AOI21_X1 U21013 ( .B1(n17809), .B2(n17871), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17820) );
  AOI21_X1 U21014 ( .B1(n17812), .B2(n17811), .A(n17810), .ZN(n18131) );
  AOI22_X1 U21015 ( .A1(n17839), .A2(n18131), .B1(n18186), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17818) );
  AOI21_X1 U21016 ( .B1(n17815), .B2(n17814), .A(n17813), .ZN(n18132) );
  AOI22_X1 U21017 ( .A1(n17863), .A2(n18132), .B1(n17816), .B2(n17844), .ZN(
        n17817) );
  OAI211_X1 U21018 ( .C1(n17820), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        P3_U2825) );
  AOI21_X1 U21019 ( .B1(n17823), .B2(n17822), .A(n17821), .ZN(n18142) );
  AOI22_X1 U21020 ( .A1(n17839), .A2(n18142), .B1(n18186), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17834) );
  AOI21_X1 U21021 ( .B1(n17826), .B2(n17825), .A(n17824), .ZN(n18136) );
  AOI21_X1 U21022 ( .B1(n17829), .B2(n17828), .A(n17827), .ZN(n17849) );
  OAI22_X1 U21023 ( .A1(n17867), .A2(n17831), .B1(n17849), .B2(n17830), .ZN(
        n17832) );
  AOI21_X1 U21024 ( .B1(n17863), .B2(n18136), .A(n17832), .ZN(n17833) );
  OAI211_X1 U21025 ( .C1(n18488), .C2(n17835), .A(n17834), .B(n17833), .ZN(
        P3_U2826) );
  AOI21_X1 U21026 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17871), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17848) );
  AOI21_X1 U21027 ( .B1(n17838), .B2(n17837), .A(n17836), .ZN(n18149) );
  AOI22_X1 U21028 ( .A1(n17839), .A2(n18149), .B1(n18186), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17847) );
  OAI21_X1 U21029 ( .B1(n17842), .B2(n17841), .A(n17840), .ZN(n17843) );
  XNOR2_X1 U21030 ( .A(n17843), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18148) );
  AOI22_X1 U21031 ( .A1(n17863), .A2(n18148), .B1(n17845), .B2(n17844), .ZN(
        n17846) );
  OAI211_X1 U21032 ( .C1(n17849), .C2(n17848), .A(n17847), .B(n17846), .ZN(
        P3_U2827) );
  INV_X1 U21033 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17857) );
  AOI21_X1 U21034 ( .B1(n9843), .B2(n17851), .A(n17850), .ZN(n18166) );
  NOR2_X1 U21035 ( .A1(n18184), .A2(n18723), .ZN(n18155) );
  XNOR2_X1 U21036 ( .A(n17853), .B(n17852), .ZN(n18170) );
  OAI22_X1 U21037 ( .A1(n17867), .A2(n17854), .B1(n17875), .B2(n18170), .ZN(
        n17855) );
  AOI211_X1 U21038 ( .C1(n17863), .C2(n18166), .A(n18155), .B(n17855), .ZN(
        n17856) );
  OAI221_X1 U21039 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18488), .C1(
        n17857), .C2(n17871), .A(n17856), .ZN(P3_U2828) );
  AOI21_X1 U21040 ( .B1(n17860), .B2(n17868), .A(n17858), .ZN(n18175) );
  NAND2_X1 U21041 ( .A1(n18818), .A2(n17859), .ZN(n17861) );
  XNOR2_X1 U21042 ( .A(n17861), .B(n17860), .ZN(n18181) );
  OAI22_X1 U21043 ( .A1(n18181), .A2(n17875), .B1(n18184), .B2(n20926), .ZN(
        n17862) );
  AOI21_X1 U21044 ( .B1(n17863), .B2(n18175), .A(n17862), .ZN(n17864) );
  OAI221_X1 U21045 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17867), .C1(
        n17866), .C2(n17865), .A(n17864), .ZN(P3_U2829) );
  OAI21_X1 U21046 ( .B1(n17869), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17868), .ZN(n18189) );
  INV_X1 U21047 ( .A(n18189), .ZN(n18191) );
  NAND3_X1 U21048 ( .A1(n18800), .A2(n17871), .A3(n17870), .ZN(n17872) );
  AOI22_X1 U21049 ( .A1(n18186), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17872), .ZN(n17873) );
  OAI221_X1 U21050 ( .B1(n18191), .B2(n17875), .C1(n18189), .C2(n17874), .A(
        n17873), .ZN(P3_U2830) );
  AOI22_X1 U21051 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18178), .B1(
        n18186), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17890) );
  NOR3_X1 U21052 ( .A1(n17894), .A2(n17876), .A3(n17892), .ZN(n17888) );
  INV_X1 U21053 ( .A(n17877), .ZN(n17885) );
  INV_X1 U21054 ( .A(n18095), .ZN(n18158) );
  NOR2_X1 U21055 ( .A1(n18082), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18160) );
  AOI21_X1 U21056 ( .B1(n18095), .B2(n17878), .A(n18160), .ZN(n17919) );
  OAI21_X1 U21057 ( .B1(n18158), .B2(n17879), .A(n17919), .ZN(n17901) );
  INV_X1 U21058 ( .A(n18041), .ZN(n18063) );
  AOI22_X1 U21059 ( .A1(n18642), .A2(n20775), .B1(n18663), .B2(n17880), .ZN(
        n17882) );
  OAI211_X1 U21060 ( .C1(n17883), .C2(n18063), .A(n17882), .B(n17881), .ZN(
        n17884) );
  AOI211_X1 U21061 ( .C1(n18630), .C2(n17885), .A(n17901), .B(n17884), .ZN(
        n17896) );
  OAI21_X1 U21062 ( .B1(n18665), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17896), .ZN(n17886) );
  OAI221_X1 U21063 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17888), 
        .C1(n17887), .C2(n17886), .A(n18182), .ZN(n17889) );
  OAI211_X1 U21064 ( .C1(n17891), .C2(n18110), .A(n17890), .B(n17889), .ZN(
        P3_U2835) );
  INV_X1 U21065 ( .A(n17892), .ZN(n17930) );
  NAND2_X1 U21066 ( .A1(n17893), .A2(n17930), .ZN(n17895) );
  AOI221_X1 U21067 ( .B1(n17896), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n17895), .C2(n17894), .A(n18176), .ZN(n17897) );
  AOI21_X1 U21068 ( .B1(n18178), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17897), .ZN(n17899) );
  OAI211_X1 U21069 ( .C1(n17900), .C2(n18110), .A(n17899), .B(n17898), .ZN(
        P3_U2836) );
  OAI21_X1 U21070 ( .B1(n17902), .B2(n17901), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17903) );
  OAI21_X1 U21071 ( .B1(n17905), .B2(n17904), .A(n17903), .ZN(n17906) );
  AOI22_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18178), .B1(
        n18182), .B2(n17906), .ZN(n17908) );
  OAI211_X1 U21073 ( .C1(n17909), .C2(n18110), .A(n17908), .B(n17907), .ZN(
        n17910) );
  AOI21_X1 U21074 ( .B1(n18150), .B2(n17911), .A(n17910), .ZN(n17912) );
  OAI21_X1 U21075 ( .B1(n17914), .B2(n17913), .A(n17912), .ZN(P3_U2837) );
  NAND2_X1 U21076 ( .A1(n18182), .A2(n17915), .ZN(n17969) );
  AOI22_X1 U21077 ( .A1(n18186), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18089), 
        .B2(n17916), .ZN(n17927) );
  INV_X1 U21078 ( .A(n18630), .ZN(n18062) );
  AOI21_X1 U21079 ( .B1(n18041), .B2(n17917), .A(n18178), .ZN(n17918) );
  OAI211_X1 U21080 ( .C1(n17920), .C2(n18062), .A(n17919), .B(n17918), .ZN(
        n17925) );
  INV_X1 U21081 ( .A(n17921), .ZN(n17923) );
  AOI211_X1 U21082 ( .C1(n18661), .C2(n17923), .A(n17922), .B(n17925), .ZN(
        n17924) );
  NOR2_X1 U21083 ( .A1(n18186), .A2(n17924), .ZN(n17929) );
  OAI211_X1 U21084 ( .C1(n18100), .C2(n17925), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17929), .ZN(n17926) );
  OAI211_X1 U21085 ( .C1(n17928), .C2(n17969), .A(n17927), .B(n17926), .ZN(
        P3_U2838) );
  OAI221_X1 U21086 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17930), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18141), .A(n17929), .ZN(
        n17931) );
  OAI211_X1 U21087 ( .C1(n17933), .C2(n18110), .A(n17932), .B(n17931), .ZN(
        P3_U2839) );
  INV_X1 U21088 ( .A(n17969), .ZN(n17972) );
  AOI22_X1 U21089 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18182), .B1(
        n17938), .B2(n17972), .ZN(n17950) );
  NAND2_X1 U21090 ( .A1(n18062), .A2(n18063), .ZN(n18067) );
  INV_X1 U21091 ( .A(n18067), .ZN(n17979) );
  OAI21_X1 U21092 ( .B1(n17977), .B2(n17963), .A(n18642), .ZN(n17934) );
  OAI221_X1 U21093 ( .B1(n18644), .B2(n17935), .C1(n18644), .C2(n17951), .A(
        n17934), .ZN(n17962) );
  AOI21_X1 U21094 ( .B1(n18642), .B2(n17936), .A(n17962), .ZN(n17937) );
  OAI21_X1 U21095 ( .B1(n17938), .B2(n17979), .A(n17937), .ZN(n17956) );
  INV_X1 U21096 ( .A(n17939), .ZN(n17954) );
  AOI22_X1 U21097 ( .A1(n18630), .A2(n17940), .B1(n18041), .B2(n12724), .ZN(
        n17952) );
  OAI21_X1 U21098 ( .B1(n17942), .B2(n18663), .A(n17941), .ZN(n17943) );
  OAI211_X1 U21099 ( .C1(n17954), .C2(n18644), .A(n17952), .B(n17943), .ZN(
        n17944) );
  AOI211_X1 U21100 ( .C1(n17999), .C2(n17945), .A(n17956), .B(n17944), .ZN(
        n17949) );
  AOI22_X1 U21101 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18178), .B1(
        n18089), .B2(n17946), .ZN(n17948) );
  OAI211_X1 U21102 ( .C1(n17950), .C2(n17949), .A(n17948), .B(n17947), .ZN(
        P3_U2840) );
  NOR2_X1 U21103 ( .A1(n18661), .A2(n18663), .ZN(n18177) );
  NAND2_X1 U21104 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17997), .ZN(
        n18021) );
  NOR2_X1 U21105 ( .A1(n17986), .A2(n18021), .ZN(n18001) );
  AOI21_X1 U21106 ( .B1(n17951), .B2(n18001), .A(n18082), .ZN(n17953) );
  NAND2_X1 U21107 ( .A1(n18182), .A2(n17952), .ZN(n18002) );
  NOR2_X1 U21108 ( .A1(n17953), .A2(n18002), .ZN(n17964) );
  OAI21_X1 U21109 ( .B1(n17954), .B2(n18177), .A(n17964), .ZN(n17955) );
  OAI21_X1 U21110 ( .B1(n17956), .B2(n17955), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17960) );
  AOI22_X1 U21111 ( .A1(n18089), .A2(n17958), .B1(n17972), .B2(n17957), .ZN(
        n17959) );
  OAI221_X1 U21112 ( .B1(n18186), .B2(n17960), .C1(n18184), .C2(n18756), .A(
        n17959), .ZN(P3_U2841) );
  AOI22_X1 U21113 ( .A1(n18186), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18089), 
        .B2(n17961), .ZN(n17968) );
  AOI21_X1 U21114 ( .B1(n17963), .B2(n18067), .A(n17962), .ZN(n17965) );
  AOI21_X1 U21115 ( .B1(n17965), .B2(n17964), .A(n18186), .ZN(n17973) );
  NOR3_X1 U21116 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18177), .A3(
        n18836), .ZN(n17966) );
  OAI21_X1 U21117 ( .B1(n17973), .B2(n17966), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17967) );
  OAI211_X1 U21118 ( .C1(n17970), .C2(n17969), .A(n17968), .B(n17967), .ZN(
        P3_U2842) );
  AOI22_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17973), .B1(
        n17972), .B2(n17971), .ZN(n17975) );
  OAI211_X1 U21120 ( .C1(n17976), .C2(n18110), .A(n17975), .B(n17974), .ZN(
        P3_U2843) );
  NOR3_X1 U21121 ( .A1(n18160), .A2(n17977), .A3(n18003), .ZN(n17978) );
  OAI22_X1 U21122 ( .A1(n17980), .A2(n17979), .B1(n18158), .B2(n17978), .ZN(
        n17981) );
  AOI211_X1 U21123 ( .C1(n18661), .C2(n17982), .A(n18002), .B(n17981), .ZN(
        n17992) );
  AOI221_X1 U21124 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17992), 
        .C1(n18158), .C2(n17992), .A(n18186), .ZN(n17988) );
  INV_X1 U21125 ( .A(n18137), .ZN(n18161) );
  INV_X1 U21126 ( .A(n18138), .ZN(n17983) );
  OAI22_X1 U21127 ( .A1(n18161), .A2(n18644), .B1(n18165), .B2(n17983), .ZN(
        n18147) );
  NAND2_X1 U21128 ( .A1(n17984), .A2(n18147), .ZN(n18120) );
  OAI21_X1 U21129 ( .B1(n18010), .B2(n18120), .A(n17985), .ZN(n18050) );
  NAND2_X1 U21130 ( .A1(n18182), .A2(n18050), .ZN(n18093) );
  NOR2_X1 U21131 ( .A1(n17986), .A2(n18093), .ZN(n18004) );
  AOI22_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17988), .B1(
        n18004), .B2(n17987), .ZN(n17990) );
  OAI211_X1 U21133 ( .C1(n18110), .C2(n17991), .A(n17990), .B(n17989), .ZN(
        P3_U2844) );
  NOR2_X1 U21134 ( .A1(n18186), .A2(n17992), .ZN(n17993) );
  AOI22_X1 U21135 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17993), .B1(
        n18186), .B2(P3_REIP_REG_17__SCAN_IN), .ZN(n17995) );
  INV_X1 U21136 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20905) );
  NAND3_X1 U21137 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18004), .A3(
        n20905), .ZN(n17994) );
  OAI211_X1 U21138 ( .C1(n17996), .C2(n18110), .A(n17995), .B(n17994), .ZN(
        P3_U2845) );
  OAI22_X1 U21139 ( .A1(n18665), .A2(n17997), .B1(n18085), .B2(n18644), .ZN(
        n18066) );
  AOI21_X1 U21140 ( .B1(n17999), .B2(n17998), .A(n18066), .ZN(n18000) );
  OAI211_X1 U21141 ( .C1(n18001), .C2(n18082), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18000), .ZN(n18011) );
  OAI221_X1 U21142 ( .B1(n18002), .B2(n18100), .C1(n18002), .C2(n18011), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U21143 ( .A1(n18089), .A2(n18005), .B1(n18004), .B2(n18003), .ZN(
        n18006) );
  OAI221_X1 U21144 ( .B1(n18186), .B2(n18007), .C1(n18184), .C2(n18747), .A(
        n18006), .ZN(P3_U2846) );
  NOR3_X1 U21145 ( .A1(n18009), .A2(n18008), .A3(n18190), .ZN(n18016) );
  NOR3_X1 U21146 ( .A1(n18010), .A2(n18120), .A3(n18026), .ZN(n18031) );
  OAI221_X1 U21147 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18031), .A(n18011), .ZN(
        n18013) );
  NAND2_X1 U21148 ( .A1(n18041), .A2(n12724), .ZN(n18012) );
  AOI221_X1 U21149 ( .B1(n18014), .B2(n18013), .C1(n18012), .C2(n18013), .A(
        n18176), .ZN(n18015) );
  AOI211_X1 U21150 ( .C1(n18017), .C2(n18089), .A(n18016), .B(n18015), .ZN(
        n18019) );
  OAI211_X1 U21151 ( .C1(n18141), .C2(n18020), .A(n18019), .B(n18018), .ZN(
        P3_U2847) );
  INV_X1 U21152 ( .A(n18066), .ZN(n18025) );
  INV_X1 U21153 ( .A(n18021), .ZN(n18081) );
  AOI21_X1 U21154 ( .B1(n18022), .B2(n18081), .A(n18082), .ZN(n18040) );
  AOI211_X1 U21155 ( .C1(n18661), .C2(n18023), .A(n18040), .B(n18029), .ZN(
        n18024) );
  OAI211_X1 U21156 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18177), .A(
        n18025), .B(n18024), .ZN(n18027) );
  OAI221_X1 U21157 ( .B1(n18027), .B2(n18642), .C1(n18027), .C2(n18026), .A(
        n18182), .ZN(n18028) );
  OAI21_X1 U21158 ( .B1(n18141), .B2(n18029), .A(n18028), .ZN(n18030) );
  OAI21_X1 U21159 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18031), .A(
        n18030), .ZN(n18037) );
  OAI22_X1 U21160 ( .A1(n18033), .A2(n18110), .B1(n18190), .B2(n18032), .ZN(
        n18034) );
  AOI21_X1 U21161 ( .B1(n18107), .B2(n18035), .A(n18034), .ZN(n18036) );
  OAI211_X1 U21162 ( .C1(n18184), .C2(n18744), .A(n18037), .B(n18036), .ZN(
        P3_U2848) );
  AOI22_X1 U21163 ( .A1(n18186), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18089), 
        .B2(n18038), .ZN(n18047) );
  AOI22_X1 U21164 ( .A1(n18661), .A2(n18039), .B1(n18642), .B2(n18068), .ZN(
        n18069) );
  AOI211_X1 U21165 ( .C1(n18041), .C2(n17694), .A(n18040), .B(n18066), .ZN(
        n18042) );
  OAI211_X1 U21166 ( .C1(n18043), .C2(n18062), .A(n18069), .B(n18042), .ZN(
        n18049) );
  AOI21_X1 U21167 ( .B1(n18642), .B2(n18044), .A(n18059), .ZN(n18053) );
  OAI21_X1 U21168 ( .B1(n18076), .B2(n18053), .A(n18182), .ZN(n18045) );
  OAI211_X1 U21169 ( .C1(n18049), .C2(n18045), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18184), .ZN(n18046) );
  OAI211_X1 U21170 ( .C1(n18093), .C2(n18048), .A(n18047), .B(n18046), .ZN(
        P3_U2849) );
  INV_X1 U21171 ( .A(n18049), .ZN(n18054) );
  AOI21_X1 U21172 ( .B1(n18051), .B2(n18050), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18052) );
  AOI211_X1 U21173 ( .C1(n18054), .C2(n18053), .A(n18052), .B(n18176), .ZN(
        n18055) );
  AOI211_X1 U21174 ( .C1(n18089), .C2(n18057), .A(n18056), .B(n18055), .ZN(
        n18058) );
  OAI21_X1 U21175 ( .B1(n18059), .B2(n18141), .A(n18058), .ZN(P3_U2850) );
  AOI22_X1 U21176 ( .A1(n18186), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18089), 
        .B2(n18060), .ZN(n18072) );
  OAI22_X1 U21177 ( .A1(n16384), .A2(n18063), .B1(n18062), .B2(n18061), .ZN(
        n18064) );
  NOR2_X1 U21178 ( .A1(n18176), .A2(n18064), .ZN(n18084) );
  OAI221_X1 U21179 ( .B1(n18082), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18082), .C2(n18081), .A(n18084), .ZN(n18065) );
  AOI211_X1 U21180 ( .C1(n18068), .C2(n18067), .A(n18066), .B(n18065), .ZN(
        n18075) );
  OAI211_X1 U21181 ( .C1(n18082), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18069), .B(n18075), .ZN(n18070) );
  NAND3_X1 U21182 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18184), .A3(
        n18070), .ZN(n18071) );
  OAI211_X1 U21183 ( .C1(n18073), .C2(n18093), .A(n18072), .B(n18071), .ZN(
        P3_U2851) );
  AOI221_X1 U21184 ( .B1(n18076), .B2(n18075), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18075), .A(n18074), .ZN(
        n18078) );
  NOR3_X1 U21185 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18092), .A3(
        n18093), .ZN(n18077) );
  AOI221_X1 U21186 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18186), .C1(n18078), 
        .C2(n18184), .A(n18077), .ZN(n18079) );
  OAI21_X1 U21187 ( .B1(n18080), .B2(n18110), .A(n18079), .ZN(P3_U2852) );
  AOI211_X1 U21188 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18082), .A(
        n18158), .B(n18081), .ZN(n18087) );
  OAI21_X1 U21189 ( .B1(n18094), .B2(n18099), .A(n18642), .ZN(n18083) );
  OAI211_X1 U21190 ( .C1(n18085), .C2(n18644), .A(n18084), .B(n18083), .ZN(
        n18086) );
  OAI21_X1 U21191 ( .B1(n18087), .B2(n18086), .A(n18184), .ZN(n18091) );
  AOI22_X1 U21192 ( .A1(n18186), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18089), 
        .B2(n18088), .ZN(n18090) );
  OAI221_X1 U21193 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18093), .C1(
        n18092), .C2(n18091), .A(n18090), .ZN(P3_U2853) );
  NOR3_X1 U21194 ( .A1(n18176), .A2(n18099), .A3(n18120), .ZN(n18104) );
  AOI22_X1 U21195 ( .A1(n18661), .A2(n18096), .B1(n18095), .B2(n18094), .ZN(
        n18098) );
  INV_X1 U21196 ( .A(n18160), .ZN(n18097) );
  NAND2_X1 U21197 ( .A1(n18098), .A2(n18097), .ZN(n18121) );
  AOI21_X1 U21198 ( .B1(n18100), .B2(n18099), .A(n18121), .ZN(n18119) );
  OAI21_X1 U21199 ( .B1(n18119), .B2(n18171), .A(n18141), .ZN(n18102) );
  NOR2_X1 U21200 ( .A1(n18184), .A2(n18734), .ZN(n18101) );
  AOI221_X1 U21201 ( .B1(n18104), .B2(n18103), .C1(n18102), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18101), .ZN(n18109) );
  AOI22_X1 U21202 ( .A1(n18107), .A2(n18106), .B1(n18150), .B2(n18105), .ZN(
        n18108) );
  OAI211_X1 U21203 ( .C1(n18111), .C2(n18110), .A(n18109), .B(n18108), .ZN(
        P3_U2854) );
  INV_X1 U21204 ( .A(n18120), .ZN(n18112) );
  OAI221_X1 U21205 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18112), .A(n18182), .ZN(
        n18118) );
  AOI21_X1 U21206 ( .B1(n18178), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18113), .ZN(n18117) );
  AOI22_X1 U21207 ( .A1(n18174), .A2(n18115), .B1(n18150), .B2(n18114), .ZN(
        n18116) );
  OAI211_X1 U21208 ( .C1(n18119), .C2(n18118), .A(n18117), .B(n18116), .ZN(
        P3_U2855) );
  NOR2_X1 U21209 ( .A1(n18176), .A2(n18120), .ZN(n18125) );
  INV_X1 U21210 ( .A(n18121), .ZN(n18122) );
  OAI21_X1 U21211 ( .B1(n18122), .B2(n18176), .A(n18141), .ZN(n18130) );
  AOI221_X1 U21212 ( .B1(n18125), .B2(n18124), .C1(n18130), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18123), .ZN(n18129) );
  AOI22_X1 U21213 ( .A1(n18174), .A2(n18127), .B1(n18150), .B2(n18126), .ZN(
        n18128) );
  NAND2_X1 U21214 ( .A1(n18129), .A2(n18128), .ZN(P3_U2856) );
  NAND4_X1 U21215 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n18182), .A4(n18147), .ZN(
        n18135) );
  AOI22_X1 U21216 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18130), .B1(
        n18186), .B2(P3_REIP_REG_5__SCAN_IN), .ZN(n18134) );
  AOI22_X1 U21217 ( .A1(n18174), .A2(n18132), .B1(n18150), .B2(n18131), .ZN(
        n18133) );
  OAI211_X1 U21218 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18135), .A(
        n18134), .B(n18133), .ZN(P3_U2857) );
  NAND3_X1 U21219 ( .A1(n18182), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18147), .ZN(n18146) );
  AOI22_X1 U21220 ( .A1(n18186), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18174), 
        .B2(n18136), .ZN(n18145) );
  OAI22_X1 U21221 ( .A1(n18158), .A2(n18138), .B1(n18644), .B2(n18137), .ZN(
        n18139) );
  NOR3_X1 U21222 ( .A1(n18160), .A2(n18140), .A3(n18139), .ZN(n18154) );
  OAI21_X1 U21223 ( .B1(n18154), .B2(n18171), .A(n18141), .ZN(n18143) );
  AOI22_X1 U21224 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18143), .B1(
        n18150), .B2(n18142), .ZN(n18144) );
  OAI211_X1 U21225 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18146), .A(
        n18145), .B(n18144), .ZN(P3_U2858) );
  OAI21_X1 U21226 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18147), .A(
        n18182), .ZN(n18153) );
  AOI22_X1 U21227 ( .A1(n18186), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18174), 
        .B2(n18148), .ZN(n18152) );
  AOI22_X1 U21228 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18178), .B1(
        n18150), .B2(n18149), .ZN(n18151) );
  OAI211_X1 U21229 ( .C1(n18154), .C2(n18153), .A(n18152), .B(n18151), .ZN(
        P3_U2859) );
  AOI21_X1 U21230 ( .B1(n18178), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18155), .ZN(n18169) );
  NAND2_X1 U21231 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18156), .ZN(
        n18164) );
  NAND2_X1 U21232 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18157) );
  OAI22_X1 U21233 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18158), .B1(
        n18644), .B2(n18157), .ZN(n18159) );
  OAI21_X1 U21234 ( .B1(n18160), .B2(n18159), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18163) );
  NAND2_X1 U21235 ( .A1(n18661), .A2(n18161), .ZN(n18162) );
  OAI211_X1 U21236 ( .C1(n18165), .C2(n18164), .A(n18163), .B(n18162), .ZN(
        n18167) );
  AOI22_X1 U21237 ( .A1(n18182), .A2(n18167), .B1(n18174), .B2(n18166), .ZN(
        n18168) );
  OAI211_X1 U21238 ( .C1(n18190), .C2(n18170), .A(n18169), .B(n18168), .ZN(
        P3_U2860) );
  NOR2_X1 U21239 ( .A1(n18184), .A2(n20926), .ZN(n18173) );
  AOI211_X1 U21240 ( .C1(n18665), .C2(n18818), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18171), .ZN(n18172) );
  AOI211_X1 U21241 ( .C1(n18175), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        n18180) );
  NOR3_X1 U21242 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18177), .A3(
        n18176), .ZN(n18183) );
  OAI21_X1 U21243 ( .B1(n18178), .B2(n18183), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18179) );
  OAI211_X1 U21244 ( .C1(n18181), .C2(n18190), .A(n18180), .B(n18179), .ZN(
        P3_U2861) );
  AOI21_X1 U21245 ( .B1(n18665), .B2(n18182), .A(n18818), .ZN(n18185) );
  AOI221_X1 U21246 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18186), .C1(n18185), 
        .C2(n18184), .A(n18183), .ZN(n18187) );
  OAI221_X1 U21247 ( .B1(n18191), .B2(n18190), .C1(n18189), .C2(n18188), .A(
        n18187), .ZN(P3_U2862) );
  AOI21_X1 U21248 ( .B1(n18194), .B2(n18193), .A(n18192), .ZN(n18688) );
  INV_X1 U21249 ( .A(n18371), .ZN(n18240) );
  OAI21_X1 U21250 ( .B1(n18688), .B2(n18240), .A(n18199), .ZN(n18195) );
  OAI221_X1 U21251 ( .B1(n18668), .B2(n18842), .C1(n18668), .C2(n18199), .A(
        n18195), .ZN(P3_U2863) );
  INV_X1 U21252 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18677) );
  NOR2_X1 U21253 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18674), .ZN(
        n18373) );
  NAND2_X1 U21254 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18674), .ZN(
        n18418) );
  INV_X1 U21255 ( .A(n18418), .ZN(n18464) );
  NOR2_X1 U21256 ( .A1(n18373), .A2(n18464), .ZN(n18197) );
  OAI22_X1 U21257 ( .A1(n18198), .A2(n18677), .B1(n18197), .B2(n18196), .ZN(
        P3_U2866) );
  NOR2_X1 U21258 ( .A1(n18678), .A2(n18199), .ZN(P3_U2867) );
  NAND2_X1 U21259 ( .A1(n18575), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18579) );
  NOR2_X1 U21260 ( .A1(n18677), .A2(n18348), .ZN(n18573) );
  NAND2_X1 U21261 ( .A1(n18573), .A2(n18668), .ZN(n18559) );
  NAND2_X1 U21262 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18575), .ZN(n18545) );
  INV_X1 U21263 ( .A(n18545), .ZN(n18571) );
  NAND2_X1 U21264 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20932), .ZN(
        n18419) );
  NAND2_X1 U21265 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18512) );
  NOR2_X2 U21266 ( .A1(n18419), .A2(n18512), .ZN(n18612) );
  NOR2_X2 U21267 ( .A1(n18486), .A2(n18200), .ZN(n18570) );
  NAND2_X1 U21268 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18573), .ZN(
        n18617) );
  NAND2_X1 U21269 ( .A1(n20932), .A2(n18668), .ZN(n18670) );
  NAND2_X1 U21270 ( .A1(n18674), .A2(n18677), .ZN(n18260) );
  NOR2_X2 U21271 ( .A1(n18670), .A2(n18260), .ZN(n18296) );
  INV_X1 U21272 ( .A(n18296), .ZN(n18303) );
  AOI21_X1 U21273 ( .B1(n18617), .B2(n18303), .A(n18569), .ZN(n18234) );
  AOI22_X1 U21274 ( .A1(n18571), .A2(n18612), .B1(n18570), .B2(n18234), .ZN(
        n18205) );
  INV_X1 U21275 ( .A(n18612), .ZN(n18628) );
  NAND2_X1 U21276 ( .A1(n18559), .A2(n18628), .ZN(n18542) );
  OAI21_X1 U21277 ( .B1(n18668), .B2(n18789), .A(n18305), .ZN(n18441) );
  AOI21_X1 U21278 ( .B1(n18617), .B2(n18303), .A(n18441), .ZN(n18262) );
  AOI21_X1 U21279 ( .B1(n18575), .B2(n18542), .A(n18262), .ZN(n18237) );
  NOR2_X1 U21280 ( .A1(n18202), .A2(n18201), .ZN(n18228) );
  INV_X1 U21281 ( .A(n18228), .ZN(n18235) );
  NOR2_X2 U21282 ( .A1(n18203), .A2(n18235), .ZN(n18576) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18237), .B1(
        n18576), .B2(n18296), .ZN(n18204) );
  OAI211_X1 U21284 ( .C1(n18579), .C2(n18559), .A(n18205), .B(n18204), .ZN(
        P3_U2868) );
  NAND2_X1 U21285 ( .A1(n18575), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18521) );
  AND2_X1 U21286 ( .A1(n18305), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18580) );
  NAND2_X1 U21287 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18575), .ZN(n18586) );
  INV_X1 U21288 ( .A(n18586), .ZN(n18518) );
  AOI22_X1 U21289 ( .A1(n18580), .A2(n18234), .B1(n18518), .B2(n18612), .ZN(
        n18208) );
  NOR2_X2 U21290 ( .A1(n18206), .A2(n18235), .ZN(n18582) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18237), .B1(
        n18582), .B2(n18296), .ZN(n18207) );
  OAI211_X1 U21292 ( .C1(n18521), .C2(n18559), .A(n18208), .B(n18207), .ZN(
        P3_U2869) );
  NAND2_X1 U21293 ( .A1(n18228), .A2(n18209), .ZN(n18592) );
  NOR2_X2 U21294 ( .A1(n18486), .A2(n18210), .ZN(n18587) );
  NOR2_X2 U21295 ( .A1(n18488), .A2(n18211), .ZN(n18589) );
  INV_X1 U21296 ( .A(n18559), .ZN(n18562) );
  AOI22_X1 U21297 ( .A1(n18587), .A2(n18234), .B1(n18589), .B2(n18562), .ZN(
        n18213) );
  AND2_X1 U21298 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18575), .ZN(n18588) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18237), .B1(
        n18588), .B2(n18612), .ZN(n18212) );
  OAI211_X1 U21300 ( .C1(n18592), .C2(n18303), .A(n18213), .B(n18212), .ZN(
        P3_U2870) );
  NAND2_X1 U21301 ( .A1(n18228), .A2(n18214), .ZN(n18598) );
  NOR2_X2 U21302 ( .A1(n18215), .A2(n18488), .ZN(n18594) );
  AND2_X1 U21303 ( .A1(n18305), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18593) );
  AOI22_X1 U21304 ( .A1(n18594), .A2(n18612), .B1(n18593), .B2(n18234), .ZN(
        n18217) );
  NOR2_X2 U21305 ( .A1(n18488), .A2(n15118), .ZN(n18595) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18237), .B1(
        n18595), .B2(n18562), .ZN(n18216) );
  OAI211_X1 U21307 ( .C1(n18598), .C2(n18303), .A(n18217), .B(n18216), .ZN(
        P3_U2871) );
  OR2_X1 U21308 ( .A1(n18235), .A2(n18218), .ZN(n18604) );
  NOR2_X2 U21309 ( .A1(n18488), .A2(n18219), .ZN(n18600) );
  NOR2_X2 U21310 ( .A1(n18486), .A2(n18220), .ZN(n18599) );
  AOI22_X1 U21311 ( .A1(n18600), .A2(n18562), .B1(n18599), .B2(n18234), .ZN(
        n18222) );
  AND2_X1 U21312 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18575), .ZN(n18601) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18237), .B1(
        n18601), .B2(n18612), .ZN(n18221) );
  OAI211_X1 U21314 ( .C1(n18604), .C2(n18303), .A(n18222), .B(n18221), .ZN(
        P3_U2872) );
  NAND2_X1 U21315 ( .A1(n18228), .A2(n18223), .ZN(n18610) );
  NOR2_X2 U21316 ( .A1(n19200), .A2(n18488), .ZN(n18607) );
  NOR2_X2 U21317 ( .A1(n18486), .A2(n18224), .ZN(n18606) );
  AOI22_X1 U21318 ( .A1(n18607), .A2(n18612), .B1(n18606), .B2(n18234), .ZN(
        n18226) );
  NOR2_X2 U21319 ( .A1(n18488), .A2(n15107), .ZN(n18605) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18237), .B1(
        n18605), .B2(n18562), .ZN(n18225) );
  OAI211_X1 U21321 ( .C1(n18610), .C2(n18303), .A(n18226), .B(n18225), .ZN(
        P3_U2873) );
  NAND2_X1 U21322 ( .A1(n18228), .A2(n18227), .ZN(n18618) );
  NOR2_X2 U21323 ( .A1(n20757), .A2(n18488), .ZN(n18614) );
  NOR2_X2 U21324 ( .A1(n18229), .A2(n18486), .ZN(n18611) );
  AOI22_X1 U21325 ( .A1(n18614), .A2(n18612), .B1(n18611), .B2(n18234), .ZN(
        n18231) );
  NOR2_X2 U21326 ( .A1(n19208), .A2(n18488), .ZN(n18613) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18237), .B1(
        n18613), .B2(n18562), .ZN(n18230) );
  OAI211_X1 U21328 ( .C1(n18618), .C2(n18303), .A(n18231), .B(n18230), .ZN(
        P3_U2874) );
  NAND2_X1 U21329 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18575), .ZN(n18629) );
  NOR2_X1 U21330 ( .A1(n18488), .A2(n18232), .ZN(n18622) );
  NOR2_X2 U21331 ( .A1(n18233), .A2(n18486), .ZN(n18620) );
  AOI22_X1 U21332 ( .A1(n18622), .A2(n18612), .B1(n18620), .B2(n18234), .ZN(
        n18239) );
  NOR2_X2 U21333 ( .A1(n18236), .A2(n18235), .ZN(n18624) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18237), .B1(
        n18624), .B2(n18296), .ZN(n18238) );
  OAI211_X1 U21335 ( .C1(n18629), .C2(n18559), .A(n18239), .B(n18238), .ZN(
        P3_U2875) );
  INV_X1 U21336 ( .A(n18579), .ZN(n18538) );
  INV_X1 U21337 ( .A(n18617), .ZN(n18623) );
  OR2_X1 U21338 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18569), .ZN(
        n18511) );
  NOR2_X1 U21339 ( .A1(n18260), .A2(n18511), .ZN(n18256) );
  AOI22_X1 U21340 ( .A1(n18538), .A2(n18623), .B1(n18570), .B2(n18256), .ZN(
        n18242) );
  INV_X1 U21341 ( .A(n18260), .ZN(n18281) );
  NOR2_X1 U21342 ( .A1(n18486), .A2(n18240), .ZN(n18572) );
  AND2_X1 U21343 ( .A1(n20932), .A2(n18572), .ZN(n18513) );
  AOI22_X1 U21344 ( .A1(n18575), .A2(n18573), .B1(n18281), .B2(n18513), .ZN(
        n18257) );
  NOR2_X2 U21345 ( .A1(n18260), .A2(n18419), .ZN(n18322) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18257), .B1(
        n18322), .B2(n18576), .ZN(n18241) );
  OAI211_X1 U21347 ( .C1(n18545), .C2(n18559), .A(n18242), .B(n18241), .ZN(
        P3_U2876) );
  INV_X1 U21348 ( .A(n18521), .ZN(n18581) );
  AOI22_X1 U21349 ( .A1(n18581), .A2(n18623), .B1(n18580), .B2(n18256), .ZN(
        n18244) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18257), .B1(
        n18322), .B2(n18582), .ZN(n18243) );
  OAI211_X1 U21351 ( .C1(n18586), .C2(n18559), .A(n18244), .B(n18243), .ZN(
        P3_U2877) );
  INV_X1 U21352 ( .A(n18322), .ZN(n18255) );
  AOI22_X1 U21353 ( .A1(n18588), .A2(n18562), .B1(n18587), .B2(n18256), .ZN(
        n18246) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18257), .B1(
        n18589), .B2(n18623), .ZN(n18245) );
  OAI211_X1 U21355 ( .C1(n18255), .C2(n18592), .A(n18246), .B(n18245), .ZN(
        P3_U2878) );
  AOI22_X1 U21356 ( .A1(n18594), .A2(n18562), .B1(n18593), .B2(n18256), .ZN(
        n18248) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18257), .B1(
        n18595), .B2(n18623), .ZN(n18247) );
  OAI211_X1 U21358 ( .C1(n18255), .C2(n18598), .A(n18248), .B(n18247), .ZN(
        P3_U2879) );
  AOI22_X1 U21359 ( .A1(n18600), .A2(n18623), .B1(n18599), .B2(n18256), .ZN(
        n18250) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18257), .B1(
        n18601), .B2(n18562), .ZN(n18249) );
  OAI211_X1 U21361 ( .C1(n18255), .C2(n18604), .A(n18250), .B(n18249), .ZN(
        P3_U2880) );
  AOI22_X1 U21362 ( .A1(n18606), .A2(n18256), .B1(n18605), .B2(n18623), .ZN(
        n18252) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18257), .B1(
        n18607), .B2(n18562), .ZN(n18251) );
  OAI211_X1 U21364 ( .C1(n18255), .C2(n18610), .A(n18252), .B(n18251), .ZN(
        P3_U2881) );
  AOI22_X1 U21365 ( .A1(n18613), .A2(n18623), .B1(n18611), .B2(n18256), .ZN(
        n18254) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18257), .B1(
        n18614), .B2(n18562), .ZN(n18253) );
  OAI211_X1 U21367 ( .C1(n18255), .C2(n18618), .A(n18254), .B(n18253), .ZN(
        P3_U2882) );
  INV_X1 U21368 ( .A(n18622), .ZN(n18567) );
  INV_X1 U21369 ( .A(n18629), .ZN(n18561) );
  AOI22_X1 U21370 ( .A1(n18561), .A2(n18623), .B1(n18620), .B2(n18256), .ZN(
        n18259) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18257), .B1(
        n18322), .B2(n18624), .ZN(n18258) );
  OAI211_X1 U21372 ( .C1(n18567), .C2(n18559), .A(n18259), .B(n18258), .ZN(
        P3_U2883) );
  NOR2_X1 U21373 ( .A1(n20932), .A2(n18260), .ZN(n18326) );
  NAND2_X1 U21374 ( .A1(n18326), .A2(n18668), .ZN(n18347) );
  INV_X1 U21375 ( .A(n18347), .ZN(n18340) );
  NOR2_X1 U21376 ( .A1(n18340), .A2(n18322), .ZN(n18304) );
  NOR2_X1 U21377 ( .A1(n18569), .A2(n18304), .ZN(n18277) );
  AOI22_X1 U21378 ( .A1(n18538), .A2(n18296), .B1(n18570), .B2(n18277), .ZN(
        n18264) );
  INV_X1 U21379 ( .A(n18441), .ZN(n18539) );
  INV_X1 U21380 ( .A(n18304), .ZN(n18261) );
  AOI22_X1 U21381 ( .A1(n18541), .A2(n18262), .B1(n18539), .B2(n18261), .ZN(
        n18278) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18278), .B1(
        n18340), .B2(n18576), .ZN(n18263) );
  OAI211_X1 U21383 ( .C1(n18545), .C2(n18617), .A(n18264), .B(n18263), .ZN(
        P3_U2884) );
  AOI22_X1 U21384 ( .A1(n18581), .A2(n18296), .B1(n18580), .B2(n18277), .ZN(
        n18266) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18278), .B1(
        n18340), .B2(n18582), .ZN(n18265) );
  OAI211_X1 U21386 ( .C1(n18586), .C2(n18617), .A(n18266), .B(n18265), .ZN(
        P3_U2885) );
  AOI22_X1 U21387 ( .A1(n18588), .A2(n18623), .B1(n18587), .B2(n18277), .ZN(
        n18268) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18278), .B1(
        n18589), .B2(n18296), .ZN(n18267) );
  OAI211_X1 U21389 ( .C1(n18347), .C2(n18592), .A(n18268), .B(n18267), .ZN(
        P3_U2886) );
  AOI22_X1 U21390 ( .A1(n18595), .A2(n18296), .B1(n18593), .B2(n18277), .ZN(
        n18270) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18278), .B1(
        n18594), .B2(n18623), .ZN(n18269) );
  OAI211_X1 U21392 ( .C1(n18347), .C2(n18598), .A(n18270), .B(n18269), .ZN(
        P3_U2887) );
  AOI22_X1 U21393 ( .A1(n18600), .A2(n18296), .B1(n18599), .B2(n18277), .ZN(
        n18272) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18278), .B1(
        n18601), .B2(n18623), .ZN(n18271) );
  OAI211_X1 U21395 ( .C1(n18347), .C2(n18604), .A(n18272), .B(n18271), .ZN(
        P3_U2888) );
  AOI22_X1 U21396 ( .A1(n18607), .A2(n18623), .B1(n18606), .B2(n18277), .ZN(
        n18274) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18278), .B1(
        n18605), .B2(n18296), .ZN(n18273) );
  OAI211_X1 U21398 ( .C1(n18347), .C2(n18610), .A(n18274), .B(n18273), .ZN(
        P3_U2889) );
  AOI22_X1 U21399 ( .A1(n18614), .A2(n18623), .B1(n18611), .B2(n18277), .ZN(
        n18276) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18278), .B1(
        n18613), .B2(n18296), .ZN(n18275) );
  OAI211_X1 U21401 ( .C1(n18347), .C2(n18618), .A(n18276), .B(n18275), .ZN(
        P3_U2890) );
  AOI22_X1 U21402 ( .A1(n18561), .A2(n18296), .B1(n18620), .B2(n18277), .ZN(
        n18280) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18278), .B1(
        n18340), .B2(n18624), .ZN(n18279) );
  OAI211_X1 U21404 ( .C1(n18567), .C2(n18617), .A(n18280), .B(n18279), .ZN(
        P3_U2891) );
  NAND2_X1 U21405 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18326), .ZN(
        n18370) );
  INV_X1 U21406 ( .A(n18370), .ZN(n18363) );
  INV_X1 U21407 ( .A(n18541), .ZN(n18443) );
  AOI21_X1 U21408 ( .B1(n20932), .B2(n18443), .A(n18486), .ZN(n18372) );
  OAI211_X1 U21409 ( .C1(n18789), .C2(n18363), .A(n18281), .B(n18372), .ZN(
        n18300) );
  INV_X1 U21410 ( .A(n18300), .ZN(n18285) );
  INV_X1 U21411 ( .A(n18326), .ZN(n18282) );
  NOR2_X1 U21412 ( .A1(n18569), .A2(n18282), .ZN(n18299) );
  AOI22_X1 U21413 ( .A1(n18571), .A2(n18296), .B1(n18570), .B2(n18299), .ZN(
        n18284) );
  AOI22_X1 U21414 ( .A1(n18363), .A2(n18576), .B1(n18322), .B2(n18538), .ZN(
        n18283) );
  OAI211_X1 U21415 ( .C1(n18285), .C2(n20872), .A(n18284), .B(n18283), .ZN(
        P3_U2892) );
  AOI22_X1 U21416 ( .A1(n18322), .A2(n18581), .B1(n18580), .B2(n18299), .ZN(
        n18287) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18300), .B1(
        n18363), .B2(n18582), .ZN(n18286) );
  OAI211_X1 U21418 ( .C1(n18586), .C2(n18303), .A(n18287), .B(n18286), .ZN(
        P3_U2893) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18300), .B1(
        n18587), .B2(n18299), .ZN(n18289) );
  AOI22_X1 U21420 ( .A1(n18322), .A2(n18589), .B1(n18588), .B2(n18296), .ZN(
        n18288) );
  OAI211_X1 U21421 ( .C1(n18370), .C2(n18592), .A(n18289), .B(n18288), .ZN(
        P3_U2894) );
  AOI22_X1 U21422 ( .A1(n18322), .A2(n18595), .B1(n18593), .B2(n18299), .ZN(
        n18291) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18300), .B1(
        n18594), .B2(n18296), .ZN(n18290) );
  OAI211_X1 U21424 ( .C1(n18370), .C2(n18598), .A(n18291), .B(n18290), .ZN(
        P3_U2895) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18300), .B1(
        n18599), .B2(n18299), .ZN(n18293) );
  AOI22_X1 U21426 ( .A1(n18322), .A2(n18600), .B1(n18601), .B2(n18296), .ZN(
        n18292) );
  OAI211_X1 U21427 ( .C1(n18370), .C2(n18604), .A(n18293), .B(n18292), .ZN(
        P3_U2896) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18300), .B1(
        n18606), .B2(n18299), .ZN(n18295) );
  AOI22_X1 U21429 ( .A1(n18322), .A2(n18605), .B1(n18607), .B2(n18296), .ZN(
        n18294) );
  OAI211_X1 U21430 ( .C1(n18370), .C2(n18610), .A(n18295), .B(n18294), .ZN(
        P3_U2897) );
  AOI22_X1 U21431 ( .A1(n18322), .A2(n18613), .B1(n18611), .B2(n18299), .ZN(
        n18298) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18300), .B1(
        n18614), .B2(n18296), .ZN(n18297) );
  OAI211_X1 U21433 ( .C1(n18370), .C2(n18618), .A(n18298), .B(n18297), .ZN(
        P3_U2898) );
  AOI22_X1 U21434 ( .A1(n18322), .A2(n18561), .B1(n18620), .B2(n18299), .ZN(
        n18302) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18300), .B1(
        n18363), .B2(n18624), .ZN(n18301) );
  OAI211_X1 U21436 ( .C1(n18567), .C2(n18303), .A(n18302), .B(n18301), .ZN(
        P3_U2899) );
  INV_X1 U21437 ( .A(n18373), .ZN(n18327) );
  NOR2_X2 U21438 ( .A1(n18670), .A2(n18327), .ZN(n18387) );
  INV_X1 U21439 ( .A(n18387), .ZN(n18394) );
  AOI21_X1 U21440 ( .B1(n18394), .B2(n18370), .A(n18569), .ZN(n18321) );
  AOI22_X1 U21441 ( .A1(n18322), .A2(n18571), .B1(n18570), .B2(n18321), .ZN(
        n18308) );
  AOI221_X1 U21442 ( .B1(n18304), .B2(n18370), .C1(n18443), .C2(n18370), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18306) );
  OAI21_X1 U21443 ( .B1(n18387), .B2(n18306), .A(n18305), .ZN(n18323) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18323), .B1(
        n18387), .B2(n18576), .ZN(n18307) );
  OAI211_X1 U21445 ( .C1(n18347), .C2(n18579), .A(n18308), .B(n18307), .ZN(
        P3_U2900) );
  AOI22_X1 U21446 ( .A1(n18322), .A2(n18518), .B1(n18321), .B2(n18580), .ZN(
        n18310) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18323), .B1(
        n18387), .B2(n18582), .ZN(n18309) );
  OAI211_X1 U21448 ( .C1(n18347), .C2(n18521), .A(n18310), .B(n18309), .ZN(
        P3_U2901) );
  AOI22_X1 U21449 ( .A1(n18340), .A2(n18589), .B1(n18321), .B2(n18587), .ZN(
        n18312) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18323), .B1(
        n18322), .B2(n18588), .ZN(n18311) );
  OAI211_X1 U21451 ( .C1(n18394), .C2(n18592), .A(n18312), .B(n18311), .ZN(
        P3_U2902) );
  AOI22_X1 U21452 ( .A1(n18340), .A2(n18595), .B1(n18321), .B2(n18593), .ZN(
        n18314) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18323), .B1(
        n18322), .B2(n18594), .ZN(n18313) );
  OAI211_X1 U21454 ( .C1(n18394), .C2(n18598), .A(n18314), .B(n18313), .ZN(
        P3_U2903) );
  AOI22_X1 U21455 ( .A1(n18340), .A2(n18600), .B1(n18321), .B2(n18599), .ZN(
        n18316) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18323), .B1(
        n18322), .B2(n18601), .ZN(n18315) );
  OAI211_X1 U21457 ( .C1(n18394), .C2(n18604), .A(n18316), .B(n18315), .ZN(
        P3_U2904) );
  AOI22_X1 U21458 ( .A1(n18340), .A2(n18605), .B1(n18321), .B2(n18606), .ZN(
        n18318) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18323), .B1(
        n18322), .B2(n18607), .ZN(n18317) );
  OAI211_X1 U21460 ( .C1(n18394), .C2(n18610), .A(n18318), .B(n18317), .ZN(
        P3_U2905) );
  AOI22_X1 U21461 ( .A1(n18340), .A2(n18613), .B1(n18321), .B2(n18611), .ZN(
        n18320) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18323), .B1(
        n18322), .B2(n18614), .ZN(n18319) );
  OAI211_X1 U21463 ( .C1(n18394), .C2(n18618), .A(n18320), .B(n18319), .ZN(
        P3_U2906) );
  AOI22_X1 U21464 ( .A1(n18322), .A2(n18622), .B1(n18321), .B2(n18620), .ZN(
        n18325) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18323), .B1(
        n18387), .B2(n18624), .ZN(n18324) );
  OAI211_X1 U21466 ( .C1(n18347), .C2(n18629), .A(n18325), .B(n18324), .ZN(
        P3_U2907) );
  NOR2_X1 U21467 ( .A1(n18327), .A2(n18511), .ZN(n18343) );
  AOI22_X1 U21468 ( .A1(n18340), .A2(n18571), .B1(n18570), .B2(n18343), .ZN(
        n18329) );
  AOI22_X1 U21469 ( .A1(n18575), .A2(n18326), .B1(n18373), .B2(n18513), .ZN(
        n18344) );
  NOR2_X2 U21470 ( .A1(n18327), .A2(n18419), .ZN(n18413) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18344), .B1(
        n18576), .B2(n18413), .ZN(n18328) );
  OAI211_X1 U21472 ( .C1(n18370), .C2(n18579), .A(n18329), .B(n18328), .ZN(
        P3_U2908) );
  AOI22_X1 U21473 ( .A1(n18363), .A2(n18581), .B1(n18580), .B2(n18343), .ZN(
        n18331) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18344), .B1(
        n18582), .B2(n18413), .ZN(n18330) );
  OAI211_X1 U21475 ( .C1(n18347), .C2(n18586), .A(n18331), .B(n18330), .ZN(
        P3_U2909) );
  INV_X1 U21476 ( .A(n18413), .ZN(n18401) );
  AOI22_X1 U21477 ( .A1(n18363), .A2(n18589), .B1(n18587), .B2(n18343), .ZN(
        n18333) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18344), .B1(
        n18340), .B2(n18588), .ZN(n18332) );
  OAI211_X1 U21479 ( .C1(n18592), .C2(n18401), .A(n18333), .B(n18332), .ZN(
        P3_U2910) );
  AOI22_X1 U21480 ( .A1(n18363), .A2(n18595), .B1(n18593), .B2(n18343), .ZN(
        n18335) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18344), .B1(
        n18340), .B2(n18594), .ZN(n18334) );
  OAI211_X1 U21482 ( .C1(n18598), .C2(n18401), .A(n18335), .B(n18334), .ZN(
        P3_U2911) );
  AOI22_X1 U21483 ( .A1(n18363), .A2(n18600), .B1(n18599), .B2(n18343), .ZN(
        n18337) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18344), .B1(
        n18340), .B2(n18601), .ZN(n18336) );
  OAI211_X1 U21485 ( .C1(n18604), .C2(n18401), .A(n18337), .B(n18336), .ZN(
        P3_U2912) );
  AOI22_X1 U21486 ( .A1(n18363), .A2(n18605), .B1(n18606), .B2(n18343), .ZN(
        n18339) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18344), .B1(
        n18340), .B2(n18607), .ZN(n18338) );
  OAI211_X1 U21488 ( .C1(n18610), .C2(n18401), .A(n18339), .B(n18338), .ZN(
        P3_U2913) );
  AOI22_X1 U21489 ( .A1(n18340), .A2(n18614), .B1(n18611), .B2(n18343), .ZN(
        n18342) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18344), .B1(
        n18363), .B2(n18613), .ZN(n18341) );
  OAI211_X1 U21491 ( .C1(n18618), .C2(n18401), .A(n18342), .B(n18341), .ZN(
        P3_U2914) );
  AOI22_X1 U21492 ( .A1(n18363), .A2(n18561), .B1(n18620), .B2(n18343), .ZN(
        n18346) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18344), .B1(
        n18624), .B2(n18413), .ZN(n18345) );
  OAI211_X1 U21494 ( .C1(n18347), .C2(n18567), .A(n18346), .B(n18345), .ZN(
        P3_U2915) );
  NOR2_X1 U21495 ( .A1(n18348), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18417) );
  INV_X1 U21496 ( .A(n18417), .ZN(n18374) );
  NOR2_X2 U21497 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18374), .ZN(
        n18433) );
  NOR2_X1 U21498 ( .A1(n18413), .A2(n18433), .ZN(n18349) );
  NOR2_X1 U21499 ( .A1(n18569), .A2(n18349), .ZN(n18366) );
  AOI22_X1 U21500 ( .A1(n18387), .A2(n18538), .B1(n18570), .B2(n18366), .ZN(
        n18352) );
  INV_X1 U21501 ( .A(n18349), .ZN(n18395) );
  NAND2_X1 U21502 ( .A1(n18394), .A2(n18370), .ZN(n18350) );
  OAI221_X1 U21503 ( .B1(n18395), .B2(n18541), .C1(n18395), .C2(n18350), .A(
        n18539), .ZN(n18367) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18367), .B1(
        n18576), .B2(n18433), .ZN(n18351) );
  OAI211_X1 U21505 ( .C1(n18370), .C2(n18545), .A(n18352), .B(n18351), .ZN(
        P3_U2916) );
  AOI22_X1 U21506 ( .A1(n18387), .A2(n18581), .B1(n18580), .B2(n18366), .ZN(
        n18354) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18367), .B1(
        n18582), .B2(n18433), .ZN(n18353) );
  OAI211_X1 U21508 ( .C1(n18370), .C2(n18586), .A(n18354), .B(n18353), .ZN(
        P3_U2917) );
  INV_X1 U21509 ( .A(n18433), .ZN(n18440) );
  AOI22_X1 U21510 ( .A1(n18363), .A2(n18588), .B1(n18587), .B2(n18366), .ZN(
        n18356) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18367), .B1(
        n18387), .B2(n18589), .ZN(n18355) );
  OAI211_X1 U21512 ( .C1(n18592), .C2(n18440), .A(n18356), .B(n18355), .ZN(
        P3_U2918) );
  AOI22_X1 U21513 ( .A1(n18363), .A2(n18594), .B1(n18593), .B2(n18366), .ZN(
        n18358) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18367), .B1(
        n18387), .B2(n18595), .ZN(n18357) );
  OAI211_X1 U21515 ( .C1(n18598), .C2(n18440), .A(n18358), .B(n18357), .ZN(
        P3_U2919) );
  AOI22_X1 U21516 ( .A1(n18363), .A2(n18601), .B1(n18599), .B2(n18366), .ZN(
        n18360) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18367), .B1(
        n18387), .B2(n18600), .ZN(n18359) );
  OAI211_X1 U21518 ( .C1(n18604), .C2(n18440), .A(n18360), .B(n18359), .ZN(
        P3_U2920) );
  AOI22_X1 U21519 ( .A1(n18363), .A2(n18607), .B1(n18606), .B2(n18366), .ZN(
        n18362) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18367), .B1(
        n18387), .B2(n18605), .ZN(n18361) );
  OAI211_X1 U21521 ( .C1(n18610), .C2(n18440), .A(n18362), .B(n18361), .ZN(
        P3_U2921) );
  AOI22_X1 U21522 ( .A1(n18387), .A2(n18613), .B1(n18611), .B2(n18366), .ZN(
        n18365) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18367), .B1(
        n18363), .B2(n18614), .ZN(n18364) );
  OAI211_X1 U21524 ( .C1(n18618), .C2(n18440), .A(n18365), .B(n18364), .ZN(
        P3_U2922) );
  AOI22_X1 U21525 ( .A1(n18387), .A2(n18561), .B1(n18620), .B2(n18366), .ZN(
        n18369) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18367), .B1(
        n18624), .B2(n18433), .ZN(n18368) );
  OAI211_X1 U21527 ( .C1(n18370), .C2(n18567), .A(n18369), .B(n18368), .ZN(
        P3_U2923) );
  NAND3_X1 U21528 ( .A1(n18373), .A2(n18372), .A3(n18371), .ZN(n18391) );
  NOR2_X1 U21529 ( .A1(n18569), .A2(n18374), .ZN(n18390) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18391), .B1(
        n18570), .B2(n18390), .ZN(n18376) );
  NOR2_X2 U21531 ( .A1(n18668), .A2(n18374), .ZN(n18460) );
  AOI22_X1 U21532 ( .A1(n18387), .A2(n18571), .B1(n18576), .B2(n18460), .ZN(
        n18375) );
  OAI211_X1 U21533 ( .C1(n18579), .C2(n18401), .A(n18376), .B(n18375), .ZN(
        P3_U2924) );
  AOI22_X1 U21534 ( .A1(n18387), .A2(n18518), .B1(n18580), .B2(n18390), .ZN(
        n18378) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18391), .B1(
        n18582), .B2(n18460), .ZN(n18377) );
  OAI211_X1 U21536 ( .C1(n18521), .C2(n18401), .A(n18378), .B(n18377), .ZN(
        P3_U2925) );
  INV_X1 U21537 ( .A(n18460), .ZN(n18424) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18391), .B1(
        n18587), .B2(n18390), .ZN(n18380) );
  AOI22_X1 U21539 ( .A1(n18387), .A2(n18588), .B1(n18589), .B2(n18413), .ZN(
        n18379) );
  OAI211_X1 U21540 ( .C1(n18592), .C2(n18424), .A(n18380), .B(n18379), .ZN(
        P3_U2926) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18391), .B1(
        n18593), .B2(n18390), .ZN(n18382) );
  AOI22_X1 U21542 ( .A1(n18387), .A2(n18594), .B1(n18595), .B2(n18413), .ZN(
        n18381) );
  OAI211_X1 U21543 ( .C1(n18598), .C2(n18424), .A(n18382), .B(n18381), .ZN(
        P3_U2927) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18391), .B1(
        n18599), .B2(n18390), .ZN(n18384) );
  AOI22_X1 U21545 ( .A1(n18387), .A2(n18601), .B1(n18600), .B2(n18413), .ZN(
        n18383) );
  OAI211_X1 U21546 ( .C1(n18604), .C2(n18424), .A(n18384), .B(n18383), .ZN(
        P3_U2928) );
  AOI22_X1 U21547 ( .A1(n18606), .A2(n18390), .B1(n18605), .B2(n18413), .ZN(
        n18386) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18391), .B1(
        n18387), .B2(n18607), .ZN(n18385) );
  OAI211_X1 U21549 ( .C1(n18610), .C2(n18424), .A(n18386), .B(n18385), .ZN(
        P3_U2929) );
  AOI22_X1 U21550 ( .A1(n18613), .A2(n18413), .B1(n18611), .B2(n18390), .ZN(
        n18389) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18391), .B1(
        n18387), .B2(n18614), .ZN(n18388) );
  OAI211_X1 U21552 ( .C1(n18618), .C2(n18424), .A(n18389), .B(n18388), .ZN(
        P3_U2930) );
  AOI22_X1 U21553 ( .A1(n18561), .A2(n18413), .B1(n18620), .B2(n18390), .ZN(
        n18393) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18391), .B1(
        n18624), .B2(n18460), .ZN(n18392) );
  OAI211_X1 U21555 ( .C1(n18394), .C2(n18567), .A(n18393), .B(n18392), .ZN(
        P3_U2931) );
  NOR2_X2 U21556 ( .A1(n18670), .A2(n18418), .ZN(n18482) );
  INV_X1 U21557 ( .A(n18482), .ZN(n18470) );
  NAND2_X1 U21558 ( .A1(n18424), .A2(n18470), .ZN(n18396) );
  INV_X1 U21559 ( .A(n18396), .ZN(n18442) );
  NOR2_X1 U21560 ( .A1(n18569), .A2(n18442), .ZN(n18412) );
  AOI22_X1 U21561 ( .A1(n18571), .A2(n18413), .B1(n18570), .B2(n18412), .ZN(
        n18398) );
  OAI221_X1 U21562 ( .B1(n18396), .B2(n18541), .C1(n18396), .C2(n18395), .A(
        n18539), .ZN(n18414) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18414), .B1(
        n18576), .B2(n18482), .ZN(n18397) );
  OAI211_X1 U21564 ( .C1(n18579), .C2(n18440), .A(n18398), .B(n18397), .ZN(
        P3_U2932) );
  AOI22_X1 U21565 ( .A1(n18581), .A2(n18433), .B1(n18580), .B2(n18412), .ZN(
        n18400) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18414), .B1(
        n18582), .B2(n18482), .ZN(n18399) );
  OAI211_X1 U21567 ( .C1(n18586), .C2(n18401), .A(n18400), .B(n18399), .ZN(
        P3_U2933) );
  AOI22_X1 U21568 ( .A1(n18587), .A2(n18412), .B1(n18589), .B2(n18433), .ZN(
        n18403) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18414), .B1(
        n18588), .B2(n18413), .ZN(n18402) );
  OAI211_X1 U21570 ( .C1(n18592), .C2(n18470), .A(n18403), .B(n18402), .ZN(
        P3_U2934) );
  AOI22_X1 U21571 ( .A1(n18595), .A2(n18433), .B1(n18593), .B2(n18412), .ZN(
        n18405) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18414), .B1(
        n18594), .B2(n18413), .ZN(n18404) );
  OAI211_X1 U21573 ( .C1(n18598), .C2(n18470), .A(n18405), .B(n18404), .ZN(
        P3_U2935) );
  AOI22_X1 U21574 ( .A1(n18600), .A2(n18433), .B1(n18599), .B2(n18412), .ZN(
        n18407) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18414), .B1(
        n18601), .B2(n18413), .ZN(n18406) );
  OAI211_X1 U21576 ( .C1(n18604), .C2(n18470), .A(n18407), .B(n18406), .ZN(
        P3_U2936) );
  AOI22_X1 U21577 ( .A1(n18607), .A2(n18413), .B1(n18606), .B2(n18412), .ZN(
        n18409) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18414), .B1(
        n18605), .B2(n18433), .ZN(n18408) );
  OAI211_X1 U21579 ( .C1(n18610), .C2(n18470), .A(n18409), .B(n18408), .ZN(
        P3_U2937) );
  AOI22_X1 U21580 ( .A1(n18614), .A2(n18413), .B1(n18611), .B2(n18412), .ZN(
        n18411) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18414), .B1(
        n18613), .B2(n18433), .ZN(n18410) );
  OAI211_X1 U21582 ( .C1(n18618), .C2(n18470), .A(n18411), .B(n18410), .ZN(
        P3_U2938) );
  AOI22_X1 U21583 ( .A1(n18622), .A2(n18413), .B1(n18620), .B2(n18412), .ZN(
        n18416) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18414), .B1(
        n18624), .B2(n18482), .ZN(n18415) );
  OAI211_X1 U21585 ( .C1(n18629), .C2(n18440), .A(n18416), .B(n18415), .ZN(
        P3_U2939) );
  NOR2_X1 U21586 ( .A1(n18511), .A2(n18418), .ZN(n18436) );
  AOI22_X1 U21587 ( .A1(n18538), .A2(n18460), .B1(n18570), .B2(n18436), .ZN(
        n18421) );
  AOI22_X1 U21588 ( .A1(n18575), .A2(n18417), .B1(n18513), .B2(n18464), .ZN(
        n18437) );
  NOR2_X2 U21589 ( .A1(n18419), .A2(n18418), .ZN(n18507) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18437), .B1(
        n18576), .B2(n18507), .ZN(n18420) );
  OAI211_X1 U21591 ( .C1(n18545), .C2(n18440), .A(n18421), .B(n18420), .ZN(
        P3_U2940) );
  AOI22_X1 U21592 ( .A1(n18580), .A2(n18436), .B1(n18518), .B2(n18433), .ZN(
        n18423) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18437), .B1(
        n18582), .B2(n18507), .ZN(n18422) );
  OAI211_X1 U21594 ( .C1(n18521), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2941) );
  INV_X1 U21595 ( .A(n18507), .ZN(n18495) );
  AOI22_X1 U21596 ( .A1(n18587), .A2(n18436), .B1(n18589), .B2(n18460), .ZN(
        n18426) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18437), .B1(
        n18588), .B2(n18433), .ZN(n18425) );
  OAI211_X1 U21598 ( .C1(n18592), .C2(n18495), .A(n18426), .B(n18425), .ZN(
        P3_U2942) );
  AOI22_X1 U21599 ( .A1(n18594), .A2(n18433), .B1(n18593), .B2(n18436), .ZN(
        n18428) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18437), .B1(
        n18595), .B2(n18460), .ZN(n18427) );
  OAI211_X1 U21601 ( .C1(n18598), .C2(n18495), .A(n18428), .B(n18427), .ZN(
        P3_U2943) );
  AOI22_X1 U21602 ( .A1(n18601), .A2(n18433), .B1(n18599), .B2(n18436), .ZN(
        n18430) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18437), .B1(
        n18600), .B2(n18460), .ZN(n18429) );
  OAI211_X1 U21604 ( .C1(n18604), .C2(n18495), .A(n18430), .B(n18429), .ZN(
        P3_U2944) );
  AOI22_X1 U21605 ( .A1(n18607), .A2(n18433), .B1(n18606), .B2(n18436), .ZN(
        n18432) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18437), .B1(
        n18605), .B2(n18460), .ZN(n18431) );
  OAI211_X1 U21607 ( .C1(n18610), .C2(n18495), .A(n18432), .B(n18431), .ZN(
        P3_U2945) );
  AOI22_X1 U21608 ( .A1(n18614), .A2(n18433), .B1(n18611), .B2(n18436), .ZN(
        n18435) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18437), .B1(
        n18613), .B2(n18460), .ZN(n18434) );
  OAI211_X1 U21610 ( .C1(n18618), .C2(n18495), .A(n18435), .B(n18434), .ZN(
        P3_U2946) );
  AOI22_X1 U21611 ( .A1(n18561), .A2(n18460), .B1(n18620), .B2(n18436), .ZN(
        n18439) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18437), .B1(
        n18624), .B2(n18507), .ZN(n18438) );
  OAI211_X1 U21613 ( .C1(n18567), .C2(n18440), .A(n18439), .B(n18438), .ZN(
        P3_U2947) );
  NAND2_X1 U21614 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18464), .ZN(
        n18465) );
  NOR2_X2 U21615 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18465), .ZN(
        n18530) );
  NOR2_X1 U21616 ( .A1(n18507), .A2(n18530), .ZN(n18489) );
  NOR2_X1 U21617 ( .A1(n18569), .A2(n18489), .ZN(n18459) );
  AOI22_X1 U21618 ( .A1(n18571), .A2(n18460), .B1(n18570), .B2(n18459), .ZN(
        n18446) );
  AOI221_X1 U21619 ( .B1(n18489), .B2(n18443), .C1(n18489), .C2(n18442), .A(
        n18441), .ZN(n18444) );
  INV_X1 U21620 ( .A(n18444), .ZN(n18461) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18461), .B1(
        n18576), .B2(n18530), .ZN(n18445) );
  OAI211_X1 U21622 ( .C1(n18579), .C2(n18470), .A(n18446), .B(n18445), .ZN(
        P3_U2948) );
  AOI22_X1 U21623 ( .A1(n18580), .A2(n18459), .B1(n18518), .B2(n18460), .ZN(
        n18448) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18461), .B1(
        n18582), .B2(n18530), .ZN(n18447) );
  OAI211_X1 U21625 ( .C1(n18521), .C2(n18470), .A(n18448), .B(n18447), .ZN(
        P3_U2949) );
  INV_X1 U21626 ( .A(n18530), .ZN(n18536) );
  AOI22_X1 U21627 ( .A1(n18587), .A2(n18459), .B1(n18589), .B2(n18482), .ZN(
        n18450) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18461), .B1(
        n18588), .B2(n18460), .ZN(n18449) );
  OAI211_X1 U21629 ( .C1(n18592), .C2(n18536), .A(n18450), .B(n18449), .ZN(
        P3_U2950) );
  AOI22_X1 U21630 ( .A1(n18594), .A2(n18460), .B1(n18593), .B2(n18459), .ZN(
        n18452) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18461), .B1(
        n18595), .B2(n18482), .ZN(n18451) );
  OAI211_X1 U21632 ( .C1(n18598), .C2(n18536), .A(n18452), .B(n18451), .ZN(
        P3_U2951) );
  AOI22_X1 U21633 ( .A1(n18601), .A2(n18460), .B1(n18599), .B2(n18459), .ZN(
        n18454) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18461), .B1(
        n18600), .B2(n18482), .ZN(n18453) );
  OAI211_X1 U21635 ( .C1(n18604), .C2(n18536), .A(n18454), .B(n18453), .ZN(
        P3_U2952) );
  AOI22_X1 U21636 ( .A1(n18606), .A2(n18459), .B1(n18605), .B2(n18482), .ZN(
        n18456) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18461), .B1(
        n18607), .B2(n18460), .ZN(n18455) );
  OAI211_X1 U21638 ( .C1(n18610), .C2(n18536), .A(n18456), .B(n18455), .ZN(
        P3_U2953) );
  AOI22_X1 U21639 ( .A1(n18613), .A2(n18482), .B1(n18611), .B2(n18459), .ZN(
        n18458) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18461), .B1(
        n18614), .B2(n18460), .ZN(n18457) );
  OAI211_X1 U21641 ( .C1(n18618), .C2(n18536), .A(n18458), .B(n18457), .ZN(
        P3_U2954) );
  AOI22_X1 U21642 ( .A1(n18622), .A2(n18460), .B1(n18620), .B2(n18459), .ZN(
        n18463) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18461), .B1(
        n18624), .B2(n18530), .ZN(n18462) );
  OAI211_X1 U21644 ( .C1(n18629), .C2(n18470), .A(n18463), .B(n18462), .ZN(
        P3_U2955) );
  NOR2_X1 U21645 ( .A1(n18569), .A2(n18465), .ZN(n18481) );
  AOI22_X1 U21646 ( .A1(n18538), .A2(n18507), .B1(n18570), .B2(n18481), .ZN(
        n18467) );
  INV_X1 U21647 ( .A(n18465), .ZN(n18515) );
  AOI22_X1 U21648 ( .A1(n18575), .A2(n18464), .B1(n18572), .B2(n18515), .ZN(
        n18483) );
  NOR2_X2 U21649 ( .A1(n18668), .A2(n18465), .ZN(n18556) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18483), .B1(
        n18576), .B2(n18556), .ZN(n18466) );
  OAI211_X1 U21651 ( .C1(n18545), .C2(n18470), .A(n18467), .B(n18466), .ZN(
        P3_U2956) );
  AOI22_X1 U21652 ( .A1(n18581), .A2(n18507), .B1(n18580), .B2(n18481), .ZN(
        n18469) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18483), .B1(
        n18582), .B2(n18556), .ZN(n18468) );
  OAI211_X1 U21654 ( .C1(n18586), .C2(n18470), .A(n18469), .B(n18468), .ZN(
        P3_U2957) );
  INV_X1 U21655 ( .A(n18556), .ZN(n18566) );
  AOI22_X1 U21656 ( .A1(n18587), .A2(n18481), .B1(n18589), .B2(n18507), .ZN(
        n18472) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18483), .B1(
        n18588), .B2(n18482), .ZN(n18471) );
  OAI211_X1 U21658 ( .C1(n18592), .C2(n18566), .A(n18472), .B(n18471), .ZN(
        P3_U2958) );
  AOI22_X1 U21659 ( .A1(n18595), .A2(n18507), .B1(n18593), .B2(n18481), .ZN(
        n18474) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18483), .B1(
        n18594), .B2(n18482), .ZN(n18473) );
  OAI211_X1 U21661 ( .C1(n18598), .C2(n18566), .A(n18474), .B(n18473), .ZN(
        P3_U2959) );
  AOI22_X1 U21662 ( .A1(n18600), .A2(n18507), .B1(n18599), .B2(n18481), .ZN(
        n18476) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18483), .B1(
        n18601), .B2(n18482), .ZN(n18475) );
  OAI211_X1 U21664 ( .C1(n18604), .C2(n18566), .A(n18476), .B(n18475), .ZN(
        P3_U2960) );
  AOI22_X1 U21665 ( .A1(n18606), .A2(n18481), .B1(n18605), .B2(n18507), .ZN(
        n18478) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18483), .B1(
        n18607), .B2(n18482), .ZN(n18477) );
  OAI211_X1 U21667 ( .C1(n18610), .C2(n18566), .A(n18478), .B(n18477), .ZN(
        P3_U2961) );
  AOI22_X1 U21668 ( .A1(n18614), .A2(n18482), .B1(n18611), .B2(n18481), .ZN(
        n18480) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18483), .B1(
        n18613), .B2(n18507), .ZN(n18479) );
  OAI211_X1 U21670 ( .C1(n18618), .C2(n18566), .A(n18480), .B(n18479), .ZN(
        P3_U2962) );
  AOI22_X1 U21671 ( .A1(n18622), .A2(n18482), .B1(n18620), .B2(n18481), .ZN(
        n18485) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18483), .B1(
        n18624), .B2(n18556), .ZN(n18484) );
  OAI211_X1 U21673 ( .C1(n18629), .C2(n18495), .A(n18485), .B(n18484), .ZN(
        P3_U2963) );
  NOR2_X2 U21674 ( .A1(n18670), .A2(n18512), .ZN(n18621) );
  INV_X1 U21675 ( .A(n18621), .ZN(n18585) );
  NAND2_X1 U21676 ( .A1(n18566), .A2(n18585), .ZN(n18540) );
  INV_X1 U21677 ( .A(n18540), .ZN(n18487) );
  NOR2_X1 U21678 ( .A1(n18569), .A2(n18487), .ZN(n18506) );
  AOI22_X1 U21679 ( .A1(n18571), .A2(n18507), .B1(n18570), .B2(n18506), .ZN(
        n18492) );
  OAI22_X1 U21680 ( .A1(n18489), .A2(n18488), .B1(n18487), .B2(n18486), .ZN(
        n18490) );
  OAI21_X1 U21681 ( .B1(n18621), .B2(n18789), .A(n18490), .ZN(n18508) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18508), .B1(
        n18576), .B2(n18621), .ZN(n18491) );
  OAI211_X1 U21683 ( .C1(n18579), .C2(n18536), .A(n18492), .B(n18491), .ZN(
        P3_U2964) );
  AOI22_X1 U21684 ( .A1(n18581), .A2(n18530), .B1(n18580), .B2(n18506), .ZN(
        n18494) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18508), .B1(
        n18582), .B2(n18621), .ZN(n18493) );
  OAI211_X1 U21686 ( .C1(n18586), .C2(n18495), .A(n18494), .B(n18493), .ZN(
        P3_U2965) );
  AOI22_X1 U21687 ( .A1(n18588), .A2(n18507), .B1(n18587), .B2(n18506), .ZN(
        n18497) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18508), .B1(
        n18589), .B2(n18530), .ZN(n18496) );
  OAI211_X1 U21689 ( .C1(n18592), .C2(n18585), .A(n18497), .B(n18496), .ZN(
        P3_U2966) );
  AOI22_X1 U21690 ( .A1(n18595), .A2(n18530), .B1(n18593), .B2(n18506), .ZN(
        n18499) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18508), .B1(
        n18594), .B2(n18507), .ZN(n18498) );
  OAI211_X1 U21692 ( .C1(n18598), .C2(n18585), .A(n18499), .B(n18498), .ZN(
        P3_U2967) );
  AOI22_X1 U21693 ( .A1(n18600), .A2(n18530), .B1(n18599), .B2(n18506), .ZN(
        n18501) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18508), .B1(
        n18601), .B2(n18507), .ZN(n18500) );
  OAI211_X1 U21695 ( .C1(n18604), .C2(n18585), .A(n18501), .B(n18500), .ZN(
        P3_U2968) );
  AOI22_X1 U21696 ( .A1(n18607), .A2(n18507), .B1(n18606), .B2(n18506), .ZN(
        n18503) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18508), .B1(
        n18605), .B2(n18530), .ZN(n18502) );
  OAI211_X1 U21698 ( .C1(n18610), .C2(n18585), .A(n18503), .B(n18502), .ZN(
        P3_U2969) );
  AOI22_X1 U21699 ( .A1(n18614), .A2(n18507), .B1(n18611), .B2(n18506), .ZN(
        n18505) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18508), .B1(
        n18613), .B2(n18530), .ZN(n18504) );
  OAI211_X1 U21701 ( .C1(n18618), .C2(n18585), .A(n18505), .B(n18504), .ZN(
        P3_U2970) );
  AOI22_X1 U21702 ( .A1(n18622), .A2(n18507), .B1(n18620), .B2(n18506), .ZN(
        n18510) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18508), .B1(
        n18624), .B2(n18621), .ZN(n18509) );
  OAI211_X1 U21704 ( .C1(n18629), .C2(n18536), .A(n18510), .B(n18509), .ZN(
        P3_U2971) );
  NOR2_X1 U21705 ( .A1(n18512), .A2(n18511), .ZN(n18574) );
  AOI22_X1 U21706 ( .A1(n18538), .A2(n18556), .B1(n18570), .B2(n18574), .ZN(
        n18517) );
  INV_X1 U21707 ( .A(n18512), .ZN(n18514) );
  AOI22_X1 U21708 ( .A1(n18575), .A2(n18515), .B1(n18514), .B2(n18513), .ZN(
        n18533) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18533), .B1(
        n18576), .B2(n18612), .ZN(n18516) );
  OAI211_X1 U21710 ( .C1(n18545), .C2(n18536), .A(n18517), .B(n18516), .ZN(
        P3_U2972) );
  AOI22_X1 U21711 ( .A1(n18580), .A2(n18574), .B1(n18518), .B2(n18530), .ZN(
        n18520) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18533), .B1(
        n18582), .B2(n18612), .ZN(n18519) );
  OAI211_X1 U21713 ( .C1(n18521), .C2(n18566), .A(n18520), .B(n18519), .ZN(
        P3_U2973) );
  AOI22_X1 U21714 ( .A1(n18587), .A2(n18574), .B1(n18589), .B2(n18556), .ZN(
        n18523) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18533), .B1(
        n18588), .B2(n18530), .ZN(n18522) );
  OAI211_X1 U21716 ( .C1(n18592), .C2(n18628), .A(n18523), .B(n18522), .ZN(
        P3_U2974) );
  AOI22_X1 U21717 ( .A1(n18595), .A2(n18556), .B1(n18593), .B2(n18574), .ZN(
        n18525) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18533), .B1(
        n18594), .B2(n18530), .ZN(n18524) );
  OAI211_X1 U21719 ( .C1(n18598), .C2(n18628), .A(n18525), .B(n18524), .ZN(
        P3_U2975) );
  AOI22_X1 U21720 ( .A1(n18600), .A2(n18556), .B1(n18599), .B2(n18574), .ZN(
        n18527) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18533), .B1(
        n18601), .B2(n18530), .ZN(n18526) );
  OAI211_X1 U21722 ( .C1(n18604), .C2(n18628), .A(n18527), .B(n18526), .ZN(
        P3_U2976) );
  AOI22_X1 U21723 ( .A1(n18606), .A2(n18574), .B1(n18605), .B2(n18556), .ZN(
        n18529) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18533), .B1(
        n18607), .B2(n18530), .ZN(n18528) );
  OAI211_X1 U21725 ( .C1(n18610), .C2(n18628), .A(n18529), .B(n18528), .ZN(
        P3_U2977) );
  AOI22_X1 U21726 ( .A1(n18614), .A2(n18530), .B1(n18611), .B2(n18574), .ZN(
        n18532) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18533), .B1(
        n18613), .B2(n18556), .ZN(n18531) );
  OAI211_X1 U21728 ( .C1(n18618), .C2(n18628), .A(n18532), .B(n18531), .ZN(
        P3_U2978) );
  AOI22_X1 U21729 ( .A1(n18561), .A2(n18556), .B1(n18620), .B2(n18574), .ZN(
        n18535) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18533), .B1(
        n18624), .B2(n18612), .ZN(n18534) );
  OAI211_X1 U21731 ( .C1(n18567), .C2(n18536), .A(n18535), .B(n18534), .ZN(
        P3_U2979) );
  INV_X1 U21732 ( .A(n18542), .ZN(n18537) );
  NOR2_X1 U21733 ( .A1(n18569), .A2(n18537), .ZN(n18560) );
  AOI22_X1 U21734 ( .A1(n18538), .A2(n18621), .B1(n18570), .B2(n18560), .ZN(
        n18544) );
  OAI221_X1 U21735 ( .B1(n18542), .B2(n18541), .C1(n18542), .C2(n18540), .A(
        n18539), .ZN(n18563) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18563), .B1(
        n18576), .B2(n18562), .ZN(n18543) );
  OAI211_X1 U21737 ( .C1(n18545), .C2(n18566), .A(n18544), .B(n18543), .ZN(
        P3_U2980) );
  AOI22_X1 U21738 ( .A1(n18581), .A2(n18621), .B1(n18580), .B2(n18560), .ZN(
        n18547) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18563), .B1(
        n18582), .B2(n18562), .ZN(n18546) );
  OAI211_X1 U21740 ( .C1(n18586), .C2(n18566), .A(n18547), .B(n18546), .ZN(
        P3_U2981) );
  AOI22_X1 U21741 ( .A1(n18587), .A2(n18560), .B1(n18589), .B2(n18621), .ZN(
        n18549) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18563), .B1(
        n18588), .B2(n18556), .ZN(n18548) );
  OAI211_X1 U21743 ( .C1(n18592), .C2(n18559), .A(n18549), .B(n18548), .ZN(
        P3_U2982) );
  AOI22_X1 U21744 ( .A1(n18594), .A2(n18556), .B1(n18593), .B2(n18560), .ZN(
        n18551) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18563), .B1(
        n18595), .B2(n18621), .ZN(n18550) );
  OAI211_X1 U21746 ( .C1(n18598), .C2(n18559), .A(n18551), .B(n18550), .ZN(
        P3_U2983) );
  AOI22_X1 U21747 ( .A1(n18601), .A2(n18556), .B1(n18599), .B2(n18560), .ZN(
        n18553) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18563), .B1(
        n18600), .B2(n18621), .ZN(n18552) );
  OAI211_X1 U21749 ( .C1(n18604), .C2(n18559), .A(n18553), .B(n18552), .ZN(
        P3_U2984) );
  AOI22_X1 U21750 ( .A1(n18607), .A2(n18556), .B1(n18606), .B2(n18560), .ZN(
        n18555) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18563), .B1(
        n18605), .B2(n18621), .ZN(n18554) );
  OAI211_X1 U21752 ( .C1(n18610), .C2(n18559), .A(n18555), .B(n18554), .ZN(
        P3_U2985) );
  AOI22_X1 U21753 ( .A1(n18614), .A2(n18556), .B1(n18611), .B2(n18560), .ZN(
        n18558) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18563), .B1(
        n18613), .B2(n18621), .ZN(n18557) );
  OAI211_X1 U21755 ( .C1(n18618), .C2(n18559), .A(n18558), .B(n18557), .ZN(
        P3_U2986) );
  AOI22_X1 U21756 ( .A1(n18561), .A2(n18621), .B1(n18620), .B2(n18560), .ZN(
        n18565) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18563), .B1(
        n18624), .B2(n18562), .ZN(n18564) );
  OAI211_X1 U21758 ( .C1(n18567), .C2(n18566), .A(n18565), .B(n18564), .ZN(
        P3_U2987) );
  INV_X1 U21759 ( .A(n18573), .ZN(n18568) );
  NOR2_X1 U21760 ( .A1(n18569), .A2(n18568), .ZN(n18619) );
  AOI22_X1 U21761 ( .A1(n18571), .A2(n18621), .B1(n18570), .B2(n18619), .ZN(
        n18578) );
  AOI22_X1 U21762 ( .A1(n18575), .A2(n18574), .B1(n18573), .B2(n18572), .ZN(
        n18625) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18625), .B1(
        n18576), .B2(n18623), .ZN(n18577) );
  OAI211_X1 U21764 ( .C1(n18579), .C2(n18628), .A(n18578), .B(n18577), .ZN(
        P3_U2988) );
  AOI22_X1 U21765 ( .A1(n18581), .A2(n18612), .B1(n18580), .B2(n18619), .ZN(
        n18584) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18625), .B1(
        n18582), .B2(n18623), .ZN(n18583) );
  OAI211_X1 U21767 ( .C1(n18586), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2989) );
  AOI22_X1 U21768 ( .A1(n18588), .A2(n18621), .B1(n18587), .B2(n18619), .ZN(
        n18591) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18625), .B1(
        n18589), .B2(n18612), .ZN(n18590) );
  OAI211_X1 U21770 ( .C1(n18592), .C2(n18617), .A(n18591), .B(n18590), .ZN(
        P3_U2990) );
  AOI22_X1 U21771 ( .A1(n18594), .A2(n18621), .B1(n18593), .B2(n18619), .ZN(
        n18597) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18625), .B1(
        n18595), .B2(n18612), .ZN(n18596) );
  OAI211_X1 U21773 ( .C1(n18598), .C2(n18617), .A(n18597), .B(n18596), .ZN(
        P3_U2991) );
  AOI22_X1 U21774 ( .A1(n18600), .A2(n18612), .B1(n18599), .B2(n18619), .ZN(
        n18603) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18625), .B1(
        n18601), .B2(n18621), .ZN(n18602) );
  OAI211_X1 U21776 ( .C1(n18604), .C2(n18617), .A(n18603), .B(n18602), .ZN(
        P3_U2992) );
  AOI22_X1 U21777 ( .A1(n18606), .A2(n18619), .B1(n18605), .B2(n18612), .ZN(
        n18609) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18625), .B1(
        n18607), .B2(n18621), .ZN(n18608) );
  OAI211_X1 U21779 ( .C1(n18610), .C2(n18617), .A(n18609), .B(n18608), .ZN(
        P3_U2993) );
  AOI22_X1 U21780 ( .A1(n18613), .A2(n18612), .B1(n18611), .B2(n18619), .ZN(
        n18616) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18625), .B1(
        n18614), .B2(n18621), .ZN(n18615) );
  OAI211_X1 U21782 ( .C1(n18618), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        P3_U2994) );
  AOI22_X1 U21783 ( .A1(n18622), .A2(n18621), .B1(n18620), .B2(n18619), .ZN(
        n18627) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18625), .B1(
        n18624), .B2(n18623), .ZN(n18626) );
  OAI211_X1 U21785 ( .C1(n18629), .C2(n18628), .A(n18627), .B(n18626), .ZN(
        P3_U2995) );
  NOR2_X1 U21786 ( .A1(n18661), .A2(n18630), .ZN(n18633) );
  OAI222_X1 U21787 ( .A1(n18636), .A2(n18635), .B1(n18634), .B2(n18633), .C1(
        n18632), .C2(n18631), .ZN(n18832) );
  OAI21_X1 U21788 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18637), .ZN(n18638) );
  OAI211_X1 U21789 ( .C1(n18640), .C2(n18662), .A(n18639), .B(n18638), .ZN(
        n18683) );
  INV_X1 U21790 ( .A(n18641), .ZN(n18653) );
  AOI21_X1 U21791 ( .B1(n18663), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18642), .ZN(n18666) );
  OAI22_X1 U21792 ( .A1(n18644), .A2(n18653), .B1(n18643), .B2(n18666), .ZN(
        n18645) );
  AND2_X1 U21793 ( .A1(n20947), .A2(n18645), .ZN(n18795) );
  AOI22_X1 U21794 ( .A1(n18648), .A2(n18647), .B1(n9801), .B2(n18646), .ZN(
        n18652) );
  NAND2_X1 U21795 ( .A1(n18649), .A2(n18652), .ZN(n18656) );
  AND2_X1 U21796 ( .A1(n18650), .A2(n9801), .ZN(n18651) );
  AOI21_X1 U21797 ( .B1(n18652), .B2(n18651), .A(n18658), .ZN(n18654) );
  AOI211_X1 U21798 ( .C1(n18821), .C2(n18656), .A(n18654), .B(n18653), .ZN(
        n18791) );
  AOI21_X1 U21799 ( .B1(n18791), .B2(n18662), .A(n20947), .ZN(n18655) );
  AOI21_X1 U21800 ( .B1(n18662), .B2(n18795), .A(n18655), .ZN(n18681) );
  AND3_X1 U21801 ( .A1(n18657), .A2(n18656), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18660) );
  AOI211_X1 U21802 ( .C1(n12634), .C2(n18807), .A(n18666), .B(n18658), .ZN(
        n18659) );
  AOI211_X1 U21803 ( .C1(n18661), .C2(n18801), .A(n18660), .B(n18659), .ZN(
        n18804) );
  AOI22_X1 U21804 ( .A1(n18672), .A2(n18807), .B1(n18804), .B2(n18662), .ZN(
        n18676) );
  NOR2_X1 U21805 ( .A1(n18664), .A2(n18663), .ZN(n18667) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18665), .B1(
        n18667), .B2(n18821), .ZN(n18816) );
  OAI22_X1 U21807 ( .A1(n18667), .A2(n18808), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18666), .ZN(n18813) );
  OR3_X1 U21808 ( .A1(n18816), .A2(n20932), .A3(n18668), .ZN(n18669) );
  AOI22_X1 U21809 ( .A1(n18816), .A2(n20932), .B1(n18813), .B2(n18669), .ZN(
        n18671) );
  OAI21_X1 U21810 ( .B1(n18672), .B2(n18671), .A(n18670), .ZN(n18675) );
  AND2_X1 U21811 ( .A1(n18676), .A2(n18675), .ZN(n18673) );
  OAI221_X1 U21812 ( .B1(n18676), .B2(n18675), .C1(n18674), .C2(n18673), .A(
        n18678), .ZN(n18680) );
  AOI21_X1 U21813 ( .B1(n18678), .B2(n18677), .A(n18676), .ZN(n18679) );
  AOI222_X1 U21814 ( .A1(n18681), .A2(n18680), .B1(n18681), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18680), .C2(n18679), .ZN(
        n18682) );
  NOR4_X1 U21815 ( .A1(n18684), .A2(n18832), .A3(n18683), .A4(n18682), .ZN(
        n18693) );
  NAND2_X1 U21816 ( .A1(n18837), .A2(n18845), .ZN(n18700) );
  AOI221_X1 U21817 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18700), 
        .C1(n18685), .C2(n18700), .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18691) );
  NOR2_X1 U21818 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18844), .ZN(n18695) );
  OAI211_X1 U21819 ( .C1(n18687), .C2(n18686), .A(n18699), .B(n18693), .ZN(
        n18696) );
  NAND2_X1 U21820 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18696), .ZN(n18787) );
  NOR4_X1 U21821 ( .A1(n18689), .A2(n18695), .A3(n18688), .A4(n18787), .ZN(
        n18690) );
  OAI22_X1 U21822 ( .A1(n18693), .A2(n18692), .B1(n18691), .B2(n18690), .ZN(
        P3_U2996) );
  AOI21_X1 U21823 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18695), .A(n18694), 
        .ZN(n18702) );
  INV_X1 U21824 ( .A(n18695), .ZN(n18697) );
  OAI211_X1 U21825 ( .C1(n18699), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        n18701) );
  OAI211_X1 U21826 ( .C1(n18702), .C2(n18800), .A(n18701), .B(n18700), .ZN(
        P3_U2997) );
  AND3_X1 U21827 ( .A1(n18702), .A2(n18839), .A3(n18788), .ZN(P3_U2998) );
  AND2_X1 U21828 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18783), .ZN(
        P3_U2999) );
  AND2_X1 U21829 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18783), .ZN(
        P3_U3000) );
  AND2_X1 U21830 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18783), .ZN(
        P3_U3001) );
  INV_X1 U21831 ( .A(P3_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20781) );
  NOR2_X1 U21832 ( .A1(n20781), .A2(n18786), .ZN(P3_U3002) );
  AND2_X1 U21833 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18783), .ZN(
        P3_U3003) );
  AND2_X1 U21834 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18783), .ZN(
        P3_U3004) );
  AND2_X1 U21835 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18783), .ZN(
        P3_U3005) );
  AND2_X1 U21836 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18783), .ZN(
        P3_U3006) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18783), .ZN(
        P3_U3007) );
  INV_X1 U21838 ( .A(P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20911) );
  NOR2_X1 U21839 ( .A1(n20911), .A2(n18786), .ZN(P3_U3008) );
  AND2_X1 U21840 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18703), .ZN(
        P3_U3009) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18703), .ZN(
        P3_U3010) );
  INV_X1 U21842 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20935) );
  NOR2_X1 U21843 ( .A1(n20935), .A2(n18786), .ZN(P3_U3011) );
  AND2_X1 U21844 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18703), .ZN(
        P3_U3012) );
  AND2_X1 U21845 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18703), .ZN(
        P3_U3013) );
  AND2_X1 U21846 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18703), .ZN(
        P3_U3014) );
  AND2_X1 U21847 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18783), .ZN(
        P3_U3015) );
  INV_X1 U21848 ( .A(P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20948) );
  NOR2_X1 U21849 ( .A1(n20948), .A2(n18786), .ZN(P3_U3016) );
  AND2_X1 U21850 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18783), .ZN(
        P3_U3017) );
  INV_X1 U21851 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20910) );
  NOR2_X1 U21852 ( .A1(n20910), .A2(n18786), .ZN(P3_U3018) );
  AND2_X1 U21853 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18783), .ZN(
        P3_U3019) );
  AND2_X1 U21854 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18783), .ZN(
        P3_U3020) );
  AND2_X1 U21855 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18783), .ZN(P3_U3021) );
  AND2_X1 U21856 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18783), .ZN(P3_U3022) );
  AND2_X1 U21857 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18783), .ZN(P3_U3023) );
  AND2_X1 U21858 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18783), .ZN(P3_U3024) );
  AND2_X1 U21859 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18783), .ZN(P3_U3025) );
  AND2_X1 U21860 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18783), .ZN(P3_U3026) );
  AND2_X1 U21861 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18783), .ZN(P3_U3027) );
  AND2_X1 U21862 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18783), .ZN(P3_U3028) );
  NAND2_X1 U21863 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n18710) );
  NOR2_X1 U21864 ( .A1(n18721), .A2(n20594), .ZN(n18717) );
  INV_X1 U21865 ( .A(n18717), .ZN(n18704) );
  AND3_X1 U21866 ( .A1(n18710), .A2(n18704), .A3(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18707) );
  NAND2_X1 U21867 ( .A1(n18837), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18715) );
  INV_X1 U21868 ( .A(n18715), .ZN(n18713) );
  OAI21_X1 U21869 ( .B1(n18713), .B2(n18719), .A(n18721), .ZN(n18706) );
  NAND3_X1 U21870 ( .A1(NA), .A2(n18719), .A3(n18705), .ZN(n18714) );
  OAI211_X1 U21871 ( .C1(n18848), .C2(n18707), .A(n18706), .B(n18714), .ZN(
        P3_U3029) );
  OAI21_X1 U21872 ( .B1(n18708), .B2(n20594), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18709) );
  OAI21_X1 U21873 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n18710), .A(n18709), 
        .ZN(n18711) );
  AOI22_X1 U21874 ( .A1(n18837), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18711), .ZN(n18712) );
  NAND2_X1 U21875 ( .A1(n18712), .A2(n18833), .ZN(P3_U3030) );
  AOI21_X1 U21876 ( .B1(n18719), .B2(n18714), .A(n18713), .ZN(n18720) );
  OAI22_X1 U21877 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18715), .ZN(n18716) );
  OAI22_X1 U21878 ( .A1(n18717), .A2(n18716), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18718) );
  OAI22_X1 U21879 ( .A1(n18720), .A2(n18721), .B1(n18719), .B2(n18718), .ZN(
        P3_U3031) );
  OAI222_X1 U21880 ( .A1(n20926), .A2(n18776), .B1(n18722), .B2(n18848), .C1(
        n18723), .C2(n18772), .ZN(P3_U3032) );
  OAI222_X1 U21881 ( .A1(n18772), .A2(n18725), .B1(n18724), .B2(n18848), .C1(
        n18723), .C2(n18776), .ZN(P3_U3033) );
  OAI222_X1 U21882 ( .A1(n18772), .A2(n18727), .B1(n18726), .B2(n18848), .C1(
        n18725), .C2(n18776), .ZN(P3_U3034) );
  OAI222_X1 U21883 ( .A1(n18772), .A2(n20797), .B1(n18728), .B2(n18848), .C1(
        n18727), .C2(n18776), .ZN(P3_U3035) );
  OAI222_X1 U21884 ( .A1(n20797), .A2(n18776), .B1(n20793), .B2(n18848), .C1(
        n18729), .C2(n18772), .ZN(P3_U3036) );
  OAI222_X1 U21885 ( .A1(n18772), .A2(n18731), .B1(n18730), .B2(n18848), .C1(
        n18729), .C2(n18776), .ZN(P3_U3037) );
  OAI222_X1 U21886 ( .A1(n18772), .A2(n18734), .B1(n18732), .B2(n18848), .C1(
        n18731), .C2(n18776), .ZN(P3_U3038) );
  OAI222_X1 U21887 ( .A1(n18734), .A2(n18776), .B1(n18733), .B2(n18848), .C1(
        n18735), .C2(n18772), .ZN(P3_U3039) );
  OAI222_X1 U21888 ( .A1(n18772), .A2(n18736), .B1(n20920), .B2(n18848), .C1(
        n18735), .C2(n18776), .ZN(P3_U3040) );
  OAI222_X1 U21889 ( .A1(n18772), .A2(n18737), .B1(n20803), .B2(n18848), .C1(
        n18736), .C2(n18776), .ZN(P3_U3041) );
  OAI222_X1 U21890 ( .A1(n18772), .A2(n18740), .B1(n18738), .B2(n18848), .C1(
        n18737), .C2(n18776), .ZN(P3_U3042) );
  OAI222_X1 U21891 ( .A1(n18740), .A2(n18776), .B1(n18739), .B2(n18848), .C1(
        n18741), .C2(n18772), .ZN(P3_U3043) );
  OAI222_X1 U21892 ( .A1(n18772), .A2(n18744), .B1(n18742), .B2(n18848), .C1(
        n18741), .C2(n18776), .ZN(P3_U3044) );
  OAI222_X1 U21893 ( .A1(n18744), .A2(n18776), .B1(n18743), .B2(n18848), .C1(
        n18745), .C2(n18772), .ZN(P3_U3045) );
  OAI222_X1 U21894 ( .A1(n18772), .A2(n18747), .B1(n18746), .B2(n18848), .C1(
        n18745), .C2(n18776), .ZN(P3_U3046) );
  OAI222_X1 U21895 ( .A1(n18772), .A2(n18750), .B1(n18748), .B2(n18848), .C1(
        n18747), .C2(n18776), .ZN(P3_U3047) );
  OAI222_X1 U21896 ( .A1(n18750), .A2(n18776), .B1(n18749), .B2(n18848), .C1(
        n20902), .C2(n18772), .ZN(P3_U3048) );
  OAI222_X1 U21897 ( .A1(n20902), .A2(n18776), .B1(n18751), .B2(n18848), .C1(
        n18752), .C2(n18772), .ZN(P3_U3049) );
  OAI222_X1 U21898 ( .A1(n18772), .A2(n18754), .B1(n18753), .B2(n18848), .C1(
        n18752), .C2(n18776), .ZN(P3_U3050) );
  OAI222_X1 U21899 ( .A1(n18772), .A2(n18756), .B1(n18755), .B2(n18848), .C1(
        n18754), .C2(n18776), .ZN(P3_U3051) );
  OAI222_X1 U21900 ( .A1(n18772), .A2(n18758), .B1(n18757), .B2(n18848), .C1(
        n18756), .C2(n18776), .ZN(P3_U3052) );
  OAI222_X1 U21901 ( .A1(n18772), .A2(n18760), .B1(n18759), .B2(n18848), .C1(
        n18758), .C2(n18776), .ZN(P3_U3053) );
  OAI222_X1 U21902 ( .A1(n18772), .A2(n18762), .B1(n18761), .B2(n18848), .C1(
        n18760), .C2(n18776), .ZN(P3_U3054) );
  OAI222_X1 U21903 ( .A1(n18772), .A2(n20745), .B1(n18763), .B2(n18848), .C1(
        n18762), .C2(n18776), .ZN(P3_U3055) );
  INV_X1 U21904 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18765) );
  OAI222_X1 U21905 ( .A1(n18772), .A2(n18765), .B1(n18764), .B2(n18848), .C1(
        n20745), .C2(n18776), .ZN(P3_U3056) );
  OAI222_X1 U21906 ( .A1(n18772), .A2(n18767), .B1(n18766), .B2(n18848), .C1(
        n18765), .C2(n18776), .ZN(P3_U3057) );
  INV_X1 U21907 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18769) );
  OAI222_X1 U21908 ( .A1(n18772), .A2(n18769), .B1(n20891), .B2(n18848), .C1(
        n18767), .C2(n18776), .ZN(P3_U3058) );
  OAI222_X1 U21909 ( .A1(n18769), .A2(n18776), .B1(n18768), .B2(n18848), .C1(
        n18770), .C2(n18772), .ZN(P3_U3059) );
  OAI222_X1 U21910 ( .A1(n18772), .A2(n18775), .B1(n18771), .B2(n18848), .C1(
        n18770), .C2(n18776), .ZN(P3_U3060) );
  OAI222_X1 U21911 ( .A1(n18776), .A2(n18775), .B1(n18774), .B2(n18848), .C1(
        n18773), .C2(n18772), .ZN(P3_U3061) );
  INV_X1 U21912 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18777) );
  AOI22_X1 U21913 ( .A1(n18848), .A2(n20791), .B1(n18777), .B2(n18849), .ZN(
        P3_U3274) );
  INV_X1 U21914 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18825) );
  INV_X1 U21915 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U21916 ( .A1(n18848), .A2(n18825), .B1(n20730), .B2(n18849), .ZN(
        P3_U3275) );
  INV_X1 U21917 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18778) );
  AOI22_X1 U21918 ( .A1(n18848), .A2(n18779), .B1(n18778), .B2(n18849), .ZN(
        P3_U3276) );
  INV_X1 U21919 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18828) );
  INV_X1 U21920 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18780) );
  AOI22_X1 U21921 ( .A1(n18848), .A2(n18828), .B1(n18780), .B2(n18849), .ZN(
        P3_U3277) );
  INV_X1 U21922 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18782) );
  INV_X1 U21923 ( .A(n18784), .ZN(n18781) );
  AOI21_X1 U21924 ( .B1(n18783), .B2(n18782), .A(n18781), .ZN(P3_U3280) );
  OAI21_X1 U21925 ( .B1(n18786), .B2(n18785), .A(n18784), .ZN(P3_U3281) );
  INV_X1 U21926 ( .A(n18787), .ZN(n18790) );
  OAI21_X1 U21927 ( .B1(n18790), .B2(n18789), .A(n18788), .ZN(P3_U3282) );
  NOR2_X1 U21928 ( .A1(n18791), .A2(n18803), .ZN(n18792) );
  INV_X1 U21929 ( .A(n18819), .ZN(n18822) );
  NOR2_X1 U21930 ( .A1(n18792), .A2(n18822), .ZN(n18797) );
  INV_X1 U21931 ( .A(n18793), .ZN(n18794) );
  AOI22_X1 U21932 ( .A1(n18817), .A2(n18795), .B1(n18815), .B2(n18794), .ZN(
        n18796) );
  OAI22_X1 U21933 ( .A1(n20947), .A2(n18797), .B1(n18822), .B2(n18796), .ZN(
        P3_U3285) );
  AOI22_X1 U21934 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18799), .B2(n18798), .ZN(
        n18809) );
  NOR2_X1 U21935 ( .A1(n18800), .A2(n18818), .ZN(n18810) );
  INV_X1 U21936 ( .A(n18815), .ZN(n18802) );
  OAI22_X1 U21937 ( .A1(n18804), .A2(n18803), .B1(n18802), .B2(n18801), .ZN(
        n18805) );
  AOI21_X1 U21938 ( .B1(n18809), .B2(n18810), .A(n18805), .ZN(n18806) );
  AOI22_X1 U21939 ( .A1(n18822), .A2(n18807), .B1(n18806), .B2(n18819), .ZN(
        P3_U3288) );
  INV_X1 U21940 ( .A(n18808), .ZN(n18812) );
  INV_X1 U21941 ( .A(n18809), .ZN(n18811) );
  AOI222_X1 U21942 ( .A1(n18813), .A2(n18817), .B1(n18815), .B2(n18812), .C1(
        n18811), .C2(n18810), .ZN(n18814) );
  AOI22_X1 U21943 ( .A1(n18822), .A2(n12634), .B1(n18814), .B2(n18819), .ZN(
        P3_U3289) );
  AOI222_X1 U21944 ( .A1(n18818), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18817), 
        .B2(n18816), .C1(n18821), .C2(n18815), .ZN(n18820) );
  AOI22_X1 U21945 ( .A1(n18822), .A2(n18821), .B1(n18820), .B2(n18819), .ZN(
        P3_U3290) );
  AOI21_X1 U21946 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18823) );
  AOI22_X1 U21947 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18823), .B2(n20926), .ZN(n18826) );
  AOI22_X1 U21948 ( .A1(n18829), .A2(n18826), .B1(n18825), .B2(n18824), .ZN(
        P3_U3292) );
  OAI21_X1 U21949 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18829), .ZN(n18827) );
  OAI21_X1 U21950 ( .B1(n18829), .B2(n18828), .A(n18827), .ZN(P3_U3293) );
  INV_X1 U21951 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18830) );
  AOI22_X1 U21952 ( .A1(n18848), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18830), 
        .B2(n18849), .ZN(P3_U3294) );
  MUX2_X1 U21953 ( .A(P3_MORE_REG_SCAN_IN), .B(n18832), .S(n18831), .Z(
        P3_U3295) );
  INV_X1 U21954 ( .A(n18833), .ZN(n18834) );
  OAI21_X1 U21955 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18835), .A(n18834), 
        .ZN(n18838) );
  AOI211_X1 U21956 ( .C1(n18854), .C2(n18838), .A(n18837), .B(n18836), .ZN(
        n18841) );
  OAI21_X1 U21957 ( .B1(n18841), .B2(n18840), .A(n18839), .ZN(n18847) );
  AOI21_X1 U21958 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18842), .ZN(n18843) );
  AOI211_X1 U21959 ( .C1(n18845), .C2(n18844), .A(n18843), .B(n18853), .ZN(
        n18846) );
  MUX2_X1 U21960 ( .A(n18847), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18846), 
        .Z(P3_U3296) );
  OAI22_X1 U21961 ( .A1(n18849), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18848), .ZN(n18850) );
  INV_X1 U21962 ( .A(n18850), .ZN(P3_U3297) );
  NOR2_X1 U21963 ( .A1(n18851), .A2(n18853), .ZN(n18855) );
  INV_X1 U21964 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18852) );
  AOI22_X1 U21965 ( .A1(n18854), .A2(n18853), .B1(n18855), .B2(n18852), .ZN(
        P3_U3298) );
  INV_X1 U21966 ( .A(n18855), .ZN(n18857) );
  OAI21_X1 U21967 ( .B1(n18857), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18856), 
        .ZN(n18858) );
  INV_X1 U21968 ( .A(n18858), .ZN(P3_U3299) );
  INV_X1 U21969 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18860) );
  INV_X1 U21970 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18859) );
  INV_X1 U21971 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19802) );
  NAND2_X1 U21972 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19802), .ZN(n19790) );
  AOI22_X1 U21973 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19790), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n18860), .ZN(n19851) );
  OAI21_X1 U21974 ( .B1(n18860), .B2(n18859), .A(n19783), .ZN(P2_U2815) );
  INV_X1 U21975 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19791) );
  OR2_X1 U21976 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19791), .ZN(n19898) );
  INV_X2 U21977 ( .A(n19898), .ZN(n19901) );
  AOI21_X1 U21978 ( .B1(n19802), .B2(n18860), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18861) );
  AOI22_X1 U21979 ( .A1(n19901), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18861), 
        .B2(n19898), .ZN(P2_U2817) );
  OAI21_X1 U21980 ( .B1(n19795), .B2(BS16), .A(n19851), .ZN(n19849) );
  OAI21_X1 U21981 ( .B1(n19851), .B2(n19666), .A(n19849), .ZN(P2_U2818) );
  AND2_X1 U21982 ( .A1(n18863), .A2(n18862), .ZN(n19896) );
  OAI21_X1 U21983 ( .B1(n19896), .B2(n18865), .A(n18864), .ZN(P2_U2819) );
  NOR4_X1 U21984 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18875) );
  NOR4_X1 U21985 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18874) );
  AOI211_X1 U21986 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18866) );
  INV_X1 U21987 ( .A(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20809) );
  INV_X1 U21988 ( .A(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20713) );
  NAND3_X1 U21989 ( .A1(n18866), .A2(n20809), .A3(n20713), .ZN(n18872) );
  NOR4_X1 U21990 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18870) );
  NOR4_X1 U21991 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n18869) );
  NOR4_X1 U21992 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18868) );
  NOR4_X1 U21993 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18867) );
  NAND4_X1 U21994 ( .A1(n18870), .A2(n18869), .A3(n18868), .A4(n18867), .ZN(
        n18871) );
  NOR4_X1 U21995 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n18872), .A4(n18871), .ZN(n18873) );
  NAND3_X1 U21996 ( .A1(n18875), .A2(n18874), .A3(n18873), .ZN(n18881) );
  NOR2_X1 U21997 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18881), .ZN(n18876) );
  INV_X1 U21998 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U21999 ( .A1(n18876), .A2(n18997), .B1(n18881), .B2(n19847), .ZN(
        P2_U2820) );
  OR3_X1 U22000 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18880) );
  INV_X1 U22001 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U22002 ( .A1(n18876), .A2(n18880), .B1(n18881), .B2(n19845), .ZN(
        P2_U2821) );
  INV_X1 U22003 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19850) );
  NAND2_X1 U22004 ( .A1(n18876), .A2(n19850), .ZN(n18879) );
  INV_X1 U22005 ( .A(n18881), .ZN(n18882) );
  OAI21_X1 U22006 ( .B1(n18997), .B2(n12971), .A(n18882), .ZN(n18877) );
  OAI21_X1 U22007 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18882), .A(n18877), 
        .ZN(n18878) );
  OAI221_X1 U22008 ( .B1(n18879), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18879), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18878), .ZN(P2_U2822) );
  INV_X1 U22009 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20839) );
  OAI221_X1 U22010 ( .B1(n18882), .B2(n20839), .C1(n18881), .C2(n18880), .A(
        n18879), .ZN(P2_U2823) );
  AOI22_X1 U22011 ( .A1(n18884), .A2(n19002), .B1(n19007), .B2(n18883), .ZN(
        n18892) );
  AOI211_X1 U22012 ( .C1(n18886), .C2(n9834), .A(n18885), .B(n12836), .ZN(
        n18890) );
  AOI22_X1 U22013 ( .A1(n18887), .A2(n20703), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19012), .ZN(n18888) );
  OAI211_X1 U22014 ( .C1(n19822), .C2(n20697), .A(n18888), .B(n18970), .ZN(
        n18889) );
  AOI211_X1 U22015 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n20694), .A(n18890), .B(
        n18889), .ZN(n18891) );
  NAND2_X1 U22016 ( .A1(n18892), .A2(n18891), .ZN(P2_U2836) );
  INV_X1 U22017 ( .A(n18901), .ZN(n18895) );
  INV_X1 U22018 ( .A(n18947), .ZN(n19011) );
  AOI22_X1 U22019 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19012), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n20694), .ZN(n18893) );
  OAI211_X1 U22020 ( .C1(n20697), .C2(n19819), .A(n18893), .B(n18933), .ZN(
        n18894) );
  AOI21_X1 U22021 ( .B1(n18895), .B2(n19011), .A(n18894), .ZN(n18896) );
  OAI21_X1 U22022 ( .B1(n18897), .B2(n19005), .A(n18896), .ZN(n18898) );
  AOI21_X1 U22023 ( .B1(n18899), .B2(n19007), .A(n18898), .ZN(n18904) );
  OAI211_X1 U22024 ( .C1(n18902), .C2(n18901), .A(n19009), .B(n18900), .ZN(
        n18903) );
  OAI211_X1 U22025 ( .C1(n20698), .C2(n18905), .A(n18904), .B(n18903), .ZN(
        P2_U2838) );
  OAI22_X1 U22026 ( .A1(n18907), .A2(n19005), .B1(n18906), .B2(n18981), .ZN(
        n18908) );
  AOI211_X1 U22027 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18986), .A(n18985), 
        .B(n18908), .ZN(n18916) );
  NOR2_X1 U22028 ( .A1(n10032), .A2(n18909), .ZN(n18910) );
  XNOR2_X1 U22029 ( .A(n18911), .B(n18910), .ZN(n18914) );
  OAI22_X1 U22030 ( .A1(n19069), .A2(n20698), .B1(n20705), .B2(n18912), .ZN(
        n18913) );
  AOI21_X1 U22031 ( .B1(n18914), .B2(n19009), .A(n18913), .ZN(n18915) );
  OAI211_X1 U22032 ( .C1(n18999), .C2(n18917), .A(n18916), .B(n18915), .ZN(
        P2_U2840) );
  INV_X1 U22033 ( .A(n18918), .ZN(n18926) );
  INV_X1 U22034 ( .A(n18919), .ZN(n18924) );
  INV_X1 U22035 ( .A(n18928), .ZN(n18922) );
  AOI22_X1 U22036 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n20694), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19012), .ZN(n18920) );
  OAI211_X1 U22037 ( .C1(n20697), .C2(n15298), .A(n18920), .B(n18933), .ZN(
        n18921) );
  AOI21_X1 U22038 ( .B1(n18922), .B2(n19011), .A(n18921), .ZN(n18923) );
  OAI21_X1 U22039 ( .B1(n18924), .B2(n19005), .A(n18923), .ZN(n18925) );
  AOI21_X1 U22040 ( .B1(n18926), .B2(n19007), .A(n18925), .ZN(n18931) );
  OAI21_X1 U22041 ( .B1(n18929), .B2(n18928), .A(n18927), .ZN(n18930) );
  OAI211_X1 U22042 ( .C1(n20698), .C2(n19074), .A(n18931), .B(n18930), .ZN(
        P2_U2842) );
  INV_X1 U22043 ( .A(n18932), .ZN(n18940) );
  AOI22_X1 U22044 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n20694), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19012), .ZN(n18934) );
  OAI211_X1 U22045 ( .C1(n20697), .C2(n19811), .A(n18934), .B(n18933), .ZN(
        n18935) );
  AOI21_X1 U22046 ( .B1(n19002), .B2(n18936), .A(n18935), .ZN(n18937) );
  OAI21_X1 U22047 ( .B1(n18938), .B2(n19005), .A(n18937), .ZN(n18939) );
  AOI21_X1 U22048 ( .B1(n18940), .B2(n19007), .A(n18939), .ZN(n18945) );
  NOR2_X1 U22049 ( .A1(n10032), .A2(n12836), .ZN(n18942) );
  OAI211_X1 U22050 ( .C1(n18943), .C2(n18946), .A(n18942), .B(n18941), .ZN(
        n18944) );
  OAI211_X1 U22051 ( .C1(n18947), .C2(n18946), .A(n18945), .B(n18944), .ZN(
        P2_U2844) );
  NAND2_X1 U22052 ( .A1(n13659), .A2(n18948), .ZN(n18950) );
  XOR2_X1 U22053 ( .A(n18950), .B(n18949), .Z(n18958) );
  INV_X1 U22054 ( .A(n18951), .ZN(n18952) );
  AOI22_X1 U22055 ( .A1(n18952), .A2(n20703), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n20694), .ZN(n18953) );
  OAI211_X1 U22056 ( .C1(n12298), .C2(n20697), .A(n18953), .B(n18933), .ZN(
        n18956) );
  INV_X1 U22057 ( .A(n19033), .ZN(n18954) );
  OAI22_X1 U22058 ( .A1(n18954), .A2(n20705), .B1(n20698), .B2(n19084), .ZN(
        n18955) );
  AOI211_X1 U22059 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19012), .A(
        n18956), .B(n18955), .ZN(n18957) );
  OAI21_X1 U22060 ( .B1(n18958), .B2(n12836), .A(n18957), .ZN(P2_U2845) );
  NOR2_X1 U22061 ( .A1(n10032), .A2(n18959), .ZN(n18960) );
  XOR2_X1 U22062 ( .A(n18961), .B(n18960), .Z(n18969) );
  AOI22_X1 U22063 ( .A1(n18962), .A2(n20703), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19012), .ZN(n18963) );
  OAI211_X1 U22064 ( .C1(n15329), .C2(n20697), .A(n18963), .B(n18933), .ZN(
        n18967) );
  INV_X1 U22065 ( .A(n18964), .ZN(n18965) );
  OAI22_X1 U22066 ( .A1(n18965), .A2(n20705), .B1(n20698), .B2(n19087), .ZN(
        n18966) );
  AOI211_X1 U22067 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n20694), .A(n18967), .B(
        n18966), .ZN(n18968) );
  OAI21_X1 U22068 ( .B1(n12836), .B2(n18969), .A(n18968), .ZN(P2_U2846) );
  OAI21_X1 U22069 ( .B1(n10734), .B2(n20697), .A(n18970), .ZN(n18973) );
  OAI22_X1 U22070 ( .A1(n18971), .A2(n19005), .B1(n18999), .B2(n13266), .ZN(
        n18972) );
  AOI211_X1 U22071 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19012), .A(
        n18973), .B(n18972), .ZN(n18980) );
  NAND2_X1 U22072 ( .A1(n10012), .A2(n18974), .ZN(n18975) );
  XNOR2_X1 U22073 ( .A(n18976), .B(n18975), .ZN(n18978) );
  AOI22_X1 U22074 ( .A1(n18978), .A2(n19009), .B1(n19007), .B2(n18977), .ZN(
        n18979) );
  OAI211_X1 U22075 ( .C1(n20698), .C2(n19093), .A(n18980), .B(n18979), .ZN(
        P2_U2849) );
  INV_X1 U22076 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18996) );
  OAI22_X1 U22077 ( .A1(n18983), .A2(n19005), .B1(n18982), .B2(n18981), .ZN(
        n18984) );
  AOI211_X1 U22078 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18986), .A(n18985), .B(
        n18984), .ZN(n18995) );
  NOR2_X1 U22079 ( .A1(n10032), .A2(n18987), .ZN(n18989) );
  XNOR2_X1 U22080 ( .A(n18990), .B(n18989), .ZN(n18993) );
  OAI22_X1 U22081 ( .A1(n19101), .A2(n20698), .B1(n20705), .B2(n18991), .ZN(
        n18992) );
  AOI21_X1 U22082 ( .B1(n18993), .B2(n19009), .A(n18992), .ZN(n18994) );
  OAI211_X1 U22083 ( .C1(n18999), .C2(n18996), .A(n18995), .B(n18994), .ZN(
        P2_U2850) );
  OAI22_X1 U22084 ( .A1(n18999), .A2(n18998), .B1(n18997), .B2(n20697), .ZN(
        n19000) );
  AOI21_X1 U22085 ( .B1(n19002), .B2(n19001), .A(n19000), .ZN(n19003) );
  OAI21_X1 U22086 ( .B1(n19005), .B2(n19004), .A(n19003), .ZN(n19006) );
  AOI21_X1 U22087 ( .B1(n19008), .B2(n19007), .A(n19006), .ZN(n19015) );
  AOI22_X1 U22088 ( .A1(n19010), .A2(n19009), .B1(n19444), .B2(n20707), .ZN(
        n19014) );
  OAI21_X1 U22089 ( .B1(n19012), .B2(n19011), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19013) );
  NAND3_X1 U22090 ( .A1(n19015), .A2(n19014), .A3(n19013), .ZN(P2_U2855) );
  OR2_X1 U22091 ( .A1(n13942), .A2(n19016), .ZN(n19017) );
  NAND2_X1 U22092 ( .A1(n13869), .A2(n19017), .ZN(n19062) );
  INV_X1 U22093 ( .A(n19062), .ZN(n19019) );
  AOI22_X1 U22094 ( .A1(n19019), .A2(n19018), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19052), .ZN(n19020) );
  OAI21_X1 U22095 ( .B1(n19052), .B2(n19021), .A(n19020), .ZN(P2_U2871) );
  AOI21_X1 U22096 ( .B1(n19024), .B2(n19023), .A(n19022), .ZN(n19027) );
  INV_X1 U22097 ( .A(n19025), .ZN(n19026) );
  NOR3_X1 U22098 ( .A1(n19027), .A2(n19026), .A3(n19041), .ZN(n19028) );
  AOI21_X1 U22099 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19052), .A(n19028), .ZN(
        n19029) );
  OAI21_X1 U22100 ( .B1(n19030), .B2(n19052), .A(n19029), .ZN(P2_U2873) );
  INV_X1 U22101 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19036) );
  AOI21_X1 U22102 ( .B1(n19032), .B2(n19031), .A(n19041), .ZN(n19034) );
  AOI22_X1 U22103 ( .A1(n19034), .A2(n13720), .B1(n19033), .B2(n19048), .ZN(
        n19035) );
  OAI21_X1 U22104 ( .B1(n19048), .B2(n19036), .A(n19035), .ZN(P2_U2877) );
  AND2_X1 U22105 ( .A1(n9755), .A2(n19037), .ZN(n19039) );
  NAND2_X1 U22106 ( .A1(n19039), .A2(n19038), .ZN(n19042) );
  AOI211_X1 U22107 ( .C1(n19043), .C2(n19042), .A(n19041), .B(n19040), .ZN(
        n19044) );
  AOI21_X1 U22108 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19052), .A(n19044), .ZN(
        n19045) );
  OAI21_X1 U22109 ( .B1(n19046), .B2(n19052), .A(n19045), .ZN(P2_U2879) );
  OAI22_X1 U22110 ( .A1(n19105), .A2(n19041), .B1(n19048), .B2(n19047), .ZN(
        n19049) );
  INV_X1 U22111 ( .A(n19049), .ZN(n19050) );
  OAI21_X1 U22112 ( .B1(n19052), .B2(n19051), .A(n19050), .ZN(P2_U2883) );
  INV_X1 U22113 ( .A(n19061), .ZN(n19055) );
  OAI22_X1 U22114 ( .A1(n19053), .A2(n19063), .B1(n19055), .B2(n19054), .ZN(
        n19056) );
  INV_X1 U22115 ( .A(n19056), .ZN(n19058) );
  AOI22_X1 U22116 ( .A1(n19060), .A2(BUF2_REG_31__SCAN_IN), .B1(n19119), .B2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n19057) );
  NAND2_X1 U22117 ( .A1(n19058), .A2(n19057), .ZN(P2_U2888) );
  AOI22_X1 U22118 ( .A1(n19059), .A2(n19185), .B1(n19119), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19068) );
  AOI22_X1 U22119 ( .A1(n19061), .A2(BUF1_REG_16__SCAN_IN), .B1(n19060), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19067) );
  OAI22_X1 U22120 ( .A1(n19064), .A2(n19063), .B1(n19124), .B2(n19062), .ZN(
        n19065) );
  INV_X1 U22121 ( .A(n19065), .ZN(n19066) );
  NAND3_X1 U22122 ( .A1(n19068), .A2(n19067), .A3(n19066), .ZN(P2_U2903) );
  INV_X1 U22123 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19135) );
  OAI222_X1 U22124 ( .A1(n19095), .A2(n19135), .B1(n19128), .B2(n19070), .C1(
        n19069), .C2(n19102), .ZN(P2_U2904) );
  AOI22_X1 U22125 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19119), .B1(n19071), 
        .B2(n19096), .ZN(n19072) );
  OAI21_X1 U22126 ( .B1(n19102), .B2(n19073), .A(n19072), .ZN(P2_U2905) );
  INV_X1 U22127 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19139) );
  OAI222_X1 U22128 ( .A1(n19095), .A2(n19139), .B1(n19075), .B2(n19128), .C1(
        n19074), .C2(n19102), .ZN(P2_U2906) );
  INV_X1 U22129 ( .A(n19076), .ZN(n19079) );
  AOI22_X1 U22130 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19119), .B1(n19077), 
        .B2(n19096), .ZN(n19078) );
  OAI21_X1 U22131 ( .B1(n19102), .B2(n19079), .A(n19078), .ZN(P2_U2907) );
  INV_X1 U22132 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19143) );
  OAI222_X1 U22133 ( .A1(n19095), .A2(n19143), .B1(n19081), .B2(n19128), .C1(
        n19080), .C2(n19102), .ZN(P2_U2908) );
  AOI22_X1 U22134 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19119), .B1(n19082), 
        .B2(n19096), .ZN(n19083) );
  OAI21_X1 U22135 ( .B1(n19102), .B2(n19084), .A(n19083), .ZN(P2_U2909) );
  AOI22_X1 U22136 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19119), .B1(n19085), .B2(
        n19096), .ZN(n19086) );
  OAI21_X1 U22137 ( .B1(n19102), .B2(n19087), .A(n19086), .ZN(P2_U2910) );
  INV_X1 U22138 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19149) );
  OAI222_X1 U22139 ( .A1(n19095), .A2(n19149), .B1(n19089), .B2(n19128), .C1(
        n19088), .C2(n19102), .ZN(P2_U2911) );
  INV_X1 U22140 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19151) );
  INV_X1 U22141 ( .A(n19090), .ZN(n19091) );
  OAI222_X1 U22142 ( .A1(n19095), .A2(n19151), .B1(n19092), .B2(n19128), .C1(
        n19091), .C2(n19102), .ZN(P2_U2912) );
  INV_X1 U22143 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20888) );
  OAI222_X1 U22144 ( .A1(n19095), .A2(n20888), .B1(n19094), .B2(n19128), .C1(
        n19093), .C2(n19102), .ZN(P2_U2913) );
  AOI22_X1 U22145 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19119), .B1(n19203), .B2(
        n19096), .ZN(n19100) );
  AOI21_X1 U22146 ( .B1(n20699), .B2(n19866), .A(n19097), .ZN(n19114) );
  XNOR2_X1 U22147 ( .A(n19445), .B(n19861), .ZN(n19113) );
  NOR2_X1 U22148 ( .A1(n19114), .A2(n19113), .ZN(n19112) );
  AOI21_X1 U22149 ( .B1(n19445), .B2(n19861), .A(n19112), .ZN(n19098) );
  NOR2_X1 U22150 ( .A1(n19098), .A2(n19103), .ZN(n19104) );
  OR3_X1 U22151 ( .A1(n19104), .A2(n19105), .A3(n19124), .ZN(n19099) );
  OAI211_X1 U22152 ( .C1(n19102), .C2(n19101), .A(n19100), .B(n19099), .ZN(
        P2_U2914) );
  AOI22_X1 U22153 ( .A1(n19120), .A2(n19103), .B1(n19119), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19109) );
  XOR2_X1 U22154 ( .A(n19105), .B(n19104), .Z(n19107) );
  NAND2_X1 U22155 ( .A1(n19107), .A2(n19106), .ZN(n19108) );
  OAI211_X1 U22156 ( .C1(n19110), .C2(n19128), .A(n19109), .B(n19108), .ZN(
        P2_U2915) );
  INV_X1 U22157 ( .A(n19861), .ZN(n19111) );
  AOI22_X1 U22158 ( .A1(n19111), .A2(n19120), .B1(n19119), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19117) );
  AOI21_X1 U22159 ( .B1(n19114), .B2(n19113), .A(n19112), .ZN(n19115) );
  OR2_X1 U22160 ( .A1(n19115), .A2(n19124), .ZN(n19116) );
  OAI211_X1 U22161 ( .C1(n19118), .C2(n19128), .A(n19117), .B(n19116), .ZN(
        P2_U2916) );
  AOI22_X1 U22162 ( .A1(n19879), .A2(n19120), .B1(n19119), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19127) );
  AOI21_X1 U22163 ( .B1(n19123), .B2(n19122), .A(n19121), .ZN(n19125) );
  OR2_X1 U22164 ( .A1(n19125), .A2(n19124), .ZN(n19126) );
  OAI211_X1 U22165 ( .C1(n19129), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        P2_U2918) );
  NOR2_X1 U22166 ( .A1(n19152), .A2(n19130), .ZN(P2_U2920) );
  INV_X1 U22167 ( .A(n19131), .ZN(n19132) );
  AOI22_X1 U22168 ( .A1(n19132), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19167), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n19133) );
  OAI21_X1 U22169 ( .B1(n20783), .B2(n19152), .A(n19133), .ZN(P2_U2933) );
  AOI22_X1 U22170 ( .A1(n19167), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U22171 ( .B1(n19170), .B2(n19135), .A(n19134), .ZN(P2_U2936) );
  AOI22_X1 U22172 ( .A1(n19167), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19136) );
  OAI21_X1 U22173 ( .B1(n19170), .B2(n19137), .A(n19136), .ZN(P2_U2937) );
  AOI22_X1 U22174 ( .A1(n19167), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19138) );
  OAI21_X1 U22175 ( .B1(n19170), .B2(n19139), .A(n19138), .ZN(P2_U2938) );
  AOI22_X1 U22176 ( .A1(n19167), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22177 ( .B1(n19170), .B2(n19141), .A(n19140), .ZN(P2_U2939) );
  AOI22_X1 U22178 ( .A1(n19167), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22179 ( .B1(n19170), .B2(n19143), .A(n19142), .ZN(P2_U2940) );
  AOI22_X1 U22180 ( .A1(n19167), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19144) );
  OAI21_X1 U22181 ( .B1(n19170), .B2(n19145), .A(n19144), .ZN(P2_U2941) );
  AOI22_X1 U22182 ( .A1(n19167), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19146) );
  OAI21_X1 U22183 ( .B1(n19170), .B2(n19147), .A(n19146), .ZN(P2_U2942) );
  AOI22_X1 U22184 ( .A1(n19167), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19148) );
  OAI21_X1 U22185 ( .B1(n19170), .B2(n19149), .A(n19148), .ZN(P2_U2943) );
  AOI22_X1 U22186 ( .A1(n19167), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U22187 ( .B1(n19170), .B2(n19151), .A(n19150), .ZN(P2_U2944) );
  INV_X1 U22188 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n19153) );
  OAI222_X1 U22189 ( .A1(n19153), .A2(n19156), .B1(n20888), .B2(n19170), .C1(
        n20749), .C2(n19152), .ZN(P2_U2945) );
  INV_X1 U22190 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U22191 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19154), .B1(n19157), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n19155) );
  OAI21_X1 U22192 ( .B1(n20718), .B2(n19156), .A(n19155), .ZN(P2_U2946) );
  INV_X1 U22193 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19159) );
  AOI22_X1 U22194 ( .A1(n19167), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19157), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22195 ( .B1(n19170), .B2(n19159), .A(n19158), .ZN(P2_U2947) );
  INV_X1 U22196 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19161) );
  AOI22_X1 U22197 ( .A1(n19167), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19160) );
  OAI21_X1 U22198 ( .B1(n19170), .B2(n19161), .A(n19160), .ZN(P2_U2948) );
  AOI22_X1 U22199 ( .A1(n19167), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19162) );
  OAI21_X1 U22200 ( .B1(n19170), .B2(n19163), .A(n19162), .ZN(P2_U2949) );
  INV_X1 U22201 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19165) );
  AOI22_X1 U22202 ( .A1(n19167), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19164) );
  OAI21_X1 U22203 ( .B1(n19170), .B2(n19165), .A(n19164), .ZN(P2_U2950) );
  INV_X1 U22204 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19169) );
  AOI22_X1 U22205 ( .A1(n19167), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19166), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19168) );
  OAI21_X1 U22206 ( .B1(n19170), .B2(n19169), .A(n19168), .ZN(P2_U2951) );
  INV_X1 U22207 ( .A(n20693), .ZN(n19171) );
  OAI22_X1 U22208 ( .A1(n19174), .A2(n19173), .B1(n19172), .B2(n19171), .ZN(
        n19175) );
  INV_X1 U22209 ( .A(n19175), .ZN(n19178) );
  NAND2_X1 U22210 ( .A1(n13180), .A2(n19176), .ZN(n19177) );
  OAI211_X1 U22211 ( .C1(n19180), .C2(n19179), .A(n19178), .B(n19177), .ZN(
        n19181) );
  INV_X1 U22212 ( .A(n19181), .ZN(n19183) );
  OAI211_X1 U22213 ( .C1(n19184), .C2(n12760), .A(n19183), .B(n19182), .ZN(
        P2_U3012) );
  AOI22_X1 U22214 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19213), .ZN(n19735) );
  INV_X1 U22215 ( .A(n19735), .ZN(n19623) );
  AND2_X1 U22216 ( .A1(n19216), .A2(n10243), .ZN(n19724) );
  AOI22_X1 U22217 ( .A1(n19777), .A2(n19623), .B1(n19190), .B2(n19724), .ZN(
        n19189) );
  AND2_X1 U22218 ( .A1(n19621), .A2(n19185), .ZN(n19725) );
  OAI22_X2 U22219 ( .A1(n19187), .A2(n19223), .B1(n19186), .B2(n19221), .ZN(
        n19732) );
  AOI22_X1 U22220 ( .A1(n19725), .A2(n19224), .B1(n19262), .B2(n19732), .ZN(
        n19188) );
  OAI211_X1 U22221 ( .C1(n19228), .C2(n20885), .A(n19189), .B(n19188), .ZN(
        P2_U3048) );
  INV_X1 U22222 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19195) );
  INV_X1 U22223 ( .A(n19741), .ZN(n19554) );
  AND2_X1 U22224 ( .A1(n19216), .A2(n13143), .ZN(n19736) );
  AOI22_X1 U22225 ( .A1(n19777), .A2(n19554), .B1(n19190), .B2(n19736), .ZN(
        n19194) );
  AND2_X1 U22226 ( .A1(n19191), .A2(n19621), .ZN(n19737) );
  OAI22_X2 U22227 ( .A1(n19192), .A2(n19223), .B1(n13875), .B2(n19221), .ZN(
        n19738) );
  AOI22_X1 U22228 ( .A1(n19737), .A2(n19224), .B1(n19262), .B2(n19738), .ZN(
        n19193) );
  OAI211_X1 U22229 ( .C1(n19228), .C2(n19195), .A(n19194), .B(n19193), .ZN(
        P2_U3049) );
  NAND2_X1 U22230 ( .A1(n19216), .A2(n10236), .ZN(n19685) );
  OAI22_X1 U22231 ( .A1(n19218), .A2(n19747), .B1(n19217), .B2(n19685), .ZN(
        n19196) );
  INV_X1 U22232 ( .A(n19196), .ZN(n19199) );
  AND2_X1 U22233 ( .A1(n19621), .A2(n19197), .ZN(n19743) );
  AOI22_X1 U22234 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19213), .ZN(n19686) );
  AOI22_X1 U22235 ( .A1(n19743), .A2(n19224), .B1(n19262), .B2(n19744), .ZN(
        n19198) );
  OAI211_X1 U22236 ( .C1(n19228), .C2(n13187), .A(n19199), .B(n19198), .ZN(
        P2_U3050) );
  OAI22_X1 U22237 ( .A1(n19201), .A2(n19223), .B1(n19200), .B2(n19221), .ZN(
        n19565) );
  NAND2_X1 U22238 ( .A1(n19216), .A2(n12214), .ZN(n19700) );
  OAI22_X1 U22239 ( .A1(n19218), .A2(n19765), .B1(n19217), .B2(n19700), .ZN(
        n19202) );
  INV_X1 U22240 ( .A(n19202), .ZN(n19205) );
  AND2_X1 U22241 ( .A1(n19203), .A2(n19621), .ZN(n19761) );
  AOI22_X1 U22242 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19213), .ZN(n19701) );
  INV_X1 U22243 ( .A(n19701), .ZN(n19762) );
  AOI22_X1 U22244 ( .A1(n19761), .A2(n19224), .B1(n19262), .B2(n19762), .ZN(
        n19204) );
  OAI211_X1 U22245 ( .C1(n19228), .C2(n13259), .A(n19205), .B(n19204), .ZN(
        P2_U3053) );
  INV_X1 U22246 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19212) );
  AND2_X1 U22247 ( .A1(n19216), .A2(n10216), .ZN(n19766) );
  INV_X1 U22248 ( .A(n19766), .ZN(n19705) );
  OAI22_X1 U22249 ( .A1(n19218), .A2(n19771), .B1(n19217), .B2(n19705), .ZN(
        n19206) );
  INV_X1 U22250 ( .A(n19206), .ZN(n19211) );
  AND2_X1 U22251 ( .A1(n19207), .A2(n19621), .ZN(n19767) );
  OAI22_X2 U22252 ( .A1(n19209), .A2(n19223), .B1(n19208), .B2(n19221), .ZN(
        n19768) );
  AOI22_X1 U22253 ( .A1(n19767), .A2(n19224), .B1(n19262), .B2(n19768), .ZN(
        n19210) );
  OAI211_X1 U22254 ( .C1(n19228), .C2(n19212), .A(n19211), .B(n19210), .ZN(
        P2_U3054) );
  AOI22_X1 U22255 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19214), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19213), .ZN(n19782) );
  NAND2_X1 U22256 ( .A1(n19216), .A2(n19215), .ZN(n19711) );
  OAI22_X1 U22257 ( .A1(n19218), .A2(n9848), .B1(n19217), .B2(n19711), .ZN(
        n19219) );
  INV_X1 U22258 ( .A(n19219), .ZN(n19226) );
  AND2_X1 U22259 ( .A1(n19220), .A2(n19621), .ZN(n19774) );
  AOI22_X1 U22260 ( .A1(n19774), .A2(n19224), .B1(n19262), .B2(n19776), .ZN(
        n19225) );
  OAI211_X1 U22261 ( .C1(n19228), .C2(n19227), .A(n19226), .B(n19225), .ZN(
        P2_U3055) );
  INV_X1 U22262 ( .A(n19732), .ZN(n19679) );
  NAND2_X1 U22263 ( .A1(n19295), .A2(n19881), .ZN(n19235) );
  NOR2_X1 U22264 ( .A1(n19890), .A2(n19235), .ZN(n19238) );
  INV_X1 U22265 ( .A(n19238), .ZN(n19259) );
  NAND2_X1 U22266 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19259), .ZN(n19229) );
  NOR2_X1 U22267 ( .A1(n10483), .A2(n19229), .ZN(n19234) );
  AND2_X1 U22268 ( .A1(n19235), .A2(n19723), .ZN(n19230) );
  INV_X1 U22269 ( .A(n19725), .ZN(n19613) );
  INV_X1 U22270 ( .A(n19724), .ZN(n19662) );
  OAI22_X1 U22271 ( .A1(n19260), .A2(n19613), .B1(n19662), .B2(n19259), .ZN(
        n19231) );
  INV_X1 U22272 ( .A(n19231), .ZN(n19240) );
  NAND2_X1 U22273 ( .A1(n19445), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19420) );
  INV_X1 U22274 ( .A(n19420), .ZN(n19233) );
  NAND2_X1 U22275 ( .A1(n19233), .A2(n19232), .ZN(n19236) );
  AOI21_X1 U22276 ( .B1(n19236), .B2(n19235), .A(n19234), .ZN(n19237) );
  OAI211_X1 U22277 ( .C1(n19238), .C2(n19668), .A(n19237), .B(n19621), .ZN(
        n19263) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19623), .ZN(n19239) );
  OAI211_X1 U22279 ( .C1(n19679), .C2(n19293), .A(n19240), .B(n19239), .ZN(
        P2_U3056) );
  INV_X1 U22280 ( .A(n19738), .ZN(n19684) );
  INV_X1 U22281 ( .A(n19737), .ZN(n19626) );
  INV_X1 U22282 ( .A(n19736), .ZN(n19680) );
  OAI22_X1 U22283 ( .A1(n19260), .A2(n19626), .B1(n19680), .B2(n19259), .ZN(
        n19241) );
  INV_X1 U22284 ( .A(n19241), .ZN(n19243) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19554), .ZN(n19242) );
  OAI211_X1 U22286 ( .C1(n19684), .C2(n19293), .A(n19243), .B(n19242), .ZN(
        P2_U3057) );
  INV_X1 U22287 ( .A(n19743), .ZN(n19630) );
  OAI22_X1 U22288 ( .A1(n19260), .A2(n19630), .B1(n19685), .B2(n19259), .ZN(
        n19244) );
  INV_X1 U22289 ( .A(n19244), .ZN(n19246) );
  INV_X1 U22290 ( .A(n19747), .ZN(n19632) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19632), .ZN(n19245) );
  OAI211_X1 U22292 ( .C1(n19686), .C2(n19293), .A(n19246), .B(n19245), .ZN(
        P2_U3058) );
  INV_X1 U22293 ( .A(n19750), .ZN(n19691) );
  INV_X1 U22294 ( .A(n19748), .ZN(n19690) );
  OAI22_X1 U22295 ( .A1(n19260), .A2(n19635), .B1(n19690), .B2(n19259), .ZN(
        n19247) );
  INV_X1 U22296 ( .A(n19247), .ZN(n19249) );
  INV_X1 U22297 ( .A(n19753), .ZN(n19559) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19559), .ZN(n19248) );
  OAI211_X1 U22299 ( .C1(n19691), .C2(n19293), .A(n19249), .B(n19248), .ZN(
        P2_U3059) );
  INV_X1 U22300 ( .A(n19756), .ZN(n19696) );
  INV_X1 U22301 ( .A(n19754), .ZN(n19695) );
  OAI22_X1 U22302 ( .A1(n19260), .A2(n19639), .B1(n19695), .B2(n19259), .ZN(
        n19250) );
  INV_X1 U22303 ( .A(n19250), .ZN(n19252) );
  INV_X1 U22304 ( .A(n19759), .ZN(n19562) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19562), .ZN(n19251) );
  OAI211_X1 U22306 ( .C1(n19696), .C2(n19293), .A(n19252), .B(n19251), .ZN(
        P2_U3060) );
  INV_X1 U22307 ( .A(n19761), .ZN(n19643) );
  OAI22_X1 U22308 ( .A1(n19260), .A2(n19643), .B1(n19700), .B2(n19259), .ZN(
        n19253) );
  INV_X1 U22309 ( .A(n19253), .ZN(n19255) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19565), .ZN(n19254) );
  OAI211_X1 U22311 ( .C1(n19701), .C2(n19293), .A(n19255), .B(n19254), .ZN(
        P2_U3061) );
  INV_X1 U22312 ( .A(n19768), .ZN(n19709) );
  INV_X1 U22313 ( .A(n19767), .ZN(n19647) );
  OAI22_X1 U22314 ( .A1(n19260), .A2(n19647), .B1(n19705), .B2(n19259), .ZN(
        n19256) );
  INV_X1 U22315 ( .A(n19256), .ZN(n19258) );
  INV_X1 U22316 ( .A(n19771), .ZN(n19649) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n19649), .ZN(n19257) );
  OAI211_X1 U22318 ( .C1(n19709), .C2(n19293), .A(n19258), .B(n19257), .ZN(
        P2_U3062) );
  INV_X1 U22319 ( .A(n19776), .ZN(n19712) );
  INV_X1 U22320 ( .A(n19774), .ZN(n19654) );
  OAI22_X1 U22321 ( .A1(n19260), .A2(n19654), .B1(n19711), .B2(n19259), .ZN(
        n19261) );
  INV_X1 U22322 ( .A(n19261), .ZN(n19265) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19263), .B1(
        n19262), .B2(n9847), .ZN(n19264) );
  OAI211_X1 U22324 ( .C1(n19712), .C2(n19293), .A(n19265), .B(n19264), .ZN(
        P2_U3063) );
  NOR3_X2 U22325 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19881), .A3(
        n19266), .ZN(n19288) );
  OAI21_X1 U22326 ( .B1(n19269), .B2(n19288), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19268) );
  INV_X1 U22327 ( .A(n19520), .ZN(n19267) );
  NAND2_X1 U22328 ( .A1(n19267), .A2(n19295), .ZN(n19270) );
  NAND2_X1 U22329 ( .A1(n19268), .A2(n19270), .ZN(n19289) );
  AOI22_X1 U22330 ( .A1(n19289), .A2(n19725), .B1(n19724), .B2(n19288), .ZN(
        n19275) );
  NOR2_X2 U22331 ( .A1(n19386), .A2(n19856), .ZN(n19317) );
  INV_X1 U22332 ( .A(n19869), .ZN(n19876) );
  AOI21_X1 U22333 ( .B1(n19293), .B2(n19327), .A(n19876), .ZN(n19273) );
  AOI21_X1 U22334 ( .B1(n19269), .B2(n19668), .A(n19288), .ZN(n19271) );
  OAI21_X1 U22335 ( .B1(n19271), .B2(n19852), .A(n19270), .ZN(n19272) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19732), .ZN(n19274) );
  OAI211_X1 U22337 ( .C1(n19735), .C2(n19293), .A(n19275), .B(n19274), .ZN(
        P2_U3064) );
  AOI22_X1 U22338 ( .A1(n19289), .A2(n19737), .B1(n19736), .B2(n19288), .ZN(
        n19277) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19738), .ZN(n19276) );
  OAI211_X1 U22340 ( .C1(n19741), .C2(n19293), .A(n19277), .B(n19276), .ZN(
        P2_U3065) );
  INV_X1 U22341 ( .A(n19685), .ZN(n19742) );
  AOI22_X1 U22342 ( .A1(n19289), .A2(n19743), .B1(n19742), .B2(n19288), .ZN(
        n19279) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19744), .ZN(n19278) );
  OAI211_X1 U22344 ( .C1(n19747), .C2(n19293), .A(n19279), .B(n19278), .ZN(
        P2_U3066) );
  AOI22_X1 U22345 ( .A1(n19289), .A2(n19749), .B1(n19748), .B2(n19288), .ZN(
        n19281) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19750), .ZN(n19280) );
  OAI211_X1 U22347 ( .C1(n19753), .C2(n19293), .A(n19281), .B(n19280), .ZN(
        P2_U3067) );
  AOI22_X1 U22348 ( .A1(n19289), .A2(n19755), .B1(n19754), .B2(n19288), .ZN(
        n19283) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19756), .ZN(n19282) );
  OAI211_X1 U22350 ( .C1(n19759), .C2(n19293), .A(n19283), .B(n19282), .ZN(
        P2_U3068) );
  AOI22_X1 U22351 ( .A1(n19289), .A2(n19761), .B1(n19760), .B2(n19288), .ZN(
        n19285) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19762), .ZN(n19284) );
  OAI211_X1 U22353 ( .C1(n19765), .C2(n19293), .A(n19285), .B(n19284), .ZN(
        P2_U3069) );
  AOI22_X1 U22354 ( .A1(n19289), .A2(n19767), .B1(n19766), .B2(n19288), .ZN(
        n19287) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19768), .ZN(n19286) );
  OAI211_X1 U22356 ( .C1(n19771), .C2(n19293), .A(n19287), .B(n19286), .ZN(
        P2_U3070) );
  INV_X1 U22357 ( .A(n19711), .ZN(n19772) );
  AOI22_X1 U22358 ( .A1(n19289), .A2(n19774), .B1(n19772), .B2(n19288), .ZN(
        n19292) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19290), .B1(
        n19317), .B2(n19776), .ZN(n19291) );
  OAI211_X1 U22360 ( .C1(n9848), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U3071) );
  OAI21_X1 U22361 ( .B1(n19420), .B2(n19856), .A(n19852), .ZN(n19305) );
  NAND2_X1 U22362 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19295), .ZN(
        n19304) );
  INV_X1 U22363 ( .A(n19304), .ZN(n19294) );
  OR2_X1 U22364 ( .A1(n19305), .A2(n19294), .ZN(n19300) );
  NAND2_X1 U22365 ( .A1(n19302), .A2(n19668), .ZN(n19298) );
  NAND2_X1 U22366 ( .A1(n19296), .A2(n19295), .ZN(n19301) );
  AND2_X1 U22367 ( .A1(n19301), .A2(n19581), .ZN(n19297) );
  AOI21_X1 U22368 ( .B1(n19298), .B2(n19297), .A(n19730), .ZN(n19299) );
  INV_X1 U22369 ( .A(n19301), .ZN(n19322) );
  AOI22_X1 U22370 ( .A1(n19344), .A2(n19732), .B1(n19322), .B2(n19724), .ZN(
        n19307) );
  OAI21_X1 U22371 ( .B1(n19302), .B2(n19322), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19303) );
  OAI21_X1 U22372 ( .B1(n19305), .B2(n19304), .A(n19303), .ZN(n19323) );
  AOI22_X1 U22373 ( .A1(n19725), .A2(n19323), .B1(n19317), .B2(n19623), .ZN(
        n19306) );
  OAI211_X1 U22374 ( .C1(n19308), .C2(n20951), .A(n19307), .B(n19306), .ZN(
        P2_U3072) );
  AOI22_X1 U22375 ( .A1(n19344), .A2(n19738), .B1(n19322), .B2(n19736), .ZN(
        n19310) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19324), .B1(
        n19737), .B2(n19323), .ZN(n19309) );
  OAI211_X1 U22377 ( .C1(n19741), .C2(n19327), .A(n19310), .B(n19309), .ZN(
        P2_U3073) );
  AOI22_X1 U22378 ( .A1(n19344), .A2(n19744), .B1(n19322), .B2(n19742), .ZN(
        n19312) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19324), .B1(
        n19743), .B2(n19323), .ZN(n19311) );
  OAI211_X1 U22380 ( .C1(n19747), .C2(n19327), .A(n19312), .B(n19311), .ZN(
        P2_U3074) );
  AOI22_X1 U22381 ( .A1(n19317), .A2(n19559), .B1(n19748), .B2(n19322), .ZN(
        n19314) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19324), .B1(
        n19749), .B2(n19323), .ZN(n19313) );
  OAI211_X1 U22383 ( .C1(n19691), .C2(n19356), .A(n19314), .B(n19313), .ZN(
        P2_U3075) );
  AOI22_X1 U22384 ( .A1(n19317), .A2(n19562), .B1(n19754), .B2(n19322), .ZN(
        n19316) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19324), .B1(
        n19755), .B2(n19323), .ZN(n19315) );
  OAI211_X1 U22386 ( .C1(n19696), .C2(n19356), .A(n19316), .B(n19315), .ZN(
        P2_U3076) );
  AOI22_X1 U22387 ( .A1(n19317), .A2(n19565), .B1(n19322), .B2(n19760), .ZN(
        n19319) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19324), .B1(
        n19761), .B2(n19323), .ZN(n19318) );
  OAI211_X1 U22389 ( .C1(n19701), .C2(n19356), .A(n19319), .B(n19318), .ZN(
        P2_U3077) );
  AOI22_X1 U22390 ( .A1(n19344), .A2(n19768), .B1(n19322), .B2(n19766), .ZN(
        n19321) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19324), .B1(
        n19767), .B2(n19323), .ZN(n19320) );
  OAI211_X1 U22392 ( .C1(n19771), .C2(n19327), .A(n19321), .B(n19320), .ZN(
        P2_U3078) );
  AOI22_X1 U22393 ( .A1(n19344), .A2(n19776), .B1(n19322), .B2(n19772), .ZN(
        n19326) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19324), .B1(
        n19774), .B2(n19323), .ZN(n19325) );
  OAI211_X1 U22395 ( .C1(n9848), .C2(n19327), .A(n19326), .B(n19325), .ZN(
        P2_U3079) );
  NOR2_X1 U22396 ( .A1(n19328), .A2(n19389), .ZN(n19586) );
  NAND2_X1 U22397 ( .A1(n19586), .A2(n19864), .ZN(n19330) );
  OR2_X1 U22398 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19330), .ZN(n19329) );
  NAND2_X1 U22399 ( .A1(n19864), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19415) );
  NOR2_X1 U22400 ( .A1(n19447), .A2(n19415), .ZN(n19351) );
  NOR3_X1 U22401 ( .A1(n10492), .A2(n19351), .A3(n19723), .ZN(n19331) );
  AOI21_X1 U22402 ( .B1(n19723), .B2(n19329), .A(n19331), .ZN(n19352) );
  AOI22_X1 U22403 ( .A1(n19352), .A2(n19725), .B1(n19724), .B2(n19351), .ZN(
        n19337) );
  INV_X1 U22404 ( .A(n19330), .ZN(n19335) );
  AOI21_X1 U22405 ( .B1(n19356), .B2(n19378), .A(n19666), .ZN(n19334) );
  INV_X1 U22406 ( .A(n19351), .ZN(n19332) );
  AOI211_X1 U22407 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19332), .A(n19730), 
        .B(n19331), .ZN(n19333) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19353), .B1(
        n19380), .B2(n19732), .ZN(n19336) );
  OAI211_X1 U22409 ( .C1(n19735), .C2(n19356), .A(n19337), .B(n19336), .ZN(
        P2_U3080) );
  AOI22_X1 U22410 ( .A1(n19352), .A2(n19737), .B1(n19736), .B2(n19351), .ZN(
        n19339) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19353), .B1(
        n19344), .B2(n19554), .ZN(n19338) );
  OAI211_X1 U22412 ( .C1(n19684), .C2(n19378), .A(n19339), .B(n19338), .ZN(
        P2_U3081) );
  AOI22_X1 U22413 ( .A1(n19352), .A2(n19743), .B1(n19742), .B2(n19351), .ZN(
        n19341) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19353), .B1(
        n19380), .B2(n19744), .ZN(n19340) );
  OAI211_X1 U22415 ( .C1(n19747), .C2(n19356), .A(n19341), .B(n19340), .ZN(
        P2_U3082) );
  AOI22_X1 U22416 ( .A1(n19352), .A2(n19749), .B1(n19748), .B2(n19351), .ZN(
        n19343) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19353), .B1(
        n19380), .B2(n19750), .ZN(n19342) );
  OAI211_X1 U22418 ( .C1(n19753), .C2(n19356), .A(n19343), .B(n19342), .ZN(
        P2_U3083) );
  AOI22_X1 U22419 ( .A1(n19352), .A2(n19755), .B1(n19754), .B2(n19351), .ZN(
        n19346) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19353), .B1(
        n19344), .B2(n19562), .ZN(n19345) );
  OAI211_X1 U22421 ( .C1(n19696), .C2(n19378), .A(n19346), .B(n19345), .ZN(
        P2_U3084) );
  AOI22_X1 U22422 ( .A1(n19352), .A2(n19761), .B1(n19760), .B2(n19351), .ZN(
        n19348) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19353), .B1(
        n19380), .B2(n19762), .ZN(n19347) );
  OAI211_X1 U22424 ( .C1(n19765), .C2(n19356), .A(n19348), .B(n19347), .ZN(
        P2_U3085) );
  AOI22_X1 U22425 ( .A1(n19352), .A2(n19767), .B1(n19766), .B2(n19351), .ZN(
        n19350) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19353), .B1(
        n19380), .B2(n19768), .ZN(n19349) );
  OAI211_X1 U22427 ( .C1(n19771), .C2(n19356), .A(n19350), .B(n19349), .ZN(
        P2_U3086) );
  AOI22_X1 U22428 ( .A1(n19352), .A2(n19774), .B1(n19772), .B2(n19351), .ZN(
        n19355) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19353), .B1(
        n19380), .B2(n19776), .ZN(n19354) );
  OAI211_X1 U22430 ( .C1(n9848), .C2(n19356), .A(n19355), .B(n19354), .ZN(
        P2_U3087) );
  NOR2_X1 U22431 ( .A1(n19415), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19360) );
  INV_X1 U22432 ( .A(n19360), .ZN(n19362) );
  NOR2_X1 U22433 ( .A1(n19890), .A2(n19362), .ZN(n19379) );
  AOI22_X1 U22434 ( .A1(n19387), .A2(n19732), .B1(n19379), .B2(n19724), .ZN(
        n19365) );
  OAI21_X1 U22435 ( .B1(n19608), .B2(n19420), .A(n19852), .ZN(n19363) );
  INV_X1 U22436 ( .A(n19379), .ZN(n19357) );
  OAI211_X1 U22437 ( .C1(n19358), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19357), 
        .B(n19581), .ZN(n19359) );
  OAI211_X1 U22438 ( .C1(n19363), .C2(n19360), .A(n19621), .B(n19359), .ZN(
        n19382) );
  OAI21_X1 U22439 ( .B1(n10537), .B2(n19379), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19361) );
  OAI21_X1 U22440 ( .B1(n19363), .B2(n19362), .A(n19361), .ZN(n19381) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19382), .B1(
        n19725), .B2(n19381), .ZN(n19364) );
  OAI211_X1 U22442 ( .C1(n19735), .C2(n19378), .A(n19365), .B(n19364), .ZN(
        P2_U3088) );
  AOI22_X1 U22443 ( .A1(n19387), .A2(n19738), .B1(n19379), .B2(n19736), .ZN(
        n19367) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19382), .B1(
        n19737), .B2(n19381), .ZN(n19366) );
  OAI211_X1 U22445 ( .C1(n19741), .C2(n19378), .A(n19367), .B(n19366), .ZN(
        P2_U3089) );
  AOI22_X1 U22446 ( .A1(n19387), .A2(n19744), .B1(n19379), .B2(n19742), .ZN(
        n19369) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19382), .B1(
        n19743), .B2(n19381), .ZN(n19368) );
  OAI211_X1 U22448 ( .C1(n19747), .C2(n19378), .A(n19369), .B(n19368), .ZN(
        P2_U3090) );
  AOI22_X1 U22449 ( .A1(n19387), .A2(n19750), .B1(n19748), .B2(n19379), .ZN(
        n19371) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19382), .B1(
        n19749), .B2(n19381), .ZN(n19370) );
  OAI211_X1 U22451 ( .C1(n19753), .C2(n19378), .A(n19371), .B(n19370), .ZN(
        P2_U3091) );
  AOI22_X1 U22452 ( .A1(n19380), .A2(n19562), .B1(n19754), .B2(n19379), .ZN(
        n19373) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19382), .B1(
        n19755), .B2(n19381), .ZN(n19372) );
  OAI211_X1 U22454 ( .C1(n19696), .C2(n19413), .A(n19373), .B(n19372), .ZN(
        P2_U3092) );
  AOI22_X1 U22455 ( .A1(n19380), .A2(n19565), .B1(n19379), .B2(n19760), .ZN(
        n19375) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19382), .B1(
        n19761), .B2(n19381), .ZN(n19374) );
  OAI211_X1 U22457 ( .C1(n19701), .C2(n19413), .A(n19375), .B(n19374), .ZN(
        P2_U3093) );
  AOI22_X1 U22458 ( .A1(n19387), .A2(n19768), .B1(n19379), .B2(n19766), .ZN(
        n19377) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19382), .B1(
        n19767), .B2(n19381), .ZN(n19376) );
  OAI211_X1 U22460 ( .C1(n19771), .C2(n19378), .A(n19377), .B(n19376), .ZN(
        P2_U3094) );
  AOI22_X1 U22461 ( .A1(n19380), .A2(n9847), .B1(n19379), .B2(n19772), .ZN(
        n19384) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19382), .B1(
        n19774), .B2(n19381), .ZN(n19383) );
  OAI211_X1 U22463 ( .C1(n19712), .C2(n19413), .A(n19384), .B(n19383), .ZN(
        P2_U3095) );
  INV_X1 U22464 ( .A(n19415), .ZN(n19388) );
  NAND3_X1 U22465 ( .A1(n19389), .A2(n19668), .A3(n19388), .ZN(n19385) );
  NOR3_X2 U22466 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19719), .ZN(n19408) );
  NOR3_X1 U22467 ( .A1(n10488), .A2(n19408), .A3(n19723), .ZN(n19390) );
  AOI21_X1 U22468 ( .B1(n19723), .B2(n19385), .A(n19390), .ZN(n19409) );
  AOI22_X1 U22469 ( .A1(n19409), .A2(n19725), .B1(n19724), .B2(n19408), .ZN(
        n19395) );
  OAI21_X1 U22470 ( .B1(n19387), .B2(n19440), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19392) );
  NAND2_X1 U22471 ( .A1(n19389), .A2(n19388), .ZN(n19391) );
  AOI211_X1 U22472 ( .C1(n19392), .C2(n19391), .A(n19730), .B(n19390), .ZN(
        n19393) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19732), .ZN(n19394) );
  OAI211_X1 U22474 ( .C1(n19735), .C2(n19413), .A(n19395), .B(n19394), .ZN(
        P2_U3096) );
  AOI22_X1 U22475 ( .A1(n19409), .A2(n19737), .B1(n19736), .B2(n19408), .ZN(
        n19397) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19738), .ZN(n19396) );
  OAI211_X1 U22477 ( .C1(n19741), .C2(n19413), .A(n19397), .B(n19396), .ZN(
        P2_U3097) );
  AOI22_X1 U22478 ( .A1(n19409), .A2(n19743), .B1(n19742), .B2(n19408), .ZN(
        n19399) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19744), .ZN(n19398) );
  OAI211_X1 U22480 ( .C1(n19747), .C2(n19413), .A(n19399), .B(n19398), .ZN(
        P2_U3098) );
  AOI22_X1 U22481 ( .A1(n19409), .A2(n19749), .B1(n19748), .B2(n19408), .ZN(
        n19401) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19750), .ZN(n19400) );
  OAI211_X1 U22483 ( .C1(n19753), .C2(n19413), .A(n19401), .B(n19400), .ZN(
        P2_U3099) );
  AOI22_X1 U22484 ( .A1(n19409), .A2(n19755), .B1(n19754), .B2(n19408), .ZN(
        n19403) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19756), .ZN(n19402) );
  OAI211_X1 U22486 ( .C1(n19759), .C2(n19413), .A(n19403), .B(n19402), .ZN(
        P2_U3100) );
  AOI22_X1 U22487 ( .A1(n19409), .A2(n19761), .B1(n19760), .B2(n19408), .ZN(
        n19405) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19762), .ZN(n19404) );
  OAI211_X1 U22489 ( .C1(n19765), .C2(n19413), .A(n19405), .B(n19404), .ZN(
        P2_U3101) );
  AOI22_X1 U22490 ( .A1(n19409), .A2(n19767), .B1(n19766), .B2(n19408), .ZN(
        n19407) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19768), .ZN(n19406) );
  OAI211_X1 U22492 ( .C1(n19771), .C2(n19413), .A(n19407), .B(n19406), .ZN(
        P2_U3102) );
  AOI22_X1 U22493 ( .A1(n19409), .A2(n19774), .B1(n19772), .B2(n19408), .ZN(
        n19412) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19410), .B1(
        n19440), .B2(n19776), .ZN(n19411) );
  OAI211_X1 U22495 ( .C1(n9848), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P2_U3103) );
  NOR2_X1 U22496 ( .A1(n19719), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19424) );
  INV_X1 U22497 ( .A(n19424), .ZN(n19418) );
  NOR2_X1 U22498 ( .A1(n19547), .A2(n19415), .ZN(n19453) );
  OR2_X1 U22499 ( .A1(n19453), .A2(n19723), .ZN(n19416) );
  NOR2_X1 U22500 ( .A1(n10493), .A2(n19416), .ZN(n19422) );
  AOI211_X2 U22501 ( .C1(n19418), .C2(n19723), .A(n19417), .B(n19422), .ZN(
        n19439) );
  AOI22_X1 U22502 ( .A1(n19439), .A2(n19725), .B1(n19453), .B2(n19724), .ZN(
        n19426) );
  NOR2_X1 U22503 ( .A1(n19420), .A2(n19419), .ZN(n19853) );
  OAI21_X1 U22504 ( .B1(n19453), .B2(n19668), .A(n19621), .ZN(n19421) );
  NOR2_X1 U22505 ( .A1(n19422), .A2(n19421), .ZN(n19423) );
  OAI21_X1 U22506 ( .B1(n19424), .B2(n19853), .A(n19423), .ZN(n19441) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19623), .ZN(n19425) );
  OAI211_X1 U22508 ( .C1(n19679), .C2(n19478), .A(n19426), .B(n19425), .ZN(
        P2_U3104) );
  AOI22_X1 U22509 ( .A1(n19439), .A2(n19737), .B1(n19453), .B2(n19736), .ZN(
        n19428) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19554), .ZN(n19427) );
  OAI211_X1 U22511 ( .C1(n19684), .C2(n19478), .A(n19428), .B(n19427), .ZN(
        P2_U3105) );
  AOI22_X1 U22512 ( .A1(n19439), .A2(n19743), .B1(n19453), .B2(n19742), .ZN(
        n19430) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19632), .ZN(n19429) );
  OAI211_X1 U22514 ( .C1(n19686), .C2(n19478), .A(n19430), .B(n19429), .ZN(
        P2_U3106) );
  AOI22_X1 U22515 ( .A1(n19439), .A2(n19749), .B1(n19748), .B2(n19453), .ZN(
        n19432) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19559), .ZN(n19431) );
  OAI211_X1 U22517 ( .C1(n19691), .C2(n19478), .A(n19432), .B(n19431), .ZN(
        P2_U3107) );
  AOI22_X1 U22518 ( .A1(n19439), .A2(n19755), .B1(n19754), .B2(n19453), .ZN(
        n19434) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19562), .ZN(n19433) );
  OAI211_X1 U22520 ( .C1(n19696), .C2(n19478), .A(n19434), .B(n19433), .ZN(
        P2_U3108) );
  AOI22_X1 U22521 ( .A1(n19439), .A2(n19761), .B1(n19453), .B2(n19760), .ZN(
        n19436) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19565), .ZN(n19435) );
  OAI211_X1 U22523 ( .C1(n19701), .C2(n19478), .A(n19436), .B(n19435), .ZN(
        P2_U3109) );
  AOI22_X1 U22524 ( .A1(n19439), .A2(n19767), .B1(n19453), .B2(n19766), .ZN(
        n19438) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n19649), .ZN(n19437) );
  OAI211_X1 U22526 ( .C1(n19709), .C2(n19478), .A(n19438), .B(n19437), .ZN(
        P2_U3110) );
  AOI22_X1 U22527 ( .A1(n19439), .A2(n19774), .B1(n19453), .B2(n19772), .ZN(
        n19443) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19441), .B1(
        n19440), .B2(n9847), .ZN(n19442) );
  OAI211_X1 U22529 ( .C1(n19712), .C2(n19478), .A(n19443), .B(n19442), .ZN(
        P2_U3111) );
  INV_X1 U22530 ( .A(n19661), .ZN(n19446) );
  NAND2_X1 U22531 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19871), .ZN(
        n19546) );
  NOR2_X1 U22532 ( .A1(n19447), .A2(n19546), .ZN(n19473) );
  AOI22_X1 U22533 ( .A1(n19503), .A2(n19732), .B1(n19473), .B2(n19724), .ZN(
        n19458) );
  INV_X1 U22534 ( .A(n19478), .ZN(n19448) );
  OAI21_X1 U22535 ( .B1(n19503), .B2(n19448), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19449) );
  NAND2_X1 U22536 ( .A1(n19449), .A2(n19852), .ZN(n19456) );
  NOR2_X1 U22537 ( .A1(n19456), .A2(n19453), .ZN(n19450) );
  AOI211_X1 U22538 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19451), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19450), .ZN(n19452) );
  NOR2_X1 U22539 ( .A1(n19453), .A2(n19473), .ZN(n19455) );
  OAI21_X1 U22540 ( .B1(n9699), .B2(n19473), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19454) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19475), .B1(
        n19725), .B2(n19474), .ZN(n19457) );
  OAI211_X1 U22542 ( .C1(n19735), .C2(n19478), .A(n19458), .B(n19457), .ZN(
        P2_U3112) );
  AOI22_X1 U22543 ( .A1(n19503), .A2(n19738), .B1(n19473), .B2(n19736), .ZN(
        n19460) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19475), .B1(
        n19737), .B2(n19474), .ZN(n19459) );
  OAI211_X1 U22545 ( .C1(n19741), .C2(n19478), .A(n19460), .B(n19459), .ZN(
        P2_U3113) );
  AOI22_X1 U22546 ( .A1(n19503), .A2(n19744), .B1(n19473), .B2(n19742), .ZN(
        n19462) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19475), .B1(
        n19743), .B2(n19474), .ZN(n19461) );
  OAI211_X1 U22548 ( .C1(n19747), .C2(n19478), .A(n19462), .B(n19461), .ZN(
        P2_U3114) );
  AOI22_X1 U22549 ( .A1(n19503), .A2(n19750), .B1(n19748), .B2(n19473), .ZN(
        n19464) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19475), .B1(
        n19749), .B2(n19474), .ZN(n19463) );
  OAI211_X1 U22551 ( .C1(n19753), .C2(n19478), .A(n19464), .B(n19463), .ZN(
        P2_U3115) );
  AOI22_X1 U22552 ( .A1(n19503), .A2(n19756), .B1(n19754), .B2(n19473), .ZN(
        n19466) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19475), .B1(
        n19755), .B2(n19474), .ZN(n19465) );
  OAI211_X1 U22554 ( .C1(n19759), .C2(n19478), .A(n19466), .B(n19465), .ZN(
        P2_U3116) );
  INV_X1 U22555 ( .A(n19473), .ZN(n19467) );
  OAI22_X1 U22556 ( .A1(n19478), .A2(n19765), .B1(n19700), .B2(n19467), .ZN(
        n19468) );
  INV_X1 U22557 ( .A(n19468), .ZN(n19470) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19475), .B1(
        n19761), .B2(n19474), .ZN(n19469) );
  OAI211_X1 U22559 ( .C1(n19701), .C2(n19511), .A(n19470), .B(n19469), .ZN(
        P2_U3117) );
  AOI22_X1 U22560 ( .A1(n19503), .A2(n19768), .B1(n19473), .B2(n19766), .ZN(
        n19472) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19475), .B1(
        n19767), .B2(n19474), .ZN(n19471) );
  OAI211_X1 U22562 ( .C1(n19771), .C2(n19478), .A(n19472), .B(n19471), .ZN(
        P2_U3118) );
  AOI22_X1 U22563 ( .A1(n19503), .A2(n19776), .B1(n19772), .B2(n19473), .ZN(
        n19477) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19475), .B1(
        n19774), .B2(n19474), .ZN(n19476) );
  OAI211_X1 U22565 ( .C1(n9848), .C2(n19478), .A(n19477), .B(n19476), .ZN(
        P2_U3119) );
  NOR2_X1 U22566 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19546), .ZN(
        n19482) );
  NAND2_X1 U22567 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19482), .ZN(
        n19512) );
  INV_X1 U22568 ( .A(n19512), .ZN(n19502) );
  AOI22_X1 U22569 ( .A1(n19503), .A2(n19623), .B1(n19724), .B2(n19502), .ZN(
        n19487) );
  NAND2_X1 U22570 ( .A1(n19857), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19615) );
  OAI21_X1 U22571 ( .B1(n19615), .B2(n19479), .A(n19852), .ZN(n19485) );
  OAI211_X1 U22572 ( .C1(n19480), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19512), 
        .B(n19581), .ZN(n19481) );
  OAI211_X1 U22573 ( .C1(n19485), .C2(n19482), .A(n19621), .B(n19481), .ZN(
        n19508) );
  INV_X1 U22574 ( .A(n19482), .ZN(n19484) );
  OAI21_X1 U22575 ( .B1(n10489), .B2(n19502), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19483) );
  OAI21_X1 U22576 ( .B1(n19485), .B2(n19484), .A(n19483), .ZN(n19507) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19508), .B1(
        n19725), .B2(n19507), .ZN(n19486) );
  OAI211_X1 U22578 ( .C1(n19679), .C2(n19544), .A(n19487), .B(n19486), .ZN(
        P2_U3120) );
  OAI22_X1 U22579 ( .A1(n19544), .A2(n19684), .B1(n19680), .B2(n19512), .ZN(
        n19488) );
  INV_X1 U22580 ( .A(n19488), .ZN(n19490) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19508), .B1(
        n19737), .B2(n19507), .ZN(n19489) );
  OAI211_X1 U22582 ( .C1(n19741), .C2(n19511), .A(n19490), .B(n19489), .ZN(
        P2_U3121) );
  OAI22_X1 U22583 ( .A1(n19544), .A2(n19686), .B1(n19685), .B2(n19512), .ZN(
        n19491) );
  INV_X1 U22584 ( .A(n19491), .ZN(n19493) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19508), .B1(
        n19743), .B2(n19507), .ZN(n19492) );
  OAI211_X1 U22586 ( .C1(n19747), .C2(n19511), .A(n19493), .B(n19492), .ZN(
        P2_U3122) );
  OAI22_X1 U22587 ( .A1(n19544), .A2(n19691), .B1(n19690), .B2(n19512), .ZN(
        n19494) );
  INV_X1 U22588 ( .A(n19494), .ZN(n19496) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19508), .B1(
        n19749), .B2(n19507), .ZN(n19495) );
  OAI211_X1 U22590 ( .C1(n19753), .C2(n19511), .A(n19496), .B(n19495), .ZN(
        P2_U3123) );
  AOI22_X1 U22591 ( .A1(n19503), .A2(n19562), .B1(n19754), .B2(n19502), .ZN(
        n19498) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19508), .B1(
        n19755), .B2(n19507), .ZN(n19497) );
  OAI211_X1 U22593 ( .C1(n19696), .C2(n19544), .A(n19498), .B(n19497), .ZN(
        P2_U3124) );
  OAI22_X1 U22594 ( .A1(n19544), .A2(n19701), .B1(n19700), .B2(n19512), .ZN(
        n19499) );
  INV_X1 U22595 ( .A(n19499), .ZN(n19501) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19508), .B1(
        n19761), .B2(n19507), .ZN(n19500) );
  OAI211_X1 U22597 ( .C1(n19765), .C2(n19511), .A(n19501), .B(n19500), .ZN(
        P2_U3125) );
  AOI22_X1 U22598 ( .A1(n19503), .A2(n19649), .B1(n19766), .B2(n19502), .ZN(
        n19505) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19508), .B1(
        n19767), .B2(n19507), .ZN(n19504) );
  OAI211_X1 U22600 ( .C1(n19709), .C2(n19544), .A(n19505), .B(n19504), .ZN(
        P2_U3126) );
  OAI22_X1 U22601 ( .A1(n19544), .A2(n19712), .B1(n19711), .B2(n19512), .ZN(
        n19506) );
  INV_X1 U22602 ( .A(n19506), .ZN(n19510) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19508), .B1(
        n19774), .B2(n19507), .ZN(n19509) );
  OAI211_X1 U22604 ( .C1(n9848), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P2_U3127) );
  NAND2_X1 U22605 ( .A1(n19661), .A2(n19868), .ZN(n19536) );
  OAI221_X1 U22606 ( .B1(n19666), .B2(n19536), .C1(n19666), .C2(n19544), .A(
        n19512), .ZN(n19515) );
  OAI21_X1 U22607 ( .B1(n19513), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19581), 
        .ZN(n19514) );
  NAND2_X1 U22608 ( .A1(n19515), .A2(n19514), .ZN(n19517) );
  NOR2_X1 U22609 ( .A1(n19881), .A2(n19546), .ZN(n19549) );
  INV_X1 U22610 ( .A(n19549), .ZN(n19545) );
  NOR2_X1 U22611 ( .A1(n19545), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19539) );
  INV_X1 U22612 ( .A(n19539), .ZN(n19516) );
  NAND2_X1 U22613 ( .A1(n19517), .A2(n19516), .ZN(n19518) );
  OAI21_X1 U22614 ( .B1(n9701), .B2(n19539), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19519) );
  AOI22_X1 U22615 ( .A1(n19540), .A2(n19725), .B1(n19724), .B2(n19539), .ZN(
        n19522) );
  INV_X1 U22616 ( .A(n19544), .ZN(n19533) );
  AOI22_X1 U22617 ( .A1(n19572), .A2(n19732), .B1(n19533), .B2(n19623), .ZN(
        n19521) );
  OAI211_X1 U22618 ( .C1(n19524), .C2(n19523), .A(n19522), .B(n19521), .ZN(
        P2_U3128) );
  AOI22_X1 U22619 ( .A1(n19540), .A2(n19737), .B1(n19736), .B2(n19539), .ZN(
        n19526) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19541), .B1(
        n19572), .B2(n19738), .ZN(n19525) );
  OAI211_X1 U22621 ( .C1(n19741), .C2(n19544), .A(n19526), .B(n19525), .ZN(
        P2_U3129) );
  AOI22_X1 U22622 ( .A1(n19540), .A2(n19743), .B1(n19742), .B2(n19539), .ZN(
        n19528) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19541), .B1(
        n19572), .B2(n19744), .ZN(n19527) );
  OAI211_X1 U22624 ( .C1(n19747), .C2(n19544), .A(n19528), .B(n19527), .ZN(
        P2_U3130) );
  AOI22_X1 U22625 ( .A1(n19540), .A2(n19749), .B1(n19748), .B2(n19539), .ZN(
        n19530) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19541), .B1(
        n19572), .B2(n19750), .ZN(n19529) );
  OAI211_X1 U22627 ( .C1(n19753), .C2(n19544), .A(n19530), .B(n19529), .ZN(
        P2_U3131) );
  AOI22_X1 U22628 ( .A1(n19540), .A2(n19755), .B1(n19754), .B2(n19539), .ZN(
        n19532) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19541), .B1(
        n19572), .B2(n19756), .ZN(n19531) );
  OAI211_X1 U22630 ( .C1(n19759), .C2(n19544), .A(n19532), .B(n19531), .ZN(
        P2_U3132) );
  AOI22_X1 U22631 ( .A1(n19540), .A2(n19761), .B1(n19760), .B2(n19539), .ZN(
        n19535) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19541), .B1(
        n19533), .B2(n19565), .ZN(n19534) );
  OAI211_X1 U22633 ( .C1(n19701), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P2_U3133) );
  AOI22_X1 U22634 ( .A1(n19540), .A2(n19767), .B1(n19766), .B2(n19539), .ZN(
        n19538) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19541), .B1(
        n19572), .B2(n19768), .ZN(n19537) );
  OAI211_X1 U22636 ( .C1(n19771), .C2(n19544), .A(n19538), .B(n19537), .ZN(
        P2_U3134) );
  AOI22_X1 U22637 ( .A1(n19540), .A2(n19774), .B1(n19772), .B2(n19539), .ZN(
        n19543) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19541), .B1(
        n19572), .B2(n19776), .ZN(n19542) );
  OAI211_X1 U22639 ( .C1(n9848), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        P2_U3135) );
  OR2_X1 U22640 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19545), .ZN(n19548) );
  NOR2_X1 U22641 ( .A1(n19547), .A2(n19546), .ZN(n19570) );
  NOR3_X1 U22642 ( .A1(n10491), .A2(n19570), .A3(n19723), .ZN(n19550) );
  AOI21_X1 U22643 ( .B1(n19723), .B2(n19548), .A(n19550), .ZN(n19571) );
  AOI22_X1 U22644 ( .A1(n19571), .A2(n19725), .B1(n19724), .B2(n19570), .ZN(
        n19553) );
  NOR2_X1 U22645 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19615), .ZN(n19727) );
  AOI22_X1 U22646 ( .A1(n19868), .A2(n19727), .B1(n19882), .B2(n19549), .ZN(
        n19551) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19623), .ZN(n19552) );
  OAI211_X1 U22648 ( .C1(n19679), .C2(n19607), .A(n19553), .B(n19552), .ZN(
        P2_U3136) );
  AOI22_X1 U22649 ( .A1(n19571), .A2(n19737), .B1(n19736), .B2(n19570), .ZN(
        n19556) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19554), .ZN(n19555) );
  OAI211_X1 U22651 ( .C1(n19684), .C2(n19607), .A(n19556), .B(n19555), .ZN(
        P2_U3137) );
  AOI22_X1 U22652 ( .A1(n19571), .A2(n19743), .B1(n19742), .B2(n19570), .ZN(
        n19558) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19632), .ZN(n19557) );
  OAI211_X1 U22654 ( .C1(n19686), .C2(n19607), .A(n19558), .B(n19557), .ZN(
        P2_U3138) );
  AOI22_X1 U22655 ( .A1(n19571), .A2(n19749), .B1(n19748), .B2(n19570), .ZN(
        n19561) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19559), .ZN(n19560) );
  OAI211_X1 U22657 ( .C1(n19691), .C2(n19607), .A(n19561), .B(n19560), .ZN(
        P2_U3139) );
  AOI22_X1 U22658 ( .A1(n19571), .A2(n19755), .B1(n19754), .B2(n19570), .ZN(
        n19564) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19562), .ZN(n19563) );
  OAI211_X1 U22660 ( .C1(n19696), .C2(n19607), .A(n19564), .B(n19563), .ZN(
        P2_U3140) );
  AOI22_X1 U22661 ( .A1(n19571), .A2(n19761), .B1(n19760), .B2(n19570), .ZN(
        n19567) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19565), .ZN(n19566) );
  OAI211_X1 U22663 ( .C1(n19701), .C2(n19607), .A(n19567), .B(n19566), .ZN(
        P2_U3141) );
  AOI22_X1 U22664 ( .A1(n19571), .A2(n19767), .B1(n19766), .B2(n19570), .ZN(
        n19569) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19649), .ZN(n19568) );
  OAI211_X1 U22666 ( .C1(n19709), .C2(n19607), .A(n19569), .B(n19568), .ZN(
        P2_U3142) );
  AOI22_X1 U22667 ( .A1(n19571), .A2(n19774), .B1(n19772), .B2(n19570), .ZN(
        n19575) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n9847), .ZN(n19574) );
  OAI211_X1 U22669 ( .C1(n19712), .C2(n19607), .A(n19575), .B(n19574), .ZN(
        P2_U3143) );
  INV_X1 U22670 ( .A(n19576), .ZN(n19579) );
  INV_X1 U22671 ( .A(n19586), .ZN(n19578) );
  NAND3_X1 U22672 ( .A1(n19881), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19619) );
  NOR2_X1 U22673 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19619), .ZN(
        n19602) );
  OAI21_X1 U22674 ( .B1(n19580), .B2(n19602), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19577) );
  AOI22_X1 U22675 ( .A1(n19603), .A2(n19725), .B1(n19724), .B2(n19602), .ZN(
        n19589) );
  NAND2_X1 U22676 ( .A1(n19661), .A2(n19616), .ZN(n19660) );
  AOI21_X1 U22677 ( .B1(n19607), .B2(n19660), .A(n19666), .ZN(n19587) );
  INV_X1 U22678 ( .A(n19580), .ZN(n19583) );
  INV_X1 U22679 ( .A(n19602), .ZN(n19582) );
  OAI211_X1 U22680 ( .C1(n19583), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19582), 
        .B(n19581), .ZN(n19584) );
  AND2_X1 U22681 ( .A1(n19584), .A2(n19621), .ZN(n19585) );
  OAI211_X1 U22682 ( .C1(n19587), .C2(n19586), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19585), .ZN(n19604) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19732), .ZN(n19588) );
  OAI211_X1 U22684 ( .C1(n19735), .C2(n19607), .A(n19589), .B(n19588), .ZN(
        P2_U3144) );
  AOI22_X1 U22685 ( .A1(n19603), .A2(n19737), .B1(n19736), .B2(n19602), .ZN(
        n19591) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19738), .ZN(n19590) );
  OAI211_X1 U22687 ( .C1(n19741), .C2(n19607), .A(n19591), .B(n19590), .ZN(
        P2_U3145) );
  AOI22_X1 U22688 ( .A1(n19603), .A2(n19743), .B1(n19742), .B2(n19602), .ZN(
        n19593) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19744), .ZN(n19592) );
  OAI211_X1 U22690 ( .C1(n19747), .C2(n19607), .A(n19593), .B(n19592), .ZN(
        P2_U3146) );
  AOI22_X1 U22691 ( .A1(n19603), .A2(n19749), .B1(n19748), .B2(n19602), .ZN(
        n19595) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19750), .ZN(n19594) );
  OAI211_X1 U22693 ( .C1(n19753), .C2(n19607), .A(n19595), .B(n19594), .ZN(
        P2_U3147) );
  AOI22_X1 U22694 ( .A1(n19603), .A2(n19755), .B1(n19754), .B2(n19602), .ZN(
        n19597) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19756), .ZN(n19596) );
  OAI211_X1 U22696 ( .C1(n19759), .C2(n19607), .A(n19597), .B(n19596), .ZN(
        P2_U3148) );
  AOI22_X1 U22697 ( .A1(n19603), .A2(n19761), .B1(n19760), .B2(n19602), .ZN(
        n19599) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19762), .ZN(n19598) );
  OAI211_X1 U22699 ( .C1(n19765), .C2(n19607), .A(n19599), .B(n19598), .ZN(
        P2_U3149) );
  AOI22_X1 U22700 ( .A1(n19603), .A2(n19767), .B1(n19766), .B2(n19602), .ZN(
        n19601) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19768), .ZN(n19600) );
  OAI211_X1 U22702 ( .C1(n19771), .C2(n19607), .A(n19601), .B(n19600), .ZN(
        P2_U3150) );
  AOI22_X1 U22703 ( .A1(n19603), .A2(n19774), .B1(n19772), .B2(n19602), .ZN(
        n19606) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19604), .B1(
        n19650), .B2(n19776), .ZN(n19605) );
  OAI211_X1 U22705 ( .C1(n9848), .C2(n19607), .A(n19606), .B(n19605), .ZN(
        P2_U3151) );
  NOR2_X1 U22706 ( .A1(n19890), .A2(n19619), .ZN(n19671) );
  INV_X1 U22707 ( .A(n19671), .ZN(n19653) );
  NAND2_X1 U22708 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19653), .ZN(n19610) );
  NOR2_X1 U22709 ( .A1(n10480), .A2(n19610), .ZN(n19618) );
  INV_X1 U22710 ( .A(n19619), .ZN(n19611) );
  AOI21_X1 U22711 ( .B1(n19668), .B2(n19611), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19612) );
  OAI22_X1 U22712 ( .A1(n19655), .A2(n19613), .B1(n19662), .B2(n19653), .ZN(
        n19614) );
  INV_X1 U22713 ( .A(n19614), .ZN(n19625) );
  INV_X1 U22714 ( .A(n19615), .ZN(n19617) );
  NAND2_X1 U22715 ( .A1(n19617), .A2(n19616), .ZN(n19620) );
  AOI21_X1 U22716 ( .B1(n19620), .B2(n19619), .A(n19618), .ZN(n19622) );
  OAI211_X1 U22717 ( .C1(n19671), .C2(n19668), .A(n19622), .B(n19621), .ZN(
        n19657) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19657), .B1(
        n19650), .B2(n19623), .ZN(n19624) );
  OAI211_X1 U22719 ( .C1(n19679), .C2(n19718), .A(n19625), .B(n19624), .ZN(
        P2_U3152) );
  OAI22_X1 U22720 ( .A1(n19655), .A2(n19626), .B1(n19680), .B2(n19653), .ZN(
        n19627) );
  INV_X1 U22721 ( .A(n19627), .ZN(n19629) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19657), .B1(
        n19664), .B2(n19738), .ZN(n19628) );
  OAI211_X1 U22723 ( .C1(n19741), .C2(n19660), .A(n19629), .B(n19628), .ZN(
        P2_U3153) );
  OAI22_X1 U22724 ( .A1(n19655), .A2(n19630), .B1(n19685), .B2(n19653), .ZN(
        n19631) );
  INV_X1 U22725 ( .A(n19631), .ZN(n19634) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19657), .B1(
        n19650), .B2(n19632), .ZN(n19633) );
  OAI211_X1 U22727 ( .C1(n19686), .C2(n19718), .A(n19634), .B(n19633), .ZN(
        P2_U3154) );
  OAI22_X1 U22728 ( .A1(n19655), .A2(n19635), .B1(n19690), .B2(n19653), .ZN(
        n19636) );
  INV_X1 U22729 ( .A(n19636), .ZN(n19638) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19657), .B1(
        n19664), .B2(n19750), .ZN(n19637) );
  OAI211_X1 U22731 ( .C1(n19753), .C2(n19660), .A(n19638), .B(n19637), .ZN(
        P2_U3155) );
  OAI22_X1 U22732 ( .A1(n19655), .A2(n19639), .B1(n19695), .B2(n19653), .ZN(
        n19640) );
  INV_X1 U22733 ( .A(n19640), .ZN(n19642) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19657), .B1(
        n19664), .B2(n19756), .ZN(n19641) );
  OAI211_X1 U22735 ( .C1(n19759), .C2(n19660), .A(n19642), .B(n19641), .ZN(
        P2_U3156) );
  OAI22_X1 U22736 ( .A1(n19655), .A2(n19643), .B1(n19700), .B2(n19653), .ZN(
        n19644) );
  INV_X1 U22737 ( .A(n19644), .ZN(n19646) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19657), .B1(
        n19664), .B2(n19762), .ZN(n19645) );
  OAI211_X1 U22739 ( .C1(n19765), .C2(n19660), .A(n19646), .B(n19645), .ZN(
        P2_U3157) );
  OAI22_X1 U22740 ( .A1(n19655), .A2(n19647), .B1(n19705), .B2(n19653), .ZN(
        n19648) );
  INV_X1 U22741 ( .A(n19648), .ZN(n19652) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19657), .B1(
        n19650), .B2(n19649), .ZN(n19651) );
  OAI211_X1 U22743 ( .C1(n19709), .C2(n19718), .A(n19652), .B(n19651), .ZN(
        P2_U3158) );
  OAI22_X1 U22744 ( .A1(n19655), .A2(n19654), .B1(n19711), .B2(n19653), .ZN(
        n19656) );
  INV_X1 U22745 ( .A(n19656), .ZN(n19659) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19657), .B1(
        n19664), .B2(n19776), .ZN(n19658) );
  OAI211_X1 U22747 ( .C1(n9848), .C2(n19660), .A(n19659), .B(n19658), .ZN(
        P2_U3159) );
  NOR3_X1 U22748 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19864), .A3(
        n19719), .ZN(n19672) );
  INV_X1 U22749 ( .A(n19672), .ZN(n19710) );
  OAI22_X1 U22750 ( .A1(n19718), .A2(n19735), .B1(n19662), .B2(n19710), .ZN(
        n19663) );
  INV_X1 U22751 ( .A(n19663), .ZN(n19678) );
  NOR3_X1 U22752 ( .A1(n19673), .A2(n19672), .A3(n19723), .ZN(n19670) );
  INV_X1 U22753 ( .A(n19781), .ZN(n19665) );
  NOR2_X1 U22754 ( .A1(n19665), .A2(n19664), .ZN(n19667) );
  OAI21_X1 U22755 ( .B1(n19667), .B2(n19666), .A(n19852), .ZN(n19676) );
  AOI221_X1 U22756 ( .B1(n19668), .B2(n19676), .C1(n19668), .C2(n19671), .A(
        n19672), .ZN(n19669) );
  NOR2_X1 U22757 ( .A1(n19672), .A2(n19671), .ZN(n19675) );
  OAI21_X1 U22758 ( .B1(n19673), .B2(n19672), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19674) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19715), .B1(
        n19725), .B2(n19714), .ZN(n19677) );
  OAI211_X1 U22760 ( .C1(n19679), .C2(n19781), .A(n19678), .B(n19677), .ZN(
        P2_U3160) );
  OAI22_X1 U22761 ( .A1(n19718), .A2(n19741), .B1(n19680), .B2(n19710), .ZN(
        n19681) );
  INV_X1 U22762 ( .A(n19681), .ZN(n19683) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19715), .B1(
        n19737), .B2(n19714), .ZN(n19682) );
  OAI211_X1 U22764 ( .C1(n19684), .C2(n19781), .A(n19683), .B(n19682), .ZN(
        P2_U3161) );
  OAI22_X1 U22765 ( .A1(n19781), .A2(n19686), .B1(n19685), .B2(n19710), .ZN(
        n19687) );
  INV_X1 U22766 ( .A(n19687), .ZN(n19689) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19715), .B1(
        n19743), .B2(n19714), .ZN(n19688) );
  OAI211_X1 U22768 ( .C1(n19747), .C2(n19718), .A(n19689), .B(n19688), .ZN(
        P2_U3162) );
  OAI22_X1 U22769 ( .A1(n19781), .A2(n19691), .B1(n19690), .B2(n19710), .ZN(
        n19692) );
  INV_X1 U22770 ( .A(n19692), .ZN(n19694) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19715), .B1(
        n19749), .B2(n19714), .ZN(n19693) );
  OAI211_X1 U22772 ( .C1(n19753), .C2(n19718), .A(n19694), .B(n19693), .ZN(
        P2_U3163) );
  OAI22_X1 U22773 ( .A1(n19781), .A2(n19696), .B1(n19695), .B2(n19710), .ZN(
        n19697) );
  INV_X1 U22774 ( .A(n19697), .ZN(n19699) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19715), .B1(
        n19755), .B2(n19714), .ZN(n19698) );
  OAI211_X1 U22776 ( .C1(n19759), .C2(n19718), .A(n19699), .B(n19698), .ZN(
        P2_U3164) );
  OAI22_X1 U22777 ( .A1(n19781), .A2(n19701), .B1(n19700), .B2(n19710), .ZN(
        n19702) );
  INV_X1 U22778 ( .A(n19702), .ZN(n19704) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19715), .B1(
        n19761), .B2(n19714), .ZN(n19703) );
  OAI211_X1 U22780 ( .C1(n19765), .C2(n19718), .A(n19704), .B(n19703), .ZN(
        P2_U3165) );
  OAI22_X1 U22781 ( .A1(n19718), .A2(n19771), .B1(n19705), .B2(n19710), .ZN(
        n19706) );
  INV_X1 U22782 ( .A(n19706), .ZN(n19708) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19715), .B1(
        n19767), .B2(n19714), .ZN(n19707) );
  OAI211_X1 U22784 ( .C1(n19709), .C2(n19781), .A(n19708), .B(n19707), .ZN(
        P2_U3166) );
  OAI22_X1 U22785 ( .A1(n19781), .A2(n19712), .B1(n19711), .B2(n19710), .ZN(
        n19713) );
  INV_X1 U22786 ( .A(n19713), .ZN(n19717) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19715), .B1(
        n19774), .B2(n19714), .ZN(n19716) );
  OAI211_X1 U22788 ( .C1(n9848), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3167) );
  NOR2_X1 U22789 ( .A1(n19864), .A2(n19719), .ZN(n19726) );
  INV_X1 U22790 ( .A(n19726), .ZN(n19720) );
  OR2_X1 U22791 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19720), .ZN(n19722) );
  INV_X1 U22792 ( .A(n19721), .ZN(n19773) );
  NOR3_X1 U22793 ( .A1(n10482), .A2(n19773), .A3(n19723), .ZN(n19729) );
  AOI21_X1 U22794 ( .B1(n19723), .B2(n19722), .A(n19729), .ZN(n19775) );
  AOI22_X1 U22795 ( .A1(n19775), .A2(n19725), .B1(n19773), .B2(n19724), .ZN(
        n19734) );
  AOI22_X1 U22796 ( .A1(n19728), .A2(n19727), .B1(n19882), .B2(n19726), .ZN(
        n19731) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19732), .ZN(n19733) );
  OAI211_X1 U22798 ( .C1(n19735), .C2(n19781), .A(n19734), .B(n19733), .ZN(
        P2_U3168) );
  AOI22_X1 U22799 ( .A1(n19775), .A2(n19737), .B1(n19773), .B2(n19736), .ZN(
        n19740) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19738), .ZN(n19739) );
  OAI211_X1 U22801 ( .C1(n19741), .C2(n19781), .A(n19740), .B(n19739), .ZN(
        P2_U3169) );
  AOI22_X1 U22802 ( .A1(n19775), .A2(n19743), .B1(n19773), .B2(n19742), .ZN(
        n19746) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19744), .ZN(n19745) );
  OAI211_X1 U22804 ( .C1(n19747), .C2(n19781), .A(n19746), .B(n19745), .ZN(
        P2_U3170) );
  AOI22_X1 U22805 ( .A1(n19775), .A2(n19749), .B1(n19773), .B2(n19748), .ZN(
        n19752) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19750), .ZN(n19751) );
  OAI211_X1 U22807 ( .C1(n19753), .C2(n19781), .A(n19752), .B(n19751), .ZN(
        P2_U3171) );
  AOI22_X1 U22808 ( .A1(n19775), .A2(n19755), .B1(n19773), .B2(n19754), .ZN(
        n19758) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19756), .ZN(n19757) );
  OAI211_X1 U22810 ( .C1(n19759), .C2(n19781), .A(n19758), .B(n19757), .ZN(
        P2_U3172) );
  AOI22_X1 U22811 ( .A1(n19775), .A2(n19761), .B1(n19773), .B2(n19760), .ZN(
        n19764) );
  AOI22_X1 U22812 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19762), .ZN(n19763) );
  OAI211_X1 U22813 ( .C1(n19765), .C2(n19781), .A(n19764), .B(n19763), .ZN(
        P2_U3173) );
  AOI22_X1 U22814 ( .A1(n19775), .A2(n19767), .B1(n19773), .B2(n19766), .ZN(
        n19770) );
  AOI22_X1 U22815 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19768), .ZN(n19769) );
  OAI211_X1 U22816 ( .C1(n19771), .C2(n19781), .A(n19770), .B(n19769), .ZN(
        P2_U3174) );
  AOI22_X1 U22817 ( .A1(n19775), .A2(n19774), .B1(n19773), .B2(n19772), .ZN(
        n19780) );
  AOI22_X1 U22818 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19778), .B1(
        n19777), .B2(n19776), .ZN(n19779) );
  OAI211_X1 U22819 ( .C1(n9848), .C2(n19781), .A(n19780), .B(n19779), .ZN(
        P2_U3175) );
  AND2_X1 U22820 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19783), .ZN(
        P2_U3179) );
  AND2_X1 U22821 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19783), .ZN(
        P2_U3180) );
  AND2_X1 U22822 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19783), .ZN(
        P2_U3181) );
  NOR2_X1 U22823 ( .A1(n20809), .A2(n19851), .ZN(P2_U3182) );
  AND2_X1 U22824 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19783), .ZN(
        P2_U3183) );
  AND2_X1 U22825 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19783), .ZN(
        P2_U3184) );
  AND2_X1 U22826 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19783), .ZN(
        P2_U3185) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19783), .ZN(
        P2_U3186) );
  AND2_X1 U22828 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19783), .ZN(
        P2_U3187) );
  AND2_X1 U22829 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19783), .ZN(
        P2_U3188) );
  AND2_X1 U22830 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19783), .ZN(
        P2_U3189) );
  INV_X1 U22831 ( .A(P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(n20818) );
  NOR2_X1 U22832 ( .A1(n20818), .A2(n19851), .ZN(P2_U3190) );
  AND2_X1 U22833 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19783), .ZN(
        P2_U3191) );
  AND2_X1 U22834 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19783), .ZN(
        P2_U3192) );
  AND2_X1 U22835 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19783), .ZN(
        P2_U3193) );
  AND2_X1 U22836 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19783), .ZN(
        P2_U3194) );
  AND2_X1 U22837 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19783), .ZN(
        P2_U3195) );
  AND2_X1 U22838 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19783), .ZN(
        P2_U3196) );
  AND2_X1 U22839 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19783), .ZN(
        P2_U3197) );
  AND2_X1 U22840 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19783), .ZN(
        P2_U3198) );
  AND2_X1 U22841 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19783), .ZN(
        P2_U3199) );
  AND2_X1 U22842 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19783), .ZN(
        P2_U3200) );
  AND2_X1 U22843 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19783), .ZN(P2_U3201) );
  AND2_X1 U22844 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19783), .ZN(P2_U3202) );
  AND2_X1 U22845 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19783), .ZN(P2_U3203) );
  AND2_X1 U22846 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19783), .ZN(P2_U3204) );
  AND2_X1 U22847 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19783), .ZN(P2_U3205) );
  NOR2_X1 U22848 ( .A1(n20713), .A2(n19851), .ZN(P2_U3206) );
  AND2_X1 U22849 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19783), .ZN(P2_U3207) );
  AND2_X1 U22850 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19783), .ZN(P2_U3208) );
  NAND2_X1 U22851 ( .A1(n19793), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19796) );
  NAND3_X1 U22852 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19796), .ZN(n19785) );
  AOI211_X1 U22853 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20594), .A(
        n19795), .B(n19901), .ZN(n19784) );
  INV_X1 U22854 ( .A(NA), .ZN(n20598) );
  NOR3_X1 U22855 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .A3(n20598), .ZN(n19801) );
  AOI211_X1 U22856 ( .C1(n19802), .C2(n19785), .A(n19784), .B(n19801), .ZN(
        n19786) );
  INV_X1 U22857 ( .A(n19786), .ZN(P2_U3209) );
  AOI21_X1 U22858 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20594), .A(n19802), 
        .ZN(n19792) );
  NOR2_X1 U22859 ( .A1(n18860), .A2(n19792), .ZN(n19788) );
  AOI21_X1 U22860 ( .B1(n19788), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n19787), .ZN(n19789) );
  OAI211_X1 U22861 ( .C1(n20594), .C2(n19790), .A(n19789), .B(n19796), .ZN(
        P2_U3210) );
  NOR2_X1 U22862 ( .A1(n19802), .A2(n19791), .ZN(n19794) );
  AOI21_X1 U22863 ( .B1(n19794), .B2(n19793), .A(n19792), .ZN(n19800) );
  INV_X1 U22864 ( .A(n19795), .ZN(n19797) );
  OAI22_X1 U22865 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19797), .B1(NA), 
        .B2(n19796), .ZN(n19798) );
  OAI211_X1 U22866 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19798), .ZN(n19799) );
  OAI21_X1 U22867 ( .B1(n19801), .B2(n19800), .A(n19799), .ZN(P2_U3211) );
  OAI222_X1 U22868 ( .A1(n19842), .A2(n20696), .B1(n20721), .B2(n19901), .C1(
        n12971), .C2(n19840), .ZN(P2_U3212) );
  OAI222_X1 U22869 ( .A1(n19842), .A2(n10289), .B1(n20821), .B2(n19901), .C1(
        n20696), .C2(n19840), .ZN(P2_U3213) );
  OAI222_X1 U22870 ( .A1(n19842), .A2(n12251), .B1(n19803), .B2(n19901), .C1(
        n10289), .C2(n19840), .ZN(P2_U3214) );
  OAI222_X1 U22871 ( .A1(n19842), .A2(n10731), .B1(n19804), .B2(n19901), .C1(
        n12251), .C2(n19840), .ZN(P2_U3215) );
  OAI222_X1 U22872 ( .A1(n19842), .A2(n10734), .B1(n19805), .B2(n19901), .C1(
        n10731), .C2(n19840), .ZN(P2_U3216) );
  OAI222_X1 U22873 ( .A1(n19842), .A2(n10739), .B1(n19806), .B2(n19901), .C1(
        n10734), .C2(n19840), .ZN(P2_U3217) );
  OAI222_X1 U22874 ( .A1(n19842), .A2(n13663), .B1(n19807), .B2(n19901), .C1(
        n10739), .C2(n19840), .ZN(P2_U3218) );
  OAI222_X1 U22875 ( .A1(n19842), .A2(n15329), .B1(n19808), .B2(n19901), .C1(
        n13663), .C2(n19840), .ZN(P2_U3219) );
  OAI222_X1 U22876 ( .A1(n19842), .A2(n12298), .B1(n19809), .B2(n19901), .C1(
        n15329), .C2(n19840), .ZN(P2_U3220) );
  OAI222_X1 U22877 ( .A1(n19842), .A2(n19811), .B1(n19810), .B2(n19901), .C1(
        n12298), .C2(n19840), .ZN(P2_U3221) );
  OAI222_X1 U22878 ( .A1(n19842), .A2(n10757), .B1(n19812), .B2(n19901), .C1(
        n19811), .C2(n19840), .ZN(P2_U3222) );
  OAI222_X1 U22879 ( .A1(n19842), .A2(n15298), .B1(n19813), .B2(n19901), .C1(
        n10757), .C2(n19840), .ZN(P2_U3223) );
  OAI222_X1 U22880 ( .A1(n19842), .A2(n19815), .B1(n19814), .B2(n19901), .C1(
        n15298), .C2(n19840), .ZN(P2_U3224) );
  OAI222_X1 U22881 ( .A1(n19842), .A2(n19817), .B1(n19816), .B2(n19901), .C1(
        n19815), .C2(n19840), .ZN(P2_U3225) );
  OAI222_X1 U22882 ( .A1(n19842), .A2(n14142), .B1(n20728), .B2(n19901), .C1(
        n19817), .C2(n19840), .ZN(P2_U3226) );
  OAI222_X1 U22883 ( .A1(n19842), .A2(n19819), .B1(n19818), .B2(n19901), .C1(
        n14142), .C2(n19840), .ZN(P2_U3227) );
  OAI222_X1 U22884 ( .A1(n19842), .A2(n15245), .B1(n19820), .B2(n19901), .C1(
        n19819), .C2(n19840), .ZN(P2_U3228) );
  OAI222_X1 U22885 ( .A1(n19842), .A2(n19822), .B1(n19821), .B2(n19901), .C1(
        n15245), .C2(n19840), .ZN(P2_U3229) );
  OAI222_X1 U22886 ( .A1(n19842), .A2(n19824), .B1(n19823), .B2(n19901), .C1(
        n19822), .C2(n19840), .ZN(P2_U3230) );
  OAI222_X1 U22887 ( .A1(n19842), .A2(n19826), .B1(n19825), .B2(n19901), .C1(
        n19824), .C2(n19840), .ZN(P2_U3231) );
  OAI222_X1 U22888 ( .A1(n19842), .A2(n10788), .B1(n19827), .B2(n19901), .C1(
        n19826), .C2(n19840), .ZN(P2_U3232) );
  OAI222_X1 U22889 ( .A1(n19842), .A2(n10792), .B1(n19828), .B2(n19901), .C1(
        n10788), .C2(n19840), .ZN(P2_U3233) );
  OAI222_X1 U22890 ( .A1(n19842), .A2(n15183), .B1(n19829), .B2(n19901), .C1(
        n10792), .C2(n19840), .ZN(P2_U3234) );
  OAI222_X1 U22891 ( .A1(n19842), .A2(n19831), .B1(n19830), .B2(n19901), .C1(
        n15183), .C2(n19840), .ZN(P2_U3235) );
  OAI222_X1 U22892 ( .A1(n19842), .A2(n19833), .B1(n19832), .B2(n19901), .C1(
        n19831), .C2(n19840), .ZN(P2_U3236) );
  OAI222_X1 U22893 ( .A1(n19842), .A2(n19836), .B1(n19834), .B2(n19901), .C1(
        n19833), .C2(n19840), .ZN(P2_U3237) );
  OAI222_X1 U22894 ( .A1(n19840), .A2(n19836), .B1(n19835), .B2(n19901), .C1(
        n15146), .C2(n19842), .ZN(P2_U3238) );
  OAI222_X1 U22895 ( .A1(n19842), .A2(n19838), .B1(n19837), .B2(n19901), .C1(
        n15146), .C2(n19840), .ZN(P2_U3239) );
  OAI222_X1 U22896 ( .A1(n19842), .A2(n15131), .B1(n19839), .B2(n19901), .C1(
        n19838), .C2(n19840), .ZN(P2_U3240) );
  OAI222_X1 U22897 ( .A1(n19842), .A2(n12842), .B1(n19841), .B2(n19901), .C1(
        n15131), .C2(n19840), .ZN(P2_U3241) );
  INV_X1 U22898 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19843) );
  AOI22_X1 U22899 ( .A1(n19901), .A2(n20839), .B1(n19843), .B2(n19898), .ZN(
        P2_U3585) );
  MUX2_X1 U22900 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19901), .Z(P2_U3586) );
  INV_X1 U22901 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U22902 ( .A1(n19901), .A2(n19845), .B1(n19844), .B2(n19898), .ZN(
        P2_U3587) );
  INV_X1 U22903 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U22904 ( .A1(n19901), .A2(n19847), .B1(n19846), .B2(n19898), .ZN(
        P2_U3588) );
  OAI21_X1 U22905 ( .B1(n19851), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19849), 
        .ZN(n19848) );
  INV_X1 U22906 ( .A(n19848), .ZN(P2_U3591) );
  OAI21_X1 U22907 ( .B1(n19851), .B2(n19850), .A(n19849), .ZN(P2_U3592) );
  NAND2_X1 U22908 ( .A1(n19853), .A2(n19852), .ZN(n19860) );
  NAND3_X1 U22909 ( .A1(n19877), .A2(n19854), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19855) );
  NAND2_X1 U22910 ( .A1(n19855), .A2(n19872), .ZN(n19865) );
  OAI21_X1 U22911 ( .B1(n19856), .B2(n19876), .A(n19865), .ZN(n19858) );
  NAND2_X1 U22912 ( .A1(n19858), .A2(n19857), .ZN(n19859) );
  OAI211_X1 U22913 ( .C1(n19861), .C2(n19668), .A(n19860), .B(n19859), .ZN(
        n19862) );
  INV_X1 U22914 ( .A(n19862), .ZN(n19863) );
  AOI22_X1 U22915 ( .A1(n19891), .A2(n19864), .B1(n19863), .B2(n19888), .ZN(
        P2_U3602) );
  OAI22_X1 U22916 ( .A1(n19866), .A2(n19865), .B1(n20699), .B2(n19668), .ZN(
        n19867) );
  AOI21_X1 U22917 ( .B1(n19869), .B2(n19868), .A(n19867), .ZN(n19870) );
  AOI22_X1 U22918 ( .A1(n19891), .A2(n19871), .B1(n19870), .B2(n19888), .ZN(
        P2_U3603) );
  INV_X1 U22919 ( .A(n19872), .ZN(n19883) );
  AND2_X1 U22920 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19873) );
  OR3_X1 U22921 ( .A1(n19874), .A2(n19883), .A3(n19873), .ZN(n19875) );
  OAI21_X1 U22922 ( .B1(n19877), .B2(n19876), .A(n19875), .ZN(n19878) );
  AOI21_X1 U22923 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19879), .A(n19878), 
        .ZN(n19880) );
  AOI22_X1 U22924 ( .A1(n19891), .A2(n19881), .B1(n19880), .B2(n19888), .ZN(
        P2_U3604) );
  OAI21_X1 U22925 ( .B1(n19884), .B2(n19883), .A(n19882), .ZN(n19885) );
  AOI21_X1 U22926 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(n19889) );
  AOI22_X1 U22927 ( .A1(n19891), .A2(n19890), .B1(n19889), .B2(n19888), .ZN(
        P2_U3605) );
  INV_X1 U22928 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19892) );
  AOI22_X1 U22929 ( .A1(n19901), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19892), 
        .B2(n19898), .ZN(P2_U3608) );
  OAI21_X1 U22930 ( .B1(n19895), .B2(n19894), .A(n19893), .ZN(n19897) );
  MUX2_X1 U22931 ( .A(P2_MORE_REG_SCAN_IN), .B(n19897), .S(n19896), .Z(
        P2_U3609) );
  INV_X1 U22932 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19899) );
  AOI22_X1 U22933 ( .A1(n19901), .A2(n19900), .B1(n19899), .B2(n19898), .ZN(
        P2_U3611) );
  INV_X1 U22934 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19902) );
  OAI21_X1 U22935 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n19902), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20601) );
  INV_X1 U22936 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20592) );
  OAI21_X1 U22937 ( .B1(n20601), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20689), .ZN(
        n19903) );
  INV_X1 U22938 ( .A(n19903), .ZN(P1_U2802) );
  NOR2_X1 U22939 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19905) );
  OAI21_X1 U22940 ( .B1(n19905), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20689), .ZN(
        n19904) );
  OAI21_X1 U22941 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20689), .A(n19904), 
        .ZN(P1_U2804) );
  NAND2_X1 U22942 ( .A1(n20601), .A2(n20689), .ZN(n20664) );
  INV_X1 U22943 ( .A(n20664), .ZN(n20668) );
  OAI21_X1 U22944 ( .B1(BS16), .B2(n19905), .A(n20668), .ZN(n20666) );
  OAI21_X1 U22945 ( .B1(n20668), .B2(n20321), .A(n20666), .ZN(P1_U2805) );
  OAI21_X1 U22946 ( .B1(n19908), .B2(n19907), .A(n19906), .ZN(P1_U2806) );
  NOR4_X1 U22947 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19912) );
  NOR4_X1 U22948 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19911) );
  NOR4_X1 U22949 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19910) );
  NOR4_X1 U22950 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19909) );
  NAND4_X1 U22951 ( .A1(n19912), .A2(n19911), .A3(n19910), .A4(n19909), .ZN(
        n19918) );
  NOR4_X1 U22952 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19916) );
  AOI211_X1 U22953 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_11__SCAN_IN), .B(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19915) );
  NOR4_X1 U22954 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19914) );
  NOR4_X1 U22955 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19913) );
  NAND4_X1 U22956 ( .A1(n19916), .A2(n19915), .A3(n19914), .A4(n19913), .ZN(
        n19917) );
  NOR2_X1 U22957 ( .A1(n19918), .A2(n19917), .ZN(n20673) );
  INV_X1 U22958 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20661) );
  NOR3_X1 U22959 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19920) );
  OAI21_X1 U22960 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19920), .A(n20673), .ZN(
        n19919) );
  OAI21_X1 U22961 ( .B1(n20673), .B2(n20661), .A(n19919), .ZN(P1_U2807) );
  INV_X1 U22962 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20669) );
  INV_X1 U22963 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20667) );
  AOI21_X1 U22964 ( .B1(n20669), .B2(n20667), .A(n19920), .ZN(n19921) );
  INV_X1 U22965 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20658) );
  INV_X1 U22966 ( .A(n20673), .ZN(n20675) );
  AOI22_X1 U22967 ( .A1(n20673), .A2(n19921), .B1(n20658), .B2(n20675), .ZN(
        P1_U2808) );
  NAND2_X1 U22968 ( .A1(n19949), .A2(n19924), .ZN(n19944) );
  OAI21_X1 U22969 ( .B1(n19996), .B2(n19922), .A(n19982), .ZN(n19926) );
  OAI22_X1 U22970 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19924), .B1(n20010), 
        .B2(n19923), .ZN(n19925) );
  AOI211_X1 U22971 ( .C1(P1_EBX_REG_9__SCAN_IN), .C2(n20006), .A(n19926), .B(
        n19925), .ZN(n19931) );
  INV_X1 U22972 ( .A(n19927), .ZN(n19929) );
  AOI22_X1 U22973 ( .A1(n19929), .A2(n19959), .B1(n20013), .B2(n19928), .ZN(
        n19930) );
  OAI211_X1 U22974 ( .C1(n20624), .C2(n19944), .A(n19931), .B(n19930), .ZN(
        P1_U2831) );
  NOR3_X1 U22975 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19933), .A3(n19932), .ZN(
        n19938) );
  OAI21_X1 U22976 ( .B1(n19996), .B2(n20950), .A(n19982), .ZN(n19934) );
  AOI21_X1 U22977 ( .B1(n20006), .B2(P1_EBX_REG_8__SCAN_IN), .A(n19934), .ZN(
        n19935) );
  OAI21_X1 U22978 ( .B1(n19936), .B2(n20010), .A(n19935), .ZN(n19937) );
  AOI211_X1 U22979 ( .C1(n19939), .C2(n19959), .A(n19938), .B(n19937), .ZN(
        n19940) );
  INV_X1 U22980 ( .A(n19940), .ZN(n19941) );
  AOI21_X1 U22981 ( .B1(n19942), .B2(n20013), .A(n19941), .ZN(n19943) );
  OAI21_X1 U22982 ( .B1(n20622), .B2(n19944), .A(n19943), .ZN(P1_U2832) );
  OAI21_X1 U22983 ( .B1(n19996), .B2(n11672), .A(n19982), .ZN(n19947) );
  NAND3_X1 U22984 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n19964), .ZN(n19948) );
  OAI22_X1 U22985 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19948), .B1(n20010), 
        .B2(n19945), .ZN(n19946) );
  AOI211_X1 U22986 ( .C1(P1_EBX_REG_7__SCAN_IN), .C2(n20006), .A(n19947), .B(
        n19946), .ZN(n19952) );
  AND2_X1 U22987 ( .A1(n19949), .A2(n19948), .ZN(n19958) );
  AOI22_X1 U22988 ( .A1(n19950), .A2(n19959), .B1(n19958), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n19951) );
  OAI211_X1 U22989 ( .C1(n19953), .C2(n19991), .A(n19952), .B(n19951), .ZN(
        P1_U2833) );
  NAND2_X1 U22990 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19964), .ZN(n19955) );
  AOI22_X1 U22991 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20006), .B1(n19993), .B2(
        n9831), .ZN(n19954) );
  OAI21_X1 U22992 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19955), .A(n19954), .ZN(
        n19956) );
  AOI211_X1 U22993 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19957), .B(n19956), .ZN(n19961) );
  AOI22_X1 U22994 ( .A1(n20018), .A2(n19959), .B1(n19958), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n19960) );
  OAI211_X1 U22995 ( .C1(n19962), .C2(n19991), .A(n19961), .B(n19960), .ZN(
        P1_U2834) );
  AOI22_X1 U22996 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20006), .B1(n19964), .B2(
        n13766), .ZN(n19970) );
  INV_X1 U22997 ( .A(n20017), .ZN(n19987) );
  NOR2_X1 U22998 ( .A1(n19964), .A2(n19963), .ZN(n19988) );
  AOI22_X1 U22999 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20014), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n19988), .ZN(n19965) );
  OAI211_X1 U23000 ( .C1(n19966), .C2(n20010), .A(n19982), .B(n19965), .ZN(
        n19967) );
  AOI21_X1 U23001 ( .B1(n19968), .B2(n19987), .A(n19967), .ZN(n19969) );
  OAI211_X1 U23002 ( .C1(n19971), .C2(n19991), .A(n19970), .B(n19969), .ZN(
        P1_U2835) );
  INV_X1 U23003 ( .A(n19972), .ZN(n19975) );
  INV_X1 U23004 ( .A(n19973), .ZN(n19974) );
  OAI21_X1 U23005 ( .B1(n19976), .B2(n19975), .A(n19974), .ZN(n19978) );
  AND2_X1 U23006 ( .A1(n19978), .A2(n19977), .ZN(n20077) );
  NOR3_X1 U23007 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19980), .A3(n19979), .ZN(
        n19986) );
  AOI22_X1 U23008 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20014), .B1(
        n19981), .B2(n20007), .ZN(n19983) );
  OAI211_X1 U23009 ( .C1(n19984), .C2(n20846), .A(n19983), .B(n19982), .ZN(
        n19985) );
  AOI211_X1 U23010 ( .C1(n20077), .C2(n19993), .A(n19986), .B(n19985), .ZN(
        n19990) );
  AOI22_X1 U23011 ( .A1(n19988), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n20061), 
        .B2(n19987), .ZN(n19989) );
  OAI211_X1 U23012 ( .C1(n20065), .C2(n19991), .A(n19990), .B(n19989), .ZN(
        P1_U2836) );
  AOI21_X1 U23013 ( .B1(n20005), .B2(n20669), .A(n19992), .ZN(n20004) );
  INV_X1 U23014 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20612) );
  AOI22_X1 U23015 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(n20006), .B1(n19993), .B2(
        n20099), .ZN(n20003) );
  INV_X1 U23016 ( .A(n13519), .ZN(n20124) );
  NAND3_X1 U23017 ( .A1(n20005), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n20612), 
        .ZN(n19994) );
  OAI21_X1 U23018 ( .B1(n19996), .B2(n19995), .A(n19994), .ZN(n19997) );
  AOI21_X1 U23019 ( .B1(n20124), .B2(n20007), .A(n19997), .ZN(n19998) );
  OAI21_X1 U23020 ( .B1(n19999), .B2(n20017), .A(n19998), .ZN(n20000) );
  AOI21_X1 U23021 ( .B1(n20001), .B2(n20013), .A(n20000), .ZN(n20002) );
  OAI211_X1 U23022 ( .C1(n20004), .C2(n20612), .A(n20003), .B(n20002), .ZN(
        P1_U2838) );
  AOI22_X1 U23023 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20006), .B1(n20005), .B2(
        n20669), .ZN(n20016) );
  INV_X1 U23024 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20069) );
  INV_X1 U23025 ( .A(n20007), .ZN(n20008) );
  OAI222_X1 U23026 ( .A1(n20011), .A2(n20010), .B1(n20009), .B2(n20669), .C1(
        n20436), .C2(n20008), .ZN(n20012) );
  AOI221_X1 U23027 ( .B1(n20014), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C1(
        n20013), .C2(n20069), .A(n20012), .ZN(n20015) );
  OAI211_X1 U23028 ( .C1(n20017), .C2(n20075), .A(n20016), .B(n20015), .ZN(
        P1_U2839) );
  AOI22_X1 U23029 ( .A1(n20018), .A2(n12893), .B1(n20021), .B2(n9831), .ZN(
        n20019) );
  OAI21_X1 U23030 ( .B1(n20023), .B2(n20020), .A(n20019), .ZN(P1_U2866) );
  AOI22_X1 U23031 ( .A1(n20061), .A2(n12893), .B1(n20021), .B2(n20077), .ZN(
        n20022) );
  OAI21_X1 U23032 ( .B1(n20023), .B2(n20846), .A(n20022), .ZN(P1_U2868) );
  AOI22_X1 U23033 ( .A1(n20036), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20024) );
  OAI21_X1 U23034 ( .B1(n20025), .B2(n20045), .A(n20024), .ZN(P1_U2921) );
  AOI22_X1 U23035 ( .A1(P1_EAX_REG_14__SCAN_IN), .A2(n20035), .B1(n20036), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20026) );
  OAI21_X1 U23036 ( .B1(n20731), .B2(n20044), .A(n20026), .ZN(P1_U2922) );
  AOI22_X1 U23037 ( .A1(n20036), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20027) );
  OAI21_X1 U23038 ( .B1(n13403), .B2(n20045), .A(n20027), .ZN(P1_U2923) );
  AOI22_X1 U23039 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n20035), .B1(n20036), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20028) );
  OAI21_X1 U23040 ( .B1(n20824), .B2(n20044), .A(n20028), .ZN(P1_U2924) );
  AOI22_X1 U23041 ( .A1(n20036), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20029) );
  OAI21_X1 U23042 ( .B1(n14216), .B2(n20045), .A(n20029), .ZN(P1_U2925) );
  AOI22_X1 U23043 ( .A1(n20036), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20030) );
  OAI21_X1 U23044 ( .B1(n13406), .B2(n20045), .A(n20030), .ZN(P1_U2926) );
  AOI22_X1 U23045 ( .A1(n20036), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U23046 ( .B1(n14106), .B2(n20045), .A(n20031), .ZN(P1_U2927) );
  AOI22_X1 U23047 ( .A1(n20036), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U23048 ( .B1(n13938), .B2(n20045), .A(n20032), .ZN(P1_U2928) );
  AOI22_X1 U23049 ( .A1(n20036), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U23050 ( .B1(n13419), .B2(n20045), .A(n20033), .ZN(P1_U2929) );
  AOI22_X1 U23051 ( .A1(n20036), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U23052 ( .B1(n13846), .B2(n20045), .A(n20034), .ZN(P1_U2930) );
  AOI222_X1 U23053 ( .A1(n20036), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20035), 
        .B2(P1_EAX_REG_5__SCAN_IN), .C1(n20038), .C2(P1_DATAO_REG_5__SCAN_IN), 
        .ZN(n20037) );
  INV_X1 U23054 ( .A(n20037), .ZN(P1_U2931) );
  AOI22_X1 U23055 ( .A1(n20036), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20039) );
  OAI21_X1 U23056 ( .B1(n13738), .B2(n20045), .A(n20039), .ZN(P1_U2932) );
  INV_X1 U23057 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n20917) );
  OAI222_X1 U23058 ( .A1(n20046), .A2(n20917), .B1(n20045), .B2(n13411), .C1(
        n20044), .C2(n20040), .ZN(P1_U2933) );
  AOI22_X1 U23059 ( .A1(n20036), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20038), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20041) );
  OAI21_X1 U23060 ( .B1(n13400), .B2(n20045), .A(n20041), .ZN(P1_U2934) );
  INV_X1 U23061 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U23062 ( .A1(n20044), .A2(n20867), .B1(n20045), .B2(n13397), .C1(
        n20046), .C2(n20042), .ZN(P1_U2935) );
  INV_X1 U23063 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n20882) );
  OAI222_X1 U23064 ( .A1(n20046), .A2(n20882), .B1(n20045), .B2(n13394), .C1(
        n20044), .C2(n20043), .ZN(P1_U2936) );
  AOI22_X1 U23065 ( .A1(n20054), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20053), .ZN(n20048) );
  NAND2_X1 U23066 ( .A1(n20048), .A2(n20047), .ZN(P1_U2961) );
  AOI22_X1 U23067 ( .A1(n20054), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20053), .ZN(n20050) );
  NAND2_X1 U23068 ( .A1(n20050), .A2(n20049), .ZN(P1_U2963) );
  AOI22_X1 U23069 ( .A1(n20054), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20053), .ZN(n20052) );
  NAND2_X1 U23070 ( .A1(n20052), .A2(n20051), .ZN(P1_U2964) );
  AOI22_X1 U23071 ( .A1(n20054), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20053), .ZN(n20056) );
  NAND2_X1 U23072 ( .A1(n20056), .A2(n20055), .ZN(P1_U2966) );
  AOI22_X1 U23073 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20064) );
  OAI21_X1 U23074 ( .B1(n20059), .B2(n20058), .A(n20057), .ZN(n20060) );
  INV_X1 U23075 ( .A(n20060), .ZN(n20078) );
  AOI22_X1 U23076 ( .A1(n20078), .A2(n20071), .B1(n20062), .B2(n20061), .ZN(
        n20063) );
  OAI211_X1 U23077 ( .C1(n20066), .C2(n20065), .A(n20064), .B(n20063), .ZN(
        P1_U2995) );
  AOI22_X1 U23078 ( .A1(n20067), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20106), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20074) );
  INV_X1 U23079 ( .A(n20068), .ZN(n20072) );
  AOI22_X1 U23080 ( .A1(n20072), .A2(n20071), .B1(n20070), .B2(n20069), .ZN(
        n20073) );
  OAI211_X1 U23081 ( .C1(n20076), .C2(n20075), .A(n20074), .B(n20073), .ZN(
        P1_U2998) );
  AOI22_X1 U23082 ( .A1(n20098), .A2(n20077), .B1(n20106), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20083) );
  AOI22_X1 U23083 ( .A1(n20078), .A2(n20103), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20089), .ZN(n20082) );
  OAI211_X1 U23084 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20080), .B(n20079), .ZN(n20081) );
  NAND3_X1 U23085 ( .A1(n20083), .A2(n20082), .A3(n20081), .ZN(P1_U3027) );
  INV_X1 U23086 ( .A(n20084), .ZN(n20085) );
  AOI21_X1 U23087 ( .B1(n20098), .B2(n20086), .A(n20085), .ZN(n20091) );
  INV_X1 U23088 ( .A(n20087), .ZN(n20088) );
  AOI22_X1 U23089 ( .A1(n20089), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20088), .B2(n20103), .ZN(n20090) );
  OAI211_X1 U23090 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20092), .A(
        n20091), .B(n20090), .ZN(P1_U3028) );
  NAND2_X1 U23091 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20095) );
  INV_X1 U23092 ( .A(n20093), .ZN(n20094) );
  OAI21_X1 U23093 ( .B1(n20095), .B2(n20107), .A(n20094), .ZN(n20096) );
  AOI22_X1 U23094 ( .A1(n20099), .A2(n20098), .B1(n20097), .B2(n20096), .ZN(
        n20112) );
  OAI21_X1 U23095 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20101), .A(
        n20100), .ZN(n20105) );
  INV_X1 U23096 ( .A(n20102), .ZN(n20104) );
  AOI22_X1 U23097 ( .A1(n20105), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20104), .B2(n20103), .ZN(n20111) );
  NAND2_X1 U23098 ( .A1(n20106), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20110) );
  NAND3_X1 U23099 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20108), .A3(
        n20107), .ZN(n20109) );
  NAND4_X1 U23100 ( .A1(n20112), .A2(n20111), .A3(n20110), .A4(n20109), .ZN(
        P1_U3029) );
  NOR2_X1 U23101 ( .A1(n20114), .A2(n20113), .ZN(P1_U3032) );
  INV_X1 U23102 ( .A(n20115), .ZN(n20116) );
  INV_X1 U23103 ( .A(n20224), .ZN(n20119) );
  INV_X1 U23104 ( .A(n20262), .ZN(n20118) );
  NOR2_X1 U23105 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20222) );
  INV_X1 U23106 ( .A(n20431), .ZN(n20120) );
  NAND2_X1 U23107 ( .A1(n20222), .A2(n20120), .ZN(n20152) );
  OAI22_X1 U23108 ( .A1(n20587), .A2(n20544), .B1(n20152), .B2(n20432), .ZN(
        n20121) );
  INV_X1 U23109 ( .A(n20121), .ZN(n20133) );
  INV_X1 U23110 ( .A(n20182), .ZN(n20122) );
  INV_X1 U23111 ( .A(n20587), .ZN(n20540) );
  OAI21_X1 U23112 ( .B1(n20122), .B2(n20540), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20123) );
  NAND2_X1 U23113 ( .A1(n20123), .A2(n20538), .ZN(n20131) );
  OR2_X1 U23114 ( .A1(n20125), .A2(n20124), .ZN(n20225) );
  NOR2_X1 U23115 ( .A1(n20225), .A2(n20488), .ZN(n20129) );
  OR2_X1 U23116 ( .A1(n20127), .A2(n20126), .ZN(n20260) );
  AOI22_X1 U23117 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20260), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20152), .ZN(n20128) );
  OAI211_X1 U23118 ( .C1(n20131), .C2(n20129), .A(n20128), .B(n20354), .ZN(
        n20155) );
  INV_X1 U23119 ( .A(n20129), .ZN(n20130) );
  OAI22_X1 U23120 ( .A1(n20131), .A2(n20130), .B1(n20359), .B2(n20260), .ZN(
        n20154) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20155), .B1(
        n20528), .B2(n20154), .ZN(n20132) );
  OAI211_X1 U23122 ( .C1(n20500), .C2(n20182), .A(n20133), .B(n20132), .ZN(
        P1_U3033) );
  OAI22_X1 U23123 ( .A1(n20587), .A2(n9858), .B1(n20152), .B2(n20447), .ZN(
        n20134) );
  INV_X1 U23124 ( .A(n20134), .ZN(n20136) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20155), .B1(
        n20546), .B2(n20154), .ZN(n20135) );
  OAI211_X1 U23126 ( .C1(n20549), .C2(n20182), .A(n20136), .B(n20135), .ZN(
        P1_U3034) );
  OAI22_X1 U23127 ( .A1(n20587), .A2(n20456), .B1(n20152), .B2(n20452), .ZN(
        n20137) );
  INV_X1 U23128 ( .A(n20137), .ZN(n20139) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20155), .B1(
        n20551), .B2(n20154), .ZN(n20138) );
  OAI211_X1 U23130 ( .C1(n20555), .C2(n20182), .A(n20139), .B(n20138), .ZN(
        P1_U3035) );
  OAI22_X1 U23131 ( .A1(n20587), .A2(n9856), .B1(n20152), .B2(n20457), .ZN(
        n20140) );
  INV_X1 U23132 ( .A(n20140), .ZN(n20142) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20155), .B1(
        n20557), .B2(n20154), .ZN(n20141) );
  OAI211_X1 U23134 ( .C1(n20560), .C2(n20182), .A(n20142), .B(n20141), .ZN(
        P1_U3036) );
  OAI22_X1 U23135 ( .A1(n20587), .A2(n20466), .B1(n20152), .B2(n20462), .ZN(
        n20143) );
  INV_X1 U23136 ( .A(n20143), .ZN(n20145) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20155), .B1(
        n20562), .B2(n20154), .ZN(n20144) );
  OAI211_X1 U23138 ( .C1(n20566), .C2(n20182), .A(n20145), .B(n20144), .ZN(
        P1_U3037) );
  OAI22_X1 U23139 ( .A1(n20587), .A2(n9854), .B1(n20152), .B2(n20467), .ZN(
        n20146) );
  INV_X1 U23140 ( .A(n20146), .ZN(n20148) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20155), .B1(
        n20568), .B2(n20154), .ZN(n20147) );
  OAI211_X1 U23142 ( .C1(n20571), .C2(n20182), .A(n20148), .B(n20147), .ZN(
        P1_U3038) );
  OAI22_X1 U23143 ( .A1(n20587), .A2(n20476), .B1(n20152), .B2(n20472), .ZN(
        n20149) );
  INV_X1 U23144 ( .A(n20149), .ZN(n20151) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20155), .B1(
        n20573), .B2(n20154), .ZN(n20150) );
  OAI211_X1 U23146 ( .C1(n9852), .C2(n20182), .A(n20151), .B(n20150), .ZN(
        P1_U3039) );
  OAI22_X1 U23147 ( .A1(n20587), .A2(n20486), .B1(n20152), .B2(n20477), .ZN(
        n20153) );
  INV_X1 U23148 ( .A(n20153), .ZN(n20157) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20155), .B1(
        n20581), .B2(n20154), .ZN(n20156) );
  OAI211_X1 U23150 ( .C1(n9850), .C2(n20182), .A(n20157), .B(n20156), .ZN(
        P1_U3040) );
  INV_X1 U23151 ( .A(n20225), .ZN(n20158) );
  NAND2_X1 U23152 ( .A1(n20222), .A2(n20524), .ZN(n20159) );
  NOR2_X1 U23153 ( .A1(n20317), .A2(n20159), .ZN(n20177) );
  AOI21_X1 U23154 ( .B1(n20158), .B2(n20318), .A(n20177), .ZN(n20160) );
  OAI22_X1 U23155 ( .A1(n20160), .A2(n20530), .B1(n20159), .B2(n20525), .ZN(
        n20178) );
  AOI22_X1 U23156 ( .A1(n20528), .A2(n20178), .B1(n20527), .B2(n20177), .ZN(
        n20164) );
  INV_X1 U23157 ( .A(n20159), .ZN(n20162) );
  OAI211_X1 U23158 ( .C1(n20224), .C2(n20321), .A(n20538), .B(n20160), .ZN(
        n20161) );
  OAI211_X1 U23159 ( .C1(n20538), .C2(n20162), .A(n20536), .B(n20161), .ZN(
        n20179) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n20539), .ZN(n20163) );
  OAI211_X1 U23161 ( .C1(n20544), .C2(n20182), .A(n20164), .B(n20163), .ZN(
        P1_U3041) );
  AOI22_X1 U23162 ( .A1(n20546), .A2(n20178), .B1(n20545), .B2(n20177), .ZN(
        n20166) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n20408), .ZN(n20165) );
  OAI211_X1 U23164 ( .C1(n9858), .C2(n20182), .A(n20166), .B(n20165), .ZN(
        P1_U3042) );
  AOI22_X1 U23165 ( .A1(n20551), .A2(n20178), .B1(n20550), .B2(n20177), .ZN(
        n20168) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n20411), .ZN(n20167) );
  OAI211_X1 U23167 ( .C1(n20456), .C2(n20182), .A(n20168), .B(n20167), .ZN(
        P1_U3043) );
  AOI22_X1 U23168 ( .A1(n20557), .A2(n20178), .B1(n20556), .B2(n20177), .ZN(
        n20170) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n20414), .ZN(n20169) );
  OAI211_X1 U23170 ( .C1(n9856), .C2(n20182), .A(n20170), .B(n20169), .ZN(
        P1_U3044) );
  AOI22_X1 U23171 ( .A1(n20562), .A2(n20178), .B1(n20561), .B2(n20177), .ZN(
        n20172) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n20303), .ZN(n20171) );
  OAI211_X1 U23173 ( .C1(n20466), .C2(n20182), .A(n20172), .B(n20171), .ZN(
        P1_U3045) );
  AOI22_X1 U23174 ( .A1(n20568), .A2(n20178), .B1(n20567), .B2(n20177), .ZN(
        n20174) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n20336), .ZN(n20173) );
  OAI211_X1 U23176 ( .C1(n9854), .C2(n20182), .A(n20174), .B(n20173), .ZN(
        P1_U3046) );
  AOI22_X1 U23177 ( .A1(n20573), .A2(n20178), .B1(n20572), .B2(n20177), .ZN(
        n20176) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n9851), .ZN(n20175) );
  OAI211_X1 U23179 ( .C1(n20476), .C2(n20182), .A(n20176), .B(n20175), .ZN(
        P1_U3047) );
  AOI22_X1 U23180 ( .A1(n20581), .A2(n20178), .B1(n20579), .B2(n20177), .ZN(
        n20181) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20179), .B1(
        n20184), .B2(n9849), .ZN(n20180) );
  OAI211_X1 U23182 ( .C1(n20486), .C2(n20182), .A(n20181), .B(n20180), .ZN(
        P1_U3048) );
  NAND2_X1 U23183 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20222), .ZN(
        n20229) );
  OR2_X1 U23184 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20229), .ZN(
        n20215) );
  OAI22_X1 U23185 ( .A1(n20253), .A2(n20500), .B1(n20215), .B2(n20432), .ZN(
        n20183) );
  INV_X1 U23186 ( .A(n20183), .ZN(n20196) );
  INV_X1 U23187 ( .A(n20253), .ZN(n20185) );
  OAI21_X1 U23188 ( .B1(n20185), .B2(n20184), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20186) );
  NAND2_X1 U23189 ( .A1(n20186), .A2(n20538), .ZN(n20194) );
  NOR2_X1 U23190 ( .A1(n20225), .A2(n20436), .ZN(n20190) );
  AOI211_X1 U23191 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20215), .A(n20188), 
        .B(n20187), .ZN(n20189) );
  INV_X1 U23192 ( .A(n20190), .ZN(n20193) );
  INV_X1 U23193 ( .A(n20191), .ZN(n20192) );
  OAI22_X1 U23194 ( .A1(n20194), .A2(n20193), .B1(n20192), .B2(n20359), .ZN(
        n20218) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20219), .B1(
        n20528), .B2(n20218), .ZN(n20195) );
  OAI211_X1 U23196 ( .C1(n20544), .C2(n20216), .A(n20196), .B(n20195), .ZN(
        P1_U3049) );
  OAI22_X1 U23197 ( .A1(n20216), .A2(n9858), .B1(n20215), .B2(n20447), .ZN(
        n20197) );
  INV_X1 U23198 ( .A(n20197), .ZN(n20199) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20219), .B1(
        n20546), .B2(n20218), .ZN(n20198) );
  OAI211_X1 U23200 ( .C1(n20549), .C2(n20253), .A(n20199), .B(n20198), .ZN(
        P1_U3050) );
  OAI22_X1 U23201 ( .A1(n20253), .A2(n20555), .B1(n20215), .B2(n20452), .ZN(
        n20200) );
  INV_X1 U23202 ( .A(n20200), .ZN(n20202) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20219), .B1(
        n20551), .B2(n20218), .ZN(n20201) );
  OAI211_X1 U23204 ( .C1(n20456), .C2(n20216), .A(n20202), .B(n20201), .ZN(
        P1_U3051) );
  OAI22_X1 U23205 ( .A1(n20216), .A2(n9856), .B1(n20215), .B2(n20457), .ZN(
        n20203) );
  INV_X1 U23206 ( .A(n20203), .ZN(n20205) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20219), .B1(
        n20557), .B2(n20218), .ZN(n20204) );
  OAI211_X1 U23208 ( .C1(n20560), .C2(n20253), .A(n20205), .B(n20204), .ZN(
        P1_U3052) );
  OAI22_X1 U23209 ( .A1(n20216), .A2(n20466), .B1(n20215), .B2(n20462), .ZN(
        n20206) );
  INV_X1 U23210 ( .A(n20206), .ZN(n20208) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20219), .B1(
        n20562), .B2(n20218), .ZN(n20207) );
  OAI211_X1 U23212 ( .C1(n20566), .C2(n20253), .A(n20208), .B(n20207), .ZN(
        P1_U3053) );
  OAI22_X1 U23213 ( .A1(n20253), .A2(n20571), .B1(n20215), .B2(n20467), .ZN(
        n20209) );
  INV_X1 U23214 ( .A(n20209), .ZN(n20211) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20219), .B1(
        n20568), .B2(n20218), .ZN(n20210) );
  OAI211_X1 U23216 ( .C1(n9854), .C2(n20216), .A(n20211), .B(n20210), .ZN(
        P1_U3054) );
  OAI22_X1 U23217 ( .A1(n20216), .A2(n20476), .B1(n20215), .B2(n20472), .ZN(
        n20212) );
  INV_X1 U23218 ( .A(n20212), .ZN(n20214) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20219), .B1(
        n20573), .B2(n20218), .ZN(n20213) );
  OAI211_X1 U23220 ( .C1(n9852), .C2(n20253), .A(n20214), .B(n20213), .ZN(
        P1_U3055) );
  OAI22_X1 U23221 ( .A1(n20216), .A2(n20486), .B1(n20215), .B2(n20477), .ZN(
        n20217) );
  INV_X1 U23222 ( .A(n20217), .ZN(n20221) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20219), .B1(
        n20581), .B2(n20218), .ZN(n20220) );
  OAI211_X1 U23224 ( .C1(n9850), .C2(n20253), .A(n20221), .B(n20220), .ZN(
        P1_U3056) );
  NAND2_X1 U23225 ( .A1(n20222), .A2(n20391), .ZN(n20252) );
  OAI22_X1 U23226 ( .A1(n20253), .A2(n20544), .B1(n20252), .B2(n20432), .ZN(
        n20223) );
  INV_X1 U23227 ( .A(n20223), .ZN(n20233) );
  AOI21_X1 U23228 ( .B1(n20224), .B2(n20389), .A(n20533), .ZN(n20230) );
  OR2_X1 U23229 ( .A1(n20225), .A2(n20519), .ZN(n20226) );
  INV_X1 U23230 ( .A(n20231), .ZN(n20228) );
  AOI21_X1 U23231 ( .B1(n20530), .B2(n20229), .A(n20396), .ZN(n20227) );
  OAI21_X1 U23232 ( .B1(n20230), .B2(n20228), .A(n20227), .ZN(n20256) );
  OAI22_X1 U23233 ( .A1(n20231), .A2(n20230), .B1(n20525), .B2(n20229), .ZN(
        n20255) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20256), .B1(
        n20528), .B2(n20255), .ZN(n20232) );
  OAI211_X1 U23235 ( .C1(n20500), .C2(n20279), .A(n20233), .B(n20232), .ZN(
        P1_U3057) );
  OAI22_X1 U23236 ( .A1(n20253), .A2(n9858), .B1(n20252), .B2(n20447), .ZN(
        n20234) );
  INV_X1 U23237 ( .A(n20234), .ZN(n20236) );
  AOI22_X1 U23238 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20256), .B1(
        n20546), .B2(n20255), .ZN(n20235) );
  OAI211_X1 U23239 ( .C1(n20549), .C2(n20279), .A(n20236), .B(n20235), .ZN(
        P1_U3058) );
  OAI22_X1 U23240 ( .A1(n20253), .A2(n20456), .B1(n20252), .B2(n20452), .ZN(
        n20237) );
  INV_X1 U23241 ( .A(n20237), .ZN(n20239) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20256), .B1(
        n20551), .B2(n20255), .ZN(n20238) );
  OAI211_X1 U23243 ( .C1(n20555), .C2(n20279), .A(n20239), .B(n20238), .ZN(
        P1_U3059) );
  OAI22_X1 U23244 ( .A1(n20253), .A2(n9856), .B1(n20252), .B2(n20457), .ZN(
        n20240) );
  INV_X1 U23245 ( .A(n20240), .ZN(n20242) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20256), .B1(
        n20557), .B2(n20255), .ZN(n20241) );
  OAI211_X1 U23247 ( .C1(n20560), .C2(n20279), .A(n20242), .B(n20241), .ZN(
        P1_U3060) );
  OAI22_X1 U23248 ( .A1(n20279), .A2(n20566), .B1(n20252), .B2(n20462), .ZN(
        n20243) );
  INV_X1 U23249 ( .A(n20243), .ZN(n20245) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20256), .B1(
        n20562), .B2(n20255), .ZN(n20244) );
  OAI211_X1 U23251 ( .C1(n20466), .C2(n20253), .A(n20245), .B(n20244), .ZN(
        P1_U3061) );
  OAI22_X1 U23252 ( .A1(n20253), .A2(n9854), .B1(n20252), .B2(n20467), .ZN(
        n20246) );
  INV_X1 U23253 ( .A(n20246), .ZN(n20248) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20256), .B1(
        n20568), .B2(n20255), .ZN(n20247) );
  OAI211_X1 U23255 ( .C1(n20571), .C2(n20279), .A(n20248), .B(n20247), .ZN(
        P1_U3062) );
  OAI22_X1 U23256 ( .A1(n20279), .A2(n9852), .B1(n20252), .B2(n20472), .ZN(
        n20249) );
  INV_X1 U23257 ( .A(n20249), .ZN(n20251) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20256), .B1(
        n20573), .B2(n20255), .ZN(n20250) );
  OAI211_X1 U23259 ( .C1(n20476), .C2(n20253), .A(n20251), .B(n20250), .ZN(
        P1_U3063) );
  OAI22_X1 U23260 ( .A1(n20253), .A2(n20486), .B1(n20252), .B2(n20477), .ZN(
        n20254) );
  INV_X1 U23261 ( .A(n20254), .ZN(n20258) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20256), .B1(
        n20581), .B2(n20255), .ZN(n20257) );
  OAI211_X1 U23263 ( .C1(n9850), .C2(n20279), .A(n20258), .B(n20257), .ZN(
        P1_U3064) );
  NAND3_X1 U23264 ( .A1(n20289), .A2(n20538), .A3(n20436), .ZN(n20259) );
  OAI21_X1 U23265 ( .B1(n20260), .B2(n20490), .A(n20259), .ZN(n20283) );
  INV_X1 U23266 ( .A(n20288), .ZN(n20261) );
  NOR2_X1 U23267 ( .A1(n20261), .A2(n20431), .ZN(n20282) );
  AOI22_X1 U23268 ( .A1(n20528), .A2(n20283), .B1(n20527), .B2(n20282), .ZN(
        n20267) );
  AOI21_X1 U23269 ( .B1(n20279), .B2(n20316), .A(n20321), .ZN(n20263) );
  AOI21_X1 U23270 ( .B1(n20289), .B2(n20436), .A(n20263), .ZN(n20264) );
  NOR2_X1 U23271 ( .A1(n20264), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20265) );
  INV_X1 U23272 ( .A(n20316), .ZN(n20276) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20285), .B1(
        n20276), .B2(n20539), .ZN(n20266) );
  OAI211_X1 U23274 ( .C1(n20544), .C2(n20279), .A(n20267), .B(n20266), .ZN(
        P1_U3065) );
  AOI22_X1 U23275 ( .A1(n20546), .A2(n20283), .B1(n20545), .B2(n20282), .ZN(
        n20269) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n9857), .ZN(n20268) );
  OAI211_X1 U23277 ( .C1(n20549), .C2(n20316), .A(n20269), .B(n20268), .ZN(
        P1_U3066) );
  AOI22_X1 U23278 ( .A1(n20551), .A2(n20283), .B1(n20550), .B2(n20282), .ZN(
        n20271) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20285), .B1(
        n20276), .B2(n20411), .ZN(n20270) );
  OAI211_X1 U23280 ( .C1(n20456), .C2(n20279), .A(n20271), .B(n20270), .ZN(
        P1_U3067) );
  AOI22_X1 U23281 ( .A1(n20557), .A2(n20283), .B1(n20556), .B2(n20282), .ZN(
        n20273) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n9855), .ZN(n20272) );
  OAI211_X1 U23283 ( .C1(n20560), .C2(n20316), .A(n20273), .B(n20272), .ZN(
        P1_U3068) );
  AOI22_X1 U23284 ( .A1(n20562), .A2(n20283), .B1(n20561), .B2(n20282), .ZN(
        n20275) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20563), .ZN(n20274) );
  OAI211_X1 U23286 ( .C1(n20566), .C2(n20316), .A(n20275), .B(n20274), .ZN(
        P1_U3069) );
  AOI22_X1 U23287 ( .A1(n20568), .A2(n20283), .B1(n20567), .B2(n20282), .ZN(
        n20278) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20285), .B1(
        n20276), .B2(n20336), .ZN(n20277) );
  OAI211_X1 U23289 ( .C1(n9854), .C2(n20279), .A(n20278), .B(n20277), .ZN(
        P1_U3070) );
  AOI22_X1 U23290 ( .A1(n20573), .A2(n20283), .B1(n20572), .B2(n20282), .ZN(
        n20281) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20574), .ZN(n20280) );
  OAI211_X1 U23292 ( .C1(n9852), .C2(n20316), .A(n20281), .B(n20280), .ZN(
        P1_U3071) );
  AOI22_X1 U23293 ( .A1(n20581), .A2(n20283), .B1(n20579), .B2(n20282), .ZN(
        n20287) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20582), .ZN(n20286) );
  OAI211_X1 U23295 ( .C1(n9850), .C2(n20316), .A(n20287), .B(n20286), .ZN(
        P1_U3072) );
  NAND2_X1 U23296 ( .A1(n20288), .A2(n20524), .ZN(n20290) );
  NOR2_X1 U23297 ( .A1(n20317), .A2(n20290), .ZN(n20310) );
  AOI21_X1 U23298 ( .B1(n20289), .B2(n20318), .A(n20310), .ZN(n20291) );
  OAI22_X1 U23299 ( .A1(n20291), .A2(n20530), .B1(n20290), .B2(n20525), .ZN(
        n20311) );
  AOI22_X1 U23300 ( .A1(n20528), .A2(n20311), .B1(n20527), .B2(n20310), .ZN(
        n20296) );
  INV_X1 U23301 ( .A(n20290), .ZN(n20294) );
  OAI211_X1 U23302 ( .C1(n20292), .C2(n20321), .A(n20538), .B(n20291), .ZN(
        n20293) );
  OAI211_X1 U23303 ( .C1(n20538), .C2(n20294), .A(n20536), .B(n20293), .ZN(
        n20313) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20539), .ZN(n20295) );
  OAI211_X1 U23305 ( .C1(n20544), .C2(n20316), .A(n20296), .B(n20295), .ZN(
        P1_U3073) );
  AOI22_X1 U23306 ( .A1(n20546), .A2(n20311), .B1(n20545), .B2(n20310), .ZN(
        n20298) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20408), .ZN(n20297) );
  OAI211_X1 U23308 ( .C1(n9858), .C2(n20316), .A(n20298), .B(n20297), .ZN(
        P1_U3074) );
  AOI22_X1 U23309 ( .A1(n20551), .A2(n20311), .B1(n20550), .B2(n20310), .ZN(
        n20300) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20411), .ZN(n20299) );
  OAI211_X1 U23311 ( .C1(n20456), .C2(n20316), .A(n20300), .B(n20299), .ZN(
        P1_U3075) );
  AOI22_X1 U23312 ( .A1(n20557), .A2(n20311), .B1(n20556), .B2(n20310), .ZN(
        n20302) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20414), .ZN(n20301) );
  OAI211_X1 U23314 ( .C1(n9856), .C2(n20316), .A(n20302), .B(n20301), .ZN(
        P1_U3076) );
  AOI22_X1 U23315 ( .A1(n20562), .A2(n20311), .B1(n20561), .B2(n20310), .ZN(
        n20305) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20303), .ZN(n20304) );
  OAI211_X1 U23317 ( .C1(n20466), .C2(n20316), .A(n20305), .B(n20304), .ZN(
        P1_U3077) );
  AOI22_X1 U23318 ( .A1(n20568), .A2(n20311), .B1(n20567), .B2(n20310), .ZN(
        n20307) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20336), .ZN(n20306) );
  OAI211_X1 U23320 ( .C1(n9854), .C2(n20316), .A(n20307), .B(n20306), .ZN(
        P1_U3078) );
  AOI22_X1 U23321 ( .A1(n20573), .A2(n20311), .B1(n20572), .B2(n20310), .ZN(
        n20309) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n9851), .ZN(n20308) );
  OAI211_X1 U23323 ( .C1(n20476), .C2(n20316), .A(n20309), .B(n20308), .ZN(
        P1_U3079) );
  AOI22_X1 U23324 ( .A1(n20581), .A2(n20311), .B1(n20579), .B2(n20310), .ZN(
        n20315) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n9849), .ZN(n20314) );
  OAI211_X1 U23326 ( .C1(n20486), .C2(n20316), .A(n20315), .B(n20314), .ZN(
        P1_U3080) );
  NAND2_X1 U23327 ( .A1(n20392), .A2(n20524), .ZN(n20319) );
  NOR2_X1 U23328 ( .A1(n20317), .A2(n20319), .ZN(n20343) );
  AOI21_X1 U23329 ( .B1(n20352), .B2(n20318), .A(n20343), .ZN(n20320) );
  OAI22_X1 U23330 ( .A1(n20320), .A2(n20530), .B1(n20319), .B2(n20525), .ZN(
        n20344) );
  AOI22_X1 U23331 ( .A1(n20528), .A2(n20344), .B1(n20527), .B2(n20343), .ZN(
        n20327) );
  INV_X1 U23332 ( .A(n20319), .ZN(n20323) );
  OAI211_X1 U23333 ( .C1(n20390), .C2(n20321), .A(n20538), .B(n20320), .ZN(
        n20322) );
  OAI211_X1 U23334 ( .C1(n20538), .C2(n20323), .A(n20536), .B(n20322), .ZN(
        n20346) );
  INV_X1 U23335 ( .A(n20324), .ZN(n20325) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20346), .B1(
        n20339), .B2(n20539), .ZN(n20326) );
  OAI211_X1 U23337 ( .C1(n20544), .C2(n20342), .A(n20327), .B(n20326), .ZN(
        P1_U3105) );
  AOI22_X1 U23338 ( .A1(n20546), .A2(n20344), .B1(n20545), .B2(n20343), .ZN(
        n20329) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20346), .B1(
        n20339), .B2(n20408), .ZN(n20328) );
  OAI211_X1 U23340 ( .C1(n9858), .C2(n20342), .A(n20329), .B(n20328), .ZN(
        P1_U3106) );
  AOI22_X1 U23341 ( .A1(n20551), .A2(n20344), .B1(n20550), .B2(n20343), .ZN(
        n20331) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20346), .B1(
        n20339), .B2(n20411), .ZN(n20330) );
  OAI211_X1 U23343 ( .C1(n20456), .C2(n20342), .A(n20331), .B(n20330), .ZN(
        P1_U3107) );
  AOI22_X1 U23344 ( .A1(n20557), .A2(n20344), .B1(n20556), .B2(n20343), .ZN(
        n20333) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20346), .B1(
        n20339), .B2(n20414), .ZN(n20332) );
  OAI211_X1 U23346 ( .C1(n9856), .C2(n20342), .A(n20333), .B(n20332), .ZN(
        P1_U3108) );
  AOI22_X1 U23347 ( .A1(n20562), .A2(n20344), .B1(n20561), .B2(n20343), .ZN(
        n20335) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20563), .ZN(n20334) );
  OAI211_X1 U23349 ( .C1(n20566), .C2(n20383), .A(n20335), .B(n20334), .ZN(
        P1_U3109) );
  AOI22_X1 U23350 ( .A1(n20568), .A2(n20344), .B1(n20567), .B2(n20343), .ZN(
        n20338) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20346), .B1(
        n20339), .B2(n20336), .ZN(n20337) );
  OAI211_X1 U23352 ( .C1(n9854), .C2(n20342), .A(n20338), .B(n20337), .ZN(
        P1_U3110) );
  AOI22_X1 U23353 ( .A1(n20573), .A2(n20344), .B1(n20572), .B2(n20343), .ZN(
        n20341) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20346), .B1(
        n20339), .B2(n9851), .ZN(n20340) );
  OAI211_X1 U23355 ( .C1(n20476), .C2(n20342), .A(n20341), .B(n20340), .ZN(
        P1_U3111) );
  AOI22_X1 U23356 ( .A1(n20581), .A2(n20344), .B1(n20579), .B2(n20343), .ZN(
        n20348) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20582), .ZN(n20347) );
  OAI211_X1 U23358 ( .C1(n9850), .C2(n20383), .A(n20348), .B(n20347), .ZN(
        P1_U3112) );
  INV_X1 U23359 ( .A(n20487), .ZN(n20349) );
  NAND2_X1 U23360 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20392), .ZN(
        n20399) );
  NOR2_X1 U23361 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20399), .ZN(
        n20355) );
  INV_X1 U23362 ( .A(n20355), .ZN(n20382) );
  OAI22_X1 U23363 ( .A1(n20430), .A2(n20500), .B1(n20382), .B2(n20432), .ZN(
        n20350) );
  INV_X1 U23364 ( .A(n20350), .ZN(n20363) );
  NAND3_X1 U23365 ( .A1(n20430), .A2(n20383), .A3(n20538), .ZN(n20351) );
  NAND2_X1 U23366 ( .A1(n20351), .A2(n20434), .ZN(n20358) );
  NAND2_X1 U23367 ( .A1(n20352), .A2(n20488), .ZN(n20360) );
  OR2_X1 U23368 ( .A1(n20353), .A2(n11318), .ZN(n20489) );
  NAND2_X1 U23369 ( .A1(n20489), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20495) );
  OAI211_X1 U23370 ( .C1(n20439), .C2(n20355), .A(n20495), .B(n20354), .ZN(
        n20356) );
  AOI21_X1 U23371 ( .B1(n20358), .B2(n20360), .A(n20356), .ZN(n20357) );
  INV_X1 U23372 ( .A(n20358), .ZN(n20361) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20386), .B1(
        n20528), .B2(n20385), .ZN(n20362) );
  OAI211_X1 U23374 ( .C1(n20544), .C2(n20383), .A(n20363), .B(n20362), .ZN(
        P1_U3113) );
  OAI22_X1 U23375 ( .A1(n20430), .A2(n20549), .B1(n20382), .B2(n20447), .ZN(
        n20364) );
  INV_X1 U23376 ( .A(n20364), .ZN(n20366) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20386), .B1(
        n20546), .B2(n20385), .ZN(n20365) );
  OAI211_X1 U23378 ( .C1(n9858), .C2(n20383), .A(n20366), .B(n20365), .ZN(
        P1_U3114) );
  OAI22_X1 U23379 ( .A1(n20383), .A2(n20456), .B1(n20382), .B2(n20452), .ZN(
        n20367) );
  INV_X1 U23380 ( .A(n20367), .ZN(n20369) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20386), .B1(
        n20551), .B2(n20385), .ZN(n20368) );
  OAI211_X1 U23382 ( .C1(n20555), .C2(n20430), .A(n20369), .B(n20368), .ZN(
        P1_U3115) );
  OAI22_X1 U23383 ( .A1(n20430), .A2(n20560), .B1(n20382), .B2(n20457), .ZN(
        n20370) );
  INV_X1 U23384 ( .A(n20370), .ZN(n20372) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20386), .B1(
        n20557), .B2(n20385), .ZN(n20371) );
  OAI211_X1 U23386 ( .C1(n9856), .C2(n20383), .A(n20372), .B(n20371), .ZN(
        P1_U3116) );
  OAI22_X1 U23387 ( .A1(n20383), .A2(n20466), .B1(n20382), .B2(n20462), .ZN(
        n20373) );
  INV_X1 U23388 ( .A(n20373), .ZN(n20375) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20386), .B1(
        n20562), .B2(n20385), .ZN(n20374) );
  OAI211_X1 U23390 ( .C1(n20566), .C2(n20430), .A(n20375), .B(n20374), .ZN(
        P1_U3117) );
  OAI22_X1 U23391 ( .A1(n20430), .A2(n20571), .B1(n20382), .B2(n20467), .ZN(
        n20376) );
  INV_X1 U23392 ( .A(n20376), .ZN(n20378) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20386), .B1(
        n20568), .B2(n20385), .ZN(n20377) );
  OAI211_X1 U23394 ( .C1(n9854), .C2(n20383), .A(n20378), .B(n20377), .ZN(
        P1_U3118) );
  OAI22_X1 U23395 ( .A1(n20383), .A2(n20476), .B1(n20382), .B2(n20472), .ZN(
        n20379) );
  INV_X1 U23396 ( .A(n20379), .ZN(n20381) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20386), .B1(
        n20573), .B2(n20385), .ZN(n20380) );
  OAI211_X1 U23398 ( .C1(n9852), .C2(n20430), .A(n20381), .B(n20380), .ZN(
        P1_U3119) );
  OAI22_X1 U23399 ( .A1(n20383), .A2(n20486), .B1(n20382), .B2(n20477), .ZN(
        n20384) );
  INV_X1 U23400 ( .A(n20384), .ZN(n20388) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20386), .B1(
        n20581), .B2(n20385), .ZN(n20387) );
  OAI211_X1 U23402 ( .C1(n9850), .C2(n20430), .A(n20388), .B(n20387), .ZN(
        P1_U3120) );
  NAND2_X1 U23403 ( .A1(n20390), .A2(n20389), .ZN(n20394) );
  NAND2_X1 U23404 ( .A1(n20392), .A2(n20391), .ZN(n20401) );
  OAI21_X1 U23405 ( .B1(n20393), .B2(n20519), .A(n20401), .ZN(n20398) );
  AOI21_X1 U23406 ( .B1(n20395), .B2(n20394), .A(n20398), .ZN(n20397) );
  AOI211_X1 U23407 ( .C1(n20530), .C2(n20399), .A(n20397), .B(n20396), .ZN(
        n20407) );
  INV_X1 U23408 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20727) );
  INV_X1 U23409 ( .A(n20398), .ZN(n20400) );
  OAI22_X1 U23410 ( .A1(n20400), .A2(n20530), .B1(n20399), .B2(n20525), .ZN(
        n20425) );
  INV_X1 U23411 ( .A(n20401), .ZN(n20424) );
  AOI22_X1 U23412 ( .A1(n20528), .A2(n20425), .B1(n20527), .B2(n20424), .ZN(
        n20406) );
  INV_X1 U23413 ( .A(n20402), .ZN(n20403) );
  INV_X1 U23414 ( .A(n20485), .ZN(n20426) );
  INV_X1 U23415 ( .A(n20430), .ZN(n20421) );
  AOI22_X1 U23416 ( .A1(n20426), .A2(n20539), .B1(n20421), .B2(n20497), .ZN(
        n20405) );
  OAI211_X1 U23417 ( .C1(n20407), .C2(n20727), .A(n20406), .B(n20405), .ZN(
        P1_U3121) );
  AOI22_X1 U23418 ( .A1(n20546), .A2(n20425), .B1(n20545), .B2(n20424), .ZN(
        n20410) );
  INV_X1 U23419 ( .A(n20407), .ZN(n20427) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20408), .ZN(n20409) );
  OAI211_X1 U23421 ( .C1(n9858), .C2(n20430), .A(n20410), .B(n20409), .ZN(
        P1_U3122) );
  AOI22_X1 U23422 ( .A1(n20551), .A2(n20425), .B1(n20550), .B2(n20424), .ZN(
        n20413) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20411), .ZN(n20412) );
  OAI211_X1 U23424 ( .C1(n20456), .C2(n20430), .A(n20413), .B(n20412), .ZN(
        P1_U3123) );
  AOI22_X1 U23425 ( .A1(n20557), .A2(n20425), .B1(n20556), .B2(n20424), .ZN(
        n20416) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n20414), .ZN(n20415) );
  OAI211_X1 U23427 ( .C1(n9856), .C2(n20430), .A(n20416), .B(n20415), .ZN(
        P1_U3124) );
  AOI22_X1 U23428 ( .A1(n20562), .A2(n20425), .B1(n20561), .B2(n20424), .ZN(
        n20418) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20427), .B1(
        n20421), .B2(n20563), .ZN(n20417) );
  OAI211_X1 U23430 ( .C1(n20566), .C2(n20485), .A(n20418), .B(n20417), .ZN(
        P1_U3125) );
  AOI22_X1 U23431 ( .A1(n20568), .A2(n20425), .B1(n20567), .B2(n20424), .ZN(
        n20420) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20427), .B1(
        n20421), .B2(n9853), .ZN(n20419) );
  OAI211_X1 U23433 ( .C1(n20571), .C2(n20485), .A(n20420), .B(n20419), .ZN(
        P1_U3126) );
  AOI22_X1 U23434 ( .A1(n20573), .A2(n20425), .B1(n20572), .B2(n20424), .ZN(
        n20423) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20427), .B1(
        n20421), .B2(n20574), .ZN(n20422) );
  OAI211_X1 U23436 ( .C1(n9852), .C2(n20485), .A(n20423), .B(n20422), .ZN(
        P1_U3127) );
  AOI22_X1 U23437 ( .A1(n20581), .A2(n20425), .B1(n20579), .B2(n20424), .ZN(
        n20429) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20427), .B1(
        n20426), .B2(n9849), .ZN(n20428) );
  OAI211_X1 U23439 ( .C1(n20486), .C2(n20430), .A(n20429), .B(n20428), .ZN(
        P1_U3128) );
  OR2_X1 U23440 ( .A1(n20431), .A2(n20523), .ZN(n20478) );
  OAI22_X1 U23441 ( .A1(n20479), .A2(n20500), .B1(n20478), .B2(n20432), .ZN(
        n20433) );
  INV_X1 U23442 ( .A(n20433), .ZN(n20446) );
  INV_X1 U23443 ( .A(n20478), .ZN(n20440) );
  NAND3_X1 U23444 ( .A1(n20485), .A2(n20538), .A3(n20479), .ZN(n20435) );
  NAND2_X1 U23445 ( .A1(n20435), .A2(n20434), .ZN(n20441) );
  NAND2_X1 U23446 ( .A1(n20522), .A2(n20436), .ZN(n20443) );
  INV_X1 U23447 ( .A(n20437), .ZN(n20442) );
  AOI22_X1 U23448 ( .A1(n20441), .A2(n20443), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20442), .ZN(n20438) );
  OAI211_X1 U23449 ( .C1(n20440), .C2(n20439), .A(n20494), .B(n20438), .ZN(
        n20482) );
  INV_X1 U23450 ( .A(n20441), .ZN(n20444) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20482), .B1(
        n20528), .B2(n20481), .ZN(n20445) );
  OAI211_X1 U23452 ( .C1(n20544), .C2(n20485), .A(n20446), .B(n20445), .ZN(
        P1_U3129) );
  OAI22_X1 U23453 ( .A1(n20479), .A2(n20549), .B1(n20478), .B2(n20447), .ZN(
        n20448) );
  INV_X1 U23454 ( .A(n20448), .ZN(n20450) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20482), .B1(
        n20546), .B2(n20481), .ZN(n20449) );
  OAI211_X1 U23456 ( .C1(n9858), .C2(n20485), .A(n20450), .B(n20449), .ZN(
        P1_U3130) );
  OAI22_X1 U23457 ( .A1(n20479), .A2(n20555), .B1(n20478), .B2(n20452), .ZN(
        n20453) );
  INV_X1 U23458 ( .A(n20453), .ZN(n20455) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20482), .B1(
        n20551), .B2(n20481), .ZN(n20454) );
  OAI211_X1 U23460 ( .C1(n20456), .C2(n20485), .A(n20455), .B(n20454), .ZN(
        P1_U3131) );
  OAI22_X1 U23461 ( .A1(n20479), .A2(n20560), .B1(n20478), .B2(n20457), .ZN(
        n20458) );
  INV_X1 U23462 ( .A(n20458), .ZN(n20460) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20482), .B1(
        n20557), .B2(n20481), .ZN(n20459) );
  OAI211_X1 U23464 ( .C1(n9856), .C2(n20485), .A(n20460), .B(n20459), .ZN(
        P1_U3132) );
  OAI22_X1 U23465 ( .A1(n20479), .A2(n20566), .B1(n20478), .B2(n20462), .ZN(
        n20463) );
  INV_X1 U23466 ( .A(n20463), .ZN(n20465) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20482), .B1(
        n20562), .B2(n20481), .ZN(n20464) );
  OAI211_X1 U23468 ( .C1(n20466), .C2(n20485), .A(n20465), .B(n20464), .ZN(
        P1_U3133) );
  OAI22_X1 U23469 ( .A1(n20479), .A2(n20571), .B1(n20478), .B2(n20467), .ZN(
        n20468) );
  INV_X1 U23470 ( .A(n20468), .ZN(n20470) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20482), .B1(
        n20568), .B2(n20481), .ZN(n20469) );
  OAI211_X1 U23472 ( .C1(n9854), .C2(n20485), .A(n20470), .B(n20469), .ZN(
        P1_U3134) );
  OAI22_X1 U23473 ( .A1(n20479), .A2(n9852), .B1(n20478), .B2(n20472), .ZN(
        n20473) );
  INV_X1 U23474 ( .A(n20473), .ZN(n20475) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20482), .B1(
        n20573), .B2(n20481), .ZN(n20474) );
  OAI211_X1 U23476 ( .C1(n20476), .C2(n20485), .A(n20475), .B(n20474), .ZN(
        P1_U3135) );
  OAI22_X1 U23477 ( .A1(n20479), .A2(n9850), .B1(n20478), .B2(n20477), .ZN(
        n20480) );
  INV_X1 U23478 ( .A(n20480), .ZN(n20484) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20482), .B1(
        n20581), .B2(n20481), .ZN(n20483) );
  OAI211_X1 U23480 ( .C1(n20486), .C2(n20485), .A(n20484), .B(n20483), .ZN(
        P1_U3136) );
  NAND2_X1 U23481 ( .A1(n20522), .A2(n20488), .ZN(n20492) );
  OAI22_X1 U23482 ( .A1(n20492), .A2(n20530), .B1(n20490), .B2(n20489), .ZN(
        n20514) );
  NOR3_X2 U23483 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20524), .A3(
        n20523), .ZN(n20513) );
  AOI22_X1 U23484 ( .A1(n20528), .A2(n20514), .B1(n20527), .B2(n20513), .ZN(
        n20499) );
  OAI21_X1 U23485 ( .B1(n20583), .B2(n20515), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20493) );
  AOI21_X1 U23486 ( .B1(n20493), .B2(n20492), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20496) );
  AOI22_X1 U23487 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20515), .B2(n20497), .ZN(n20498) );
  OAI211_X1 U23488 ( .C1(n20500), .C2(n20543), .A(n20499), .B(n20498), .ZN(
        P1_U3145) );
  AOI22_X1 U23489 ( .A1(n20546), .A2(n20514), .B1(n20545), .B2(n20513), .ZN(
        n20502) );
  AOI22_X1 U23490 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20515), .B2(n9857), .ZN(n20501) );
  OAI211_X1 U23491 ( .C1(n20549), .C2(n20543), .A(n20502), .B(n20501), .ZN(
        P1_U3146) );
  AOI22_X1 U23492 ( .A1(n20551), .A2(n20514), .B1(n20550), .B2(n20513), .ZN(
        n20504) );
  AOI22_X1 U23493 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20515), .B2(n20552), .ZN(n20503) );
  OAI211_X1 U23494 ( .C1(n20555), .C2(n20543), .A(n20504), .B(n20503), .ZN(
        P1_U3147) );
  AOI22_X1 U23495 ( .A1(n20557), .A2(n20514), .B1(n20556), .B2(n20513), .ZN(
        n20506) );
  AOI22_X1 U23496 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n20515), .B2(n9855), .ZN(n20505) );
  OAI211_X1 U23497 ( .C1(n20560), .C2(n20543), .A(n20506), .B(n20505), .ZN(
        P1_U3148) );
  AOI22_X1 U23498 ( .A1(n20562), .A2(n20514), .B1(n20561), .B2(n20513), .ZN(
        n20508) );
  AOI22_X1 U23499 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n20515), .B2(n20563), .ZN(n20507) );
  OAI211_X1 U23500 ( .C1(n20566), .C2(n20543), .A(n20508), .B(n20507), .ZN(
        P1_U3149) );
  AOI22_X1 U23501 ( .A1(n20568), .A2(n20514), .B1(n20567), .B2(n20513), .ZN(
        n20510) );
  AOI22_X1 U23502 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20515), .B2(n9853), .ZN(n20509) );
  OAI211_X1 U23503 ( .C1(n20571), .C2(n20543), .A(n20510), .B(n20509), .ZN(
        P1_U3150) );
  AOI22_X1 U23504 ( .A1(n20573), .A2(n20514), .B1(n20572), .B2(n20513), .ZN(
        n20512) );
  AOI22_X1 U23505 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n20515), .B2(n20574), .ZN(n20511) );
  OAI211_X1 U23506 ( .C1(n9852), .C2(n20543), .A(n20512), .B(n20511), .ZN(
        P1_U3151) );
  AOI22_X1 U23507 ( .A1(n20581), .A2(n20514), .B1(n20579), .B2(n20513), .ZN(
        n20518) );
  AOI22_X1 U23508 ( .A1(n20516), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20515), .B2(n20582), .ZN(n20517) );
  OAI211_X1 U23509 ( .C1(n9850), .C2(n20543), .A(n20518), .B(n20517), .ZN(
        P1_U3152) );
  INV_X1 U23510 ( .A(n20519), .ZN(n20521) );
  NOR2_X1 U23511 ( .A1(n20520), .A2(n20523), .ZN(n20578) );
  AOI21_X1 U23512 ( .B1(n20522), .B2(n20521), .A(n20578), .ZN(n20532) );
  NOR2_X1 U23513 ( .A1(n20524), .A2(n20523), .ZN(n20537) );
  INV_X1 U23514 ( .A(n20537), .ZN(n20526) );
  OAI22_X1 U23515 ( .A1(n20532), .A2(n20530), .B1(n20526), .B2(n20525), .ZN(
        n20580) );
  AOI22_X1 U23516 ( .A1(n20528), .A2(n20580), .B1(n20527), .B2(n20578), .ZN(
        n20542) );
  INV_X1 U23517 ( .A(n20529), .ZN(n20531) );
  NOR2_X1 U23518 ( .A1(n20531), .A2(n20530), .ZN(n20534) );
  OAI21_X1 U23519 ( .B1(n20534), .B2(n20533), .A(n20532), .ZN(n20535) );
  OAI211_X1 U23520 ( .C1(n20538), .C2(n20537), .A(n20536), .B(n20535), .ZN(
        n20584) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20584), .B1(
        n20540), .B2(n20539), .ZN(n20541) );
  OAI211_X1 U23522 ( .C1(n20544), .C2(n20543), .A(n20542), .B(n20541), .ZN(
        P1_U3153) );
  AOI22_X1 U23523 ( .A1(n20546), .A2(n20580), .B1(n20545), .B2(n20578), .ZN(
        n20548) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n9857), .ZN(n20547) );
  OAI211_X1 U23525 ( .C1(n20549), .C2(n20587), .A(n20548), .B(n20547), .ZN(
        P1_U3154) );
  AOI22_X1 U23526 ( .A1(n20551), .A2(n20580), .B1(n20550), .B2(n20578), .ZN(
        n20554) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20552), .ZN(n20553) );
  OAI211_X1 U23528 ( .C1(n20555), .C2(n20587), .A(n20554), .B(n20553), .ZN(
        P1_U3155) );
  AOI22_X1 U23529 ( .A1(n20557), .A2(n20580), .B1(n20556), .B2(n20578), .ZN(
        n20559) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n9855), .ZN(n20558) );
  OAI211_X1 U23531 ( .C1(n20560), .C2(n20587), .A(n20559), .B(n20558), .ZN(
        P1_U3156) );
  AOI22_X1 U23532 ( .A1(n20562), .A2(n20580), .B1(n20561), .B2(n20578), .ZN(
        n20565) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20563), .ZN(n20564) );
  OAI211_X1 U23534 ( .C1(n20566), .C2(n20587), .A(n20565), .B(n20564), .ZN(
        P1_U3157) );
  AOI22_X1 U23535 ( .A1(n20568), .A2(n20580), .B1(n20567), .B2(n20578), .ZN(
        n20570) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n9853), .ZN(n20569) );
  OAI211_X1 U23537 ( .C1(n20571), .C2(n20587), .A(n20570), .B(n20569), .ZN(
        P1_U3158) );
  AOI22_X1 U23538 ( .A1(n20573), .A2(n20580), .B1(n20572), .B2(n20578), .ZN(
        n20576) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20574), .ZN(n20575) );
  OAI211_X1 U23540 ( .C1(n9852), .C2(n20587), .A(n20576), .B(n20575), .ZN(
        P1_U3159) );
  AOI22_X1 U23541 ( .A1(n20581), .A2(n20580), .B1(n20579), .B2(n20578), .ZN(
        n20586) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20582), .ZN(n20585) );
  OAI211_X1 U23543 ( .C1(n9850), .C2(n20587), .A(n20586), .B(n20585), .ZN(
        P1_U3160) );
  NOR2_X1 U23544 ( .A1(n20589), .A2(n20684), .ZN(n20591) );
  NAND2_X1 U23545 ( .A1(n20591), .A2(n20590), .ZN(P1_U3163) );
  AND2_X1 U23546 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20664), .ZN(
        P1_U3164) );
  AND2_X1 U23547 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20664), .ZN(
        P1_U3165) );
  AND2_X1 U23548 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20664), .ZN(
        P1_U3166) );
  AND2_X1 U23549 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20664), .ZN(
        P1_U3167) );
  AND2_X1 U23550 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20664), .ZN(
        P1_U3168) );
  AND2_X1 U23551 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20664), .ZN(
        P1_U3169) );
  AND2_X1 U23552 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20664), .ZN(
        P1_U3170) );
  AND2_X1 U23553 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20664), .ZN(
        P1_U3171) );
  AND2_X1 U23554 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20664), .ZN(
        P1_U3172) );
  AND2_X1 U23555 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20664), .ZN(
        P1_U3173) );
  INV_X1 U23556 ( .A(P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20866) );
  NOR2_X1 U23557 ( .A1(n20668), .A2(n20866), .ZN(P1_U3174) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20664), .ZN(
        P1_U3175) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20664), .ZN(
        P1_U3176) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20664), .ZN(
        P1_U3177) );
  INV_X1 U23561 ( .A(P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20901) );
  NOR2_X1 U23562 ( .A1(n20668), .A2(n20901), .ZN(P1_U3178) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20664), .ZN(
        P1_U3179) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20664), .ZN(
        P1_U3180) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20664), .ZN(
        P1_U3181) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20664), .ZN(
        P1_U3182) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20664), .ZN(
        P1_U3183) );
  INV_X1 U23568 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20852) );
  NOR2_X1 U23569 ( .A1(n20668), .A2(n20852), .ZN(P1_U3184) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20664), .ZN(
        P1_U3185) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20664), .ZN(P1_U3186) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20664), .ZN(P1_U3187) );
  AND2_X1 U23573 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20664), .ZN(P1_U3188) );
  AND2_X1 U23574 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20664), .ZN(P1_U3189) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20664), .ZN(P1_U3190) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20664), .ZN(P1_U3191) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20664), .ZN(P1_U3192) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20664), .ZN(P1_U3193) );
  AOI21_X1 U23579 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20593), .A(n20592), 
        .ZN(n20599) );
  INV_X1 U23580 ( .A(n20689), .ZN(n20688) );
  INV_X1 U23581 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20605) );
  NOR2_X1 U23582 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20595) );
  OAI22_X1 U23583 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20598), .B1(n20595), 
        .B2(n20594), .ZN(n20596) );
  NOR2_X1 U23584 ( .A1(n20605), .A2(n20596), .ZN(n20597) );
  OAI22_X1 U23585 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20599), .B1(n20688), 
        .B2(n20597), .ZN(P1_U3194) );
  NAND2_X1 U23586 ( .A1(n20598), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20602) );
  AOI221_X1 U23587 ( .B1(n20609), .B2(n20605), .C1(n20609), .C2(n20602), .A(
        n20599), .ZN(n20600) );
  INV_X1 U23588 ( .A(n20600), .ZN(n20608) );
  OAI21_X1 U23589 ( .B1(n20603), .B2(n20602), .A(n20601), .ZN(n20604) );
  OAI211_X1 U23590 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20605), .A(HOLD), .B(
        n20604), .ZN(n20606) );
  OAI221_X1 U23591 ( .B1(n20608), .B2(NA), .C1(n20608), .C2(n20607), .A(n20606), .ZN(P1_U3196) );
  NAND2_X1 U23592 ( .A1(n20688), .A2(n20609), .ZN(n20655) );
  INV_X1 U23593 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20610) );
  NAND2_X1 U23594 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20688), .ZN(n20651) );
  OAI222_X1 U23595 ( .A1(n20655), .A2(n20612), .B1(n20610), .B2(n20688), .C1(
        n20669), .C2(n20651), .ZN(P1_U3197) );
  INV_X1 U23596 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20611) );
  OAI222_X1 U23597 ( .A1(n20651), .A2(n20612), .B1(n20611), .B2(n20688), .C1(
        n20614), .C2(n20655), .ZN(P1_U3198) );
  OAI222_X1 U23598 ( .A1(n20651), .A2(n20614), .B1(n20613), .B2(n20688), .C1(
        n20615), .C2(n20655), .ZN(P1_U3199) );
  INV_X1 U23599 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20616) );
  OAI222_X1 U23600 ( .A1(n20655), .A2(n13766), .B1(n20616), .B2(n20688), .C1(
        n20615), .C2(n20651), .ZN(P1_U3200) );
  INV_X1 U23601 ( .A(n20655), .ZN(n20649) );
  AOI22_X1 U23602 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20689), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20649), .ZN(n20617) );
  OAI21_X1 U23603 ( .B1(n13766), .B2(n20651), .A(n20617), .ZN(P1_U3201) );
  INV_X1 U23604 ( .A(n20651), .ZN(n20653) );
  AOI22_X1 U23605 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20689), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20653), .ZN(n20618) );
  OAI21_X1 U23606 ( .B1(n20620), .B2(n20655), .A(n20618), .ZN(P1_U3202) );
  INV_X1 U23607 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20619) );
  OAI222_X1 U23608 ( .A1(n20651), .A2(n20620), .B1(n20619), .B2(n20688), .C1(
        n20622), .C2(n20655), .ZN(P1_U3203) );
  INV_X1 U23609 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20621) );
  OAI222_X1 U23610 ( .A1(n20651), .A2(n20622), .B1(n20621), .B2(n20688), .C1(
        n20624), .C2(n20655), .ZN(P1_U3204) );
  INV_X1 U23611 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20623) );
  OAI222_X1 U23612 ( .A1(n20651), .A2(n20624), .B1(n20623), .B2(n20688), .C1(
        n14812), .C2(n20655), .ZN(P1_U3205) );
  INV_X1 U23613 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20625) );
  OAI222_X1 U23614 ( .A1(n20655), .A2(n14888), .B1(n20625), .B2(n20688), .C1(
        n14812), .C2(n20651), .ZN(P1_U3206) );
  AOI22_X1 U23615 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20689), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20649), .ZN(n20626) );
  OAI21_X1 U23616 ( .B1(n14888), .B2(n20651), .A(n20626), .ZN(P1_U3207) );
  AOI22_X1 U23617 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20689), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20653), .ZN(n20627) );
  OAI21_X1 U23618 ( .B1(n20629), .B2(n20655), .A(n20627), .ZN(P1_U3208) );
  INV_X1 U23619 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20628) );
  OAI222_X1 U23620 ( .A1(n20651), .A2(n20629), .B1(n20628), .B2(n20688), .C1(
        n20630), .C2(n20655), .ZN(P1_U3209) );
  INV_X1 U23621 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20887) );
  OAI222_X1 U23622 ( .A1(n20655), .A2(n20796), .B1(n20887), .B2(n20688), .C1(
        n20630), .C2(n20651), .ZN(P1_U3210) );
  INV_X1 U23623 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20631) );
  OAI222_X1 U23624 ( .A1(n20655), .A2(n20633), .B1(n20631), .B2(n20688), .C1(
        n20796), .C2(n20651), .ZN(P1_U3211) );
  AOI22_X1 U23625 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20689), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20649), .ZN(n20632) );
  OAI21_X1 U23626 ( .B1(n20633), .B2(n20651), .A(n20632), .ZN(P1_U3212) );
  AOI22_X1 U23627 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20689), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20653), .ZN(n20634) );
  OAI21_X1 U23628 ( .B1(n14771), .B2(n20655), .A(n20634), .ZN(P1_U3213) );
  INV_X1 U23629 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20635) );
  OAI222_X1 U23630 ( .A1(n20651), .A2(n14771), .B1(n20635), .B2(n20688), .C1(
        n20636), .C2(n20655), .ZN(P1_U3214) );
  INV_X1 U23631 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20637) );
  OAI222_X1 U23632 ( .A1(n20655), .A2(n20639), .B1(n20637), .B2(n20688), .C1(
        n20636), .C2(n20651), .ZN(P1_U3215) );
  INV_X1 U23633 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20638) );
  OAI222_X1 U23634 ( .A1(n20651), .A2(n20639), .B1(n20638), .B2(n20688), .C1(
        n14873), .C2(n20655), .ZN(P1_U3216) );
  INV_X1 U23635 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20640) );
  OAI222_X1 U23636 ( .A1(n20651), .A2(n14873), .B1(n20640), .B2(n20688), .C1(
        n14761), .C2(n20655), .ZN(P1_U3217) );
  INV_X1 U23637 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20957) );
  OAI222_X1 U23638 ( .A1(n20651), .A2(n14761), .B1(n20957), .B2(n20688), .C1(
        n20837), .C2(n20655), .ZN(P1_U3218) );
  AOI22_X1 U23639 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20649), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20689), .ZN(n20641) );
  OAI21_X1 U23640 ( .B1(n20837), .B2(n20651), .A(n20641), .ZN(P1_U3219) );
  AOI22_X1 U23641 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20653), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20689), .ZN(n20642) );
  OAI21_X1 U23642 ( .B1(n20644), .B2(n20655), .A(n20642), .ZN(P1_U3220) );
  AOI22_X1 U23643 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20649), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20689), .ZN(n20643) );
  OAI21_X1 U23644 ( .B1(n20644), .B2(n20651), .A(n20643), .ZN(P1_U3221) );
  AOI22_X1 U23645 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20653), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20689), .ZN(n20645) );
  OAI21_X1 U23646 ( .B1(n20647), .B2(n20655), .A(n20645), .ZN(P1_U3222) );
  AOI22_X1 U23647 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20649), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20689), .ZN(n20646) );
  OAI21_X1 U23648 ( .B1(n20647), .B2(n20651), .A(n20646), .ZN(P1_U3223) );
  AOI22_X1 U23649 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20653), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20689), .ZN(n20648) );
  OAI21_X1 U23650 ( .B1(n20652), .B2(n20655), .A(n20648), .ZN(P1_U3224) );
  AOI22_X1 U23651 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20649), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20689), .ZN(n20650) );
  OAI21_X1 U23652 ( .B1(n20652), .B2(n20651), .A(n20650), .ZN(P1_U3225) );
  AOI22_X1 U23653 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20653), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20689), .ZN(n20654) );
  OAI21_X1 U23654 ( .B1(n20656), .B2(n20655), .A(n20654), .ZN(P1_U3226) );
  INV_X1 U23655 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20657) );
  AOI22_X1 U23656 ( .A1(n20688), .A2(n20658), .B1(n20657), .B2(n20689), .ZN(
        P1_U3458) );
  INV_X1 U23657 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20671) );
  INV_X1 U23658 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20659) );
  AOI22_X1 U23659 ( .A1(n20688), .A2(n20671), .B1(n20659), .B2(n20689), .ZN(
        P1_U3459) );
  INV_X1 U23660 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20660) );
  AOI22_X1 U23661 ( .A1(n20688), .A2(n20661), .B1(n20660), .B2(n20689), .ZN(
        P1_U3460) );
  INV_X1 U23662 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20676) );
  INV_X1 U23663 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20662) );
  AOI22_X1 U23664 ( .A1(n20688), .A2(n20676), .B1(n20662), .B2(n20689), .ZN(
        P1_U3461) );
  INV_X1 U23665 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20665) );
  INV_X1 U23666 ( .A(n20666), .ZN(n20663) );
  AOI21_X1 U23667 ( .B1(n20665), .B2(n20664), .A(n20663), .ZN(P1_U3464) );
  OAI21_X1 U23668 ( .B1(n20668), .B2(n20667), .A(n20666), .ZN(P1_U3465) );
  AOI21_X1 U23669 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20670) );
  AOI22_X1 U23670 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20670), .B2(n20669), .ZN(n20672) );
  AOI22_X1 U23671 ( .A1(n20673), .A2(n20672), .B1(n20671), .B2(n20675), .ZN(
        P1_U3481) );
  NOR2_X1 U23672 ( .A1(n20675), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U23673 ( .A1(n20676), .A2(n20675), .B1(n13254), .B2(n20674), .ZN(
        P1_U3482) );
  AOI22_X1 U23674 ( .A1(n20688), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20746), 
        .B2(n20689), .ZN(P1_U3483) );
  OAI21_X1 U23675 ( .B1(n20677), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20679) );
  OAI22_X1 U23676 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20680), .B1(n20679), 
        .B2(n20678), .ZN(n20687) );
  AOI211_X1 U23677 ( .C1(n20684), .C2(n20683), .A(n20682), .B(n20681), .ZN(
        n20686) );
  NAND2_X1 U23678 ( .A1(n20686), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20685) );
  OAI21_X1 U23679 ( .B1(n20687), .B2(n20686), .A(n20685), .ZN(P1_U3485) );
  OAI22_X1 U23680 ( .A1(n20689), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20688), .ZN(n20690) );
  INV_X1 U23681 ( .A(n20690), .ZN(P1_U3486) );
  NAND2_X1 U23682 ( .A1(n10012), .A2(n20691), .ZN(n20692) );
  XOR2_X1 U23683 ( .A(n20693), .B(n20692), .Z(n20710) );
  AOI22_X1 U23684 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n20694), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19012), .ZN(n20695) );
  OAI21_X1 U23685 ( .B1(n20697), .B2(n20696), .A(n20695), .ZN(n20701) );
  NOR2_X1 U23686 ( .A1(n20699), .A2(n20698), .ZN(n20700) );
  AOI211_X1 U23687 ( .C1(n20703), .C2(n20702), .A(n20701), .B(n20700), .ZN(
        n20704) );
  OAI21_X1 U23688 ( .B1(n13197), .B2(n20705), .A(n20704), .ZN(n20706) );
  AOI21_X1 U23689 ( .B1(n20708), .B2(n20707), .A(n20706), .ZN(n20709) );
  OAI21_X1 U23690 ( .B1(n20710), .B2(n12836), .A(n20709), .ZN(n20971) );
  INV_X1 U23691 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n20712) );
  AOI22_X1 U23692 ( .A1(n20713), .A2(keyinput51), .B1(n20712), .B2(keyinput116), .ZN(n20711) );
  OAI221_X1 U23693 ( .B1(n20713), .B2(keyinput51), .C1(n20712), .C2(
        keyinput116), .A(n20711), .ZN(n20725) );
  INV_X1 U23694 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20715) );
  AOI22_X1 U23695 ( .A1(n20716), .A2(keyinput110), .B1(n20715), .B2(keyinput94), .ZN(n20714) );
  OAI221_X1 U23696 ( .B1(n20716), .B2(keyinput110), .C1(n20715), .C2(
        keyinput94), .A(n20714), .ZN(n20724) );
  AOI22_X1 U23697 ( .A1(n20719), .A2(keyinput52), .B1(keyinput3), .B2(n20718), 
        .ZN(n20717) );
  OAI221_X1 U23698 ( .B1(n20719), .B2(keyinput52), .C1(n20718), .C2(keyinput3), 
        .A(n20717), .ZN(n20723) );
  AOI22_X1 U23699 ( .A1(n20721), .A2(keyinput115), .B1(keyinput25), .B2(n13403), .ZN(n20720) );
  OAI221_X1 U23700 ( .B1(n20721), .B2(keyinput115), .C1(n13403), .C2(
        keyinput25), .A(n20720), .ZN(n20722) );
  NOR4_X1 U23701 ( .A1(n20725), .A2(n20724), .A3(n20723), .A4(n20722), .ZN(
        n20773) );
  AOI22_X1 U23702 ( .A1(n20728), .A2(keyinput23), .B1(keyinput125), .B2(n20727), .ZN(n20726) );
  OAI221_X1 U23703 ( .B1(n20728), .B2(keyinput23), .C1(n20727), .C2(
        keyinput125), .A(n20726), .ZN(n20741) );
  AOI22_X1 U23704 ( .A1(n20731), .A2(keyinput103), .B1(keyinput88), .B2(n20730), .ZN(n20729) );
  OAI221_X1 U23705 ( .B1(n20731), .B2(keyinput103), .C1(n20730), .C2(
        keyinput88), .A(n20729), .ZN(n20740) );
  AOI22_X1 U23706 ( .A1(n20734), .A2(keyinput32), .B1(n20733), .B2(keyinput93), 
        .ZN(n20732) );
  OAI221_X1 U23707 ( .B1(n20734), .B2(keyinput32), .C1(n20733), .C2(keyinput93), .A(n20732), .ZN(n20739) );
  AOI22_X1 U23708 ( .A1(n20737), .A2(keyinput19), .B1(keyinput98), .B2(n20736), 
        .ZN(n20735) );
  OAI221_X1 U23709 ( .B1(n20737), .B2(keyinput19), .C1(n20736), .C2(keyinput98), .A(n20735), .ZN(n20738) );
  NOR4_X1 U23710 ( .A1(n20741), .A2(n20740), .A3(n20739), .A4(n20738), .ZN(
        n20772) );
  AOI22_X1 U23711 ( .A1(n13373), .A2(keyinput5), .B1(keyinput126), .B2(n20743), 
        .ZN(n20742) );
  OAI221_X1 U23712 ( .B1(n13373), .B2(keyinput5), .C1(n20743), .C2(keyinput126), .A(n20742), .ZN(n20755) );
  AOI22_X1 U23713 ( .A1(n20746), .A2(keyinput14), .B1(n20745), .B2(keyinput81), 
        .ZN(n20744) );
  OAI221_X1 U23714 ( .B1(n20746), .B2(keyinput14), .C1(n20745), .C2(keyinput81), .A(n20744), .ZN(n20754) );
  AOI22_X1 U23715 ( .A1(n20749), .A2(keyinput2), .B1(n20748), .B2(keyinput122), 
        .ZN(n20747) );
  OAI221_X1 U23716 ( .B1(n20749), .B2(keyinput2), .C1(n20748), .C2(keyinput122), .A(n20747), .ZN(n20753) );
  INV_X1 U23717 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U23718 ( .A1(n13337), .A2(keyinput41), .B1(keyinput127), .B2(n20751), .ZN(n20750) );
  OAI221_X1 U23719 ( .B1(n13337), .B2(keyinput41), .C1(n20751), .C2(
        keyinput127), .A(n20750), .ZN(n20752) );
  NOR4_X1 U23720 ( .A1(n20755), .A2(n20754), .A3(n20753), .A4(n20752), .ZN(
        n20771) );
  INV_X1 U23721 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20758) );
  AOI22_X1 U23722 ( .A1(n20758), .A2(keyinput43), .B1(keyinput62), .B2(n20757), 
        .ZN(n20756) );
  OAI221_X1 U23723 ( .B1(n20758), .B2(keyinput43), .C1(n20757), .C2(keyinput62), .A(n20756), .ZN(n20769) );
  AOI22_X1 U23724 ( .A1(n20761), .A2(keyinput27), .B1(n20760), .B2(keyinput97), 
        .ZN(n20759) );
  OAI221_X1 U23725 ( .B1(n20761), .B2(keyinput27), .C1(n20760), .C2(keyinput97), .A(n20759), .ZN(n20768) );
  INV_X1 U23726 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20763) );
  AOI22_X1 U23727 ( .A1(n13346), .A2(keyinput79), .B1(keyinput89), .B2(n20763), 
        .ZN(n20762) );
  OAI221_X1 U23728 ( .B1(n13346), .B2(keyinput79), .C1(n20763), .C2(keyinput89), .A(n20762), .ZN(n20767) );
  AOI22_X1 U23729 ( .A1(n20765), .A2(keyinput92), .B1(n11898), .B2(keyinput123), .ZN(n20764) );
  OAI221_X1 U23730 ( .B1(n20765), .B2(keyinput92), .C1(n11898), .C2(
        keyinput123), .A(n20764), .ZN(n20766) );
  NOR4_X1 U23731 ( .A1(n20769), .A2(n20768), .A3(n20767), .A4(n20766), .ZN(
        n20770) );
  NAND4_X1 U23732 ( .A1(n20773), .A2(n20772), .A3(n20771), .A4(n20770), .ZN(
        n20969) );
  AOI22_X1 U23733 ( .A1(n20776), .A2(keyinput28), .B1(keyinput113), .B2(n20775), .ZN(n20774) );
  OAI221_X1 U23734 ( .B1(n20776), .B2(keyinput28), .C1(n20775), .C2(
        keyinput113), .A(n20774), .ZN(n20787) );
  INV_X1 U23735 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U23736 ( .A1(n20779), .A2(keyinput36), .B1(n20778), .B2(keyinput80), 
        .ZN(n20777) );
  OAI221_X1 U23737 ( .B1(n20779), .B2(keyinput36), .C1(n20778), .C2(keyinput80), .A(n20777), .ZN(n20786) );
  AOI22_X1 U23738 ( .A1(n12022), .A2(keyinput100), .B1(keyinput16), .B2(n20781), .ZN(n20780) );
  OAI221_X1 U23739 ( .B1(n12022), .B2(keyinput100), .C1(n20781), .C2(
        keyinput16), .A(n20780), .ZN(n20785) );
  AOI22_X1 U23740 ( .A1(n20783), .A2(keyinput117), .B1(n20983), .B2(
        keyinput112), .ZN(n20782) );
  OAI221_X1 U23741 ( .B1(n20783), .B2(keyinput117), .C1(n20983), .C2(
        keyinput112), .A(n20782), .ZN(n20784) );
  NOR4_X1 U23742 ( .A1(n20787), .A2(n20786), .A3(n20785), .A4(n20784), .ZN(
        n20835) );
  INV_X1 U23743 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U23744 ( .A1(n20789), .A2(keyinput70), .B1(n20984), .B2(keyinput73), 
        .ZN(n20788) );
  OAI221_X1 U23745 ( .B1(n20789), .B2(keyinput70), .C1(n20984), .C2(keyinput73), .A(n20788), .ZN(n20801) );
  AOI22_X1 U23746 ( .A1(n13406), .A2(keyinput0), .B1(keyinput20), .B2(n20791), 
        .ZN(n20790) );
  OAI221_X1 U23747 ( .B1(n13406), .B2(keyinput0), .C1(n20791), .C2(keyinput20), 
        .A(n20790), .ZN(n20800) );
  INV_X1 U23748 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20794) );
  AOI22_X1 U23749 ( .A1(n20794), .A2(keyinput4), .B1(keyinput72), .B2(n20793), 
        .ZN(n20792) );
  OAI221_X1 U23750 ( .B1(n20794), .B2(keyinput4), .C1(n20793), .C2(keyinput72), 
        .A(n20792), .ZN(n20799) );
  AOI22_X1 U23751 ( .A1(n20797), .A2(keyinput78), .B1(n20796), .B2(keyinput26), 
        .ZN(n20795) );
  OAI221_X1 U23752 ( .B1(n20797), .B2(keyinput78), .C1(n20796), .C2(keyinput26), .A(n20795), .ZN(n20798) );
  NOR4_X1 U23753 ( .A1(n20801), .A2(n20800), .A3(n20799), .A4(n20798), .ZN(
        n20834) );
  AOI22_X1 U23754 ( .A1(n20804), .A2(keyinput45), .B1(keyinput68), .B2(n20803), 
        .ZN(n20802) );
  OAI221_X1 U23755 ( .B1(n20804), .B2(keyinput45), .C1(n20803), .C2(keyinput68), .A(n20802), .ZN(n20816) );
  AOI22_X1 U23756 ( .A1(n20807), .A2(keyinput31), .B1(keyinput53), .B2(n20806), 
        .ZN(n20805) );
  OAI221_X1 U23757 ( .B1(n20807), .B2(keyinput31), .C1(n20806), .C2(keyinput53), .A(n20805), .ZN(n20815) );
  INV_X1 U23758 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20985) );
  AOI22_X1 U23759 ( .A1(n20985), .A2(keyinput46), .B1(keyinput67), .B2(n20809), 
        .ZN(n20808) );
  OAI221_X1 U23760 ( .B1(n20985), .B2(keyinput46), .C1(n20809), .C2(keyinput67), .A(n20808), .ZN(n20814) );
  INV_X1 U23761 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20812) );
  AOI22_X1 U23762 ( .A1(n20812), .A2(keyinput37), .B1(keyinput34), .B2(n20811), 
        .ZN(n20810) );
  OAI221_X1 U23763 ( .B1(n20812), .B2(keyinput37), .C1(n20811), .C2(keyinput34), .A(n20810), .ZN(n20813) );
  NOR4_X1 U23764 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        n20833) );
  INV_X1 U23765 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20819) );
  AOI22_X1 U23766 ( .A1(n20819), .A2(keyinput11), .B1(keyinput104), .B2(n20818), .ZN(n20817) );
  OAI221_X1 U23767 ( .B1(n20819), .B2(keyinput11), .C1(n20818), .C2(
        keyinput104), .A(n20817), .ZN(n20831) );
  AOI22_X1 U23768 ( .A1(n20821), .A2(keyinput121), .B1(keyinput118), .B2(
        n11402), .ZN(n20820) );
  OAI221_X1 U23769 ( .B1(n20821), .B2(keyinput121), .C1(n11402), .C2(
        keyinput118), .A(n20820), .ZN(n20830) );
  AOI22_X1 U23770 ( .A1(n20824), .A2(keyinput17), .B1(n20823), .B2(keyinput95), 
        .ZN(n20822) );
  OAI221_X1 U23771 ( .B1(n20824), .B2(keyinput17), .C1(n20823), .C2(keyinput95), .A(n20822), .ZN(n20829) );
  INV_X1 U23772 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20826) );
  AOI22_X1 U23773 ( .A1(n20827), .A2(keyinput108), .B1(n20826), .B2(keyinput49), .ZN(n20825) );
  OAI221_X1 U23774 ( .B1(n20827), .B2(keyinput108), .C1(n20826), .C2(
        keyinput49), .A(n20825), .ZN(n20828) );
  NOR4_X1 U23775 ( .A1(n20831), .A2(n20830), .A3(n20829), .A4(n20828), .ZN(
        n20832) );
  NAND4_X1 U23776 ( .A1(n20835), .A2(n20834), .A3(n20833), .A4(n20832), .ZN(
        n20968) );
  AOI22_X1 U23777 ( .A1(n14761), .A2(keyinput15), .B1(n20837), .B2(keyinput85), 
        .ZN(n20836) );
  OAI221_X1 U23778 ( .B1(n14761), .B2(keyinput15), .C1(n20837), .C2(keyinput85), .A(n20836), .ZN(n20850) );
  AOI22_X1 U23779 ( .A1(n20840), .A2(keyinput69), .B1(keyinput8), .B2(n20839), 
        .ZN(n20838) );
  OAI221_X1 U23780 ( .B1(n20840), .B2(keyinput69), .C1(n20839), .C2(keyinput8), 
        .A(n20838), .ZN(n20849) );
  INV_X1 U23781 ( .A(DATAI_8_), .ZN(n20842) );
  AOI22_X1 U23782 ( .A1(n20843), .A2(keyinput35), .B1(n20842), .B2(keyinput6), 
        .ZN(n20841) );
  OAI221_X1 U23783 ( .B1(n20843), .B2(keyinput35), .C1(n20842), .C2(keyinput6), 
        .A(n20841), .ZN(n20848) );
  INV_X1 U23784 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U23785 ( .A1(n20846), .A2(keyinput87), .B1(n20845), .B2(keyinput119), .ZN(n20844) );
  OAI221_X1 U23786 ( .B1(n20846), .B2(keyinput87), .C1(n20845), .C2(
        keyinput119), .A(n20844), .ZN(n20847) );
  NOR4_X1 U23787 ( .A1(n20850), .A2(n20849), .A3(n20848), .A4(n20847), .ZN(
        n20899) );
  AOI22_X1 U23788 ( .A1(n20853), .A2(keyinput106), .B1(keyinput7), .B2(n20852), 
        .ZN(n20851) );
  OAI221_X1 U23789 ( .B1(n20853), .B2(keyinput106), .C1(n20852), .C2(keyinput7), .A(n20851), .ZN(n20864) );
  AOI22_X1 U23790 ( .A1(n15329), .A2(keyinput63), .B1(keyinput38), .B2(n20855), 
        .ZN(n20854) );
  OAI221_X1 U23791 ( .B1(n15329), .B2(keyinput63), .C1(n20855), .C2(keyinput38), .A(n20854), .ZN(n20863) );
  INV_X1 U23792 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U23793 ( .A1(n20858), .A2(keyinput48), .B1(keyinput101), .B2(n20857), .ZN(n20856) );
  OAI221_X1 U23794 ( .B1(n20858), .B2(keyinput48), .C1(n20857), .C2(
        keyinput101), .A(n20856), .ZN(n20862) );
  INV_X1 U23795 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n20860) );
  AOI22_X1 U23796 ( .A1(n20860), .A2(keyinput102), .B1(n10788), .B2(keyinput44), .ZN(n20859) );
  OAI221_X1 U23797 ( .B1(n20860), .B2(keyinput102), .C1(n10788), .C2(
        keyinput44), .A(n20859), .ZN(n20861) );
  NOR4_X1 U23798 ( .A1(n20864), .A2(n20863), .A3(n20862), .A4(n20861), .ZN(
        n20898) );
  AOI22_X1 U23799 ( .A1(n20867), .A2(keyinput61), .B1(keyinput30), .B2(n20866), 
        .ZN(n20865) );
  OAI221_X1 U23800 ( .B1(n20867), .B2(keyinput61), .C1(n20866), .C2(keyinput30), .A(n20865), .ZN(n20879) );
  AOI22_X1 U23801 ( .A1(n14113), .A2(keyinput22), .B1(keyinput91), .B2(n20869), 
        .ZN(n20868) );
  OAI221_X1 U23802 ( .B1(n14113), .B2(keyinput22), .C1(n20869), .C2(keyinput91), .A(n20868), .ZN(n20878) );
  AOI22_X1 U23803 ( .A1(n20872), .A2(keyinput65), .B1(n20871), .B2(keyinput33), 
        .ZN(n20870) );
  OAI221_X1 U23804 ( .B1(n20872), .B2(keyinput65), .C1(n20871), .C2(keyinput33), .A(n20870), .ZN(n20877) );
  INV_X1 U23805 ( .A(DATAI_10_), .ZN(n20875) );
  AOI22_X1 U23806 ( .A1(n20875), .A2(keyinput75), .B1(keyinput64), .B2(n20874), 
        .ZN(n20873) );
  OAI221_X1 U23807 ( .B1(n20875), .B2(keyinput75), .C1(n20874), .C2(keyinput64), .A(n20873), .ZN(n20876) );
  NOR4_X1 U23808 ( .A1(n20879), .A2(n20878), .A3(n20877), .A4(n20876), .ZN(
        n20897) );
  INV_X1 U23809 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U23810 ( .A1(n20882), .A2(keyinput40), .B1(n20881), .B2(keyinput10), 
        .ZN(n20880) );
  OAI221_X1 U23811 ( .B1(n20882), .B2(keyinput40), .C1(n20881), .C2(keyinput10), .A(n20880), .ZN(n20895) );
  AOI22_X1 U23812 ( .A1(n20885), .A2(keyinput47), .B1(keyinput1), .B2(n20884), 
        .ZN(n20883) );
  OAI221_X1 U23813 ( .B1(n20885), .B2(keyinput47), .C1(n20884), .C2(keyinput1), 
        .A(n20883), .ZN(n20894) );
  AOI22_X1 U23814 ( .A1(n20888), .A2(keyinput96), .B1(keyinput71), .B2(n20887), 
        .ZN(n20886) );
  OAI221_X1 U23815 ( .B1(n20888), .B2(keyinput96), .C1(n20887), .C2(keyinput71), .A(n20886), .ZN(n20893) );
  AOI22_X1 U23816 ( .A1(n20891), .A2(keyinput105), .B1(n20890), .B2(
        keyinput111), .ZN(n20889) );
  OAI221_X1 U23817 ( .B1(n20891), .B2(keyinput105), .C1(n20890), .C2(
        keyinput111), .A(n20889), .ZN(n20892) );
  NOR4_X1 U23818 ( .A1(n20895), .A2(n20894), .A3(n20893), .A4(n20892), .ZN(
        n20896) );
  NAND4_X1 U23819 ( .A1(n20899), .A2(n20898), .A3(n20897), .A4(n20896), .ZN(
        n20967) );
  AOI22_X1 U23820 ( .A1(n20902), .A2(keyinput42), .B1(keyinput90), .B2(n20901), 
        .ZN(n20900) );
  OAI221_X1 U23821 ( .B1(n20902), .B2(keyinput42), .C1(n20901), .C2(keyinput90), .A(n20900), .ZN(n20915) );
  AOI22_X1 U23822 ( .A1(n20905), .A2(keyinput114), .B1(keyinput77), .B2(n20904), .ZN(n20903) );
  OAI221_X1 U23823 ( .B1(n20905), .B2(keyinput114), .C1(n20904), .C2(
        keyinput77), .A(n20903), .ZN(n20914) );
  INV_X1 U23824 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n20908) );
  AOI22_X1 U23825 ( .A1(n20911), .A2(keyinput82), .B1(keyinput83), .B2(n20910), 
        .ZN(n20909) );
  OAI221_X1 U23826 ( .B1(n20911), .B2(keyinput82), .C1(n20910), .C2(keyinput83), .A(n20909), .ZN(n20912) );
  NOR4_X1 U23827 ( .A1(n20915), .A2(n20914), .A3(n20913), .A4(n20912), .ZN(
        n20965) );
  INV_X1 U23828 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20918) );
  AOI22_X1 U23829 ( .A1(n20918), .A2(keyinput29), .B1(keyinput124), .B2(n20917), .ZN(n20916) );
  OAI221_X1 U23830 ( .B1(n20918), .B2(keyinput29), .C1(n20917), .C2(
        keyinput124), .A(n20916), .ZN(n20930) );
  AOI22_X1 U23831 ( .A1(n20921), .A2(keyinput74), .B1(keyinput109), .B2(n20920), .ZN(n20919) );
  OAI221_X1 U23832 ( .B1(n20921), .B2(keyinput74), .C1(n20920), .C2(
        keyinput109), .A(n20919), .ZN(n20929) );
  INV_X1 U23833 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n20923) );
  AOI22_X1 U23834 ( .A1(n20986), .A2(keyinput86), .B1(keyinput107), .B2(n20923), .ZN(n20922) );
  OAI221_X1 U23835 ( .B1(n20986), .B2(keyinput86), .C1(n20923), .C2(
        keyinput107), .A(n20922), .ZN(n20928) );
  AOI22_X1 U23836 ( .A1(n20926), .A2(keyinput54), .B1(keyinput84), .B2(n20925), 
        .ZN(n20924) );
  OAI221_X1 U23837 ( .B1(n20926), .B2(keyinput54), .C1(n20925), .C2(keyinput84), .A(n20924), .ZN(n20927) );
  NOR4_X1 U23838 ( .A1(n20930), .A2(n20929), .A3(n20928), .A4(n20927), .ZN(
        n20964) );
  INV_X1 U23839 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20933) );
  AOI22_X1 U23840 ( .A1(n20933), .A2(keyinput99), .B1(keyinput13), .B2(n20932), 
        .ZN(n20931) );
  OAI221_X1 U23841 ( .B1(n20933), .B2(keyinput99), .C1(n20932), .C2(keyinput13), .A(n20931), .ZN(n20945) );
  AOI22_X1 U23842 ( .A1(n20936), .A2(keyinput58), .B1(keyinput76), .B2(n20935), 
        .ZN(n20934) );
  OAI221_X1 U23843 ( .B1(n20936), .B2(keyinput58), .C1(n20935), .C2(keyinput76), .A(n20934), .ZN(n20944) );
  AOI22_X1 U23844 ( .A1(n20939), .A2(keyinput50), .B1(n20938), .B2(keyinput60), 
        .ZN(n20937) );
  OAI221_X1 U23845 ( .B1(n20939), .B2(keyinput50), .C1(n20938), .C2(keyinput60), .A(n20937), .ZN(n20943) );
  AOI22_X1 U23846 ( .A1(n20941), .A2(keyinput18), .B1(n12298), .B2(keyinput55), 
        .ZN(n20940) );
  OAI221_X1 U23847 ( .B1(n20941), .B2(keyinput18), .C1(n12298), .C2(keyinput55), .A(n20940), .ZN(n20942) );
  NOR4_X1 U23848 ( .A1(n20945), .A2(n20944), .A3(n20943), .A4(n20942), .ZN(
        n20963) );
  AOI22_X1 U23849 ( .A1(n20948), .A2(keyinput21), .B1(n20947), .B2(keyinput59), 
        .ZN(n20946) );
  OAI221_X1 U23850 ( .B1(n20948), .B2(keyinput21), .C1(n20947), .C2(keyinput59), .A(n20946), .ZN(n20961) );
  AOI22_X1 U23851 ( .A1(n20951), .A2(keyinput12), .B1(keyinput9), .B2(n20950), 
        .ZN(n20949) );
  OAI221_X1 U23852 ( .B1(n20951), .B2(keyinput12), .C1(n20950), .C2(keyinput9), 
        .A(n20949), .ZN(n20960) );
  INV_X1 U23853 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20954) );
  AOI22_X1 U23854 ( .A1(n20954), .A2(keyinput39), .B1(keyinput24), .B2(n20953), 
        .ZN(n20952) );
  OAI221_X1 U23855 ( .B1(n20954), .B2(keyinput39), .C1(n20953), .C2(keyinput24), .A(n20952), .ZN(n20959) );
  AOI22_X1 U23856 ( .A1(n20957), .A2(keyinput57), .B1(n20956), .B2(keyinput120), .ZN(n20955) );
  OAI221_X1 U23857 ( .B1(n20957), .B2(keyinput57), .C1(n20956), .C2(
        keyinput120), .A(n20955), .ZN(n20958) );
  NOR4_X1 U23858 ( .A1(n20961), .A2(n20960), .A3(n20959), .A4(n20958), .ZN(
        n20962) );
  NAND4_X1 U23859 ( .A1(n20965), .A2(n20964), .A3(n20963), .A4(n20962), .ZN(
        n20966) );
  NOR4_X1 U23860 ( .A1(n20969), .A2(n20968), .A3(n20967), .A4(n20966), .ZN(
        n20970) );
  XOR2_X1 U23861 ( .A(n20971), .B(n20970), .Z(n21019) );
  NOR4_X1 U23862 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__4__SCAN_IN), .A3(P3_LWORD_REG_0__SCAN_IN), .A4(
        P3_DATAO_REG_16__SCAN_IN), .ZN(n21017) );
  NOR4_X1 U23863 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), 
        .A4(P3_DATAO_REG_0__SCAN_IN), .ZN(n21016) );
  NOR4_X1 U23864 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n20972)
         );
  NAND3_X1 U23865 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20972), .A3(n10788), 
        .ZN(n20978) );
  NOR4_X1 U23866 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A3(P3_REIP_REG_18__SCAN_IN), .A4(
        P3_CODEFETCH_REG_SCAN_IN), .ZN(n20976) );
  NOR4_X1 U23867 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .A3(P3_INSTQUEUE_REG_2__3__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20975) );
  NOR4_X1 U23868 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_EBX_REG_26__SCAN_IN), .A3(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A4(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20974) );
  NOR4_X1 U23869 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        BUF1_REG_14__SCAN_IN), .A3(P2_DATAO_REG_27__SCAN_IN), .A4(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n20973) );
  NAND4_X1 U23870 ( .A1(n20976), .A2(n20975), .A3(n20974), .A4(n20973), .ZN(
        n20977) );
  NOR4_X1 U23871 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(
        P1_EAX_REG_21__SCAN_IN), .A3(n20978), .A4(n20977), .ZN(n21015) );
  NOR4_X1 U23872 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(P1_EBX_REG_4__SCAN_IN), 
        .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(P3_LWORD_REG_3__SCAN_IN), .ZN(
        n20982) );
  NOR4_X1 U23873 ( .A1(P3_ADDRESS_REG_4__SCAN_IN), .A2(
        P3_LWORD_REG_11__SCAN_IN), .A3(P3_UWORD_REG_13__SCAN_IN), .A4(
        P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20981) );
  NOR4_X1 U23874 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(BUF1_REG_4__SCAN_IN), .A3(
        BUF1_REG_2__SCAN_IN), .A4(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20980)
         );
  NOR4_X1 U23875 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_LWORD_REG_5__SCAN_IN), .A3(P1_LWORD_REG_3__SCAN_IN), .A4(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n20979) );
  NAND4_X1 U23876 ( .A1(n20982), .A2(n20981), .A3(n20980), .A4(n20979), .ZN(
        n21013) );
  NOR4_X1 U23877 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .A3(P2_INSTQUEUE_REG_6__0__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20990) );
  NOR4_X1 U23878 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .A3(P2_INSTQUEUE_REG_4__7__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20989) );
  NOR4_X1 U23879 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        BUF1_REG_8__SCAN_IN), .A3(P1_DATAO_REG_12__SCAN_IN), .A4(n20983), .ZN(
        n20988) );
  NOR4_X1 U23880 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20986), .A3(
        n20985), .A4(n20984), .ZN(n20987) );
  NAND4_X1 U23881 ( .A1(n20990), .A2(n20989), .A3(n20988), .A4(n20987), .ZN(
        n21012) );
  NAND4_X1 U23882 ( .A1(P1_EAX_REG_10__SCAN_IN), .A2(P3_REIP_REG_5__SCAN_IN), 
        .A3(P3_DATAWIDTH_REG_28__SCAN_IN), .A4(P2_DATAO_REG_18__SCAN_IN), .ZN(
        n20994) );
  NAND4_X1 U23883 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(P1_EBX_REG_1__SCAN_IN), 
        .A3(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A4(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n20993) );
  NAND4_X1 U23884 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_REIP_REG_22__SCAN_IN), .A3(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A4(
        P1_UWORD_REG_1__SCAN_IN), .ZN(n20992) );
  NAND4_X1 U23885 ( .A1(BUF1_REG_23__SCAN_IN), .A2(P1_DATAO_REG_17__SCAN_IN), 
        .A3(P3_ADDRESS_REG_9__SCAN_IN), .A4(P2_DATAWIDTH_REG_20__SCAN_IN), 
        .ZN(n20991) );
  NOR4_X1 U23886 ( .A1(n20994), .A2(n20993), .A3(n20992), .A4(n20991), .ZN(
        n21010) );
  NAND4_X1 U23887 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_11__0__SCAN_IN), .A3(P3_BE_N_REG_2__SCAN_IN), .A4(
        P2_UWORD_REG_7__SCAN_IN), .ZN(n20998) );
  NAND4_X1 U23888 ( .A1(P2_ADDRESS_REG_0__SCAN_IN), .A2(P1_EAX_REG_13__SCAN_IN), .A3(P3_EBX_REG_4__SCAN_IN), .A4(P2_LWORD_REG_5__SCAN_IN), .ZN(n20997) );
  NAND4_X1 U23889 ( .A1(BUF2_REG_30__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(BUF1_REG_11__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20996) );
  NAND4_X1 U23890 ( .A1(BUF1_REG_13__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(P1_W_R_N_REG_SCAN_IN), .A4(P2_DATAO_REG_6__SCAN_IN), .ZN(n20995)
         );
  NOR4_X1 U23891 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n21009) );
  NAND4_X1 U23892 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__4__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), 
        .A4(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21002) );
  NAND4_X1 U23893 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(P1_DATAWIDTH_REG_17__SCAN_IN), 
        .ZN(n21001) );
  NAND4_X1 U23894 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), 
        .A4(P3_EAX_REG_1__SCAN_IN), .ZN(n21000) );
  NAND4_X1 U23895 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_REIP_REG_1__SCAN_IN), .A3(P3_ADDRESS_REG_8__SCAN_IN), .A4(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20999) );
  NOR4_X1 U23896 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21008) );
  NAND4_X1 U23897 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(
        P3_EAX_REG_28__SCAN_IN), .A3(P1_DATAO_REG_1__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21006) );
  NAND4_X1 U23898 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(DATAI_8_), .A3(
        P2_BYTEENABLE_REG_3__SCAN_IN), .A4(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n21005) );
  NAND4_X1 U23899 ( .A1(P2_EAX_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), 
        .A4(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n21004) );
  NAND4_X1 U23900 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(DATAI_10_), 
        .A3(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n21003) );
  NOR4_X1 U23901 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21007) );
  NAND4_X1 U23902 ( .A1(n21010), .A2(n21009), .A3(n21008), .A4(n21007), .ZN(
        n21011) );
  NOR3_X1 U23903 ( .A1(n21013), .A2(n21012), .A3(n21011), .ZN(n21014) );
  NAND4_X1 U23904 ( .A1(n21017), .A2(n21016), .A3(n21015), .A4(n21014), .ZN(
        n21018) );
  XNOR2_X1 U23905 ( .A(n21019), .B(n21018), .ZN(P2_U2853) );
  AND2_X1 U11593 ( .A1(n10888), .A2(n10887), .ZN(n11887) );
  CLKBUF_X1 U11165 ( .A(n10988), .Z(n11929) );
  INV_X1 U15432 ( .A(n12410), .ZN(n17174) );
  NAND2_X1 U11565 ( .A1(n15152), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14278) );
  INV_X2 U11503 ( .A(n9761), .ZN(n13143) );
  AOI21_X2 U11535 ( .B1(n12162), .B2(n12161), .A(n13026), .ZN(n12377) );
  CLKBUF_X1 U11150 ( .A(n11080), .Z(n11063) );
  CLKBUF_X1 U11163 ( .A(n11015), .Z(n11369) );
  CLKBUF_X1 U11177 ( .A(n11421), .Z(n11446) );
  CLKBUF_X1 U11181 ( .A(n11117), .Z(n9726) );
  AND2_X1 U11198 ( .A1(n10948), .A2(n9728), .ZN(n10955) );
  INV_X1 U11200 ( .A(n12172), .ZN(n10249) );
  CLKBUF_X1 U11209 ( .A(n10479), .Z(n19269) );
  CLKBUF_X1 U11247 ( .A(n11299), .Z(n9750) );
  CLKBUF_X1 U11286 ( .A(n13556), .Z(n9755) );
  CLKBUF_X1 U11359 ( .A(n10481), .Z(n15647) );
  NOR2_X1 U11472 ( .A1(n16405), .A2(n16584), .ZN(n16404) );
  CLKBUF_X1 U11510 ( .A(n14612), .Z(n14613) );
  CLKBUF_X1 U11511 ( .A(n16494), .Z(n16509) );
  AND2_X2 U11531 ( .A1(n13503), .A2(n10888), .ZN(n10988) );
  XNOR2_X1 U11555 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12872), .ZN(
        n21020) );
  CLKBUF_X1 U11562 ( .A(n10945), .Z(n13574) );
endmodule

