

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9680, n9681, n9682, n9683, n9684, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12336, n12337, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753;

  BUF_X1 U11124 ( .A(n19798), .Z(n9682) );
  NAND2_X1 U11125 ( .A1(n14548), .A2(n14550), .ZN(n20155) );
  NAND3_X1 U11126 ( .A1(n10612), .A2(n10220), .A3(n10613), .ZN(n10142) );
  XNOR2_X1 U11128 ( .A(n13851), .B(n17149), .ZN(n17145) );
  BUF_X2 U11129 ( .A(n12177), .Z(n9681) );
  INV_X1 U11130 ( .A(n19818), .ZN(n11158) );
  NAND2_X1 U11131 ( .A1(n12785), .A2(n12784), .ZN(n13394) );
  CLKBUF_X2 U11132 ( .A(n11672), .Z(n9687) );
  BUF_X2 U11133 ( .A(n11125), .Z(n11126) );
  AND3_X1 U11134 ( .A1(n18641), .A2(n9717), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18536) );
  NAND2_X1 U11135 ( .A1(n10861), .A2(n10862), .ZN(n11132) );
  BUF_X1 U11136 ( .A(n12662), .Z(n14051) );
  BUF_X2 U11137 ( .A(n11998), .Z(n18105) );
  CLKBUF_X2 U11138 ( .A(n12619), .Z(n13264) );
  NOR2_X1 U11139 ( .A1(n13911), .A2(n12632), .ZN(n12676) );
  CLKBUF_X2 U11140 ( .A(n11946), .Z(n9693) );
  AND2_X2 U11141 ( .A1(n11189), .A2(n11006), .ZN(n11250) );
  AND2_X2 U11142 ( .A1(n12463), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11244) );
  CLKBUF_X3 U11144 ( .A(n18056), .Z(n18104) );
  NOR2_X1 U11145 ( .A1(n11078), .A2(n11096), .ZN(n11079) );
  AND2_X2 U11146 ( .A1(n12316), .A2(n11006), .ZN(n11306) );
  INV_X1 U11147 ( .A(n9778), .ZN(n18112) );
  OR2_X1 U11148 ( .A1(n11923), .A2(n17750), .ZN(n18016) );
  CLKBUF_X2 U11149 ( .A(n11946), .Z(n9688) );
  OR2_X1 U11150 ( .A1(n19536), .A2(n11924), .ZN(n17988) );
  INV_X2 U11151 ( .A(n14173), .ZN(n12658) );
  NAND2_X1 U11152 ( .A1(n12163), .A2(n12161), .ZN(n11920) );
  INV_X2 U11153 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12161) );
  AND2_X2 U11155 ( .A1(n12516), .A2(n14489), .ZN(n12740) );
  AND2_X2 U11156 ( .A1(n14676), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12316) );
  AND2_X2 U11157 ( .A1(n14676), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9711) );
  AND2_X1 U11158 ( .A1(n10214), .A2(n10002), .ZN(n9750) );
  AND2_X1 U11159 ( .A1(n11391), .A2(n11611), .ZN(n11425) );
  NAND2_X1 U11160 ( .A1(n12654), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12687) );
  AND2_X2 U11161 ( .A1(n14676), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9710) );
  INV_X1 U11163 ( .A(n13454), .ZN(n12639) );
  AOI21_X1 U11164 ( .B1(n10866), .B2(n10610), .A(n10609), .ZN(n10608) );
  NAND2_X1 U11165 ( .A1(n11026), .A2(n11027), .ZN(n11836) );
  NOR2_X1 U11166 ( .A1(n18502), .A2(n18859), .ZN(n18513) );
  INV_X1 U11167 ( .A(n14055), .ZN(n15267) );
  OR2_X1 U11168 ( .A1(n15565), .A2(n13892), .ZN(n10051) );
  NAND3_X2 U11169 ( .A1(n12799), .A2(n10345), .A3(n12798), .ZN(n10298) );
  NAND2_X1 U11170 ( .A1(n9943), .A2(n13850), .ZN(n13851) );
  INV_X2 U11171 ( .A(n13754), .ZN(n11876) );
  NOR2_X1 U11173 ( .A1(n14813), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U11174 ( .A1(n9988), .A2(n9987), .ZN(n16676) );
  INV_X1 U11175 ( .A(n11836), .ZN(n19869) );
  NAND3_X1 U11176 ( .A1(n18476), .A2(n10592), .A3(n9977), .ZN(n18455) );
  NOR2_X1 U11178 ( .A1(n13950), .A2(n15893), .ZN(n15863) );
  NAND3_X1 U11179 ( .A1(n12633), .A2(n14587), .A3(n12632), .ZN(n15918) );
  CLKBUF_X2 U11180 ( .A(n9698), .Z(n19879) );
  INV_X1 U11183 ( .A(n19930), .ZN(n20403) );
  NAND2_X1 U11184 ( .A1(n18536), .A2(n17208), .ZN(n18520) );
  NOR2_X1 U11185 ( .A1(n19047), .A2(n17080), .ZN(n17133) );
  INV_X1 U11186 ( .A(n20637), .ZN(n15294) );
  AND2_X1 U11187 ( .A1(n15070), .A2(n10842), .ZN(n15012) );
  OR2_X1 U11188 ( .A1(n12601), .A2(n12600), .ZN(n14587) );
  BUF_X1 U11189 ( .A(n15437), .Z(n15438) );
  NAND2_X2 U11190 ( .A1(n11080), .A2(n11402), .ZN(n15939) );
  OAI21_X1 U11191 ( .B1(n16485), .B2(n10433), .A(n13633), .ZN(n13597) );
  OAI21_X1 U11193 ( .B1(n17045), .B2(n17044), .A(n17043), .ZN(n19897) );
  NOR2_X1 U11194 ( .A1(n20398), .A2(n20058), .ZN(n20108) );
  INV_X1 U11195 ( .A(n20295), .ZN(n20271) );
  INV_X1 U11196 ( .A(n20389), .ZN(n20339) );
  NOR2_X1 U11197 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17513), .ZN(n17496) );
  NAND2_X1 U11198 ( .A1(n17138), .A2(n10706), .ZN(n18147) );
  NOR2_X1 U11199 ( .A1(n17262), .A2(n18776), .ZN(n18684) );
  NAND2_X1 U11200 ( .A1(n9690), .A2(n18626), .ZN(n18767) );
  NAND2_X1 U11201 ( .A1(n13408), .A2(n14884), .ZN(n15269) );
  OR2_X1 U11202 ( .A1(n17101), .A2(n13970), .ZN(n15671) );
  AOI21_X1 U11203 ( .B1(n17037), .B2(n17044), .A(n17036), .ZN(n19900) );
  NAND2_X1 U11204 ( .A1(n20095), .A2(n20336), .ZN(n20154) );
  NAND2_X1 U11205 ( .A1(n20337), .A2(n20160), .ZN(n20194) );
  NAND2_X1 U11206 ( .A1(n20337), .A2(n20336), .ZN(n21750) );
  INV_X1 U11207 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20300) );
  INV_X1 U11208 ( .A(n18669), .ZN(n18687) );
  AND2_X1 U11209 ( .A1(n11628), .A2(n11115), .ZN(n13754) );
  AND2_X1 U11211 ( .A1(n16647), .A2(n16637), .ZN(n9680) );
  AND4_X4 U11212 ( .A1(n12542), .A2(n12541), .A3(n12540), .A4(n12539), .ZN(
        n20812) );
  AND4_X2 U11213 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n12541) );
  NAND2_X2 U11214 ( .A1(n10621), .A2(n11270), .ZN(n11346) );
  INV_X2 U11215 ( .A(n12210), .ZN(n10864) );
  NAND2_X2 U11216 ( .A1(n11430), .A2(n9741), .ZN(n11438) );
  INV_X2 U11217 ( .A(n11431), .ZN(n11430) );
  NAND2_X2 U11218 ( .A1(n16676), .A2(n16673), .ZN(n10075) );
  AOI211_X2 U11219 ( .C1(n15006), .C2(n15446), .A(n15005), .B(n15004), .ZN(
        n15007) );
  AND4_X2 U11220 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11038), .ZN(
        n11042) );
  NAND2_X2 U11221 ( .A1(n9974), .A2(n10417), .ZN(n11974) );
  INV_X4 U11222 ( .A(n11974), .ZN(n12075) );
  XNOR2_X2 U11223 ( .A(n13530), .B(n13529), .ZN(n15300) );
  AOI211_X2 U11224 ( .C1(n19809), .C2(n16141), .A(n16140), .B(n16139), .ZN(
        n16142) );
  NOR2_X4 U11225 ( .A1(n17584), .A2(n17659), .ZN(n18641) );
  NAND2_X1 U11227 ( .A1(n10298), .A2(n13805), .ZN(n9697) );
  NOR2_X2 U11228 ( .A1(n16844), .A2(n10556), .ZN(n16754) );
  XNOR2_X1 U11229 ( .A(n12892), .B(n12891), .ZN(n20852) );
  NAND2_X1 U11230 ( .A1(n9779), .A2(n18780), .ZN(n18416) );
  AND2_X2 U11231 ( .A1(n12154), .A2(n10764), .ZN(n9779) );
  NOR3_X2 U11232 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17737) );
  AND2_X2 U11234 ( .A1(n15008), .A2(n10391), .ZN(n14866) );
  NOR2_X4 U11235 ( .A1(n15021), .A2(n15023), .ZN(n15008) );
  BUF_X2 U11236 ( .A(n11169), .Z(n9683) );
  NOR2_X1 U11237 ( .A1(n18267), .A2(n17267), .ZN(n9684) );
  NAND2_X2 U11238 ( .A1(n10074), .A2(n11340), .ZN(n11345) );
  XNOR2_X2 U11239 ( .A(n9996), .B(n11271), .ZN(n10066) );
  XNOR2_X2 U11240 ( .A(n12134), .B(n12133), .ZN(n18711) );
  AND2_X2 U11241 ( .A1(n10664), .A2(n9807), .ZN(n12134) );
  INV_X2 U11242 ( .A(n16704), .ZN(n11180) );
  NAND2_X2 U11243 ( .A1(n9951), .A2(n9949), .ZN(n9948) );
  NOR2_X1 U11244 ( .A1(n19778), .A2(n19820), .ZN(n9686) );
  INV_X2 U11245 ( .A(n19764), .ZN(n16195) );
  NAND2_X1 U11246 ( .A1(n11380), .A2(n16811), .ZN(n16562) );
  NAND2_X1 U11247 ( .A1(n16485), .A2(n10487), .ZN(n10226) );
  AOI21_X1 U11248 ( .B1(n10143), .B2(n9680), .A(n10270), .ZN(n10380) );
  NAND2_X1 U11249 ( .A1(n10057), .A2(n10281), .ZN(n10128) );
  OR2_X1 U11250 ( .A1(n14870), .A2(n15573), .ZN(n10780) );
  NAND2_X1 U11251 ( .A1(n10219), .A2(n16661), .ZN(n10057) );
  AND2_X1 U11252 ( .A1(n9810), .A2(n16647), .ZN(n13600) );
  NAND3_X1 U11253 ( .A1(n10204), .A2(n16937), .A3(n10203), .ZN(n16647) );
  CLKBUF_X1 U11254 ( .A(n16014), .Z(n16025) );
  AND2_X1 U11255 ( .A1(n10871), .A2(n10870), .ZN(n10868) );
  AND3_X1 U11256 ( .A1(n13777), .A2(n13585), .A3(n16518), .ZN(n10871) );
  AOI21_X1 U11257 ( .B1(n9794), .B2(n10051), .A(n15621), .ZN(n10050) );
  AOI21_X1 U11258 ( .B1(n10747), .B2(n9970), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U11259 ( .A1(n20155), .A2(n20116), .ZN(n20337) );
  NAND2_X1 U11260 ( .A1(n12293), .A2(n9902), .ZN(n16305) );
  NOR2_X2 U11261 ( .A1(n14540), .A2(n14539), .ZN(n14538) );
  NAND2_X1 U11262 ( .A1(n14548), .A2(n10859), .ZN(n14653) );
  NAND2_X1 U11263 ( .A1(n15012), .A2(n14999), .ZN(n14871) );
  NOR2_X1 U11264 ( .A1(n10040), .A2(n10342), .ZN(n11176) );
  INV_X1 U11265 ( .A(n18767), .ZN(n18761) );
  OAI22_X1 U11266 ( .A1(n20202), .A2(n10343), .B1(n11165), .B2(n11289), .ZN(
        n10342) );
  OR2_X1 U11267 ( .A1(n9697), .A2(n15879), .ZN(n15552) );
  OR2_X1 U11268 ( .A1(n14522), .A2(n14523), .ZN(n12225) );
  NAND2_X1 U11269 ( .A1(n10648), .A2(n11164), .ZN(n11289) );
  OR2_X1 U11270 ( .A1(n11150), .A2(n9704), .ZN(n20391) );
  AOI21_X1 U11271 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18521), .A(
        n19455), .ZN(n18588) );
  INV_X1 U11272 ( .A(n18521), .ZN(n9690) );
  NAND2_X1 U11273 ( .A1(n11178), .A2(n10647), .ZN(n11185) );
  NAND2_X1 U11275 ( .A1(n11538), .A2(n11537), .ZN(n14655) );
  OR2_X1 U11276 ( .A1(n15118), .A2(n15119), .ZN(n15120) );
  INV_X2 U11278 ( .A(n18772), .ZN(n18728) );
  NAND2_X1 U11279 ( .A1(n19715), .A2(n18880), .ZN(n18820) );
  NOR2_X2 U11280 ( .A1(n19030), .A2(n19544), .ZN(n18880) );
  NAND2_X1 U11282 ( .A1(n10636), .A2(n12765), .ZN(n12899) );
  NAND2_X1 U11283 ( .A1(n11114), .A2(n11113), .ZN(n11142) );
  AOI21_X1 U11284 ( .B1(n11125), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11108), .ZN(n11114) );
  NOR2_X1 U11285 ( .A1(n18750), .A2(n18751), .ZN(n18749) );
  OR2_X1 U11286 ( .A1(n14580), .A2(n12659), .ZN(n13928) );
  NAND2_X1 U11287 ( .A1(n11072), .A2(n10015), .ZN(n11837) );
  INV_X1 U11288 ( .A(n12118), .ZN(n18298) );
  AND2_X1 U11289 ( .A1(n10011), .A2(n10014), .ZN(n11072) );
  NAND2_X1 U11290 ( .A1(n11078), .A2(n11829), .ZN(n11105) );
  AND2_X1 U11291 ( .A1(n12640), .A2(n13937), .ZN(n14174) );
  INV_X4 U11292 ( .A(n19879), .ZN(n13593) );
  BUF_X1 U11293 ( .A(n13522), .Z(n13518) );
  CLKBUF_X1 U11294 ( .A(n11015), .Z(n19875) );
  CLKBUF_X1 U11295 ( .A(n11081), .Z(n12213) );
  NAND2_X1 U11296 ( .A1(n11651), .A2(n11650), .ZN(n11765) );
  NAND2_X1 U11297 ( .A1(n11074), .A2(n11385), .ZN(n11402) );
  OR2_X1 U11298 ( .A1(n11074), .A2(n11385), .ZN(n11080) );
  BUF_X2 U11299 ( .A(n13432), .Z(n13522) );
  NAND2_X2 U11300 ( .A1(n9720), .A2(n10371), .ZN(n18197) );
  INV_X2 U11301 ( .A(n11378), .ZN(n13641) );
  INV_X2 U11302 ( .A(n14163), .ZN(n13433) );
  INV_X1 U11303 ( .A(n14297), .ZN(n12636) );
  CLKBUF_X2 U11304 ( .A(n11063), .Z(n14813) );
  INV_X1 U11305 ( .A(n20812), .ZN(n12632) );
  NAND2_X1 U11306 ( .A1(n13430), .A2(n12637), .ZN(n13454) );
  NAND2_X2 U11307 ( .A1(n11001), .A2(n11000), .ZN(n11064) );
  NAND2_X2 U11308 ( .A1(n14173), .A2(n20812), .ZN(n14054) );
  INV_X2 U11309 ( .A(n14566), .ZN(n13916) );
  AND4_X1 U11310 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(
        n11374) );
  MUX2_X1 U11311 ( .A(n10977), .B(n10976), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11063) );
  AND4_X1 U11312 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        n12551) );
  AND4_X1 U11313 ( .A1(n12546), .A2(n12545), .A3(n12544), .A4(n12543), .ZN(
        n12552) );
  INV_X2 U11314 ( .A(n17988), .ZN(n18113) );
  INV_X2 U11315 ( .A(n18058), .ZN(n9696) );
  AND2_X2 U11316 ( .A1(n9700), .A2(n11006), .ZN(n11222) );
  AND2_X2 U11317 ( .A1(n11190), .A2(n10954), .ZN(n11245) );
  CLKBUF_X2 U11318 ( .A(n12740), .Z(n13123) );
  BUF_X2 U11319 ( .A(n12748), .Z(n13221) );
  INV_X2 U11320 ( .A(n17988), .ZN(n18017) );
  CLKBUF_X2 U11321 ( .A(n12612), .Z(n12719) );
  INV_X2 U11323 ( .A(n18058), .ZN(n18107) );
  BUF_X2 U11324 ( .A(n12713), .Z(n13297) );
  CLKBUF_X2 U11325 ( .A(n12757), .Z(n13177) );
  CLKBUF_X2 U11326 ( .A(n12733), .Z(n13315) );
  CLKBUF_X2 U11327 ( .A(n12618), .Z(n13124) );
  NOR2_X1 U11328 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17730), .ZN(n17710) );
  AND2_X2 U11329 ( .A1(n12516), .A2(n12515), .ZN(n12713) );
  CLKBUF_X2 U11330 ( .A(n12617), .Z(n13317) );
  NAND2_X1 U11331 ( .A1(n12163), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11923) );
  AND2_X2 U11332 ( .A1(n11186), .A2(n10954), .ZN(n11043) );
  AND2_X2 U11333 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14178) );
  AND2_X1 U11334 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12515) );
  NAND3_X4 U11335 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12315) );
  OR2_X1 U11336 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17750) );
  AND2_X1 U11337 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19528) );
  NAND2_X1 U11338 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18740) );
  AND2_X1 U11339 ( .A1(n13794), .A2(n13793), .ZN(n13795) );
  AOI21_X1 U11340 ( .B1(n10711), .B2(n10710), .A(n10707), .ZN(n16494) );
  OAI21_X1 U11341 ( .B1(n16834), .B2(n17193), .A(n10339), .ZN(n10338) );
  OAI21_X1 U11342 ( .B1(n16820), .B2(n10470), .A(n10469), .ZN(n10468) );
  AND2_X1 U11343 ( .A1(n10178), .A2(n10177), .ZN(n16786) );
  OAI21_X1 U11344 ( .B1(n16820), .B2(n10413), .A(n10412), .ZN(n10623) );
  NAND2_X1 U11345 ( .A1(n10241), .A2(n16495), .ZN(n10240) );
  AND2_X1 U11346 ( .A1(n13801), .A2(n13800), .ZN(n13802) );
  AND2_X1 U11347 ( .A1(n10159), .A2(n10160), .ZN(n10158) );
  NAND2_X1 U11348 ( .A1(n10094), .A2(n9739), .ZN(n10494) );
  INV_X1 U11349 ( .A(n10161), .ZN(n16820) );
  NAND2_X1 U11350 ( .A1(n10145), .A2(n13775), .ZN(n16509) );
  NAND2_X1 U11351 ( .A1(n9852), .A2(n10223), .ZN(n13664) );
  NAND2_X1 U11352 ( .A1(n10226), .A2(n13644), .ZN(n13745) );
  OAI21_X1 U11353 ( .B1(n9791), .B2(n10502), .A(n10501), .ZN(n11596) );
  XNOR2_X1 U11354 ( .A(n14913), .B(n10555), .ZN(n10421) );
  NAND2_X1 U11355 ( .A1(n16629), .A2(n10600), .ZN(n10141) );
  AOI21_X1 U11356 ( .B1(n14914), .B2(n14926), .A(n14913), .ZN(n14935) );
  OAI21_X1 U11357 ( .B1(n16562), .B2(n17193), .A(n10471), .ZN(n10161) );
  NAND2_X1 U11358 ( .A1(n10110), .A2(n9742), .ZN(n10109) );
  NAND2_X1 U11359 ( .A1(n16629), .A2(n9776), .ZN(n16588) );
  NAND2_X1 U11360 ( .A1(n10312), .A2(n9882), .ZN(n10311) );
  NAND2_X1 U11361 ( .A1(n10004), .A2(n10869), .ZN(n16517) );
  AOI21_X1 U11362 ( .B1(n10503), .B2(n11868), .A(n16680), .ZN(n10501) );
  NAND2_X1 U11363 ( .A1(n16583), .A2(n16584), .ZN(n16582) );
  AND2_X1 U11364 ( .A1(n16510), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16500) );
  NAND2_X1 U11365 ( .A1(n16510), .A2(n9914), .ZN(n16491) );
  AOI21_X1 U11366 ( .B1(n16481), .B2(n16715), .A(n16480), .ZN(n10643) );
  AND2_X1 U11367 ( .A1(n13632), .A2(n9854), .ZN(n10593) );
  AND2_X1 U11368 ( .A1(n10308), .A2(n10307), .ZN(n15685) );
  AND3_X2 U11369 ( .A1(n10264), .A2(n10095), .A3(n9820), .ZN(n16485) );
  AND2_X1 U11370 ( .A1(n10173), .A2(n9862), .ZN(n10176) );
  NAND2_X1 U11371 ( .A1(n10380), .A2(n10737), .ZN(n11380) );
  AND2_X1 U11372 ( .A1(n10192), .A2(n10917), .ZN(n11530) );
  OAI21_X1 U11373 ( .B1(n16664), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10381), .ZN(n16953) );
  OR2_X1 U11374 ( .A1(n15966), .A2(n15965), .ZN(n16721) );
  NAND2_X1 U11375 ( .A1(n10384), .A2(n10383), .ZN(n10125) );
  NAND2_X1 U11376 ( .A1(n10912), .A2(n10914), .ZN(n10910) );
  XNOR2_X1 U11377 ( .A(n16278), .B(n16277), .ZN(n16391) );
  NAND2_X1 U11378 ( .A1(n13553), .A2(n16584), .ZN(n10872) );
  NAND2_X1 U11379 ( .A1(n10057), .A2(n11483), .ZN(n16594) );
  OR2_X1 U11380 ( .A1(n12439), .A2(n10848), .ZN(n10847) );
  AND2_X1 U11381 ( .A1(n10057), .A2(n10235), .ZN(n13553) );
  NAND2_X1 U11382 ( .A1(n10028), .A2(n10027), .ZN(n10849) );
  AND2_X1 U11383 ( .A1(n10189), .A2(n10282), .ZN(n10281) );
  AND2_X1 U11384 ( .A1(n13600), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10248) );
  NAND2_X1 U11385 ( .A1(n10099), .A2(n10299), .ZN(n10189) );
  NAND2_X1 U11386 ( .A1(n12425), .A2(n12424), .ZN(n16271) );
  XNOR2_X1 U11387 ( .A(n14983), .B(n13341), .ZN(n14876) );
  NAND2_X1 U11388 ( .A1(n12407), .A2(n10029), .ZN(n12425) );
  AND2_X1 U11389 ( .A1(n15470), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15481) );
  OAI21_X1 U11390 ( .B1(n10499), .B2(n9831), .A(n10497), .ZN(n10496) );
  CLKBUF_X1 U11391 ( .A(n15021), .Z(n15022) );
  NAND2_X1 U11392 ( .A1(n9992), .A2(n16966), .ZN(n16673) );
  AND3_X1 U11393 ( .A1(n15168), .A2(n15196), .A3(n15216), .ZN(n15197) );
  NAND2_X1 U11394 ( .A1(n10491), .A2(n16224), .ZN(n16668) );
  INV_X1 U11395 ( .A(n11346), .ZN(n10430) );
  NAND2_X1 U11396 ( .A1(n10056), .A2(n11343), .ZN(n10612) );
  NAND3_X1 U11397 ( .A1(n10377), .A2(n11346), .A3(n10376), .ZN(n16674) );
  XNOR2_X1 U11398 ( .A(n10615), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16637) );
  NAND2_X1 U11399 ( .A1(n10018), .A2(n11270), .ZN(n10017) );
  NAND2_X1 U11400 ( .A1(n9995), .A2(n10621), .ZN(n10220) );
  NAND2_X1 U11401 ( .A1(n18429), .A2(n10588), .ZN(n17216) );
  AND2_X1 U11402 ( .A1(n11343), .A2(n13750), .ZN(n10336) );
  NAND2_X1 U11403 ( .A1(n9848), .A2(n10428), .ZN(n18430) );
  XNOR2_X1 U11404 ( .A(n9965), .B(n19675), .ZN(n17260) );
  NOR2_X2 U11405 ( .A1(n17032), .A2(n20398), .ZN(n21746) );
  AND2_X1 U11406 ( .A1(n9996), .A2(n11345), .ZN(n9995) );
  NOR2_X1 U11407 ( .A1(n11345), .A2(n13750), .ZN(n10130) );
  INV_X1 U11408 ( .A(n9922), .ZN(n9921) );
  AOI22_X1 U11409 ( .A1(n18756), .A2(n18802), .B1(n18684), .B2(n18800), .ZN(
        n18469) );
  NAND2_X1 U11410 ( .A1(n20095), .A2(n20306), .ZN(n20074) );
  AND2_X1 U11411 ( .A1(n13893), .A2(n9911), .ZN(n10320) );
  INV_X1 U11412 ( .A(n14822), .ZN(n10798) );
  NOR2_X2 U11413 ( .A1(n20023), .A2(n19961), .ZN(n20019) );
  XNOR2_X1 U11414 ( .A(n13747), .B(n13645), .ZN(n13725) );
  INV_X1 U11415 ( .A(n10051), .ZN(n13893) );
  NOR2_X2 U11416 ( .A1(n19909), .A2(n20023), .ZN(n19956) );
  OR2_X1 U11417 ( .A1(n16305), .A2(n12348), .ZN(n12349) );
  INV_X1 U11418 ( .A(n10685), .ZN(n11270) );
  NAND2_X1 U11419 ( .A1(n13637), .A2(n13636), .ZN(n13747) );
  NAND2_X1 U11420 ( .A1(n20155), .A2(n20116), .ZN(n20023) );
  AND2_X1 U11421 ( .A1(n15554), .A2(n13888), .ZN(n10325) );
  AOI221_X1 U11422 ( .B1(n18818), .B2(n19544), .C1(n18817), .C2(n19544), .A(
        n18856), .ZN(n18819) );
  AND2_X1 U11423 ( .A1(n12204), .A2(n9886), .ZN(n10429) );
  NAND4_X1 U11424 ( .A1(n9978), .A2(n9805), .A3(n9980), .A4(n9979), .ZN(n10787) );
  AND2_X1 U11425 ( .A1(n10251), .A2(n10250), .ZN(n10869) );
  NOR2_X1 U11426 ( .A1(n13635), .A2(n13634), .ZN(n13637) );
  AND3_X1 U11427 ( .A1(n10121), .A2(n10124), .A3(n10122), .ZN(n10117) );
  NOR2_X1 U11428 ( .A1(n17877), .A2(n21556), .ZN(n17891) );
  NAND2_X1 U11429 ( .A1(n13746), .A2(n13540), .ZN(n13635) );
  NOR2_X1 U11430 ( .A1(n11288), .A2(n9981), .ZN(n9980) );
  AND2_X1 U11431 ( .A1(n15574), .A2(n15577), .ZN(n13891) );
  NAND3_X1 U11432 ( .A1(n11177), .A2(n11176), .A3(n11175), .ZN(n9993) );
  NAND2_X1 U11433 ( .A1(n10944), .A2(n9806), .ZN(n13561) );
  AND2_X1 U11434 ( .A1(n13859), .A2(n13858), .ZN(n14610) );
  AND2_X1 U11435 ( .A1(n10506), .A2(n16568), .ZN(n10505) );
  NAND2_X1 U11436 ( .A1(n13874), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15657) );
  AND2_X1 U11437 ( .A1(n11910), .A2(n16531), .ZN(n10944) );
  OR3_X1 U11438 ( .A1(n16764), .A2(n16755), .A3(n16511), .ZN(n13784) );
  OAI21_X1 U11439 ( .B1(n13863), .B2(n10387), .A(n12870), .ZN(n14892) );
  NOR2_X1 U11440 ( .A1(n18173), .A2(n18367), .ZN(n18169) );
  NAND2_X1 U11441 ( .A1(n12225), .A2(n12224), .ZN(n14549) );
  AND2_X1 U11442 ( .A1(n15602), .A2(n15598), .ZN(n15563) );
  OR2_X1 U11443 ( .A1(n20391), .A2(n11327), .ZN(n10124) );
  AND3_X1 U11444 ( .A1(n11180), .A2(n10333), .A3(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n9719) );
  NAND2_X1 U11445 ( .A1(n9780), .A2(n11847), .ZN(n16844) );
  AND2_X1 U11446 ( .A1(n11523), .A2(n16779), .ZN(n13547) );
  NAND2_X1 U11447 ( .A1(n18182), .A2(n9775), .ZN(n18173) );
  INV_X1 U11448 ( .A(n18626), .ZN(n18577) );
  XNOR2_X1 U11449 ( .A(n10462), .B(n12872), .ZN(n13844) );
  INV_X1 U11450 ( .A(n18187), .ZN(n18182) );
  NAND2_X1 U11451 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18699), .ZN(n18626) );
  OR2_X1 U11452 ( .A1(n11181), .A2(n9704), .ZN(n20024) );
  OR2_X1 U11453 ( .A1(n11150), .A2(n12210), .ZN(n10043) );
  OR2_X1 U11454 ( .A1(n16090), .A2(n11378), .ZN(n11523) );
  OAI21_X1 U11455 ( .B1(n10215), .B2(n14230), .A(n12229), .ZN(n12232) );
  AND2_X1 U11456 ( .A1(n11159), .A2(n11158), .ZN(n11174) );
  NAND2_X1 U11457 ( .A1(n12141), .A2(n12142), .ZN(n18693) );
  OR2_X1 U11458 ( .A1(n11845), .A2(n16984), .ZN(n16959) );
  NOR2_X1 U11459 ( .A1(n11178), .A2(n11179), .ZN(n10601) );
  AND2_X1 U11460 ( .A1(n11521), .A2(n11520), .ZN(n16104) );
  NOR2_X1 U11461 ( .A1(n9825), .A2(n11516), .ZN(n19760) );
  OR2_X1 U11462 ( .A1(n16986), .A2(n16985), .ZN(n16974) );
  NAND2_X1 U11463 ( .A1(n10590), .A2(n9975), .ZN(n18943) );
  AND2_X1 U11464 ( .A1(n11158), .A2(n17184), .ZN(n10647) );
  NOR2_X2 U11465 ( .A1(n18267), .A2(n18776), .ZN(n18669) );
  NOR2_X1 U11466 ( .A1(n15908), .A2(n10783), .ZN(n10463) );
  AND2_X1 U11467 ( .A1(n12797), .A2(n12796), .ZN(n15908) );
  NAND2_X1 U11468 ( .A1(n19564), .A2(n17220), .ZN(n18776) );
  NAND2_X2 U11469 ( .A1(n19778), .A2(n19782), .ZN(n19826) );
  XNOR2_X1 U11470 ( .A(n12777), .B(n12775), .ZN(n12891) );
  NAND2_X1 U11471 ( .A1(n11865), .A2(n14701), .ZN(n16803) );
  NAND2_X1 U11472 ( .A1(n10635), .A2(n13804), .ZN(n12777) );
  NAND2_X1 U11473 ( .A1(n10048), .A2(n11133), .ZN(n11146) );
  NAND2_X1 U11474 ( .A1(n12899), .A2(n12898), .ZN(n10635) );
  NAND2_X1 U11475 ( .A1(n11140), .A2(n11132), .ZN(n10048) );
  OR2_X1 U11476 ( .A1(n12695), .A2(n12694), .ZN(n12696) );
  OAI21_X1 U11477 ( .B1(n17184), .B2(n14230), .A(n12216), .ZN(n17009) );
  XNOR2_X1 U11478 ( .A(n12899), .B(n10915), .ZN(n20784) );
  NAND2_X1 U11479 ( .A1(n10740), .A2(n18701), .ZN(n18700) );
  INV_X2 U11480 ( .A(n15429), .ZN(n20706) );
  AND2_X1 U11481 ( .A1(n15251), .A2(n10830), .ZN(n15202) );
  NAND2_X1 U11482 ( .A1(n11157), .A2(n11155), .ZN(n17184) );
  AND2_X1 U11483 ( .A1(n13710), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13711) );
  NAND2_X1 U11484 ( .A1(n14699), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17022) );
  NAND2_X1 U11485 ( .A1(n12783), .A2(n12782), .ZN(n20913) );
  CLKBUF_X1 U11486 ( .A(n12901), .Z(n20882) );
  INV_X2 U11487 ( .A(n18322), .ZN(n18329) );
  OR2_X1 U11488 ( .A1(n18737), .A2(n10663), .ZN(n10661) );
  INV_X2 U11489 ( .A(n18397), .ZN(n18405) );
  AND2_X1 U11490 ( .A1(n19520), .A2(n10398), .ZN(n19532) );
  NAND2_X1 U11491 ( .A1(n13702), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13706) );
  NAND2_X1 U11492 ( .A1(n10156), .A2(n13395), .ZN(n14579) );
  XNOR2_X1 U11493 ( .A(n12665), .B(n12682), .ZN(n20883) );
  NAND2_X1 U11494 ( .A1(n10542), .A2(n10541), .ZN(n11626) );
  AND2_X1 U11495 ( .A1(n13700), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13702) );
  AND2_X1 U11496 ( .A1(n17396), .A2(n10693), .ZN(n17519) );
  OAI21_X1 U11497 ( .B1(n12687), .B2(n12666), .A(n12667), .ZN(n12731) );
  CLKBUF_X1 U11498 ( .A(n17396), .Z(n17723) );
  NOR2_X1 U11499 ( .A1(n18147), .A2(n10705), .ZN(n17061) );
  NAND2_X1 U11500 ( .A1(n13393), .A2(n13392), .ZN(n10156) );
  XNOR2_X1 U11501 ( .A(n10694), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17396) );
  NOR2_X2 U11502 ( .A1(n18267), .A2(n17267), .ZN(n18573) );
  OAI211_X1 U11503 ( .C1(n11876), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        n11131) );
  OR2_X1 U11504 ( .A1(n12127), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10663) );
  NAND2_X1 U11505 ( .A1(n17057), .A2(n9830), .ZN(n17138) );
  OR2_X2 U11506 ( .A1(n14046), .A2(n14347), .ZN(n14154) );
  NOR2_X1 U11507 ( .A1(n18274), .A2(n12088), .ZN(n12096) );
  AND2_X1 U11508 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12126), .ZN(
        n12127) );
  XNOR2_X1 U11509 ( .A(n12126), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18738) );
  XNOR2_X1 U11510 ( .A(n12122), .B(n19036), .ZN(n18750) );
  XNOR2_X1 U11511 ( .A(n12125), .B(n12124), .ZN(n12126) );
  NAND2_X1 U11512 ( .A1(n11073), .A2(n11072), .ZN(n11629) );
  NOR2_X1 U11513 ( .A1(n12058), .A2(n12124), .ZN(n12085) );
  NOR2_X1 U11514 ( .A1(n11471), .A2(n10893), .ZN(n10892) );
  NAND4_X1 U11515 ( .A1(n12148), .A2(n19095), .A3(n12108), .A4(n18302), .ZN(
        n18342) );
  NAND2_X1 U11516 ( .A1(n15267), .A2(n14484), .ZN(n14580) );
  INV_X1 U11517 ( .A(n21412), .ZN(n14052) );
  AND2_X1 U11518 ( .A1(n11071), .A2(n11070), .ZN(n11073) );
  INV_X1 U11519 ( .A(n18762), .ZN(n9952) );
  INV_X1 U11520 ( .A(n12195), .ZN(n19091) );
  CLKBUF_X2 U11521 ( .A(n11808), .Z(n13649) );
  NAND3_X1 U11523 ( .A1(n11941), .A2(n11940), .A3(n11939), .ZN(n12177) );
  INV_X1 U11524 ( .A(n19076), .ZN(n18302) );
  INV_X1 U11525 ( .A(n10665), .ZN(n18287) );
  INV_X2 U11526 ( .A(n11378), .ZN(n13750) );
  INV_X1 U11527 ( .A(n19715), .ZN(n18343) );
  AND2_X1 U11528 ( .A1(n12671), .A2(n14587), .ZN(n13904) );
  INV_X1 U11529 ( .A(n14179), .ZN(n14484) );
  AND2_X1 U11530 ( .A1(n12658), .A2(n14566), .ZN(n10916) );
  AND2_X1 U11531 ( .A1(n12637), .A2(n10775), .ZN(n12638) );
  OR2_X1 U11532 ( .A1(n11268), .A2(n11267), .ZN(n11684) );
  OR2_X1 U11533 ( .A1(n11339), .A2(n11338), .ZN(n11691) );
  OR2_X2 U11534 ( .A1(n12632), .A2(n17176), .ZN(n12785) );
  OR2_X1 U11535 ( .A1(n12747), .A2(n12746), .ZN(n13876) );
  OR2_X1 U11536 ( .A1(n11952), .A2(n11951), .ZN(n18156) );
  OR2_X1 U11537 ( .A1(n11237), .A2(n11236), .ZN(n11662) );
  AOI211_X1 U11538 ( .C1(n18006), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n11938), .B(n11937), .ZN(n11939) );
  INV_X2 U11539 ( .A(n14297), .ZN(n17112) );
  NOR2_X2 U11540 ( .A1(n11930), .A2(n11929), .ZN(n19715) );
  OR2_X1 U11541 ( .A1(n11312), .A2(n11311), .ZN(n11688) );
  AND4_X1 U11542 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11376) );
  NAND2_X1 U11543 ( .A1(n11014), .A2(n11013), .ZN(n11075) );
  CLKBUF_X1 U11544 ( .A(n12634), .Z(n12671) );
  NAND2_X1 U11545 ( .A1(n10947), .A2(n10949), .ZN(n14198) );
  INV_X2 U11546 ( .A(U214), .ZN(n17303) );
  AND2_X1 U11547 ( .A1(n13679), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13681) );
  NAND2_X1 U11548 ( .A1(n10535), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10536) );
  NAND2_X1 U11549 ( .A1(n11042), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11053) );
  INV_X2 U11550 ( .A(n11063), .ZN(n9691) );
  AND4_X1 U11551 ( .A1(n12606), .A2(n12605), .A3(n12604), .A4(n12603), .ZN(
        n12627) );
  AND4_X1 U11552 ( .A1(n12611), .A2(n12610), .A3(n12609), .A4(n12608), .ZN(
        n12626) );
  AND4_X1 U11553 ( .A1(n12623), .A2(n12622), .A3(n12621), .A4(n12620), .ZN(
        n12624) );
  INV_X2 U11554 ( .A(n11227), .ZN(n9712) );
  AND4_X1 U11555 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12539) );
  AND4_X1 U11556 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        n12522) );
  AND4_X1 U11557 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12625) );
  NOR2_X2 U11558 ( .A1(n15350), .A2(n15573), .ZN(n14553) );
  AND4_X1 U11559 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12542) );
  AND4_X1 U11560 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12572), .ZN(
        n12591) );
  AND4_X1 U11561 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        n12590) );
  AND4_X1 U11562 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n12540) );
  AND4_X1 U11563 ( .A1(n12570), .A2(n12569), .A3(n12568), .A4(n12567), .ZN(
        n10949) );
  AND4_X1 U11564 ( .A1(n12583), .A2(n12582), .A3(n12581), .A4(n12580), .ZN(
        n12589) );
  AND4_X1 U11565 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12588) );
  AND4_X1 U11566 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n12562) );
  AND4_X1 U11567 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n12561) );
  BUF_X2 U11568 ( .A(n12755), .Z(n12720) );
  BUF_X2 U11569 ( .A(n12607), .Z(n12754) );
  BUF_X2 U11570 ( .A(n12739), .Z(n13302) );
  INV_X1 U11571 ( .A(n17788), .ZN(n17773) );
  BUF_X2 U11572 ( .A(n11713), .Z(n12294) );
  BUF_X4 U11573 ( .A(n17806), .Z(n18106) );
  AND2_X2 U11574 ( .A1(n11190), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12330) );
  AND2_X2 U11575 ( .A1(n14489), .A2(n14178), .ZN(n12612) );
  OR3_X2 U11576 ( .A1(n19726), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19055) );
  AND2_X2 U11577 ( .A1(n14486), .A2(n14504), .ZN(n12607) );
  AND2_X2 U11578 ( .A1(n12516), .A2(n12517), .ZN(n12741) );
  AND2_X2 U11579 ( .A1(n14486), .A2(n14178), .ZN(n12757) );
  INV_X2 U11580 ( .A(n19724), .ZN(n19723) );
  AND2_X2 U11581 ( .A1(n19528), .A2(n11915), .ZN(n12071) );
  AND2_X2 U11582 ( .A1(n9709), .A2(n11006), .ZN(n12336) );
  INV_X4 U11584 ( .A(n10946), .ZN(n9692) );
  NAND2_X1 U11585 ( .A1(n12466), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11227) );
  AND2_X2 U11586 ( .A1(n12510), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14486) );
  AND2_X1 U11587 ( .A1(n12509), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10049) );
  AND2_X2 U11588 ( .A1(n10774), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14489) );
  CLKBUF_X2 U11589 ( .A(n10952), .Z(n14599) );
  AND2_X2 U11590 ( .A1(n10951), .A2(n14680), .ZN(n11189) );
  INV_X1 U11591 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10774) );
  AND2_X1 U11592 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10951) );
  INV_X1 U11593 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10953) );
  NOR2_X2 U11594 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12517) );
  INV_X1 U11595 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10952) );
  INV_X2 U11596 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n17176) );
  NAND2_X1 U11597 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19536) );
  INV_X1 U11598 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19689) );
  AOI21_X1 U11599 ( .B1(n16507), .B2(n16511), .A(n16496), .ZN(n13585) );
  NOR2_X2 U11600 ( .A1(n14380), .A2(n10828), .ZN(n14466) );
  OR2_X1 U11601 ( .A1(n11143), .A2(n11142), .ZN(n11157) );
  INV_X2 U11602 ( .A(n16004), .ZN(n12490) );
  AND2_X2 U11603 ( .A1(n11074), .A2(n11607), .ZN(n11115) );
  XNOR2_X1 U11605 ( .A(n14522), .B(n14524), .ZN(n20537) );
  NAND2_X4 U11606 ( .A1(n10537), .A2(n10536), .ZN(n11074) );
  NOR2_X1 U11607 ( .A1(n11920), .A2(n19536), .ZN(n11946) );
  NOR2_X2 U11608 ( .A1(n11101), .A2(n10243), .ZN(n11862) );
  INV_X2 U11609 ( .A(n10946), .ZN(n9695) );
  OR2_X1 U11610 ( .A1(n19536), .A2(n11923), .ZN(n10946) );
  INV_X4 U11611 ( .A(n12506), .ZN(n11544) );
  NOR2_X2 U11612 ( .A1(n16043), .A2(n16042), .ZN(n16024) );
  NAND2_X2 U11613 ( .A1(n10967), .A2(n10966), .ZN(n11055) );
  INV_X4 U11614 ( .A(n11765), .ZN(n11652) );
  NAND2_X4 U11615 ( .A1(n10298), .A2(n13805), .ZN(n13880) );
  OAI22_X2 U11616 ( .A1(n15535), .A2(n15533), .B1(n15507), .B2(n15532), .ZN(
        n15521) );
  XNOR2_X1 U11617 ( .A(n14915), .B(n12507), .ZN(n13730) );
  INV_X1 U11618 ( .A(n11064), .ZN(n9698) );
  AND2_X1 U11619 ( .A1(n14676), .A2(n14599), .ZN(n9699) );
  AND2_X1 U11620 ( .A1(n14676), .A2(n14599), .ZN(n9700) );
  AND2_X1 U11621 ( .A1(n19528), .A2(n11915), .ZN(n9701) );
  NOR2_X1 U11622 ( .A1(n11173), .A2(n17184), .ZN(n11169) );
  AND2_X2 U11623 ( .A1(n12655), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12516) );
  OAI21_X1 U11624 ( .B1(n12687), .B2(n12655), .A(n12657), .ZN(n12665) );
  INV_X2 U11625 ( .A(n11999), .ZN(n9702) );
  NOR2_X1 U11626 ( .A1(n17750), .A2(n11924), .ZN(n12040) );
  INV_X4 U11627 ( .A(n11074), .ZN(n11650) );
  NOR2_X4 U11628 ( .A1(n18520), .A2(n10688), .ZN(n17386) );
  MUX2_X2 U11629 ( .A(n13984), .B(n13768), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n19778) );
  OAI21_X1 U11630 ( .B1(n14937), .B2(n17180), .A(n13773), .ZN(n13774) );
  XNOR2_X2 U11631 ( .A(n13765), .B(n13764), .ZN(n14937) );
  AND2_X2 U11632 ( .A1(n14763), .A2(n14790), .ZN(n14789) );
  NOR2_X2 U11633 ( .A1(n14740), .A2(n14765), .ZN(n14763) );
  AND2_X4 U11634 ( .A1(n14725), .A2(n15242), .ZN(n15165) );
  NOR2_X2 U11635 ( .A1(n14723), .A2(n14724), .ZN(n14725) );
  AND2_X1 U11636 ( .A1(n10951), .A2(n14680), .ZN(n9705) );
  AND2_X2 U11637 ( .A1(n10951), .A2(n14680), .ZN(n9706) );
  INV_X4 U11638 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10954) );
  AND2_X2 U11639 ( .A1(n11186), .A2(n10954), .ZN(n9708) );
  AND2_X2 U11640 ( .A1(n11186), .A2(n10954), .ZN(n9709) );
  INV_X1 U11641 ( .A(n17788), .ZN(n9713) );
  INV_X1 U11642 ( .A(n17788), .ZN(n9714) );
  AND2_X2 U11643 ( .A1(n12467), .A2(n11006), .ZN(n11358) );
  AND2_X1 U11644 ( .A1(n10189), .A2(n10650), .ZN(n10235) );
  NOR2_X1 U11645 ( .A1(n10651), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10650) );
  AND4_X1 U11646 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11375) );
  NAND2_X1 U11647 ( .A1(n10295), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10086) );
  NOR2_X1 U11648 ( .A1(n11341), .A2(n11453), .ZN(n10085) );
  AND2_X1 U11649 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  NAND2_X1 U11650 ( .A1(n11099), .A2(n11075), .ZN(n10014) );
  NAND2_X1 U11651 ( .A1(n18197), .A2(n19076), .ZN(n12104) );
  NOR2_X1 U11652 ( .A1(n10790), .A2(n10607), .ZN(n10606) );
  NAND2_X1 U11653 ( .A1(n10273), .A2(n10272), .ZN(n10219) );
  NAND2_X1 U11654 ( .A1(n16668), .A2(n10490), .ZN(n10272) );
  NAND2_X1 U11655 ( .A1(n10575), .A2(n11482), .ZN(n10273) );
  AND2_X2 U11656 ( .A1(n10787), .A2(n9982), .ZN(n10621) );
  NAND2_X1 U11657 ( .A1(n9993), .A2(n10113), .ZN(n9983) );
  NAND2_X1 U11658 ( .A1(n10115), .A2(n10785), .ZN(n9984) );
  NOR2_X1 U11659 ( .A1(n12113), .A2(n9681), .ZN(n19524) );
  NAND2_X1 U11660 ( .A1(n18721), .A2(n12087), .ZN(n12090) );
  OAI21_X1 U11661 ( .B1(n12175), .B2(n12191), .A(n12174), .ZN(n12192) );
  INV_X1 U11662 ( .A(n15456), .ZN(n13900) );
  OAI21_X1 U11663 ( .B1(n12210), .B2(n10856), .A(n10853), .ZN(n12224) );
  NAND3_X2 U11664 ( .A1(n10039), .A2(n10038), .A3(n9836), .ZN(n16510) );
  NAND2_X1 U11665 ( .A1(n10143), .A2(n9812), .ZN(n10038) );
  NAND2_X1 U11666 ( .A1(n10248), .A2(n10076), .ZN(n10039) );
  AND2_X1 U11667 ( .A1(n10919), .A2(n10918), .ZN(n10917) );
  NAND2_X1 U11668 ( .A1(n9737), .A2(n10580), .ZN(n10918) );
  INV_X1 U11669 ( .A(n10920), .ZN(n10919) );
  OAI21_X1 U11670 ( .B1(n10922), .B2(n10921), .A(n9838), .ZN(n10920) );
  NAND2_X1 U11671 ( .A1(n10191), .A2(n9745), .ZN(n10192) );
  NAND2_X1 U11672 ( .A1(n10128), .A2(n10505), .ZN(n10191) );
  OAI211_X1 U11673 ( .C1(n14227), .C2(n11627), .A(n10540), .B(n11649), .ZN(
        n10539) );
  AND3_X1 U11674 ( .A1(n11648), .A2(n11647), .A3(n11646), .ZN(n11649) );
  NAND3_X1 U11675 ( .A1(n12008), .A2(n12007), .A3(n12006), .ZN(n17262) );
  AOI211_X1 U11676 ( .C1(n18107), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n12005), .B(n12004), .ZN(n12006) );
  INV_X1 U11677 ( .A(n17262), .ZN(n18267) );
  NAND2_X1 U11678 ( .A1(n11628), .A2(n11607), .ZN(n11091) );
  NAND2_X1 U11679 ( .A1(n20346), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10136) );
  NAND2_X1 U11680 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U11681 ( .A1(n13374), .A2(n13373), .ZN(n13379) );
  XNOR2_X1 U11682 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U11683 ( .A1(n20812), .A2(n13876), .ZN(n12766) );
  INV_X1 U11684 ( .A(n13383), .ZN(n13380) );
  OAI21_X1 U11685 ( .B1(n14051), .B2(n12660), .A(n13928), .ZN(n12664) );
  INV_X1 U11686 ( .A(n10621), .ZN(n10056) );
  NAND2_X1 U11687 ( .A1(n11621), .A2(n11623), .ZN(n10543) );
  NAND2_X1 U11688 ( .A1(n17911), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10419) );
  NOR2_X1 U11689 ( .A1(n13916), .A2(n21201), .ZN(n10680) );
  INV_X1 U11690 ( .A(n13872), .ZN(n13863) );
  AND2_X1 U11691 ( .A1(n10913), .A2(n15696), .ZN(n10467) );
  NOR2_X1 U11692 ( .A1(n10835), .A2(n15133), .ZN(n10834) );
  INV_X1 U11693 ( .A(n10837), .ZN(n10835) );
  NAND2_X1 U11694 ( .A1(n10325), .A2(n15551), .ZN(n10321) );
  NOR2_X1 U11695 ( .A1(n15153), .A2(n10838), .ZN(n10837) );
  INV_X1 U11696 ( .A(n15144), .ZN(n10838) );
  AND2_X1 U11697 ( .A1(n14163), .A2(n13528), .ZN(n13502) );
  INV_X1 U11698 ( .A(n13502), .ZN(n13520) );
  AND2_X1 U11699 ( .A1(n13914), .A2(n13913), .ZN(n13930) );
  AOI21_X1 U11700 ( .B1(n9682), .B2(n15982), .A(n10533), .ZN(n10532) );
  INV_X1 U11701 ( .A(n16490), .ZN(n10533) );
  NAND2_X1 U11702 ( .A1(n10809), .A2(n14772), .ZN(n10808) );
  INV_X1 U11703 ( .A(n14775), .ZN(n10809) );
  NOR2_X1 U11704 ( .A1(n14652), .A2(n17056), .ZN(n12230) );
  NAND2_X1 U11705 ( .A1(n12214), .A2(n12213), .ZN(n14652) );
  AND2_X1 U11706 ( .A1(n14347), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U11707 ( .A1(n10035), .A2(n10034), .ZN(n10023) );
  AND2_X1 U11708 ( .A1(n10036), .A2(n11061), .ZN(n10035) );
  OAI21_X1 U11709 ( .B1(n11837), .B2(n11105), .A(n11054), .ZN(n10036) );
  AOI22_X1 U11710 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n18112), .ZN(n10401) );
  NAND2_X1 U11711 ( .A1(n18342), .A2(n9814), .ZN(n10358) );
  INV_X1 U11712 ( .A(n18700), .ZN(n9933) );
  XNOR2_X1 U11713 ( .A(n12085), .B(n18278), .ZN(n12086) );
  INV_X1 U11714 ( .A(n12058), .ZN(n12069) );
  NAND2_X1 U11715 ( .A1(n18752), .A2(n12082), .ZN(n9942) );
  NOR3_X1 U11716 ( .A1(n10365), .A2(n10364), .A3(n10362), .ZN(n10361) );
  INV_X1 U11717 ( .A(n11959), .ZN(n10365) );
  INV_X1 U11718 ( .A(n11956), .ZN(n10364) );
  NAND2_X1 U11719 ( .A1(n12100), .A2(n18156), .ZN(n12107) );
  AND2_X1 U11720 ( .A1(n12102), .A2(n19715), .ZN(n12103) );
  AND2_X2 U11721 ( .A1(n14566), .A2(n13430), .ZN(n14163) );
  NAND2_X1 U11722 ( .A1(n13274), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13313) );
  OR2_X1 U11723 ( .A1(n14579), .A2(n14054), .ZN(n17101) );
  NAND2_X1 U11724 ( .A1(n10638), .A2(n15621), .ZN(n15462) );
  INV_X1 U11725 ( .A(n15439), .ZN(n10637) );
  INV_X1 U11726 ( .A(n20772), .ZN(n13950) );
  NAND2_X1 U11727 ( .A1(n20723), .A2(n20722), .ZN(n15893) );
  OR2_X1 U11728 ( .A1(n17102), .A2(n14055), .ZN(n14576) );
  AOI21_X1 U11729 ( .B1(n13922), .B2(n10568), .A(n20561), .ZN(n13944) );
  INV_X1 U11730 ( .A(n10569), .ZN(n10568) );
  OAI22_X1 U11731 ( .A1(n14579), .A2(n10570), .B1(n13910), .B2(n10775), .ZN(
        n10569) );
  INV_X1 U11732 ( .A(n13829), .ZN(n15907) );
  AOI21_X1 U11733 ( .B1(n19818), .B2(n12219), .A(n12218), .ZN(n14291) );
  XNOR2_X1 U11734 ( .A(n17009), .B(n12220), .ZN(n14292) );
  AND2_X1 U11735 ( .A1(n9819), .A2(n12231), .ZN(n10859) );
  NOR2_X1 U11736 ( .A1(n10459), .A2(n16266), .ZN(n10455) );
  NAND2_X1 U11737 ( .A1(n12293), .A2(n12292), .ZN(n16318) );
  NAND2_X1 U11738 ( .A1(n9789), .A2(n10825), .ZN(n10824) );
  INV_X1 U11739 ( .A(n14633), .ZN(n10825) );
  XNOR2_X1 U11740 ( .A(n13699), .B(n13698), .ZN(n13984) );
  XNOR2_X1 U11741 ( .A(n14931), .B(n13762), .ZN(n16360) );
  INV_X1 U11742 ( .A(n16742), .ZN(n10554) );
  NOR2_X1 U11743 ( .A1(n9908), .A2(n16732), .ZN(n10655) );
  NAND2_X1 U11744 ( .A1(n10271), .A2(n10096), .ZN(n10095) );
  NOR2_X1 U11745 ( .A1(n9909), .A2(n16732), .ZN(n10379) );
  AOI21_X1 U11746 ( .B1(n10606), .B2(n10604), .A(n9846), .ZN(n10603) );
  NAND2_X1 U11747 ( .A1(n10791), .A2(n10789), .ZN(n10788) );
  INV_X1 U11748 ( .A(n10606), .ZN(n10605) );
  OR2_X1 U11749 ( .A1(n11868), .A2(n11528), .ZN(n10134) );
  NAND2_X1 U11750 ( .A1(n10192), .A2(n9828), .ZN(n10503) );
  NAND2_X1 U11751 ( .A1(n16802), .A2(n9913), .ZN(n10178) );
  AOI21_X1 U11752 ( .B1(n10505), .B2(n10507), .A(n10584), .ZN(n10504) );
  NOR2_X1 U11753 ( .A1(n9764), .A2(n10651), .ZN(n10282) );
  NOR2_X1 U11754 ( .A1(n11345), .A2(n10485), .ZN(n10484) );
  NAND2_X1 U11755 ( .A1(n10199), .A2(n16621), .ZN(n16653) );
  INV_X1 U11756 ( .A(n16622), .ZN(n10199) );
  NAND2_X1 U11757 ( .A1(n10075), .A2(n16674), .ZN(n10378) );
  NAND2_X1 U11758 ( .A1(n10063), .A2(n10061), .ZN(n10295) );
  NAND2_X1 U11759 ( .A1(n10062), .A2(n11345), .ZN(n10061) );
  INV_X1 U11760 ( .A(n16674), .ZN(n10062) );
  NAND3_X1 U11761 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n11149) );
  NAND2_X1 U11762 ( .A1(n10048), .A2(n9816), .ZN(n10044) );
  NAND2_X1 U11763 ( .A1(n11626), .A2(n11625), .ZN(n14699) );
  AND2_X1 U11764 ( .A1(n20155), .A2(n17033), .ZN(n20057) );
  NAND2_X1 U11765 ( .A1(n14853), .A2(n18342), .ZN(n17381) );
  NAND2_X1 U11766 ( .A1(n17904), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n17877) );
  NOR2_X1 U11767 ( .A1(n12163), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11915) );
  NOR2_X1 U11768 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10625) );
  OAI21_X1 U11769 ( .B1(n19532), .B2(n10397), .A(n14856), .ZN(n17140) );
  AND2_X1 U11770 ( .A1(n10355), .A2(n18343), .ZN(n10397) );
  INV_X1 U11771 ( .A(n17216), .ZN(n17214) );
  NAND2_X1 U11772 ( .A1(n18943), .A2(n17077), .ZN(n12200) );
  INV_X1 U11773 ( .A(n19513), .ZN(n10351) );
  NAND2_X1 U11774 ( .A1(n17261), .A2(n19514), .ZN(n10350) );
  NAND2_X1 U11775 ( .A1(n17217), .A2(n17216), .ZN(n10231) );
  NAND2_X1 U11776 ( .A1(n12096), .A2(n12095), .ZN(n17267) );
  NAND2_X1 U11777 ( .A1(n9976), .A2(n18673), .ZN(n12201) );
  AND2_X1 U11778 ( .A1(n18607), .A2(n18910), .ZN(n10760) );
  NAND2_X1 U11779 ( .A1(n12200), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12199) );
  NAND2_X2 U11780 ( .A1(n9963), .A2(n9792), .ZN(n12154) );
  XNOR2_X1 U11781 ( .A(n12086), .B(n12128), .ZN(n18723) );
  NOR2_X1 U11782 ( .A1(n19578), .A2(n19575), .ZN(n19711) );
  OR2_X1 U11783 ( .A1(n21329), .A2(n17176), .ZN(n20561) );
  NAND2_X1 U11784 ( .A1(n11420), .A2(n10538), .ZN(n19738) );
  NAND2_X1 U11785 ( .A1(n10798), .A2(n11574), .ZN(n16337) );
  INV_X1 U11786 ( .A(n16838), .ZN(n10477) );
  INV_X1 U11787 ( .A(n17260), .ZN(n10585) );
  INV_X1 U11788 ( .A(n9946), .ZN(n9945) );
  AOI21_X1 U11789 ( .B1(n9972), .B2(n9734), .A(n17266), .ZN(n9946) );
  AND2_X1 U11790 ( .A1(n18837), .A2(n18836), .ZN(n18846) );
  NOR2_X1 U11791 ( .A1(n12210), .A2(n17056), .ZN(n10218) );
  NAND2_X1 U11792 ( .A1(n9718), .A2(n10601), .ZN(n9916) );
  NAND2_X1 U11793 ( .A1(n12210), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U11794 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10289) );
  OAI21_X1 U11795 ( .B1(n11118), .B2(n14690), .A(n11091), .ZN(n10645) );
  OAI21_X1 U11796 ( .B1(n20087), .B2(n11316), .A(n10181), .ZN(n10183) );
  NAND2_X1 U11797 ( .A1(n10864), .A2(n10182), .ZN(n10181) );
  NOR2_X1 U11798 ( .A1(n11178), .A2(n9842), .ZN(n10182) );
  NAND2_X1 U11799 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10275) );
  INV_X1 U11800 ( .A(n19902), .ZN(n10276) );
  NOR2_X1 U11801 ( .A1(n12210), .A2(n10070), .ZN(n10069) );
  INV_X1 U11802 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U11803 ( .A1(n10646), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U11804 ( .A1(n11860), .A2(n11629), .ZN(n10646) );
  AOI21_X1 U11805 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19557), .A(
        n12162), .ZN(n12164) );
  AOI21_X1 U11806 ( .B1(n13379), .B2(n13378), .A(n13377), .ZN(n13390) );
  NOR2_X1 U11807 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20783), .ZN(
        n13388) );
  INV_X1 U11808 ( .A(n15918), .ZN(n13052) );
  OR2_X1 U11809 ( .A1(n12726), .A2(n12725), .ZN(n13821) );
  AND3_X1 U11810 ( .A1(n12571), .A2(n12638), .A3(n12658), .ZN(n13902) );
  NAND2_X1 U11811 ( .A1(n11840), .A2(n11082), .ZN(n11068) );
  NAND2_X1 U11812 ( .A1(n10871), .A2(n10249), .ZN(n10867) );
  NOR2_X1 U11813 ( .A1(n16540), .A2(n13556), .ZN(n10925) );
  INV_X1 U11814 ( .A(n10649), .ZN(n10301) );
  AND3_X1 U11815 ( .A1(n10220), .A2(n16623), .A3(n10612), .ZN(n10097) );
  AND2_X1 U11816 ( .A1(n16609), .A2(n16613), .ZN(n11481) );
  AOI21_X1 U11817 ( .B1(n16214), .B2(n13750), .A(n11453), .ZN(n10649) );
  NAND2_X1 U11818 ( .A1(n10180), .A2(n11343), .ZN(n10613) );
  AND2_X1 U11819 ( .A1(n9868), .A2(n11301), .ZN(n9978) );
  INV_X1 U11820 ( .A(n10115), .ZN(n10077) );
  NAND2_X1 U11821 ( .A1(n9993), .A2(n14347), .ZN(n10008) );
  XNOR2_X1 U11822 ( .A(n11065), .B(n11064), .ZN(n11632) );
  NAND2_X1 U11823 ( .A1(n12337), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10260) );
  NAND2_X1 U11824 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10258) );
  NAND2_X1 U11825 ( .A1(n11367), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10259) );
  INV_X1 U11826 ( .A(n11187), .ZN(n10262) );
  NAND2_X1 U11827 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  NAND2_X1 U11828 ( .A1(n14264), .A2(n11075), .ZN(n10244) );
  NAND2_X1 U11829 ( .A1(n11100), .A2(n11082), .ZN(n10245) );
  NAND2_X1 U11830 ( .A1(n11396), .A2(n11395), .ZN(n11399) );
  XNOR2_X1 U11831 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U11832 ( .A1(n10665), .A2(n12118), .ZN(n12058) );
  NAND2_X1 U11833 ( .A1(n12119), .A2(n18287), .ZN(n12125) );
  NAND2_X1 U11834 ( .A1(n18762), .A2(n12118), .ZN(n12119) );
  NAND2_X1 U11835 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10369) );
  OR3_X1 U11836 ( .A1(n15085), .A2(n21373), .A3(n21374), .ZN(n15042) );
  AND2_X1 U11837 ( .A1(n14901), .A2(n9910), .ZN(n15233) );
  NAND2_X1 U11838 ( .A1(n15035), .A2(n15036), .ZN(n15021) );
  NOR2_X1 U11839 ( .A1(n13138), .A2(n10444), .ZN(n10443) );
  NAND2_X1 U11840 ( .A1(n15062), .A2(n10777), .ZN(n10776) );
  AND2_X1 U11841 ( .A1(n9765), .A2(n15113), .ZN(n10396) );
  NAND2_X1 U11842 ( .A1(n13052), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13336) );
  AND2_X1 U11843 ( .A1(n13901), .A2(n15697), .ZN(n10909) );
  INV_X1 U11844 ( .A(n15152), .ZN(n10836) );
  AND2_X1 U11845 ( .A1(n10782), .A2(n12840), .ZN(n10345) );
  NOR2_X1 U11846 ( .A1(n13804), .A2(n13853), .ZN(n13805) );
  INV_X1 U11847 ( .A(n15658), .ZN(n10712) );
  OAI21_X1 U11848 ( .B1(n10714), .B2(n15657), .A(n9844), .ZN(n10640) );
  NAND2_X1 U11849 ( .A1(n13844), .A2(n13871), .ZN(n9943) );
  OAI21_X1 U11850 ( .B1(n15911), .B2(n9920), .A(n9918), .ZN(n13809) );
  AOI21_X1 U11851 ( .B1(n13808), .B2(n13853), .A(n9919), .ZN(n9918) );
  NAND2_X1 U11852 ( .A1(n9917), .A2(n13808), .ZN(n14626) );
  NAND2_X1 U11853 ( .A1(n15911), .A2(n13871), .ZN(n9917) );
  OR2_X1 U11854 ( .A1(n12763), .A2(n12762), .ZN(n13820) );
  AND3_X1 U11855 ( .A1(n14566), .A2(n12632), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13383) );
  NAND2_X1 U11856 ( .A1(n12648), .A2(n20804), .ZN(n14179) );
  AND2_X1 U11857 ( .A1(n12780), .A2(n21259), .ZN(n21032) );
  NAND2_X1 U11858 ( .A1(n20883), .A2(n12712), .ZN(n12711) );
  INV_X1 U11859 ( .A(n12712), .ZN(n10717) );
  NOR2_X1 U11860 ( .A1(n16053), .A2(n10518), .ZN(n10517) );
  INV_X1 U11861 ( .A(n16063), .ZN(n10518) );
  INV_X1 U11862 ( .A(n13563), .ZN(n10901) );
  AND2_X1 U11863 ( .A1(n10901), .A2(n9796), .ZN(n10900) );
  INV_X1 U11864 ( .A(n13576), .ZN(n13539) );
  INV_X1 U11865 ( .A(n16670), .ZN(n10522) );
  NOR2_X1 U11866 ( .A1(n19802), .A2(n10524), .ZN(n10523) );
  INV_X1 U11867 ( .A(n16709), .ZN(n10524) );
  NAND2_X1 U11868 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U11869 ( .A1(n13582), .A2(n13583), .ZN(n13590) );
  NAND2_X1 U11870 ( .A1(n11811), .A2(n10814), .ZN(n10813) );
  INV_X1 U11871 ( .A(n16106), .ZN(n10814) );
  AND2_X1 U11872 ( .A1(n13544), .A2(n10687), .ZN(n10686) );
  NAND2_X1 U11873 ( .A1(n16595), .A2(n16888), .ZN(n10687) );
  INV_X1 U11874 ( .A(n10336), .ZN(n10335) );
  NAND2_X1 U11875 ( .A1(n11345), .A2(n10485), .ZN(n10337) );
  NAND2_X1 U11876 ( .A1(n10142), .A2(n16674), .ZN(n11341) );
  INV_X1 U11877 ( .A(n11270), .ZN(n10180) );
  AOI21_X1 U11878 ( .B1(n10056), .B2(n10130), .A(n10129), .ZN(n9997) );
  AND2_X1 U11879 ( .A1(n11474), .A2(n10167), .ZN(n10166) );
  NAND2_X1 U11880 ( .A1(n16237), .A2(n13750), .ZN(n10167) );
  OAI21_X1 U11881 ( .B1(n11618), .B2(n19879), .A(n10894), .ZN(n11471) );
  NAND2_X1 U11882 ( .A1(n19879), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10894) );
  AND2_X1 U11883 ( .A1(n19869), .A2(n11074), .ZN(n11057) );
  NAND2_X1 U11884 ( .A1(n11074), .A2(n20300), .ZN(n13619) );
  NOR2_X1 U11885 ( .A1(n11821), .A2(n10243), .ZN(n14677) );
  NAND2_X1 U11886 ( .A1(n14457), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10541) );
  OAI21_X1 U11887 ( .B1(n10544), .B2(n10543), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10542) );
  AOI21_X1 U11888 ( .B1(n11616), .B2(n9743), .A(n11402), .ZN(n10544) );
  NAND2_X1 U11889 ( .A1(n10037), .A2(n12210), .ZN(n11323) );
  NAND2_X1 U11890 ( .A1(n10333), .A2(n11180), .ZN(n20087) );
  AND2_X1 U11891 ( .A1(n11081), .A2(n11075), .ZN(n11059) );
  INV_X1 U11892 ( .A(n11923), .ZN(n10417) );
  NOR2_X1 U11893 ( .A1(n9932), .A2(n9927), .ZN(n9926) );
  NAND2_X1 U11894 ( .A1(n9693), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9929) );
  AOI21_X1 U11895 ( .B1(n18076), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(n9931), .ZN(n9930) );
  INV_X1 U11896 ( .A(n12047), .ZN(n10762) );
  INV_X1 U11897 ( .A(n18271), .ZN(n12095) );
  NAND2_X1 U11898 ( .A1(n18455), .A2(n12150), .ZN(n10232) );
  NAND2_X1 U11899 ( .A1(n18700), .A2(n12094), .ZN(n9937) );
  NAND3_X1 U11900 ( .A1(n9953), .A2(n9955), .A3(n9954), .ZN(n12122) );
  NAND2_X1 U11901 ( .A1(n18298), .A2(n10665), .ZN(n9953) );
  XNOR2_X1 U11902 ( .A(n12118), .B(n10665), .ZN(n12081) );
  AOI22_X1 U11903 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n19553), .B2(n19689), .ZN(
        n12189) );
  INV_X1 U11904 ( .A(n12104), .ZN(n10370) );
  NOR2_X1 U11905 ( .A1(n12107), .A2(n12195), .ZN(n10360) );
  INV_X1 U11906 ( .A(n19520), .ZN(n19537) );
  CLKBUF_X1 U11907 ( .A(n13396), .Z(n14061) );
  OR2_X1 U11908 ( .A1(n15117), .A2(n13419), .ZN(n15091) );
  AND2_X1 U11909 ( .A1(n9774), .A2(n9910), .ZN(n10677) );
  AND2_X1 U11910 ( .A1(n13448), .A2(n13447), .ZN(n14468) );
  AND2_X1 U11911 ( .A1(n13425), .A2(n10680), .ZN(n10679) );
  NAND2_X1 U11912 ( .A1(n14464), .A2(n14465), .ZN(n14540) );
  AND2_X1 U11913 ( .A1(n14577), .A2(n14576), .ZN(n14578) );
  INV_X1 U11914 ( .A(n13904), .ZN(n14590) );
  AND2_X1 U11915 ( .A1(n21201), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13340) );
  OR2_X1 U11916 ( .A1(n13198), .A2(n13197), .ZN(n13216) );
  NAND2_X1 U11917 ( .A1(n13049), .A2(n10435), .ZN(n13114) );
  AND2_X1 U11918 ( .A1(n10436), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10435) );
  OR2_X1 U11919 ( .A1(n15332), .A2(n15333), .ZN(n15330) );
  AND2_X1 U11920 ( .A1(n10909), .A2(n10907), .ZN(n10906) );
  INV_X1 U11921 ( .A(n10908), .ZN(n10907) );
  NOR2_X1 U11922 ( .A1(n9833), .A2(n10466), .ZN(n10465) );
  INV_X1 U11923 ( .A(n10467), .ZN(n10466) );
  AND2_X1 U11924 ( .A1(n9877), .A2(n10843), .ZN(n10842) );
  INV_X1 U11925 ( .A(n15010), .ZN(n10843) );
  NOR2_X1 U11926 ( .A1(n15734), .A2(n10567), .ZN(n15714) );
  AND2_X1 U11927 ( .A1(n15893), .A2(n15716), .ZN(n10567) );
  NAND2_X1 U11928 ( .A1(n10321), .A2(n10320), .ZN(n13897) );
  NAND2_X1 U11929 ( .A1(n10324), .A2(n10050), .ZN(n15498) );
  NAND2_X1 U11930 ( .A1(n10321), .A2(n13893), .ZN(n15544) );
  AND2_X1 U11931 ( .A1(n13494), .A2(n13493), .ZN(n15144) );
  AND2_X1 U11932 ( .A1(n13491), .A2(n13490), .ZN(n15153) );
  OR2_X1 U11933 ( .A1(n10572), .A2(n13947), .ZN(n15822) );
  NAND2_X1 U11934 ( .A1(n20772), .A2(n13949), .ZN(n10572) );
  NAND2_X1 U11935 ( .A1(n10298), .A2(n10054), .ZN(n15585) );
  AND2_X1 U11936 ( .A1(n13805), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10054) );
  NOR2_X1 U11937 ( .A1(n10831), .A2(n13481), .ZN(n10830) );
  INV_X1 U11938 ( .A(n10832), .ZN(n10831) );
  NOR2_X2 U11939 ( .A1(n17151), .A2(n10839), .ZN(n14894) );
  OR2_X1 U11940 ( .A1(n10840), .A2(n14895), .ZN(n10839) );
  NAND2_X1 U11941 ( .A1(n17144), .A2(n17145), .ZN(n17143) );
  NOR2_X1 U11942 ( .A1(n20723), .A2(n20760), .ZN(n15845) );
  AND3_X1 U11943 ( .A1(n13941), .A2(n13931), .A3(n14172), .ZN(n14180) );
  INV_X1 U11944 ( .A(n12898), .ZN(n10915) );
  AND2_X1 U11945 ( .A1(n14061), .A2(n14297), .ZN(n14495) );
  NAND2_X1 U11946 ( .A1(n10399), .A2(n15907), .ZN(n20881) );
  AND2_X1 U11947 ( .A1(n13829), .A2(n15908), .ZN(n21008) );
  INV_X1 U11948 ( .A(n20919), .ZN(n20824) );
  NOR2_X1 U11949 ( .A1(n21152), .A2(n21151), .ZN(n21261) );
  NOR2_X1 U11950 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14556), .ZN(n20919) );
  NAND2_X1 U11951 ( .A1(n13829), .A2(n12798), .ZN(n21265) );
  AOI21_X1 U11952 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21199), .A(n20824), 
        .ZN(n21272) );
  NAND2_X1 U11953 ( .A1(n10255), .A2(n10254), .ZN(n11422) );
  NAND2_X1 U11954 ( .A1(n11402), .A2(n11619), .ZN(n10254) );
  NAND2_X1 U11955 ( .A1(n11676), .A2(n11617), .ZN(n10255) );
  NAND2_X1 U11956 ( .A1(n16028), .A2(n16519), .ZN(n16010) );
  CLKBUF_X1 U11957 ( .A(n11629), .Z(n14345) );
  INV_X1 U11958 ( .A(n14702), .ZN(n14705) );
  INV_X1 U11959 ( .A(n12230), .ZN(n10450) );
  AND2_X1 U11960 ( .A1(n10857), .A2(n9891), .ZN(n10247) );
  AND2_X1 U11961 ( .A1(n11810), .A2(n11809), .ZN(n16463) );
  AOI21_X1 U11962 ( .B1(n10808), .B2(n11692), .A(n10807), .ZN(n10806) );
  INV_X1 U11963 ( .A(n14288), .ZN(n10807) );
  OR2_X1 U11964 ( .A1(n14747), .A2(n10808), .ZN(n14774) );
  NOR2_X1 U11965 ( .A1(n14227), .A2(n14345), .ZN(n14336) );
  NOR3_X1 U11966 ( .A1(n16744), .A2(n10550), .A3(n10555), .ZN(n10548) );
  NOR2_X1 U11967 ( .A1(n13768), .A2(n10555), .ZN(n10482) );
  NOR2_X2 U11968 ( .A1(n13606), .A2(n14916), .ZN(n14915) );
  AND2_X2 U11969 ( .A1(n16510), .A2(n10656), .ZN(n14913) );
  NOR3_X1 U11970 ( .A1(n9908), .A2(n14926), .A3(n16732), .ZN(n10656) );
  NAND2_X1 U11972 ( .A1(n10554), .A2(n10552), .ZN(n13653) );
  AND2_X1 U11973 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  NAND2_X1 U11974 ( .A1(n10249), .A2(n10603), .ZN(n10005) );
  OAI21_X1 U11975 ( .B1(n10128), .B2(n10106), .A(n10102), .ZN(n11909) );
  AOI21_X1 U11976 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10102) );
  INV_X1 U11977 ( .A(n10505), .ZN(n10104) );
  CLKBUF_X1 U11978 ( .A(n14822), .Z(n14834) );
  AND3_X1 U11979 ( .A1(n11792), .A2(n11791), .A3(n11790), .ZN(n14545) );
  NAND2_X1 U11980 ( .A1(n16576), .A2(n16575), .ZN(n16583) );
  INV_X1 U11981 ( .A(n13553), .ZN(n16575) );
  NAND2_X1 U11982 ( .A1(n10823), .A2(n10821), .ZN(n10820) );
  INV_X1 U11983 ( .A(n14016), .ZN(n10821) );
  OR2_X1 U11984 ( .A1(n14254), .A2(n10822), .ZN(n14285) );
  AND3_X1 U11985 ( .A1(n11710), .A2(n11709), .A3(n11708), .ZN(n14280) );
  INV_X1 U11986 ( .A(n11341), .ZN(n11342) );
  NAND2_X1 U11987 ( .A1(n10797), .A2(n14735), .ZN(n10796) );
  NAND3_X1 U11988 ( .A1(n10017), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        n10021), .ZN(n9987) );
  NAND2_X1 U11989 ( .A1(n10489), .A2(n11346), .ZN(n9992) );
  NOR2_X1 U11990 ( .A1(n11839), .A2(n11838), .ZN(n14661) );
  OR2_X1 U11991 ( .A1(n11835), .A2(n11834), .ZN(n11839) );
  NAND2_X1 U11992 ( .A1(n12211), .A2(n20300), .ZN(n12228) );
  INV_X1 U11993 ( .A(n10855), .ZN(n10852) );
  AOI22_X1 U11994 ( .A1(n10853), .A2(n10856), .B1(n10855), .B2(n14230), .ZN(
        n10851) );
  OR2_X1 U11995 ( .A1(n17009), .A2(n12221), .ZN(n12222) );
  NAND2_X1 U11996 ( .A1(n10513), .A2(n10512), .ZN(n17012) );
  NAND2_X1 U11997 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U11998 ( .A1(n14457), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10513) );
  AND2_X1 U11999 ( .A1(n11174), .A2(n10864), .ZN(n17042) );
  OR2_X1 U12000 ( .A1(n17042), .A2(n20393), .ZN(n10278) );
  NOR2_X1 U12001 ( .A1(n11185), .A2(n12210), .ZN(n20122) );
  INV_X1 U12002 ( .A(n19909), .ZN(n20160) );
  NAND2_X1 U12003 ( .A1(n11166), .A2(n10648), .ZN(n20202) );
  INV_X1 U12004 ( .A(n20202), .ZN(n11328) );
  NOR2_X1 U12005 ( .A1(n11185), .A2(n10864), .ZN(n20264) );
  INV_X1 U12006 ( .A(n20306), .ZN(n20269) );
  AND2_X1 U12007 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20341), .ZN(
        n20392) );
  INV_X1 U12008 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20338) );
  NOR2_X1 U12009 ( .A1(n9704), .A2(n11158), .ZN(n11164) );
  NAND2_X1 U12010 ( .A1(n20537), .A2(n20524), .ZN(n20398) );
  NAND2_X1 U12011 ( .A1(n15935), .A2(n16997), .ZN(n14456) );
  NOR2_X1 U12012 ( .A1(n19715), .A2(n18302), .ZN(n12147) );
  NAND2_X1 U12013 ( .A1(n17224), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10694) );
  NOR2_X1 U12014 ( .A1(n18197), .A2(n10702), .ZN(n10700) );
  NAND2_X1 U12015 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10405) );
  NAND2_X1 U12016 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U12017 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10406) );
  AOI21_X1 U12018 ( .B1(n12071), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n10403), .ZN(n10402) );
  NAND2_X1 U12019 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10400) );
  INV_X1 U12020 ( .A(n11972), .ZN(n10372) );
  OAI21_X1 U12021 ( .B1(n11969), .B2(n9962), .A(n12072), .ZN(n9957) );
  AOI21_X1 U12022 ( .B1(n9688), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(n9961), 
        .ZN(n9960) );
  NOR2_X1 U12023 ( .A1(n17817), .A2(n21634), .ZN(n9961) );
  NAND2_X1 U12024 ( .A1(n12073), .A2(n12077), .ZN(n9958) );
  NOR2_X1 U12025 ( .A1(n19095), .A2(n18156), .ZN(n19547) );
  NOR2_X1 U12026 ( .A1(n18430), .A2(n9883), .ZN(n17127) );
  NAND2_X1 U12027 ( .A1(n10427), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10426) );
  INV_X1 U12028 ( .A(n17069), .ZN(n10427) );
  NAND2_X1 U12029 ( .A1(n10426), .A2(n9797), .ZN(n10428) );
  NOR2_X1 U12030 ( .A1(n18487), .A2(n18805), .ZN(n18802) );
  NOR2_X1 U12031 ( .A1(n10743), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10742) );
  INV_X1 U12032 ( .A(n10943), .ZN(n10743) );
  AOI22_X1 U12033 ( .A1(n12154), .A2(n10763), .B1(n18816), .B2(n18820), .ZN(
        n18856) );
  AND2_X1 U12034 ( .A1(n18816), .A2(n10764), .ZN(n10763) );
  NAND2_X1 U12035 ( .A1(n12201), .A2(n12200), .ZN(n18572) );
  NOR3_X1 U12036 ( .A1(n18940), .A2(n18910), .A3(n10766), .ZN(n18605) );
  AND2_X1 U12037 ( .A1(n10354), .A2(n10358), .ZN(n10353) );
  OR2_X1 U12038 ( .A1(n10356), .A2(n12103), .ZN(n10354) );
  NAND2_X1 U12039 ( .A1(n18342), .A2(n19524), .ZN(n10356) );
  AND2_X1 U12040 ( .A1(n12144), .A2(n12145), .ZN(n10666) );
  OR2_X2 U12041 ( .A1(n18682), .A2(n10759), .ZN(n9963) );
  NAND2_X1 U12042 ( .A1(n9936), .A2(n9934), .ZN(n18689) );
  INV_X1 U12043 ( .A(n12094), .ZN(n9935) );
  NOR2_X1 U12044 ( .A1(n9941), .A2(n19026), .ZN(n9940) );
  NAND2_X1 U12045 ( .A1(n12127), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10662) );
  INV_X1 U12046 ( .A(n9942), .ZN(n9938) );
  NAND2_X1 U12047 ( .A1(n19727), .A2(n14855), .ZN(n19027) );
  NAND2_X1 U12048 ( .A1(n12114), .A2(n9728), .ZN(n19521) );
  INV_X1 U12049 ( .A(n19027), .ZN(n19544) );
  NOR2_X1 U12050 ( .A1(n10632), .A2(n10630), .ZN(n10629) );
  AOI21_X1 U12051 ( .B1(n19559), .B2(n19558), .A(n19557), .ZN(n10632) );
  OAI21_X1 U12052 ( .B1(n19559), .B2(n19558), .A(n10631), .ZN(n10630) );
  OR2_X1 U12053 ( .A1(n10628), .A2(n19709), .ZN(n10627) );
  OR2_X1 U12054 ( .A1(n19564), .A2(n19563), .ZN(n10628) );
  NAND2_X1 U12055 ( .A1(n10156), .A2(n10154), .ZN(n14384) );
  NOR2_X1 U12056 ( .A1(n9788), .A2(n10155), .ZN(n10154) );
  INV_X1 U12057 ( .A(n13395), .ZN(n10155) );
  NAND2_X1 U12058 ( .A1(n14384), .A2(n14043), .ZN(n21407) );
  NAND2_X1 U12059 ( .A1(n14886), .A2(n20585), .ZN(n15000) );
  OR2_X1 U12060 ( .A1(n15686), .A2(n20648), .ZN(n10153) );
  AOI21_X1 U12061 ( .B1(n15294), .B2(n14888), .A(n10152), .ZN(n10151) );
  INV_X1 U12062 ( .A(n14887), .ZN(n10152) );
  OR2_X1 U12063 ( .A1(n15100), .A2(n13412), .ZN(n15063) );
  AND2_X1 U12064 ( .A1(n13533), .A2(n13532), .ZN(n20627) );
  NOR2_X1 U12065 ( .A1(n15407), .A2(n14589), .ZN(n15397) );
  OR2_X1 U12066 ( .A1(n14866), .A2(n14867), .ZN(n14868) );
  INV_X1 U12067 ( .A(n13274), .ZN(n13276) );
  AND2_X2 U12068 ( .A1(n15671), .A2(n13974), .ZN(n20709) );
  INV_X1 U12069 ( .A(n20709), .ZN(n15673) );
  OR2_X1 U12070 ( .A1(n17102), .A2(n20561), .ZN(n13970) );
  NAND2_X1 U12071 ( .A1(n15691), .A2(n10563), .ZN(n15677) );
  NOR2_X1 U12072 ( .A1(n10564), .A2(n15680), .ZN(n10563) );
  NOR2_X1 U12073 ( .A1(n20761), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U12074 ( .A1(n10910), .A2(n15680), .ZN(n10307) );
  NAND2_X1 U12075 ( .A1(n10309), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10308) );
  INV_X1 U12076 ( .A(n10910), .ZN(n10309) );
  NOR2_X1 U12077 ( .A1(n15710), .A2(n10565), .ZN(n15691) );
  NOR2_X1 U12078 ( .A1(n13954), .A2(n15696), .ZN(n10565) );
  NAND2_X1 U12079 ( .A1(n10349), .A2(n10348), .ZN(n14864) );
  NAND2_X1 U12080 ( .A1(n13900), .A2(n9880), .ZN(n10348) );
  AND3_X1 U12081 ( .A1(n10573), .A2(n10571), .A3(n20772), .ZN(n13951) );
  INV_X1 U12082 ( .A(n13947), .ZN(n10571) );
  NOR3_X1 U12083 ( .A1(n15770), .A2(n13962), .A3(n10574), .ZN(n10573) );
  AND2_X1 U12084 ( .A1(n13944), .A2(n13927), .ZN(n20757) );
  OR2_X1 U12085 ( .A1(n13973), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20781) );
  INV_X1 U12086 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21199) );
  INV_X1 U12087 ( .A(n13825), .ZN(n12892) );
  INV_X1 U12088 ( .A(n14513), .ZN(n21153) );
  CLKBUF_X1 U12089 ( .A(n14171), .Z(n21152) );
  INV_X1 U12090 ( .A(n20970), .ZN(n20962) );
  INV_X1 U12091 ( .A(n14945), .ZN(n13738) );
  NOR2_X1 U12092 ( .A1(n14945), .A2(n19820), .ZN(n10509) );
  INV_X1 U12093 ( .A(n13731), .ZN(n10508) );
  INV_X1 U12094 ( .A(n13727), .ZN(n13742) );
  NAND2_X1 U12095 ( .A1(n10527), .A2(n10526), .ZN(n15946) );
  AOI21_X1 U12096 ( .B1(n10528), .B2(n19778), .A(n19778), .ZN(n10526) );
  NOR2_X1 U12097 ( .A1(n10529), .A2(n15961), .ZN(n10528) );
  AOI21_X1 U12098 ( .B1(n16370), .B2(n19794), .A(n10728), .ZN(n10727) );
  NAND2_X1 U12099 ( .A1(n15953), .A2(n15952), .ZN(n10728) );
  INV_X1 U12100 ( .A(n19813), .ZN(n19794) );
  AND2_X1 U12101 ( .A1(n19812), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19787) );
  NAND2_X1 U12102 ( .A1(n15942), .A2(n14721), .ZN(n19813) );
  AND2_X1 U12103 ( .A1(n14036), .A2(n13729), .ZN(n19819) );
  INV_X1 U12104 ( .A(n14801), .ZN(n14784) );
  INV_X1 U12105 ( .A(n16354), .ZN(n19828) );
  NOR2_X1 U12106 ( .A1(n16266), .A2(n12475), .ZN(n10456) );
  NAND2_X1 U12107 ( .A1(n10849), .A2(n16271), .ZN(n16278) );
  NAND2_X1 U12108 ( .A1(n9691), .A2(n19840), .ZN(n16441) );
  OR2_X1 U12109 ( .A1(n14816), .A2(n17038), .ZN(n16470) );
  NAND2_X1 U12110 ( .A1(n10226), .A2(n10224), .ZN(n10223) );
  NOR2_X1 U12111 ( .A1(n13647), .A2(n13643), .ZN(n10224) );
  NAND2_X1 U12112 ( .A1(n9924), .A2(n14914), .ZN(n16479) );
  AOI21_X1 U12113 ( .B1(n10242), .B2(n10789), .A(n16680), .ZN(n10236) );
  NAND2_X1 U12114 ( .A1(n16517), .A2(n16518), .ZN(n10145) );
  NOR2_X1 U12115 ( .A1(n16712), .A2(n10211), .ZN(n10210) );
  INV_X1 U12116 ( .A(n10600), .ZN(n10211) );
  OAI21_X1 U12117 ( .B1(n10546), .B2(n16712), .A(n10209), .ZN(n10208) );
  INV_X1 U12118 ( .A(n16522), .ZN(n10209) );
  INV_X1 U12119 ( .A(n10503), .ZN(n10502) );
  NAND2_X1 U12120 ( .A1(n11380), .A2(n9773), .ZN(n16559) );
  AND2_X1 U12121 ( .A1(n16588), .A2(n16697), .ZN(n10195) );
  NAND2_X1 U12122 ( .A1(n16672), .A2(n14355), .ZN(n16710) );
  INV_X1 U12123 ( .A(n16672), .ZN(n16707) );
  INV_X1 U12124 ( .A(n16710), .ZN(n16692) );
  NAND2_X1 U12125 ( .A1(n13664), .A2(n16944), .ZN(n10422) );
  XNOR2_X1 U12126 ( .A(n10252), .B(n9801), .ZN(n14936) );
  NAND2_X1 U12127 ( .A1(n16485), .A2(n14910), .ZN(n10652) );
  INV_X1 U12128 ( .A(n16479), .ZN(n10280) );
  XNOR2_X1 U12129 ( .A(n13597), .B(n13596), .ZN(n16483) );
  NAND2_X1 U12130 ( .A1(n13591), .A2(n10434), .ZN(n10433) );
  NAND2_X1 U12131 ( .A1(n16485), .A2(n10112), .ZN(n10108) );
  NAND2_X1 U12132 ( .A1(n10112), .A2(n16484), .ZN(n10111) );
  AND2_X1 U12133 ( .A1(n10926), .A2(n16993), .ZN(n10614) );
  OR2_X1 U12134 ( .A1(n16518), .A2(n10607), .ZN(n10146) );
  INV_X1 U12135 ( .A(n16499), .ZN(n10241) );
  OAI21_X1 U12136 ( .B1(n16517), .B2(n10605), .A(n10603), .ZN(n16499) );
  NAND2_X1 U12137 ( .A1(n10141), .A2(n10546), .ZN(n9967) );
  XNOR2_X1 U12138 ( .A(n16517), .B(n10604), .ZN(n10164) );
  NAND2_X1 U12139 ( .A1(n16629), .A2(n13599), .ZN(n10159) );
  NAND2_X1 U12140 ( .A1(n10178), .A2(n21524), .ZN(n10160) );
  NAND2_X1 U12141 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  INV_X1 U12142 ( .A(n10134), .ZN(n10132) );
  INV_X1 U12143 ( .A(n10917), .ZN(n10133) );
  OAI211_X1 U12144 ( .C1(n10179), .C2(n10739), .A(n10174), .B(n16779), .ZN(
        n10177) );
  NAND2_X1 U12145 ( .A1(n10175), .A2(n10738), .ZN(n10174) );
  INV_X1 U12146 ( .A(n10176), .ZN(n10175) );
  NAND2_X1 U12147 ( .A1(n10188), .A2(n10576), .ZN(n16539) );
  AOI21_X1 U12148 ( .B1(n10577), .B2(n10579), .A(n13556), .ZN(n10576) );
  NAND2_X1 U12149 ( .A1(n10414), .A2(n11381), .ZN(n10413) );
  INV_X1 U12150 ( .A(n16816), .ZN(n10412) );
  INV_X1 U12151 ( .A(n16812), .ZN(n10414) );
  NOR2_X1 U12152 ( .A1(n16809), .A2(n10930), .ZN(n16826) );
  AOI21_X1 U12153 ( .B1(n19784), .B2(n16970), .A(n16821), .ZN(n10469) );
  NAND2_X1 U12154 ( .A1(n10191), .A2(n10504), .ZN(n16555) );
  NAND2_X1 U12155 ( .A1(n10340), .A2(n16559), .ZN(n16834) );
  NAND2_X1 U12156 ( .A1(n16562), .A2(n16828), .ZN(n10340) );
  NAND2_X1 U12157 ( .A1(n16570), .A2(n10285), .ZN(n16853) );
  NAND2_X1 U12158 ( .A1(n10286), .A2(n9884), .ZN(n10285) );
  AND2_X1 U12159 ( .A1(n9777), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10598) );
  NAND2_X1 U12160 ( .A1(n16604), .A2(n16888), .ZN(n10323) );
  XNOR2_X1 U12161 ( .A(n10197), .B(n16640), .ZN(n16932) );
  NAND2_X1 U12162 ( .A1(n10198), .A2(n16650), .ZN(n10197) );
  NAND2_X1 U12163 ( .A1(n16653), .A2(n16651), .ZN(n10198) );
  NAND2_X1 U12164 ( .A1(n10381), .A2(n10332), .ZN(n13601) );
  INV_X1 U12165 ( .A(n10076), .ZN(n10332) );
  OR2_X1 U12166 ( .A1(n17009), .A2(n14156), .ZN(n17033) );
  AND4_X1 U12167 ( .A1(n12213), .A2(n14155), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20300), .ZN(n14156) );
  INV_X1 U12168 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20542) );
  INV_X1 U12169 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20533) );
  XNOR2_X1 U12170 ( .A(n17411), .B(n17410), .ZN(n17416) );
  INV_X1 U12171 ( .A(n17731), .ZN(n17763) );
  OAI22_X1 U12172 ( .A1(n17877), .A2(n10695), .B1(n18143), .B2(n10697), .ZN(
        n17887) );
  OR2_X1 U12173 ( .A1(n10697), .A2(n21556), .ZN(n10695) );
  AND2_X1 U12174 ( .A1(n18123), .A2(n17874), .ZN(n10697) );
  AND2_X1 U12175 ( .A1(n17220), .A2(n18302), .ZN(n10706) );
  NOR2_X1 U12176 ( .A1(n18196), .A2(n18356), .ZN(n18192) );
  NOR2_X1 U12177 ( .A1(n18291), .A2(n19105), .ZN(n18263) );
  NOR2_X1 U12178 ( .A1(n18238), .A2(n18281), .ZN(n18269) );
  INV_X1 U12179 ( .A(n18255), .ZN(n18297) );
  AND2_X1 U12180 ( .A1(n19547), .A2(n17142), .ZN(n18255) );
  NAND2_X1 U12181 ( .A1(n10756), .A2(n10758), .ZN(n10755) );
  INV_X1 U12182 ( .A(n17219), .ZN(n10757) );
  INV_X1 U12183 ( .A(n18684), .ZN(n18620) );
  INV_X1 U12184 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19676) );
  NAND2_X1 U12185 ( .A1(n17236), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9965) );
  AOI21_X1 U12186 ( .B1(n17258), .B2(n17257), .A(n10754), .ZN(n10753) );
  INV_X1 U12187 ( .A(n17259), .ZN(n10754) );
  NAND2_X1 U12188 ( .A1(n10229), .A2(n17218), .ZN(n10750) );
  NAND2_X1 U12189 ( .A1(n10231), .A2(n10230), .ZN(n10229) );
  NAND2_X1 U12190 ( .A1(n19675), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10230) );
  NOR2_X1 U12191 ( .A1(n19040), .A2(n18418), .ZN(n9971) );
  OAI21_X1 U12192 ( .B1(n18802), .B2(n18820), .A(n10447), .ZN(n10674) );
  NOR2_X1 U12193 ( .A1(n10675), .A2(n10448), .ZN(n10447) );
  NAND2_X1 U12194 ( .A1(n19053), .A2(n18801), .ZN(n10448) );
  NOR2_X1 U12195 ( .A1(n18800), .A2(n18942), .ZN(n10675) );
  INV_X1 U12196 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19575) );
  INV_X1 U12197 ( .A(n18970), .ZN(n18962) );
  NOR2_X1 U12198 ( .A1(n18820), .A2(n19054), .ZN(n19021) );
  AOI211_X1 U12199 ( .C1(n12187), .C2(n19514), .A(n12186), .B(n14854), .ZN(
        n12198) );
  INV_X1 U12200 ( .A(n19021), .ZN(n19062) );
  INV_X1 U12201 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19560) );
  AOI22_X1 U12202 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n11043), .ZN(n10981) );
  AOI22_X1 U12203 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U12204 ( .A1(n10297), .A2(n14198), .ZN(n12644) );
  AND2_X1 U12205 ( .A1(n10878), .A2(n10877), .ZN(n12378) );
  NAND2_X1 U12206 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10878) );
  NAND2_X1 U12207 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10877) );
  AOI21_X1 U12208 ( .B1(n12319), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A(n9770), .ZN(n12372) );
  NAND2_X1 U12209 ( .A1(n10269), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10268) );
  NAND2_X1 U12210 ( .A1(n9753), .A2(n10041), .ZN(n10078) );
  INV_X1 U12211 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12212 ( .A1(n11174), .A2(n10218), .ZN(n10217) );
  AND2_X1 U12213 ( .A1(n10341), .A2(n10041), .ZN(n10040) );
  NOR2_X1 U12214 ( .A1(n12210), .A2(n11167), .ZN(n10341) );
  AOI21_X1 U12215 ( .B1(n17042), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n10101), .ZN(n11299) );
  NOR2_X1 U12216 ( .A1(n19997), .A2(n11298), .ZN(n10101) );
  INV_X1 U12217 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U12218 ( .A1(n10059), .A2(n10058), .ZN(n9981) );
  NAND2_X1 U12219 ( .A1(n10060), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10059) );
  NAND2_X1 U12220 ( .A1(n11295), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10058) );
  INV_X1 U12221 ( .A(n10202), .ZN(n9979) );
  NOR2_X1 U12222 ( .A1(n10292), .A2(n11197), .ZN(n11216) );
  NOR2_X1 U12223 ( .A1(n11185), .A2(n10072), .ZN(n11197) );
  NAND2_X1 U12224 ( .A1(n10082), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10072) );
  OAI21_X1 U12225 ( .B1(n20202), .B2(n11200), .A(n10003), .ZN(n11201) );
  NOR2_X1 U12226 ( .A1(n11212), .A2(n10088), .ZN(n11213) );
  NAND2_X1 U12227 ( .A1(n9704), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10067) );
  AND2_X1 U12228 ( .A1(n11099), .A2(n11650), .ZN(n11829) );
  NAND2_X1 U12229 ( .A1(n11081), .A2(n11015), .ZN(n10012) );
  NAND2_X1 U12230 ( .A1(n13383), .A2(n13871), .ZN(n13375) );
  OR2_X1 U12231 ( .A1(n9864), .A2(n10560), .ZN(n10557) );
  INV_X1 U12232 ( .A(n13366), .ZN(n10561) );
  NOR2_X1 U12233 ( .A1(n10560), .A2(n10562), .ZN(n10559) );
  INV_X1 U12234 ( .A(n13370), .ZN(n10562) );
  INV_X1 U12235 ( .A(n13350), .ZN(n13360) );
  AND2_X1 U12236 ( .A1(n12823), .A2(n12822), .ZN(n12871) );
  INV_X1 U12237 ( .A(n12863), .ZN(n10634) );
  NOR2_X1 U12238 ( .A1(n10783), .A2(n12871), .ZN(n10782) );
  INV_X1 U12239 ( .A(n13808), .ZN(n9920) );
  NOR2_X1 U12240 ( .A1(n12766), .A2(n17176), .ZN(n12769) );
  INV_X1 U12241 ( .A(n12769), .ZN(n13804) );
  OR2_X1 U12242 ( .A1(n12795), .A2(n12794), .ZN(n13846) );
  AOI22_X1 U12243 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12741), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U12244 ( .A1(n10023), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10033) );
  INV_X1 U12245 ( .A(n10645), .ZN(n10644) );
  AOI21_X1 U12246 ( .B1(n12319), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n9895), .ZN(n12449) );
  AND2_X1 U12247 ( .A1(n10888), .A2(n10887), .ZN(n12444) );
  NAND2_X1 U12248 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10887) );
  NAND2_X1 U12249 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10888) );
  AND2_X1 U12250 ( .A1(n16291), .A2(n12406), .ZN(n10026) );
  AND2_X1 U12251 ( .A1(n10884), .A2(n10883), .ZN(n12415) );
  NAND2_X1 U12252 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10883) );
  NAND2_X1 U12253 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10884) );
  AND2_X1 U12254 ( .A1(n10882), .A2(n10881), .ZN(n12410) );
  NAND2_X1 U12255 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10881) );
  NAND2_X1 U12256 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10882) );
  AND2_X1 U12257 ( .A1(n10880), .A2(n10879), .ZN(n12395) );
  NAND2_X1 U12258 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10879) );
  NAND2_X1 U12259 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10880) );
  AOI21_X1 U12260 ( .B1(n12466), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A(n9897), .ZN(n12390) );
  AND2_X1 U12261 ( .A1(n10876), .A2(n10875), .ZN(n12359) );
  NAND2_X1 U12262 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10875) );
  NAND2_X1 U12263 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10876) );
  AOI21_X1 U12264 ( .B1(n12466), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(n9904), .ZN(n12354) );
  AND2_X1 U12265 ( .A1(n10874), .A2(n10873), .ZN(n12325) );
  NAND2_X1 U12266 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U12267 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10874) );
  AOI21_X1 U12268 ( .B1(n12319), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A(n9903), .ZN(n12320) );
  NOR2_X1 U12269 ( .A1(n11592), .A2(n10722), .ZN(n10721) );
  INV_X1 U12270 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U12271 ( .A1(n13543), .A2(n13554), .ZN(n10924) );
  NAND2_X1 U12272 ( .A1(n11505), .A2(n16554), .ZN(n10692) );
  AND2_X1 U12273 ( .A1(n11481), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10490) );
  NOR2_X1 U12274 ( .A1(n10786), .A2(n11282), .ZN(n10785) );
  INV_X1 U12275 ( .A(n11314), .ZN(n10786) );
  NOR2_X1 U12276 ( .A1(n10114), .A2(n11650), .ZN(n10113) );
  INV_X1 U12277 ( .A(n10785), .ZN(n10114) );
  NAND2_X1 U12278 ( .A1(n10060), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10121) );
  INV_X1 U12279 ( .A(n10183), .ZN(n10122) );
  NOR2_X1 U12280 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  NOR2_X1 U12281 ( .A1(n11205), .A2(n11326), .ZN(n10119) );
  NAND2_X1 U12282 ( .A1(n11174), .A2(n9747), .ZN(n10277) );
  NOR2_X1 U12283 ( .A1(n10266), .A2(n11318), .ZN(n10265) );
  AND2_X1 U12284 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11318) );
  NAND2_X1 U12285 ( .A1(n11328), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10137) );
  AND2_X1 U12286 ( .A1(n11124), .A2(n11132), .ZN(n10032) );
  NOR2_X1 U12287 ( .A1(n11183), .A2(n11179), .ZN(n10333) );
  AOI22_X1 U12288 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U12289 ( .A1(n11066), .A2(n19875), .ZN(n11639) );
  AND2_X1 U12290 ( .A1(n20338), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11387) );
  XNOR2_X1 U12291 ( .A(n21424), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11393) );
  INV_X1 U12292 ( .A(n12042), .ZN(n9927) );
  NAND2_X1 U12293 ( .A1(n12161), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11924) );
  NAND2_X1 U12294 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19696), .ZN(
        n11921) );
  NAND2_X1 U12295 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10363) );
  AOI21_X1 U12296 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19553), .A(
        n12160), .ZN(n12170) );
  NOR2_X1 U12297 ( .A1(n12189), .A2(n12159), .ZN(n12160) );
  AOI21_X1 U12298 ( .B1(n13390), .B2(n13389), .A(n13388), .ZN(n13402) );
  AND2_X1 U12299 ( .A1(n14867), .A2(n10391), .ZN(n10390) );
  NOR2_X1 U12300 ( .A1(n14998), .A2(n10392), .ZN(n10391) );
  INV_X1 U12301 ( .A(n15009), .ZN(n10392) );
  OR2_X1 U12302 ( .A1(n15528), .A2(n13339), .ZN(n13136) );
  OR2_X1 U12303 ( .A1(n14587), .A2(n21201), .ZN(n10928) );
  INV_X1 U12304 ( .A(n13336), .ZN(n13309) );
  AND2_X1 U12305 ( .A1(n10779), .A2(n13082), .ZN(n10778) );
  AND2_X1 U12306 ( .A1(n13046), .A2(n9901), .ZN(n10779) );
  INV_X1 U12307 ( .A(n12923), .ZN(n10445) );
  AND2_X1 U12308 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U12309 ( .A1(n15621), .A2(n15680), .ZN(n10908) );
  INV_X1 U12310 ( .A(n15026), .ZN(n10844) );
  NOR2_X1 U12311 ( .A1(n15039), .A2(n10846), .ZN(n10845) );
  INV_X1 U12312 ( .A(n15050), .ZN(n10846) );
  AND2_X1 U12313 ( .A1(n15104), .A2(n15094), .ZN(n15081) );
  NOR2_X1 U12314 ( .A1(n15230), .A2(n10833), .ZN(n10832) );
  INV_X1 U12315 ( .A(n15250), .ZN(n10833) );
  NAND2_X1 U12316 ( .A1(n10841), .A2(n9824), .ZN(n10840) );
  INV_X1 U12317 ( .A(n17152), .ZN(n10841) );
  OR2_X1 U12318 ( .A1(n12837), .A2(n12836), .ZN(n13864) );
  NAND2_X1 U12319 ( .A1(n20758), .A2(n13828), .ZN(n13837) );
  OR2_X1 U12320 ( .A1(n13907), .A2(n14198), .ZN(n10570) );
  OAI211_X1 U12321 ( .C1(n13380), .C2(n12768), .A(n12767), .B(n12766), .ZN(
        n12898) );
  AOI21_X1 U12322 ( .B1(n14513), .B2(n17176), .A(n12728), .ZN(n12890) );
  AND3_X1 U12323 ( .A1(n12774), .A2(n12773), .A3(n12772), .ZN(n12775) );
  NAND2_X1 U12324 ( .A1(n12711), .A2(n12686), .ZN(n12695) );
  NAND2_X1 U12325 ( .A1(n12693), .A2(n12692), .ZN(n12694) );
  AOI22_X1 U12326 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12607), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U12327 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12607), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12549) );
  AOI21_X1 U12328 ( .B1(n17172), .B2(n17177), .A(n17123), .ZN(n14556) );
  NOR2_X1 U12329 ( .A1(n13593), .A2(n11569), .ZN(n11486) );
  NOR2_X1 U12330 ( .A1(n9795), .A2(n16633), .ZN(n16160) );
  INV_X1 U12331 ( .A(n11444), .ZN(n11446) );
  INV_X1 U12332 ( .A(n11691), .ZN(n11428) );
  NAND2_X1 U12333 ( .A1(n19879), .A2(n11423), .ZN(n11424) );
  INV_X1 U12334 ( .A(n15992), .ZN(n10794) );
  AND2_X1 U12335 ( .A1(n10890), .A2(n10889), .ZN(n12470) );
  NAND2_X1 U12336 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10889) );
  NAND2_X1 U12337 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10890) );
  AOI21_X1 U12338 ( .B1(n12319), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(n9896), .ZN(n12462) );
  AND2_X1 U12339 ( .A1(n10818), .A2(n13623), .ZN(n10817) );
  AND2_X1 U12340 ( .A1(n10886), .A2(n10885), .ZN(n12434) );
  NAND2_X1 U12341 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10885) );
  NAND2_X1 U12342 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10886) );
  AOI21_X1 U12343 ( .B1(n12466), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(n9898), .ZN(n12429) );
  INV_X1 U12344 ( .A(n14652), .ZN(n12386) );
  INV_X1 U12345 ( .A(n16311), .ZN(n10860) );
  AND2_X1 U12346 ( .A1(n12249), .A2(n10858), .ZN(n10857) );
  INV_X1 U12347 ( .A(n16331), .ZN(n10858) );
  NOR2_X1 U12348 ( .A1(n11096), .A2(n11080), .ZN(n11828) );
  INV_X1 U12349 ( .A(n13647), .ZN(n10225) );
  NAND2_X1 U12350 ( .A1(n13689), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13688) );
  NAND2_X1 U12351 ( .A1(n13683), .A2(n9727), .ZN(n13684) );
  INV_X1 U12352 ( .A(n10031), .ZN(n9951) );
  OAI22_X1 U12353 ( .A1(n11140), .A2(n10030), .B1(n11124), .B2(n11132), .ZN(
        n10031) );
  NOR2_X1 U12354 ( .A1(n11147), .A2(n11133), .ZN(n10030) );
  NAND2_X1 U12355 ( .A1(n9950), .A2(n11147), .ZN(n9949) );
  INV_X1 U12356 ( .A(n10032), .ZN(n9950) );
  NAND2_X1 U12357 ( .A1(n13627), .A2(n10551), .ZN(n10550) );
  INV_X1 U12358 ( .A(n13766), .ZN(n10551) );
  NAND2_X1 U12359 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U12360 ( .A1(n13747), .A2(n13638), .ZN(n13640) );
  OR2_X1 U12361 ( .A1(n13637), .A2(n13636), .ZN(n13638) );
  NOR2_X1 U12362 ( .A1(n15967), .A2(n10819), .ZN(n10818) );
  INV_X1 U12363 ( .A(n13782), .ZN(n10819) );
  INV_X1 U12364 ( .A(n16507), .ZN(n10792) );
  INV_X1 U12365 ( .A(n16005), .ZN(n12489) );
  INV_X1 U12366 ( .A(n9876), .ZN(n10250) );
  NAND2_X1 U12367 ( .A1(n13561), .A2(n10870), .ZN(n10251) );
  INV_X1 U12368 ( .A(n16523), .ZN(n10870) );
  AND2_X1 U12369 ( .A1(n11904), .A2(n11589), .ZN(n10802) );
  INV_X1 U12370 ( .A(n10944), .ZN(n10921) );
  INV_X1 U12371 ( .A(n16338), .ZN(n11578) );
  INV_X1 U12372 ( .A(n10691), .ZN(n10103) );
  AOI21_X1 U12373 ( .B1(n9723), .B2(n10580), .A(n10923), .ZN(n10691) );
  NOR2_X1 U12374 ( .A1(n11505), .A2(n10584), .ZN(n10583) );
  INV_X1 U12375 ( .A(n14545), .ZN(n10826) );
  INV_X1 U12376 ( .A(n14472), .ZN(n10827) );
  AND2_X1 U12377 ( .A1(n11481), .A2(n10300), .ZN(n10299) );
  NAND2_X1 U12378 ( .A1(n16623), .A2(n10301), .ZN(n10300) );
  NAND2_X1 U12379 ( .A1(n9799), .A2(n10098), .ZN(n10100) );
  AND2_X1 U12380 ( .A1(n10220), .A2(n10612), .ZN(n10098) );
  INV_X1 U12381 ( .A(n10142), .ZN(n10064) );
  INV_X1 U12382 ( .A(n14656), .ZN(n10797) );
  OAI21_X1 U12383 ( .B1(n10168), .B2(n10172), .A(n10170), .ZN(n10020) );
  NAND2_X1 U12384 ( .A1(n9996), .A2(n10042), .ZN(n10168) );
  NAND2_X1 U12385 ( .A1(n9964), .A2(n11315), .ZN(n10489) );
  AOI21_X1 U12386 ( .B1(n11126), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11137), .ZN(n11532) );
  NAND2_X1 U12387 ( .A1(n10165), .A2(n16237), .ZN(n16682) );
  NAND2_X1 U12388 ( .A1(n11140), .A2(n10032), .ZN(n10126) );
  INV_X1 U12389 ( .A(n10126), .ZN(n10047) );
  NAND4_X1 U12390 ( .A1(n9698), .A2(n9691), .A3(n11065), .A4(n11015), .ZN(
        n11078) );
  NAND2_X1 U12391 ( .A1(n11029), .A2(n10016), .ZN(n10015) );
  NAND2_X1 U12392 ( .A1(n11070), .A2(n10784), .ZN(n10016) );
  NAND2_X1 U12393 ( .A1(n14227), .A2(n9826), .ZN(n10540) );
  NOR2_X1 U12394 ( .A1(n10262), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U12395 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_0__SCAN_IN), .A(n10511), .ZN(n17013) );
  NAND2_X1 U12396 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10511) );
  AND2_X1 U12397 ( .A1(n12215), .A2(n10854), .ZN(n10853) );
  NAND2_X1 U12398 ( .A1(n12212), .A2(n14230), .ZN(n10854) );
  NOR2_X1 U12399 ( .A1(n12215), .A2(n10856), .ZN(n10855) );
  NAND2_X1 U12400 ( .A1(n12386), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12220) );
  NAND2_X1 U12401 ( .A1(n11044), .A2(n11006), .ZN(n14596) );
  NAND2_X1 U12402 ( .A1(n11182), .A2(n10864), .ZN(n19902) );
  AND2_X1 U12403 ( .A1(n11173), .A2(n17184), .ZN(n11159) );
  INV_X1 U12404 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n21618) );
  INV_X1 U12405 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21575) );
  NAND2_X1 U12406 ( .A1(n20403), .A2(n20521), .ZN(n17039) );
  OR3_X1 U12407 ( .A1(n11405), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n17137), .ZN(n11615) );
  XNOR2_X1 U12408 ( .A(n11399), .B(n11397), .ZN(n11619) );
  AND2_X1 U12409 ( .A1(n14455), .A2(n14457), .ZN(n15935) );
  NAND2_X1 U12410 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11922) );
  NOR2_X1 U12411 ( .A1(n17817), .A2(n21618), .ZN(n10403) );
  INV_X1 U12412 ( .A(n11920), .ZN(n9973) );
  NAND2_X1 U12413 ( .A1(n17241), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17209) );
  NAND2_X1 U12414 ( .A1(n10689), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10688) );
  NOR2_X1 U12415 ( .A1(n10690), .A2(n18497), .ZN(n10689) );
  NAND2_X1 U12416 ( .A1(n17697), .A2(n17207), .ZN(n17659) );
  INV_X1 U12417 ( .A(n17072), .ZN(n9970) );
  NAND2_X1 U12418 ( .A1(n18693), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12144) );
  AND3_X1 U12419 ( .A1(n12148), .A2(n12180), .A3(n19525), .ZN(n14855) );
  INV_X1 U12420 ( .A(n19511), .ZN(n17357) );
  NAND2_X1 U12421 ( .A1(n10352), .A2(n12114), .ZN(n19523) );
  OR2_X1 U12422 ( .A1(n10357), .A2(n10358), .ZN(n10352) );
  NOR2_X1 U12423 ( .A1(n19537), .A2(n9802), .ZN(n19535) );
  NAND2_X1 U12424 ( .A1(n9803), .A2(n10367), .ZN(n12100) );
  NOR2_X1 U12425 ( .A1(n11966), .A2(n10368), .ZN(n10367) );
  OAI221_X1 U12426 ( .B1(n19575), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n19676), .A(n19678), .ZN(n19074) );
  AOI21_X1 U12427 ( .B1(n19562), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n10631) );
  NAND2_X1 U12428 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n10684) );
  NOR2_X1 U12429 ( .A1(n15042), .A2(n15017), .ZN(n15013) );
  NAND2_X1 U12430 ( .A1(n13116), .A2(n10443), .ZN(n13170) );
  NAND2_X1 U12431 ( .A1(n13420), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15085) );
  NOR2_X1 U12432 ( .A1(n15177), .A2(n13411), .ZN(n15115) );
  NAND2_X1 U12433 ( .A1(n15204), .A2(n13417), .ZN(n15117) );
  AND2_X1 U12434 ( .A1(n15233), .A2(n13415), .ZN(n15204) );
  AND2_X1 U12435 ( .A1(n10677), .A2(n13415), .ZN(n10676) );
  INV_X1 U12436 ( .A(n13414), .ZN(n10678) );
  NOR2_X1 U12437 ( .A1(n20584), .A2(n13414), .ZN(n14901) );
  AND2_X1 U12438 ( .A1(n20638), .A2(n10680), .ZN(n13533) );
  AND4_X1 U12439 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n14724) );
  INV_X1 U12440 ( .A(n15350), .ZN(n15405) );
  XNOR2_X1 U12441 ( .A(n13345), .B(n13344), .ZN(n14885) );
  OR2_X1 U12442 ( .A1(n13343), .A2(n13342), .ZN(n13345) );
  NAND2_X1 U12443 ( .A1(n13314), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13343) );
  INV_X1 U12444 ( .A(n13313), .ZN(n13314) );
  AND2_X1 U12445 ( .A1(n15008), .A2(n10388), .ZN(n14983) );
  AND2_X1 U12446 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  INV_X1 U12447 ( .A(n14985), .ZN(n10389) );
  AND2_X1 U12448 ( .A1(n13255), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13274) );
  OR2_X1 U12449 ( .A1(n13216), .A2(n21575), .ZN(n13237) );
  NAND2_X1 U12450 ( .A1(n13235), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13256) );
  INV_X1 U12451 ( .A(n13237), .ZN(n13235) );
  NAND2_X1 U12452 ( .A1(n13116), .A2(n9771), .ZN(n13198) );
  AND2_X1 U12453 ( .A1(n10396), .A2(n10395), .ZN(n10394) );
  NOR2_X1 U12454 ( .A1(n9875), .A2(n15049), .ZN(n10395) );
  AND2_X1 U12455 ( .A1(n13115), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13116) );
  INV_X1 U12456 ( .A(n13114), .ZN(n13115) );
  NAND2_X1 U12457 ( .A1(n13116), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13154) );
  NOR2_X1 U12458 ( .A1(n10440), .A2(n10437), .ZN(n10436) );
  OR2_X1 U12459 ( .A1(n15547), .A2(n13339), .ZN(n13099) );
  AND2_X1 U12460 ( .A1(n13048), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13049) );
  NAND2_X1 U12461 ( .A1(n13049), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13083) );
  NOR2_X1 U12462 ( .A1(n13028), .A2(n12961), .ZN(n12976) );
  NAND2_X1 U12463 ( .A1(n10431), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13026) );
  INV_X1 U12464 ( .A(n12960), .ZN(n10431) );
  INV_X1 U12465 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15232) );
  OR2_X1 U12466 ( .A1(n13026), .A2(n15232), .ZN(n13028) );
  NAND2_X1 U12467 ( .A1(n10432), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12960) );
  INV_X1 U12468 ( .A(n12954), .ZN(n10432) );
  NAND2_X1 U12469 ( .A1(n12939), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12954) );
  INV_X1 U12470 ( .A(n12938), .ZN(n12939) );
  AND2_X1 U12471 ( .A1(n14892), .A2(n14572), .ZN(n10393) );
  OR2_X1 U12472 ( .A1(n12865), .A2(n12864), .ZN(n12938) );
  NAND2_X1 U12473 ( .A1(n10445), .A2(n12843), .ZN(n12874) );
  AND2_X1 U12474 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12911) );
  NAND2_X1 U12475 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12911), .ZN(
        n12923) );
  AOI21_X1 U12476 ( .B1(n12889), .B2(n10387), .A(n10386), .ZN(n10385) );
  INV_X1 U12477 ( .A(n12909), .ZN(n10386) );
  NAND2_X1 U12478 ( .A1(n9847), .A2(n15455), .ZN(n10914) );
  NAND2_X1 U12479 ( .A1(n15456), .A2(n10467), .ZN(n10912) );
  NAND2_X1 U12480 ( .A1(n15070), .A2(n9877), .ZN(n15024) );
  NAND2_X1 U12481 ( .A1(n15070), .A2(n10845), .ZN(n15041) );
  NAND2_X1 U12482 ( .A1(n15070), .A2(n15050), .ZN(n15052) );
  INV_X1 U12483 ( .A(n13949), .ZN(n10574) );
  NOR2_X1 U12484 ( .A1(n15120), .A2(n15105), .ZN(n15104) );
  AND2_X1 U12485 ( .A1(n13496), .A2(n13495), .ZN(n15133) );
  INV_X1 U12486 ( .A(n13891), .ZN(n15565) );
  OR2_X1 U12487 ( .A1(n13880), .A2(n15816), .ZN(n15577) );
  AND2_X1 U12488 ( .A1(n10303), .A2(n10305), .ZN(n15587) );
  NOR2_X1 U12489 ( .A1(n10306), .A2(n10304), .ZN(n10303) );
  INV_X1 U12490 ( .A(n15600), .ZN(n10304) );
  AND2_X1 U12491 ( .A1(n13480), .A2(n13479), .ZN(n15200) );
  NAND2_X1 U12492 ( .A1(n15585), .A2(n13883), .ZN(n15604) );
  NAND2_X1 U12493 ( .A1(n15251), .A2(n15250), .ZN(n15249) );
  AND2_X1 U12494 ( .A1(n13469), .A2(n13468), .ZN(n14730) );
  INV_X1 U12495 ( .A(n10640), .ZN(n10639) );
  NAND2_X1 U12496 ( .A1(n10712), .A2(n15657), .ZN(n10642) );
  AND2_X1 U12497 ( .A1(n13467), .A2(n13466), .ZN(n14895) );
  OR2_X1 U12498 ( .A1(n17151), .A2(n10840), .ZN(n15327) );
  NAND2_X1 U12499 ( .A1(n14468), .A2(n10829), .ZN(n10828) );
  INV_X1 U12500 ( .A(n14381), .ZN(n10829) );
  AND2_X1 U12501 ( .A1(n20769), .A2(n20771), .ZN(n20723) );
  NAND2_X1 U12502 ( .A1(n13930), .A2(n13917), .ZN(n17102) );
  NAND2_X1 U12503 ( .A1(n17163), .A2(n17176), .ZN(n13973) );
  NAND2_X1 U12504 ( .A1(n14208), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14207) );
  NAND2_X1 U12505 ( .A1(n10297), .A2(n12639), .ZN(n13937) );
  AOI22_X1 U12506 ( .A1(n12771), .A2(n12708), .B1(n13383), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12709) );
  INV_X1 U12507 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14500) );
  AND3_X1 U12508 ( .A1(n14203), .A2(n14202), .A3(n14201), .ZN(n17090) );
  OR2_X1 U12509 ( .A1(n20881), .A2(n21148), .ZN(n20785) );
  INV_X1 U12510 ( .A(n12637), .ZN(n12648) );
  NOR2_X2 U12511 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21273) );
  OR3_X1 U12512 ( .A1(n21091), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14556), 
        .ZN(n20827) );
  XNOR2_X1 U12513 ( .A(n12628), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n13409) );
  INV_X1 U12514 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21332) );
  XNOR2_X1 U12515 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U12516 ( .A1(n13580), .A2(n13539), .ZN(n13746) );
  INV_X1 U12517 ( .A(n10532), .ZN(n10529) );
  NAND2_X1 U12518 ( .A1(n10733), .A2(n10732), .ZN(n10731) );
  INV_X1 U12519 ( .A(n10734), .ZN(n10733) );
  NOR2_X1 U12520 ( .A1(n15970), .A2(n10735), .ZN(n10732) );
  NAND2_X1 U12521 ( .A1(n10530), .A2(n10532), .ZN(n15954) );
  NAND2_X1 U12522 ( .A1(n10514), .A2(n19798), .ZN(n16028) );
  NOR2_X1 U12523 ( .A1(n10519), .A2(n10516), .ZN(n10515) );
  INV_X1 U12524 ( .A(n10517), .ZN(n10516) );
  NAND2_X1 U12525 ( .A1(n10898), .A2(n10901), .ZN(n10897) );
  INV_X1 U12526 ( .A(n13539), .ZN(n10898) );
  NOR2_X1 U12527 ( .A1(n10903), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10902) );
  INV_X1 U12528 ( .A(n11517), .ZN(n10903) );
  NAND2_X1 U12529 ( .A1(n11518), .A2(n9796), .ZN(n13562) );
  NAND2_X1 U12530 ( .A1(n16062), .A2(n16063), .ZN(n16050) );
  NOR2_X1 U12531 ( .A1(n16082), .A2(n13693), .ZN(n11905) );
  NAND2_X1 U12532 ( .A1(n13694), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13693) );
  NAND2_X1 U12533 ( .A1(n14018), .A2(n9732), .ZN(n11512) );
  NAND2_X1 U12534 ( .A1(n14018), .A2(n9726), .ZN(n11500) );
  NAND2_X1 U12535 ( .A1(n14018), .A2(n11488), .ZN(n11491) );
  NAND2_X1 U12536 ( .A1(n11446), .A2(n10896), .ZN(n14019) );
  AND2_X1 U12537 ( .A1(n11445), .A2(n16166), .ZN(n10896) );
  NAND2_X1 U12538 ( .A1(n16160), .A2(n16616), .ZN(n14015) );
  NOR2_X1 U12539 ( .A1(n14015), .A2(n16597), .ZN(n16147) );
  INV_X1 U12540 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n16166) );
  NAND2_X1 U12541 ( .A1(n11430), .A2(n10253), .ZN(n11444) );
  AND2_X1 U12542 ( .A1(n9741), .A2(n11439), .ZN(n10253) );
  AND3_X1 U12543 ( .A1(n16229), .A2(n10523), .A3(n16663), .ZN(n10520) );
  NAND2_X1 U12544 ( .A1(n11430), .A2(n11429), .ZN(n11437) );
  INV_X1 U12545 ( .A(n11471), .ZN(n10891) );
  CLKBUF_X1 U12546 ( .A(n11431), .Z(n11456) );
  NAND2_X1 U12547 ( .A1(n16229), .A2(n10523), .ZN(n16218) );
  AND2_X1 U12548 ( .A1(n13674), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13677) );
  INV_X1 U12549 ( .A(n12503), .ZN(n13758) );
  OR2_X1 U12550 ( .A1(n11723), .A2(n11722), .ZN(n14788) );
  NAND2_X1 U12551 ( .A1(n10458), .A2(n10460), .ZN(n10453) );
  NAND2_X1 U12552 ( .A1(n12456), .A2(n12475), .ZN(n10460) );
  INV_X1 U12553 ( .A(n16277), .ZN(n10848) );
  AND2_X2 U12554 ( .A1(n13781), .A2(n10815), .ZN(n14931) );
  AND2_X1 U12555 ( .A1(n10817), .A2(n10816), .ZN(n10815) );
  INV_X1 U12556 ( .A(n14932), .ZN(n10816) );
  AND2_X1 U12557 ( .A1(n12293), .A2(n9899), .ZN(n16313) );
  NAND2_X1 U12558 ( .A1(n10811), .A2(n16075), .ZN(n10810) );
  INV_X1 U12559 ( .A(n10813), .ZN(n10811) );
  AND3_X1 U12560 ( .A1(n11805), .A2(n11804), .A3(n11803), .ZN(n14633) );
  AND3_X1 U12561 ( .A1(n11778), .A2(n11777), .A3(n11776), .ZN(n14471) );
  NAND2_X1 U12562 ( .A1(n16485), .A2(n10222), .ZN(n10221) );
  NOR2_X1 U12563 ( .A1(n10225), .A2(n10488), .ZN(n10222) );
  NAND2_X1 U12564 ( .A1(n11895), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13696) );
  INV_X1 U12565 ( .A(n11894), .ZN(n11895) );
  INV_X1 U12566 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13695) );
  NOR2_X1 U12567 ( .A1(n13696), .A2(n13695), .ZN(n13700) );
  INV_X1 U12568 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16082) );
  AND2_X1 U12569 ( .A1(n13689), .A2(n10720), .ZN(n13694) );
  AND2_X1 U12570 ( .A1(n9729), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10720) );
  NAND2_X1 U12571 ( .A1(n13689), .A2(n9729), .ZN(n13691) );
  INV_X1 U12572 ( .A(n14833), .ZN(n11574) );
  BUF_X1 U12573 ( .A(n16329), .Z(n16335) );
  NAND2_X1 U12574 ( .A1(n13683), .A2(n9749), .ZN(n13686) );
  AND2_X1 U12575 ( .A1(n13683), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13685) );
  AND2_X1 U12576 ( .A1(n13676), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13679) );
  NOR2_X1 U12577 ( .A1(n13671), .A2(n11591), .ZN(n13674) );
  NAND2_X1 U12578 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U12579 ( .A1(n10499), .A2(n9733), .ZN(n10497) );
  INV_X1 U12580 ( .A(n13744), .ZN(n10498) );
  NAND2_X1 U12581 ( .A1(n13768), .A2(n10555), .ZN(n10483) );
  NOR2_X1 U12582 ( .A1(n16744), .A2(n10550), .ZN(n10549) );
  INV_X1 U12583 ( .A(n14909), .ZN(n10654) );
  NAND2_X1 U12584 ( .A1(n13639), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10434) );
  AND2_X1 U12585 ( .A1(n13613), .A2(n13612), .ZN(n16015) );
  AND2_X1 U12586 ( .A1(n13609), .A2(n13608), .ZN(n16042) );
  NAND2_X1 U12587 ( .A1(n10932), .A2(n10610), .ZN(n10383) );
  NAND2_X1 U12588 ( .A1(n16594), .A2(n9815), .ZN(n10384) );
  AND2_X1 U12589 ( .A1(n13599), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10600) );
  OAI21_X1 U12590 ( .B1(n9759), .B2(n10318), .A(n10317), .ZN(n10316) );
  NOR2_X1 U12591 ( .A1(n13558), .A2(n11868), .ZN(n10318) );
  NAND2_X1 U12592 ( .A1(n9759), .A2(n13550), .ZN(n10317) );
  NAND2_X1 U12594 ( .A1(n11901), .A2(n10802), .ZN(n11880) );
  AND2_X1 U12595 ( .A1(n17188), .A2(n13624), .ZN(n10556) );
  AND2_X1 U12596 ( .A1(n11901), .A2(n11904), .ZN(n11902) );
  AND2_X1 U12597 ( .A1(n9680), .A2(n10474), .ZN(n10140) );
  INV_X1 U12598 ( .A(n14807), .ZN(n10812) );
  AND2_X1 U12599 ( .A1(n10578), .A2(n10186), .ZN(n10185) );
  NAND2_X1 U12600 ( .A1(n10187), .A2(n11496), .ZN(n10186) );
  AND2_X1 U12601 ( .A1(n10579), .A2(n16547), .ZN(n10578) );
  INV_X1 U12602 ( .A(n10686), .ZN(n10187) );
  AND2_X1 U12603 ( .A1(n10582), .A2(n16547), .ZN(n10577) );
  INV_X1 U12604 ( .A(n10583), .ZN(n10582) );
  AOI21_X1 U12605 ( .B1(n10583), .B2(n10581), .A(n10580), .ZN(n10579) );
  INV_X1 U12606 ( .A(n16568), .ZN(n10581) );
  NAND2_X1 U12607 ( .A1(n10184), .A2(n11496), .ZN(n16569) );
  OR2_X1 U12608 ( .A1(n10686), .A2(n10507), .ZN(n10506) );
  INV_X1 U12609 ( .A(n16569), .ZN(n10286) );
  NAND2_X1 U12610 ( .A1(n10827), .A2(n9789), .ZN(n14632) );
  NAND2_X1 U12611 ( .A1(n16621), .A2(n16623), .ZN(n16610) );
  INV_X1 U12612 ( .A(n14280), .ZN(n11711) );
  CLKBUF_X1 U12613 ( .A(n14740), .Z(n14764) );
  AND2_X1 U12614 ( .A1(n11346), .A2(n13750), .ZN(n10205) );
  NAND2_X1 U12615 ( .A1(n11377), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16646) );
  INV_X1 U12616 ( .A(n10616), .ZN(n11377) );
  OAI211_X1 U12617 ( .C1(n10430), .C2(n13750), .A(n10337), .B(n10334), .ZN(
        n10616) );
  NAND2_X1 U12618 ( .A1(n10180), .A2(n10130), .ZN(n10144) );
  NAND2_X1 U12619 ( .A1(n9849), .A2(n9995), .ZN(n9994) );
  NAND2_X1 U12620 ( .A1(n11269), .A2(n11315), .ZN(n10377) );
  NAND2_X1 U12621 ( .A1(n11270), .A2(n11271), .ZN(n11269) );
  NAND2_X1 U12622 ( .A1(n10087), .A2(n10166), .ZN(n11480) );
  INV_X1 U12623 ( .A(n16688), .ZN(n11537) );
  INV_X1 U12624 ( .A(n16689), .ZN(n11538) );
  INV_X1 U12625 ( .A(n16803), .ZN(n14956) );
  NAND2_X1 U12626 ( .A1(n10804), .A2(n11659), .ZN(n14268) );
  NAND2_X1 U12627 ( .A1(n11060), .A2(n11643), .ZN(n11822) );
  NAND2_X1 U12628 ( .A1(n14442), .A2(n14441), .ZN(n14444) );
  NAND2_X1 U12629 ( .A1(n10864), .A2(n10601), .ZN(n19965) );
  NOR2_X1 U12630 ( .A1(n20199), .A2(n20528), .ZN(n10000) );
  INV_X1 U12631 ( .A(n19961), .ZN(n20522) );
  NOR3_X1 U12632 ( .A1(n10269), .A2(n20329), .A3(n20393), .ZN(n20299) );
  AND2_X1 U12633 ( .A1(n20537), .A2(n19998), .ZN(n20306) );
  NOR2_X2 U12634 ( .A1(n17038), .A2(n17039), .ZN(n19894) );
  NOR2_X2 U12635 ( .A1(n17040), .A2(n17039), .ZN(n19895) );
  INV_X1 U12636 ( .A(n19894), .ZN(n19888) );
  INV_X1 U12637 ( .A(n19895), .ZN(n19889) );
  INV_X1 U12638 ( .A(n20398), .ZN(n20336) );
  NAND2_X1 U12639 ( .A1(n14342), .A2(n14341), .ZN(n14715) );
  AND3_X1 U12640 ( .A1(n11615), .A2(n11619), .A3(n11598), .ZN(n11415) );
  NOR2_X1 U12641 ( .A1(n19510), .A2(n18341), .ZN(n17709) );
  NOR2_X1 U12642 ( .A1(n10703), .A2(n17492), .ZN(n10699) );
  INV_X1 U12643 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10703) );
  NOR2_X1 U12644 ( .A1(n18363), .A2(n10411), .ZN(n10410) );
  AND2_X1 U12645 ( .A1(n18154), .A2(n10409), .ZN(n10408) );
  INV_X1 U12646 ( .A(n18238), .ZN(n10409) );
  NOR2_X1 U12647 ( .A1(n10762), .A2(n10761), .ZN(n10416) );
  NOR2_X1 U12648 ( .A1(n9928), .A2(n9925), .ZN(n10415) );
  INV_X1 U12649 ( .A(n12046), .ZN(n10761) );
  NOR2_X1 U12650 ( .A1(n19573), .A2(n17357), .ZN(n18300) );
  AOI21_X1 U12651 ( .B1(n18430), .B2(n18573), .A(n18429), .ZN(n18420) );
  INV_X1 U12652 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18497) );
  NOR2_X1 U12653 ( .A1(n18520), .A2(n21610), .ZN(n18496) );
  NOR2_X1 U12654 ( .A1(n18773), .A2(n18728), .ZN(n18521) );
  NAND2_X1 U12655 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18539) );
  AND2_X1 U12656 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18663) );
  NAND2_X1 U12657 ( .A1(n18663), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18639) );
  NOR2_X1 U12658 ( .A1(n18728), .A2(n18741), .ZN(n18699) );
  NOR2_X1 U12659 ( .A1(n19715), .A2(n19573), .ZN(n17220) );
  NOR2_X1 U12660 ( .A1(n10589), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10588) );
  INV_X1 U12661 ( .A(n17074), .ZN(n10589) );
  NAND2_X1 U12662 ( .A1(n17127), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17213) );
  NAND2_X1 U12663 ( .A1(n17263), .A2(n18267), .ZN(n10423) );
  OAI21_X1 U12664 ( .B1(n18419), .B2(n10424), .A(n17262), .ZN(n9972) );
  NOR2_X1 U12665 ( .A1(n18430), .A2(n17267), .ZN(n10424) );
  INV_X1 U12666 ( .A(n18455), .ZN(n18467) );
  INV_X1 U12667 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18805) );
  INV_X1 U12668 ( .A(n18476), .ZN(n18530) );
  INV_X1 U12669 ( .A(n18513), .ZN(n9947) );
  NAND2_X1 U12670 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10765) );
  OR2_X1 U12671 ( .A1(n18863), .A2(n18985), .ZN(n18907) );
  NAND2_X1 U12672 ( .A1(n10591), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10590) );
  NAND2_X1 U12673 ( .A1(n18689), .A2(n9905), .ZN(n9975) );
  INV_X1 U12674 ( .A(n12099), .ZN(n10591) );
  NAND2_X1 U12675 ( .A1(n18713), .A2(n12092), .ZN(n10740) );
  XNOR2_X1 U12676 ( .A(n12090), .B(n12089), .ZN(n18714) );
  INV_X1 U12677 ( .A(n12091), .ZN(n12089) );
  NAND2_X1 U12678 ( .A1(n18714), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18713) );
  NOR2_X1 U12679 ( .A1(n10660), .A2(n18726), .ZN(n10659) );
  INV_X1 U12680 ( .A(n10662), .ZN(n10660) );
  NOR2_X1 U12681 ( .A1(n18749), .A2(n12123), .ZN(n18739) );
  XNOR2_X1 U12682 ( .A(n12081), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18754) );
  INV_X1 U12683 ( .A(n18820), .ZN(n19509) );
  INV_X1 U12684 ( .A(n11958), .ZN(n10366) );
  AOI21_X1 U12685 ( .B1(n12194), .B2(n12193), .A(n12192), .ZN(n19513) );
  NAND2_X1 U12686 ( .A1(n19528), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n19530) );
  INV_X1 U12687 ( .A(n19528), .ZN(n19533) );
  INV_X1 U12688 ( .A(n19521), .ZN(n10398) );
  INV_X1 U12689 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19553) );
  NOR2_X1 U12690 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19152) );
  NAND2_X1 U12691 ( .A1(n19072), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19316) );
  NOR2_X1 U12692 ( .A1(n11995), .A2(n11994), .ZN(n19076) );
  INV_X1 U12693 ( .A(n12100), .ZN(n19095) );
  INV_X1 U12694 ( .A(n18156), .ZN(n19099) );
  OR2_X1 U12695 ( .A1(n14050), .A2(n20561), .ZN(n14043) );
  AND2_X1 U12696 ( .A1(n14055), .A2(n13528), .ZN(n14980) );
  NOR3_X1 U12697 ( .A1(n15063), .A2(n9912), .A3(n10681), .ZN(n13429) );
  OR2_X1 U12698 ( .A1(n10684), .A2(n10682), .ZN(n10681) );
  NOR2_X1 U12699 ( .A1(n15063), .A2(n21373), .ZN(n15059) );
  AND2_X1 U12700 ( .A1(n15115), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15127) );
  OR2_X1 U12701 ( .A1(n15188), .A2(n13416), .ZN(n15177) );
  NAND2_X1 U12702 ( .A1(n20606), .A2(n9774), .ZN(n15266) );
  OAI21_X1 U12703 ( .B1(n20637), .B2(n15653), .A(n10441), .ZN(n14902) );
  INV_X1 U12704 ( .A(n10442), .ZN(n10441) );
  OAI22_X1 U12705 ( .A1(n20610), .A2(n14898), .B1(n20648), .B2(n15883), .ZN(
        n10442) );
  INV_X1 U12706 ( .A(n20608), .ZN(n20636) );
  NAND2_X1 U12707 ( .A1(n20606), .A2(n13410), .ZN(n20594) );
  INV_X1 U12708 ( .A(n15269), .ZN(n20601) );
  NOR2_X1 U12709 ( .A1(n21353), .A2(n20632), .ZN(n20606) );
  AND2_X1 U12710 ( .A1(n20638), .A2(n9767), .ZN(n15281) );
  NAND2_X1 U12711 ( .A1(n20638), .A2(n10679), .ZN(n20645) );
  AND2_X1 U12712 ( .A1(n20638), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20608) );
  MUX2_X1 U12713 ( .A(n14989), .B(n13528), .S(n14986), .Z(n13530) );
  AND2_X1 U12714 ( .A1(n20655), .A2(n20826), .ZN(n20650) );
  AND2_X1 U12715 ( .A1(n14165), .A2(n14295), .ZN(n20655) );
  OR2_X1 U12716 ( .A1(n14877), .A2(n15405), .ZN(n15399) );
  NOR2_X2 U12717 ( .A1(n14877), .A2(n15350), .ZN(n15401) );
  OR2_X1 U12718 ( .A1(n15324), .A2(n15323), .ZN(n15661) );
  INV_X1 U12719 ( .A(n14877), .ZN(n14591) );
  AND2_X1 U12720 ( .A1(n14584), .A2(n14583), .ZN(n14585) );
  OR2_X1 U12721 ( .A1(n14579), .A2(n14578), .ZN(n14586) );
  AND2_X1 U12722 ( .A1(n14299), .A2(n17111), .ZN(n20671) );
  INV_X2 U12723 ( .A(n20678), .ZN(n20683) );
  AND2_X1 U12724 ( .A1(n21412), .A2(n21341), .ZN(n14383) );
  INV_X1 U12725 ( .A(n15307), .ZN(n15520) );
  INV_X1 U12726 ( .A(n15573), .ZN(n20715) );
  XNOR2_X1 U12727 ( .A(n10911), .B(n14186), .ZN(n13971) );
  NAND2_X1 U12728 ( .A1(n10905), .A2(n10464), .ZN(n10911) );
  NAND2_X1 U12729 ( .A1(n15456), .A2(n10465), .ZN(n10464) );
  NOR2_X1 U12730 ( .A1(n15300), .A2(n20774), .ZN(n10327) );
  NAND2_X1 U12731 ( .A1(n10053), .A2(n10052), .ZN(n15457) );
  NAND2_X1 U12732 ( .A1(n15455), .A2(n9689), .ZN(n10052) );
  NAND2_X1 U12733 ( .A1(n15456), .A2(n15621), .ZN(n10053) );
  AND2_X1 U12734 ( .A1(n13953), .A2(n10566), .ZN(n15710) );
  NAND2_X1 U12735 ( .A1(n15714), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10566) );
  NOR2_X1 U12736 ( .A1(n15152), .A2(n15153), .ZN(n15145) );
  NAND2_X1 U12737 ( .A1(n10713), .A2(n15657), .ZN(n15649) );
  NAND2_X1 U12738 ( .A1(n15659), .A2(n15658), .ZN(n10713) );
  NAND2_X1 U12739 ( .A1(n17143), .A2(n13852), .ZN(n14612) );
  OR2_X1 U12740 ( .A1(n20755), .A2(n20754), .ZN(n14620) );
  AND2_X1 U12741 ( .A1(n13946), .A2(n13945), .ZN(n20772) );
  INV_X1 U12742 ( .A(n20784), .ZN(n13816) );
  INV_X1 U12743 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21157) );
  OR2_X1 U12744 ( .A1(n14579), .A2(n21091), .ZN(n15929) );
  NOR2_X1 U12745 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17163) );
  NAND2_X1 U12746 ( .A1(n14563), .A2(n14562), .ZN(n20849) );
  INV_X1 U12747 ( .A(n20866), .ZN(n20875) );
  INV_X1 U12748 ( .A(n20927), .ZN(n20938) );
  NAND2_X1 U12749 ( .A1(n21008), .A2(n20916), .ZN(n20970) );
  OAI21_X1 U12750 ( .B1(n12779), .B2(n21006), .A(n21272), .ZN(n21026) );
  OAI211_X1 U12751 ( .C1(n21054), .C2(n21091), .A(n21096), .B(n21037), .ZN(
        n21056) );
  INV_X1 U12752 ( .A(n21044), .ZN(n21055) );
  OR2_X1 U12753 ( .A1(n21126), .A2(n21206), .ZN(n21084) );
  OR2_X1 U12754 ( .A1(n21126), .A2(n21231), .ZN(n21133) );
  OAI211_X1 U12755 ( .C1(n21162), .C2(n21201), .A(n21236), .B(n21161), .ZN(
        n21194) );
  AOI22_X1 U12756 ( .A1(n21160), .A2(n21155), .B1(n21154), .B2(n21162), .ZN(
        n21198) );
  OR2_X1 U12757 ( .A1(n20825), .A2(n20824), .ZN(n21197) );
  INV_X1 U12758 ( .A(n21213), .ZN(n21224) );
  OAI211_X1 U12759 ( .C1(n21254), .C2(n21237), .A(n21236), .B(n21235), .ZN(
        n21256) );
  INV_X1 U12760 ( .A(n21244), .ZN(n21255) );
  AND2_X1 U12761 ( .A1(n20919), .A2(n15396), .ZN(n21264) );
  INV_X1 U12762 ( .A(n20790), .ZN(n21263) );
  AND2_X1 U12763 ( .A1(n20919), .A2(n14554), .ZN(n21280) );
  INV_X1 U12764 ( .A(n20800), .ZN(n21279) );
  INV_X1 U12765 ( .A(n21326), .ZN(n21288) );
  AND2_X1 U12766 ( .A1(n20919), .A2(n20803), .ZN(n21286) );
  AND2_X1 U12767 ( .A1(n20919), .A2(n20807), .ZN(n21294) );
  INV_X1 U12768 ( .A(n20813), .ZN(n21301) );
  AND2_X1 U12769 ( .A1(n20919), .A2(n20811), .ZN(n21300) );
  INV_X1 U12770 ( .A(n20817), .ZN(n21307) );
  INV_X1 U12771 ( .A(n20821), .ZN(n21313) );
  AND2_X1 U12772 ( .A1(n20919), .A2(n20820), .ZN(n21312) );
  OR2_X1 U12773 ( .A1(n21265), .A2(n21125), .ZN(n21326) );
  INV_X1 U12774 ( .A(n21291), .ZN(n21322) );
  INV_X1 U12775 ( .A(n21197), .ZN(n21318) );
  INV_X1 U12776 ( .A(n15929), .ZN(n17123) );
  NAND2_X1 U12777 ( .A1(n21201), .A2(n17174), .ZN(n17172) );
  INV_X1 U12778 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17174) );
  NAND2_X1 U12779 ( .A1(n17174), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21329) );
  NAND2_X1 U12780 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17177) );
  INV_X1 U12781 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21091) );
  AOI221_X1 U12782 ( .B1(n17176), .B2(n17174), .C1(n17118), .C2(n17174), .A(
        n17169), .ZN(n17175) );
  NAND2_X1 U12783 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21409) );
  NAND2_X1 U12784 ( .A1(n10531), .A2(n9682), .ZN(n15968) );
  OAI21_X1 U12785 ( .B1(n11516), .B2(n9885), .A(n10263), .ZN(n11521) );
  NAND2_X1 U12786 ( .A1(n11516), .A2(n19879), .ZN(n10263) );
  INV_X1 U12787 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n21703) );
  NAND2_X1 U12788 ( .A1(n16229), .A2(n16709), .ZN(n19799) );
  INV_X1 U12789 ( .A(n19809), .ZN(n19791) );
  XNOR2_X1 U12790 ( .A(n14292), .B(n14291), .ZN(n20524) );
  NAND2_X1 U12791 ( .A1(n11156), .A2(n10194), .ZN(n10193) );
  INV_X1 U12792 ( .A(n11154), .ZN(n10194) );
  INV_X1 U12793 ( .A(n19807), .ZN(n19774) );
  OR2_X1 U12794 ( .A1(n11789), .A2(n11788), .ZN(n14826) );
  OR2_X1 U12795 ( .A1(n11736), .A2(n11735), .ZN(n14848) );
  NAND2_X1 U12796 ( .A1(n10449), .A2(n14780), .ZN(n10025) );
  NAND2_X1 U12797 ( .A1(n16290), .A2(n10246), .ZN(n16286) );
  INV_X1 U12798 ( .A(n12293), .ZN(n16317) );
  AND2_X1 U12799 ( .A1(n19840), .A2(n14814), .ZN(n16466) );
  NAND2_X1 U12800 ( .A1(n14774), .A2(n11692), .ZN(n14289) );
  AND2_X1 U12801 ( .A1(n16475), .A2(n16441), .ZN(n19836) );
  NAND2_X1 U12802 ( .A1(n14548), .A2(n12231), .ZN(n14779) );
  NAND2_X1 U12803 ( .A1(n19840), .A2(n14265), .ZN(n19834) );
  INV_X1 U12804 ( .A(n17033), .ZN(n20116) );
  INV_X1 U12805 ( .A(n19840), .ZN(n16465) );
  INV_X1 U12806 ( .A(n16441), .ZN(n16472) );
  INV_X1 U12807 ( .A(n14360), .ZN(n14373) );
  INV_X1 U12808 ( .A(n19842), .ZN(n19860) );
  INV_X1 U12809 ( .A(n15940), .ZN(n19859) );
  NAND2_X1 U12810 ( .A1(n14229), .A2(n20450), .ZN(n19862) );
  NAND2_X1 U12811 ( .A1(n14228), .A2(n14154), .ZN(n14229) );
  NAND2_X1 U12812 ( .A1(n19862), .A2(n15940), .ZN(n19842) );
  INV_X2 U12813 ( .A(n14066), .ZN(n14151) );
  NAND2_X1 U12814 ( .A1(n14154), .A2(n14067), .ZN(n14066) );
  NOR2_X1 U12815 ( .A1(n16712), .A2(n10480), .ZN(n10479) );
  INV_X1 U12816 ( .A(n10483), .ZN(n10480) );
  NAND2_X1 U12817 ( .A1(n16493), .A2(n16715), .ZN(n10709) );
  INV_X1 U12818 ( .A(n16492), .ZN(n10708) );
  INV_X1 U12819 ( .A(n10926), .ZN(n16725) );
  NAND2_X1 U12820 ( .A1(n16802), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16543) );
  INV_X1 U12821 ( .A(n13774), .ZN(n10500) );
  NAND2_X1 U12822 ( .A1(n13745), .A2(n10495), .ZN(n10493) );
  AND2_X1 U12823 ( .A1(n10499), .A2(n13744), .ZN(n10495) );
  AND2_X1 U12824 ( .A1(n10496), .A2(n16944), .ZN(n10492) );
  NAND2_X1 U12825 ( .A1(n16993), .A2(n10483), .ZN(n10091) );
  INV_X1 U12826 ( .A(n10478), .ZN(n10092) );
  NAND2_X1 U12827 ( .A1(n9985), .A2(n13768), .ZN(n10481) );
  INV_X1 U12828 ( .A(n14913), .ZN(n9985) );
  XNOR2_X1 U12829 ( .A(n13779), .B(n13778), .ZN(n10116) );
  NAND2_X1 U12830 ( .A1(n10007), .A2(n10602), .ZN(n13779) );
  AOI21_X1 U12831 ( .B1(n10603), .B2(n10605), .A(n16498), .ZN(n10602) );
  XNOR2_X1 U12832 ( .A(n10141), .B(n10296), .ZN(n16774) );
  INV_X1 U12833 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10296) );
  INV_X1 U12834 ( .A(n11530), .ZN(n10312) );
  NAND2_X1 U12835 ( .A1(n11530), .A2(n10319), .ZN(n10313) );
  NOR2_X1 U12836 ( .A1(n9759), .A2(n11868), .ZN(n10319) );
  OR2_X1 U12837 ( .A1(n13599), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U12838 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16825), .ZN(
        n10470) );
  XNOR2_X1 U12839 ( .A(n10107), .B(n9879), .ZN(n16867) );
  NAND2_X1 U12840 ( .A1(n16582), .A2(n16586), .ZN(n10107) );
  AND2_X1 U12841 ( .A1(n16588), .A2(n16993), .ZN(n10196) );
  INV_X1 U12842 ( .A(n10295), .ZN(n10294) );
  INV_X1 U12843 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17017) );
  NOR2_X1 U12844 ( .A1(n20343), .A2(n20198), .ZN(n20521) );
  INV_X1 U12845 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U12846 ( .A1(n12228), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20528), .B2(n20338), .ZN(n12216) );
  INV_X1 U12847 ( .A(n20524), .ZN(n19998) );
  NAND2_X1 U12848 ( .A1(n12210), .A2(n14687), .ZN(n14673) );
  AND2_X1 U12849 ( .A1(n17008), .A2(n17007), .ZN(n17026) );
  AND2_X1 U12850 ( .A1(n10278), .A2(n20300), .ZN(n17035) );
  AND2_X1 U12851 ( .A1(n20057), .A2(n20522), .ZN(n19989) );
  OAI21_X1 U12852 ( .B1(n20030), .B2(n20029), .A(n20028), .ZN(n20052) );
  OAI21_X1 U12853 ( .B1(n20063), .B2(n20079), .A(n20403), .ZN(n20082) );
  INV_X1 U12854 ( .A(n20074), .ZN(n20081) );
  OR2_X1 U12855 ( .A1(n20094), .A2(n20093), .ZN(n20112) );
  AOI21_X1 U12856 ( .B1(n20393), .B2(n20089), .A(n20088), .ZN(n20111) );
  NOR2_X1 U12857 ( .A1(n20119), .A2(n10071), .ZN(n20120) );
  AND2_X1 U12858 ( .A1(n20159), .A2(n20158), .ZN(n20171) );
  NAND2_X1 U12859 ( .A1(n10001), .A2(n10000), .ZN(n20157) );
  INV_X1 U12860 ( .A(n20171), .ZN(n20191) );
  OAI21_X1 U12861 ( .B1(n20225), .B2(n20197), .A(n20196), .ZN(n20220) );
  INV_X1 U12862 ( .A(n20252), .ZN(n20260) );
  AND2_X1 U12863 ( .A1(n20237), .A2(n20236), .ZN(n20259) );
  NAND2_X1 U12864 ( .A1(n10073), .A2(n10127), .ZN(n20274) );
  NOR2_X1 U12865 ( .A1(n20290), .A2(n20528), .ZN(n10127) );
  INV_X1 U12866 ( .A(n20352), .ZN(n21741) );
  OAI22_X1 U12867 ( .A1(n19890), .A2(n19889), .B1(n21561), .B2(n19888), .ZN(
        n20331) );
  OR2_X1 U12868 ( .A1(n19891), .A2(n19879), .ZN(n20372) );
  INV_X1 U12869 ( .A(n20357), .ZN(n20409) );
  INV_X1 U12870 ( .A(n20362), .ZN(n20415) );
  INV_X1 U12871 ( .A(n20371), .ZN(n20423) );
  INV_X1 U12872 ( .A(n20367), .ZN(n20421) );
  INV_X1 U12873 ( .A(n20372), .ZN(n20427) );
  INV_X1 U12874 ( .A(n20144), .ZN(n20433) );
  INV_X1 U12875 ( .A(n20381), .ZN(n20439) );
  AND2_X1 U12876 ( .A1(n20402), .A2(n20394), .ZN(n21744) );
  INV_X1 U12877 ( .A(n20331), .ZN(n20444) );
  INV_X1 U12878 ( .A(n15934), .ZN(n20450) );
  INV_X1 U12879 ( .A(n17709), .ZN(n19728) );
  NAND2_X1 U12880 ( .A1(n17397), .A2(n17562), .ZN(n10693) );
  INV_X1 U12881 ( .A(n18663), .ZN(n18676) );
  NOR2_X2 U12882 ( .A1(n19666), .A2(n17751), .ZN(n17715) );
  INV_X1 U12883 ( .A(n17752), .ZN(n17764) );
  NOR2_X2 U12884 ( .A1(n19566), .A2(n17385), .ZN(n17736) );
  INV_X1 U12885 ( .A(n17736), .ZN(n17757) );
  NAND3_X1 U12886 ( .A1(n17655), .A2(n19728), .A3(n19571), .ZN(n17767) );
  NOR2_X1 U12887 ( .A1(n17901), .A2(n17873), .ZN(n17904) );
  AND2_X1 U12888 ( .A1(n17935), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17947) );
  AND2_X1 U12889 ( .A1(n18055), .A2(n9772), .ZN(n17985) );
  NAND2_X1 U12890 ( .A1(n18055), .A2(n9769), .ZN(n17998) );
  NOR2_X1 U12891 ( .A1(n18030), .A2(n17604), .ZN(n10698) );
  NAND2_X1 U12892 ( .A1(n18055), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n18027) );
  AND2_X1 U12893 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18068), .ZN(n18055) );
  INV_X1 U12894 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18069) );
  NOR2_X1 U12895 ( .A1(n18087), .A2(n18069), .ZN(n18068) );
  OR2_X1 U12896 ( .A1(n18102), .A2(n18072), .ZN(n18087) );
  NAND2_X1 U12897 ( .A1(n18120), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n18102) );
  NAND2_X1 U12898 ( .A1(n18182), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18181) );
  NOR2_X1 U12899 ( .A1(n10373), .A2(n10372), .ZN(n10371) );
  INV_X1 U12900 ( .A(n11973), .ZN(n10373) );
  NOR3_X1 U12901 ( .A1(n18230), .A2(n18354), .A3(n18352), .ZN(n18155) );
  NOR2_X1 U12902 ( .A1(n18348), .A2(n18223), .ZN(n18217) );
  NAND2_X1 U12903 ( .A1(n17142), .A2(n10407), .ZN(n18230) );
  NOR2_X1 U12904 ( .A1(n9768), .A2(n21640), .ZN(n10407) );
  INV_X1 U12905 ( .A(n18207), .ZN(n18229) );
  NOR2_X1 U12906 ( .A1(n18291), .A2(n9768), .ZN(n18234) );
  NAND2_X1 U12907 ( .A1(n17142), .A2(n10408), .ZN(n18239) );
  NOR2_X1 U12908 ( .A1(n12019), .A2(n12018), .ZN(n18271) );
  INV_X1 U12909 ( .A(n12131), .ZN(n18274) );
  INV_X1 U12910 ( .A(n18282), .ZN(n12124) );
  INV_X1 U12911 ( .A(n18292), .ZN(n18290) );
  NOR2_X1 U12912 ( .A1(n9959), .A2(n9958), .ZN(n12078) );
  NAND2_X1 U12913 ( .A1(n18335), .A2(n18340), .ZN(n18322) );
  NOR2_X1 U12914 ( .A1(n18341), .A2(n19567), .ZN(n18397) );
  NAND2_X1 U12915 ( .A1(n18641), .A2(n9717), .ZN(n18564) );
  AND2_X1 U12916 ( .A1(n18655), .A2(n17077), .ZN(n9722) );
  INV_X1 U12917 ( .A(n12200), .ZN(n18887) );
  NAND2_X1 U12918 ( .A1(n18641), .A2(n9721), .ZN(n18601) );
  OAI21_X1 U12919 ( .B1(n18777), .B2(n18940), .A(n10359), .ZN(n18655) );
  NAND2_X1 U12920 ( .A1(n18684), .A2(n18943), .ZN(n10359) );
  INV_X1 U12921 ( .A(n18655), .ZN(n18672) );
  INV_X1 U12922 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18703) );
  INV_X1 U12923 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18729) );
  INV_X2 U12924 ( .A(n19221), .ZN(n19455) );
  INV_X1 U12925 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18768) );
  OAI21_X2 U12926 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19710), .A(n17364), 
        .ZN(n18772) );
  NAND2_X1 U12927 ( .A1(n18429), .A2(n17074), .ZN(n17128) );
  NAND2_X1 U12928 ( .A1(n10426), .A2(n10429), .ZN(n12205) );
  INV_X1 U12929 ( .A(n10428), .ZN(n17073) );
  INV_X1 U12930 ( .A(n10747), .ZN(n18454) );
  OAI21_X1 U12931 ( .B1(n18808), .B2(n18970), .A(n10670), .ZN(n10669) );
  NAND2_X1 U12932 ( .A1(n19040), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n10670) );
  NOR2_X1 U12933 ( .A1(n18880), .A2(n18811), .ZN(n10673) );
  NOR2_X1 U12934 ( .A1(n18963), .A2(n10592), .ZN(n10672) );
  AOI21_X1 U12935 ( .B1(n18824), .B2(n18828), .A(n19054), .ZN(n10770) );
  OR2_X1 U12936 ( .A1(n18840), .A2(n10772), .ZN(n10771) );
  NAND2_X1 U12937 ( .A1(n18825), .A2(n10773), .ZN(n10772) );
  NOR2_X1 U12938 ( .A1(n18822), .A2(n18828), .ZN(n10773) );
  AOI21_X1 U12939 ( .B1(n18846), .B2(n10933), .A(n18963), .ZN(n18852) );
  INV_X1 U12940 ( .A(n10744), .ZN(n18561) );
  NAND2_X1 U12941 ( .A1(n12154), .A2(n18903), .ZN(n18606) );
  INV_X1 U12942 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18966) );
  INV_X1 U12943 ( .A(n9963), .ZN(n18681) );
  INV_X1 U12944 ( .A(n10657), .ZN(n18705) );
  AND2_X1 U12945 ( .A1(n10228), .A2(n10227), .ZN(n18722) );
  NAND2_X1 U12946 ( .A1(n18734), .A2(n19026), .ZN(n10228) );
  INV_X1 U12947 ( .A(n18734), .ZN(n10741) );
  INV_X1 U12948 ( .A(n10227), .ZN(n12083) );
  INV_X2 U12949 ( .A(n19049), .ZN(n19548) );
  INV_X1 U12950 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19072) );
  INV_X1 U12951 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19557) );
  NAND2_X1 U12952 ( .A1(n19560), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19219) );
  AOI22_X1 U12953 ( .A1(n19548), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19696), .B2(n19551), .ZN(n19691) );
  AOI211_X1 U12954 ( .C1(n19711), .C2(n19545), .A(n19075), .B(n14858), .ZN(
        n19697) );
  INV_X1 U12955 ( .A(n19711), .ZN(n19573) );
  AND2_X1 U12956 ( .A1(n10633), .A2(n10626), .ZN(n19574) );
  OR2_X1 U12957 ( .A1(n19561), .A2(n19562), .ZN(n10633) );
  NOR2_X1 U12958 ( .A1(n10629), .A2(n10627), .ZN(n10626) );
  NAND2_X1 U12959 ( .A1(n19676), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19578) );
  INV_X1 U12960 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19666) );
  CLKBUF_X1 U12961 ( .A(n19655), .Z(n19648) );
  NAND2_X1 U12962 ( .A1(n19598), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19724) );
  AND2_X2 U12963 ( .A1(n13999), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15350)
         );
  CLKBUF_X1 U12964 ( .A(n17338), .Z(n17349) );
  OAI21_X1 U12965 ( .B1(n15000), .B2(n21386), .A(n10150), .ZN(n14889) );
  AND2_X1 U12966 ( .A1(n10153), .A2(n10151), .ZN(n10150) );
  NOR3_X1 U12967 ( .A1(n15063), .A2(n9912), .A3(n21373), .ZN(n15006) );
  AOI21_X1 U12968 ( .B1(n14888), .B2(n15517), .A(n14869), .ZN(n10781) );
  NAND2_X1 U12969 ( .A1(n10328), .A2(n10326), .ZN(P1_U3000) );
  NOR2_X1 U12970 ( .A1(n10716), .A2(n10327), .ZN(n10326) );
  NAND2_X1 U12971 ( .A1(n13971), .A2(n20757), .ZN(n10328) );
  INV_X1 U12972 ( .A(n13969), .ZN(n10716) );
  OAI21_X1 U12973 ( .B1(n15685), .B2(n20775), .A(n15684), .ZN(P1_U3001) );
  OAI21_X1 U12974 ( .B1(n10509), .B2(n16242), .A(n10508), .ZN(n13743) );
  INV_X1 U12975 ( .A(n10726), .ZN(n10725) );
  OAI21_X1 U12976 ( .B1(n15945), .B2(n16238), .A(n10727), .ZN(n10726) );
  AOI21_X1 U12977 ( .B1(n19819), .B2(n12210), .A(n16253), .ZN(n16254) );
  NOR2_X1 U12978 ( .A1(n10941), .A2(n10934), .ZN(n12508) );
  INV_X1 U12979 ( .A(n16391), .ZN(n16385) );
  NAND2_X1 U12980 ( .A1(n10010), .A2(n10009), .ZN(n14525) );
  OAI211_X1 U12981 ( .C1(n15340), .C2(n14819), .A(n16361), .B(n9790), .ZN(
        n16362) );
  NAND2_X1 U12982 ( .A1(n10421), .A2(n16697), .ZN(n10374) );
  NAND2_X1 U12983 ( .A1(n14920), .A2(n14919), .ZN(n14921) );
  INV_X1 U12984 ( .A(n9923), .ZN(n16482) );
  OAI21_X1 U12985 ( .B1(n16479), .B2(n16712), .A(n10643), .ZN(n9923) );
  OAI211_X1 U12986 ( .C1(n16509), .C2(n10237), .A(n10240), .B(n10236), .ZN(
        n10239) );
  INV_X1 U12987 ( .A(n10242), .ZN(n10237) );
  INV_X1 U12988 ( .A(n10208), .ZN(n10207) );
  NAND2_X1 U12989 ( .A1(n9839), .A2(n9822), .ZN(n10206) );
  NAND2_X1 U12990 ( .A1(n10164), .A2(n11531), .ZN(n10163) );
  NAND2_X1 U12991 ( .A1(n10158), .A2(n16697), .ZN(n11597) );
  AOI21_X1 U12992 ( .B1(n16836), .B2(n16715), .A(n16560), .ZN(n10213) );
  NAND2_X1 U12993 ( .A1(n10477), .A2(n11531), .ZN(n10476) );
  INV_X1 U12994 ( .A(n10283), .ZN(n16572) );
  AOI21_X1 U12995 ( .B1(n16852), .B2(n16715), .A(n16571), .ZN(n10284) );
  NAND2_X1 U12996 ( .A1(n10323), .A2(n10195), .ZN(n16601) );
  AOI21_X1 U12997 ( .B1(n16932), .B2(n11531), .A(n16644), .ZN(n16645) );
  NAND2_X1 U12998 ( .A1(n10421), .A2(n16993), .ZN(n10420) );
  NAND2_X1 U12999 ( .A1(n14935), .A2(n16993), .ZN(n10799) );
  NAND2_X1 U13000 ( .A1(n14934), .A2(n14933), .ZN(n10801) );
  OAI211_X1 U13001 ( .C1(n16483), .C2(n17182), .A(n10279), .B(n10593), .ZN(
        P2_U3018) );
  NAND2_X1 U13002 ( .A1(n10280), .A2(n16993), .ZN(n10279) );
  NAND2_X1 U13003 ( .A1(n10710), .A2(n10614), .ZN(n16726) );
  NAND2_X1 U13004 ( .A1(n10238), .A2(n10240), .ZN(n16741) );
  NAND2_X1 U13005 ( .A1(n10147), .A2(n10242), .ZN(n10238) );
  AOI21_X1 U13006 ( .B1(n10164), .B2(n16944), .A(n9840), .ZN(n9986) );
  NAND2_X1 U13007 ( .A1(n10135), .A2(n16944), .ZN(n10139) );
  NAND2_X1 U13008 ( .A1(n10158), .A2(n16993), .ZN(n9968) );
  INV_X1 U13009 ( .A(n16775), .ZN(n16788) );
  INV_X1 U13010 ( .A(n16817), .ZN(n10624) );
  INV_X1 U13011 ( .A(n10468), .ZN(n16824) );
  INV_X1 U13012 ( .A(n10338), .ZN(n16837) );
  NOR2_X1 U13013 ( .A1(n16835), .A2(n9800), .ZN(n10339) );
  AOI21_X1 U13014 ( .B1(n17416), .B2(n17745), .A(n17415), .ZN(n17419) );
  OR2_X1 U13015 ( .A1(n17887), .A2(n17886), .ZN(n10696) );
  NOR2_X1 U13016 ( .A1(n18291), .A2(n18238), .ZN(n18262) );
  INV_X1 U13017 ( .A(n10750), .ZN(n10587) );
  NAND2_X1 U13018 ( .A1(n10755), .A2(n18669), .ZN(n10586) );
  INV_X1 U13019 ( .A(n10752), .ZN(n10751) );
  NAND2_X1 U13020 ( .A1(n10750), .A2(n10749), .ZN(n10748) );
  OAI21_X1 U13021 ( .B1(n17260), .B2(n19062), .A(n10753), .ZN(n10752) );
  NAND2_X1 U13022 ( .A1(n9945), .A2(n9971), .ZN(n9944) );
  NAND2_X1 U13023 ( .A1(n10671), .A2(n10667), .ZN(P3_U2838) );
  AND2_X1 U13024 ( .A1(n18807), .A2(n10668), .ZN(n10667) );
  OAI21_X1 U13025 ( .B1(n10674), .B2(n10673), .A(n10672), .ZN(n10671) );
  INV_X1 U13026 ( .A(n10669), .ZN(n10668) );
  INV_X1 U13027 ( .A(n10674), .ZN(n18812) );
  NAND2_X1 U13028 ( .A1(n10769), .A2(n10767), .ZN(P3_U2840) );
  AOI21_X1 U13029 ( .B1(n18826), .B2(n18962), .A(n10768), .ZN(n10767) );
  OAI21_X1 U13030 ( .B1(n18831), .B2(n10771), .A(n10770), .ZN(n10769) );
  OAI21_X1 U13031 ( .B1(n19053), .B2(n18828), .A(n18827), .ZN(n10768) );
  NAND2_X1 U13032 ( .A1(n17274), .A2(U214), .ZN(U212) );
  OR2_X2 U13033 ( .A1(n11922), .A2(n19536), .ZN(n9778) );
  AND2_X1 U13034 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9715) );
  INV_X2 U13035 ( .A(n11411), .ZN(n11217) );
  NAND2_X2 U13036 ( .A1(n9974), .A2(n9973), .ZN(n11969) );
  OR2_X1 U13037 ( .A1(n15101), .A2(n9875), .ZN(n9716) );
  INV_X1 U13038 ( .A(n9703), .ZN(n10082) );
  AND2_X1 U13039 ( .A1(n9735), .A2(n10937), .ZN(n9717) );
  AND2_X1 U13040 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9718) );
  INV_X1 U13041 ( .A(n11173), .ZN(n11178) );
  INV_X1 U13042 ( .A(n11178), .ZN(n10215) );
  AND3_X1 U13043 ( .A1(n9857), .A2(n9751), .A3(n11970), .ZN(n9720) );
  AND2_X1 U13044 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U13045 ( .A1(n11184), .A2(n9683), .ZN(n11205) );
  INV_X1 U13046 ( .A(n12040), .ZN(n11999) );
  AND2_X1 U13047 ( .A1(n10925), .A2(n10692), .ZN(n9723) );
  INV_X1 U13048 ( .A(n12212), .ZN(n10856) );
  NAND2_X1 U13049 ( .A1(n15165), .A2(n10779), .ZN(n9724) );
  NOR3_X1 U13050 ( .A1(n15063), .A2(n9912), .A3(n10684), .ZN(n9725) );
  NOR2_X1 U13051 ( .A1(n11486), .A2(n10904), .ZN(n9726) );
  AND2_X1 U13052 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U13053 ( .A1(n18689), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18688) );
  NOR3_X1 U13054 ( .A1(n15101), .A2(n9870), .A3(n15102), .ZN(n15061) );
  NAND2_X1 U13055 ( .A1(n10812), .A2(n11811), .ZN(n16105) );
  INV_X1 U13056 ( .A(n15601), .ZN(n10306) );
  AND3_X1 U13057 ( .A1(n19087), .A2(n10370), .A3(n10360), .ZN(n9728) );
  AND2_X1 U13058 ( .A1(n10721), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9729) );
  AND2_X1 U13059 ( .A1(n9726), .A2(n11499), .ZN(n9730) );
  AND2_X1 U13060 ( .A1(n9727), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9731) );
  AND2_X1 U13061 ( .A1(n9730), .A2(n11501), .ZN(n9732) );
  OR2_X1 U13062 ( .A1(n13646), .A2(n10555), .ZN(n9733) );
  AND2_X1 U13063 ( .A1(n10423), .A2(n17261), .ZN(n9734) );
  AND2_X1 U13064 ( .A1(n9721), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9735) );
  AND3_X1 U13065 ( .A1(n17223), .A2(n9858), .A3(n9969), .ZN(n9736) );
  AND2_X1 U13066 ( .A1(n10944), .A2(n10925), .ZN(n9737) );
  AND4_X1 U13067 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(
        n9738) );
  AND2_X1 U13068 ( .A1(n13752), .A2(n9733), .ZN(n9739) );
  AND3_X1 U13069 ( .A1(n10797), .A2(n11548), .A3(n14735), .ZN(n9740) );
  AND2_X1 U13070 ( .A1(n11436), .A2(n11429), .ZN(n9741) );
  BUF_X2 U13071 ( .A(n12732), .Z(n12749) );
  AND2_X1 U13072 ( .A1(n16487), .A2(n13591), .ZN(n9742) );
  AND2_X1 U13073 ( .A1(n11615), .A2(n11619), .ZN(n9743) );
  INV_X1 U13074 ( .A(n12154), .ZN(n18940) );
  AND2_X1 U13075 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9744) );
  AND2_X1 U13076 ( .A1(n9851), .A2(n10504), .ZN(n9745) );
  AND2_X1 U13077 ( .A1(n18688), .A2(n9798), .ZN(n9746) );
  AND2_X1 U13078 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U13079 ( .A1(n10201), .A2(n11258), .ZN(n10685) );
  INV_X1 U13080 ( .A(n10685), .ZN(n9996) );
  AND2_X1 U13081 ( .A1(n15456), .A2(n15696), .ZN(n9748) );
  AND2_X1 U13082 ( .A1(n9731), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9749) );
  AND3_X1 U13083 ( .A1(n10596), .A2(n13604), .A3(n10594), .ZN(n10547) );
  OR2_X1 U13084 ( .A1(n15974), .A2(n11378), .ZN(n16486) );
  AND4_X1 U13085 ( .A1(n10402), .A2(n10401), .A3(n11971), .A4(n10400), .ZN(
        n9751) );
  OAI21_X1 U13086 ( .B1(n16629), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10599), .ZN(n10486) );
  AND2_X1 U13087 ( .A1(n19818), .A2(n17184), .ZN(n9752) );
  AND3_X1 U13088 ( .A1(n11726), .A2(n11725), .A3(n11724), .ZN(n14257) );
  AND2_X1 U13089 ( .A1(n10082), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9753) );
  AND2_X1 U13090 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9754)
         );
  AND2_X1 U13091 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n9755)
         );
  NAND2_X1 U13092 ( .A1(n10430), .A2(n9818), .ZN(n13603) );
  INV_X1 U13093 ( .A(n13603), .ZN(n10270) );
  INV_X1 U13094 ( .A(n11149), .ZN(n11183) );
  AND2_X1 U13095 ( .A1(n10146), .A2(n10793), .ZN(n9756) );
  AND2_X1 U13096 ( .A1(n9752), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n9757)
         );
  AND2_X1 U13097 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U13098 ( .A1(n13560), .A2(n13551), .ZN(n9759) );
  INV_X1 U13099 ( .A(n13750), .ZN(n10485) );
  NAND2_X1 U13100 ( .A1(n11457), .A2(n10895), .ZN(n11459) );
  OR2_X1 U13101 ( .A1(n13706), .A2(n15997), .ZN(n9760) );
  OR3_X1 U13102 ( .A1(n13706), .A2(n10734), .A3(n15970), .ZN(n9761) );
  AND2_X1 U13103 ( .A1(n16612), .A2(n16625), .ZN(n9762) );
  NAND2_X1 U13104 ( .A1(n16507), .A2(n16511), .ZN(n10793) );
  INV_X1 U13105 ( .A(n10793), .ZN(n10789) );
  AND2_X1 U13106 ( .A1(n12489), .A2(n10794), .ZN(n9763) );
  NOR2_X1 U13107 ( .A1(n16595), .A2(n16888), .ZN(n9764) );
  AND2_X1 U13108 ( .A1(n10778), .A2(n9900), .ZN(n9765) );
  AND2_X1 U13109 ( .A1(n9763), .A2(n13790), .ZN(n9766) );
  AND2_X1 U13110 ( .A1(n10679), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U13111 ( .A1(n10408), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n9768) );
  AND2_X1 U13112 ( .A1(n10698), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n9769) );
  AND2_X1 U13113 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9770) );
  INV_X1 U13114 ( .A(n16266), .ZN(n10461) );
  AND2_X1 U13115 ( .A1(n10443), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9771) );
  NOR2_X1 U13116 ( .A1(n10766), .A2(n10765), .ZN(n10764) );
  AND2_X1 U13117 ( .A1(n9769), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n9772) );
  AND2_X1 U13118 ( .A1(n16811), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9773) );
  NOR2_X2 U13119 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20528) );
  AND2_X1 U13120 ( .A1(n10678), .A2(n13410), .ZN(n9774) );
  AND2_X1 U13121 ( .A1(n10410), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U13122 ( .A1(n9773), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10475) );
  AND2_X1 U13123 ( .A1(n16885), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9776) );
  AND2_X1 U13124 ( .A1(n9776), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9777) );
  INV_X1 U13125 ( .A(n9687), .ZN(n13621) );
  NOR2_X1 U13126 ( .A1(n11924), .A2(n11921), .ZN(n12070) );
  AND2_X2 U13127 ( .A1(n12516), .A2(n14486), .ZN(n12718) );
  AND2_X2 U13128 ( .A1(n12515), .A2(n14178), .ZN(n12734) );
  NAND2_X1 U13129 ( .A1(n11480), .A2(n11479), .ZN(n10575) );
  INV_X1 U13130 ( .A(n10065), .ZN(n10157) );
  INV_X1 U13131 ( .A(n14198), .ZN(n20804) );
  NOR2_X2 U13132 ( .A1(n16959), .A2(n11846), .ZN(n9780) );
  AND2_X1 U13133 ( .A1(n16062), .A2(n10517), .ZN(n9781) );
  INV_X1 U13134 ( .A(n18342), .ZN(n10355) );
  NAND2_X1 U13135 ( .A1(n15165), .A2(n10396), .ZN(n15101) );
  AND2_X1 U13136 ( .A1(n15165), .A2(n10394), .ZN(n15035) );
  XNOR2_X1 U13137 ( .A(n16294), .B(n12404), .ZN(n16281) );
  OR3_X1 U13138 ( .A1(n18520), .A2(n21610), .A3(n10690), .ZN(n9782) );
  AND2_X1 U13139 ( .A1(n10849), .A2(n16272), .ZN(n9783) );
  AND2_X1 U13140 ( .A1(n15165), .A2(n13046), .ZN(n9784) );
  NAND2_X1 U13141 ( .A1(n17935), .A2(n10700), .ZN(n10704) );
  AND2_X1 U13142 ( .A1(n18182), .A2(n10410), .ZN(n9785) );
  AND2_X1 U13143 ( .A1(n15165), .A2(n10778), .ZN(n9786) );
  OR2_X1 U13144 ( .A1(n15101), .A2(n15102), .ZN(n9787) );
  OR2_X1 U13145 ( .A1(n14051), .A2(n20561), .ZN(n9788) );
  NAND2_X1 U13146 ( .A1(n10294), .A2(n10293), .ZN(n16664) );
  AND2_X1 U13147 ( .A1(n11779), .A2(n10826), .ZN(n9789) );
  AND2_X1 U13148 ( .A1(n15165), .A2(n9765), .ZN(n15112) );
  OR2_X1 U13149 ( .A1(n16360), .A2(n16441), .ZN(n9790) );
  NOR2_X1 U13150 ( .A1(n11530), .A2(n11528), .ZN(n9791) );
  NAND3_X1 U13151 ( .A1(n10449), .A2(n14549), .A3(n14780), .ZN(n14548) );
  OR2_X1 U13152 ( .A1(n12140), .A2(n12144), .ZN(n9792) );
  AND2_X1 U13153 ( .A1(n11102), .A2(n10644), .ZN(n9793) );
  AND2_X1 U13154 ( .A1(n18641), .A2(n9735), .ZN(n17395) );
  NAND2_X1 U13155 ( .A1(n19689), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10446) );
  INV_X1 U13156 ( .A(n10446), .ZN(n9974) );
  INV_X2 U13157 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11006) );
  AND2_X1 U13158 ( .A1(n15543), .A2(n10938), .ZN(n9794) );
  OR2_X1 U13159 ( .A1(n16182), .A2(n16641), .ZN(n9795) );
  AND2_X1 U13160 ( .A1(n10330), .A2(n10329), .ZN(n15659) );
  AND2_X1 U13161 ( .A1(n10902), .A2(n16316), .ZN(n9796) );
  AND2_X1 U13162 ( .A1(n10429), .A2(n18445), .ZN(n9797) );
  OAI21_X1 U13163 ( .B1(n16569), .B2(n10582), .A(n10579), .ZN(n16546) );
  AND2_X1 U13164 ( .A1(n12099), .A2(n10759), .ZN(n9798) );
  AND2_X1 U13165 ( .A1(n13601), .A2(n16647), .ZN(n16636) );
  INV_X1 U13166 ( .A(n12113), .ZN(n19087) );
  INV_X1 U13167 ( .A(n19778), .ZN(n19798) );
  AND2_X1 U13168 ( .A1(n10613), .A2(n16214), .ZN(n9799) );
  AND2_X1 U13169 ( .A1(n16836), .A2(n16970), .ZN(n9800) );
  AND2_X1 U13170 ( .A1(n14912), .A2(n14911), .ZN(n9801) );
  AND2_X1 U13171 ( .A1(n19546), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9802) );
  AND4_X1 U13172 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n9803) );
  AND4_X1 U13173 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n9804) );
  AND4_X1 U13174 ( .A1(n11300), .A2(n11299), .A3(n11293), .A4(n11294), .ZN(
        n9805) );
  AND3_X1 U13175 ( .A1(n13559), .A2(n13558), .A3(n13560), .ZN(n9806) );
  NAND2_X1 U13176 ( .A1(n13605), .A2(n13607), .ZN(n13606) );
  NAND2_X1 U13177 ( .A1(n10193), .A2(n11141), .ZN(n19818) );
  AND2_X1 U13178 ( .A1(n13677), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13676) );
  NAND2_X1 U13179 ( .A1(n10744), .A2(n18673), .ZN(n18476) );
  NAND2_X1 U13180 ( .A1(n9804), .A2(n9738), .ZN(n11653) );
  OR2_X1 U13181 ( .A1(n12130), .A2(n12128), .ZN(n9807) );
  AND4_X1 U13182 ( .A1(n11373), .A2(n11372), .A3(n11371), .A4(n11370), .ZN(
        n9808) );
  AND2_X1 U13183 ( .A1(n11656), .A2(n11663), .ZN(n9809) );
  AND2_X1 U13184 ( .A1(n16637), .A2(n13602), .ZN(n9810) );
  AND2_X1 U13185 ( .A1(n10554), .A2(n10549), .ZN(n9811) );
  INV_X1 U13186 ( .A(n11118), .ZN(n10618) );
  AND3_X1 U13187 ( .A1(n9810), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16647), .ZN(n9812) );
  AND3_X1 U13188 ( .A1(n11123), .A2(n11127), .A3(n11122), .ZN(n11133) );
  AND2_X1 U13189 ( .A1(n16073), .A2(n16970), .ZN(n9813) );
  NAND2_X1 U13190 ( .A1(n10989), .A2(n10988), .ZN(n11062) );
  NOR2_X1 U13191 ( .A1(n19715), .A2(n12148), .ZN(n9814) );
  AND2_X1 U13192 ( .A1(n10932), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9815) );
  AND2_X1 U13193 ( .A1(n11148), .A2(n11133), .ZN(n9816) );
  OR2_X1 U13194 ( .A1(n14297), .A2(n13409), .ZN(n9817) );
  AND2_X1 U13195 ( .A1(n11343), .A2(n11435), .ZN(n9818) );
  NAND2_X1 U13196 ( .A1(n12232), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9819) );
  NAND3_X1 U13197 ( .A1(n10608), .A2(n13588), .A3(n10611), .ZN(n9820) );
  OR2_X1 U13198 ( .A1(n11103), .A2(n17017), .ZN(n9821) );
  INV_X1 U13199 ( .A(n18756), .ZN(n18777) );
  AND2_X1 U13200 ( .A1(n16629), .A2(n10210), .ZN(n9822) );
  INV_X1 U13201 ( .A(n13643), .ZN(n13644) );
  AND3_X1 U13202 ( .A1(n10313), .A2(n10316), .A3(n10311), .ZN(n9823) );
  OR3_X1 U13203 ( .A1(n16116), .A2(n11378), .A3(n16828), .ZN(n16553) );
  AND2_X1 U13204 ( .A1(n13463), .A2(n14618), .ZN(n9824) );
  NOR2_X1 U13205 ( .A1(n14807), .A2(n10810), .ZN(n11818) );
  AND2_X1 U13206 ( .A1(n11510), .A2(n11509), .ZN(n9825) );
  AND2_X1 U13207 ( .A1(n11622), .A2(n11635), .ZN(n9826) );
  OR2_X1 U13208 ( .A1(n13593), .A2(n11511), .ZN(n9827) );
  AND2_X1 U13209 ( .A1(n10917), .A2(n11529), .ZN(n9828) );
  AND2_X1 U13210 ( .A1(n17773), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n9829) );
  OR2_X1 U13211 ( .A1(n17058), .A2(n17059), .ZN(n9830) );
  AND2_X1 U13212 ( .A1(n9733), .A2(n10498), .ZN(n9831) );
  NOR2_X1 U13213 ( .A1(n14652), .A2(n19874), .ZN(n12215) );
  AND3_X1 U13214 ( .A1(n13988), .A2(n13987), .A3(n13986), .ZN(n9832) );
  AND2_X1 U13215 ( .A1(n10908), .A2(n15680), .ZN(n9833) );
  INV_X1 U13216 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21718) );
  OR2_X1 U13217 ( .A1(n10225), .A2(n13644), .ZN(n9834) );
  INV_X1 U13218 ( .A(n10546), .ZN(n10545) );
  NAND2_X1 U13219 ( .A1(n10547), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10546) );
  AND2_X1 U13220 ( .A1(n12490), .A2(n9763), .ZN(n9835) );
  NAND2_X1 U13221 ( .A1(n10378), .A2(n10142), .ZN(n11344) );
  INV_X1 U13222 ( .A(n10488), .ZN(n10487) );
  OAI21_X1 U13223 ( .B1(n14910), .B2(n13639), .A(n14911), .ZN(n10488) );
  NAND2_X1 U13224 ( .A1(n10595), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9836) );
  AND4_X1 U13225 ( .A1(n11194), .A2(n11193), .A3(n11192), .A4(n11191), .ZN(
        n9837) );
  INV_X1 U13226 ( .A(n13752), .ZN(n10499) );
  INV_X1 U13227 ( .A(n11345), .ZN(n11343) );
  AND2_X1 U13228 ( .A1(n11525), .A2(n11524), .ZN(n9838) );
  AND2_X1 U13229 ( .A1(n10547), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9839) );
  INV_X1 U13230 ( .A(n16487), .ZN(n10112) );
  OR2_X1 U13231 ( .A1(n16761), .A2(n16762), .ZN(n9840) );
  INV_X1 U13232 ( .A(n14054), .ZN(n10297) );
  NAND2_X1 U13233 ( .A1(n12490), .A2(n12489), .ZN(n15991) );
  NAND2_X1 U13234 ( .A1(n14018), .A2(n9730), .ZN(n9841) );
  OR2_X1 U13235 ( .A1(n11179), .A2(n11317), .ZN(n9842) );
  AND2_X1 U13236 ( .A1(n10558), .A2(n10557), .ZN(n9843) );
  AND3_X1 U13237 ( .A1(n11739), .A2(n11738), .A3(n11737), .ZN(n14283) );
  AND2_X1 U13238 ( .A1(n11074), .A2(n11385), .ZN(n11617) );
  INV_X1 U13239 ( .A(n10923), .ZN(n10922) );
  OAI21_X1 U13240 ( .B1(n16540), .B2(n10924), .A(n13546), .ZN(n10923) );
  NAND2_X1 U13241 ( .A1(n15647), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9844) );
  INV_X1 U13242 ( .A(n10106), .ZN(n10105) );
  NAND2_X1 U13243 ( .A1(n10504), .A2(n9723), .ZN(n10106) );
  INV_X1 U13244 ( .A(n10869), .ZN(n10249) );
  AND2_X1 U13245 ( .A1(n15470), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9845) );
  NAND2_X1 U13246 ( .A1(n13776), .A2(n10788), .ZN(n9846) );
  AND2_X1 U13247 ( .A1(n15462), .A2(n10909), .ZN(n9847) );
  AND2_X1 U13248 ( .A1(n10747), .A2(n10745), .ZN(n9848) );
  OAI211_X1 U13249 ( .C1(n10192), .C2(n10134), .A(n10503), .B(n10131), .ZN(
        n10135) );
  AND2_X1 U13250 ( .A1(n10621), .A2(n10485), .ZN(n9849) );
  INV_X1 U13251 ( .A(n10823), .ZN(n10822) );
  NOR2_X1 U13252 ( .A1(n14257), .A2(n14283), .ZN(n10823) );
  AND2_X1 U13253 ( .A1(n14653), .A2(n10857), .ZN(n9850) );
  AND2_X1 U13254 ( .A1(n9737), .A2(n16553), .ZN(n9851) );
  AND2_X1 U13255 ( .A1(n10221), .A2(n9834), .ZN(n9852) );
  NAND2_X1 U13256 ( .A1(n16491), .A2(n16719), .ZN(n10710) );
  AND2_X1 U13257 ( .A1(n15987), .A2(n13616), .ZN(n13781) );
  NAND2_X1 U13258 ( .A1(n12078), .A2(n12079), .ZN(n18762) );
  OR2_X1 U13259 ( .A1(n13769), .A2(n13768), .ZN(n9853) );
  OR2_X1 U13260 ( .A1(n12038), .A2(n12039), .ZN(n10665) );
  INV_X1 U13261 ( .A(n11185), .ZN(n10041) );
  OR2_X1 U13262 ( .A1(n16274), .A2(n17185), .ZN(n9854) );
  AOI21_X1 U13263 ( .B1(n15564), .B2(n13891), .A(n13886), .ZN(n15554) );
  OR2_X1 U13264 ( .A1(n12138), .A2(n12137), .ZN(n9855) );
  AND2_X2 U13265 ( .A1(n12319), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11367) );
  AND2_X1 U13266 ( .A1(n13657), .A2(n13656), .ZN(n9856) );
  AND3_X1 U13267 ( .A1(n10406), .A2(n10405), .A3(n10404), .ZN(n9857) );
  NAND2_X1 U13268 ( .A1(n10792), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10791) );
  INV_X1 U13269 ( .A(n10791), .ZN(n10790) );
  NAND2_X1 U13270 ( .A1(n13781), .A2(n10817), .ZN(n13648) );
  NAND2_X1 U13271 ( .A1(n13683), .A2(n9731), .ZN(n10730) );
  OR2_X1 U13272 ( .A1(n17222), .A2(n18620), .ZN(n9858) );
  NAND2_X1 U13273 ( .A1(n11518), .A2(n10902), .ZN(n9859) );
  AND2_X1 U13274 ( .A1(n9732), .A2(n9827), .ZN(n9860) );
  AND2_X1 U13275 ( .A1(n17270), .A2(n18411), .ZN(n9861) );
  OR2_X1 U13276 ( .A1(n13603), .A2(n10475), .ZN(n9862) );
  INV_X1 U13277 ( .A(n13852), .ZN(n10715) );
  AND2_X1 U13278 ( .A1(n12843), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9863) );
  NAND2_X1 U13279 ( .A1(n13380), .A2(n13398), .ZN(n9864) );
  AND2_X1 U13280 ( .A1(n11574), .A2(n11578), .ZN(n9865) );
  AND2_X1 U13281 ( .A1(n13761), .A2(n10500), .ZN(n9866) );
  AND2_X1 U13282 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U13283 ( .A1(n20264), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n9868) );
  INV_X1 U13284 ( .A(n13376), .ZN(n10560) );
  INV_X1 U13285 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18565) );
  INV_X1 U13286 ( .A(n13604), .ZN(n10595) );
  NAND2_X1 U13287 ( .A1(n10270), .A2(n13602), .ZN(n13604) );
  INV_X1 U13288 ( .A(n13879), .ZN(n10714) );
  NOR2_X2 U13289 ( .A1(n19891), .A2(n11602), .ZN(n9869) );
  INV_X1 U13290 ( .A(n19039), .ZN(n19054) );
  NAND2_X1 U13291 ( .A1(n15075), .A2(n15097), .ZN(n9870) );
  NAND2_X1 U13292 ( .A1(n15251), .A2(n10832), .ZN(n15199) );
  NOR2_X1 U13293 ( .A1(n14807), .A2(n10813), .ZN(n16076) );
  AND2_X1 U13294 ( .A1(n20638), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n9871) );
  OR2_X1 U13295 ( .A1(n14254), .A2(n14257), .ZN(n14255) );
  AND2_X1 U13296 ( .A1(n20606), .A2(n10677), .ZN(n9872) );
  NAND2_X1 U13297 ( .A1(n10827), .A2(n11779), .ZN(n14470) );
  INV_X1 U13298 ( .A(n16518), .ZN(n10604) );
  AND2_X1 U13299 ( .A1(n16069), .A2(n11527), .ZN(n11528) );
  INV_X1 U13300 ( .A(n11205), .ZN(n10269) );
  NOR2_X1 U13301 ( .A1(n13706), .A2(n10734), .ZN(n9873) );
  NAND3_X1 U13302 ( .A1(n11457), .A2(n10895), .A3(n10891), .ZN(n9874) );
  OR2_X1 U13303 ( .A1(n10776), .A2(n9870), .ZN(n9875) );
  NOR2_X1 U13304 ( .A1(n14655), .A2(n14656), .ZN(n14654) );
  NAND2_X1 U13305 ( .A1(n13880), .A2(n15850), .ZN(n15601) );
  NAND2_X1 U13306 ( .A1(n14653), .A2(n12249), .ZN(n14804) );
  NAND2_X1 U13307 ( .A1(n10836), .A2(n10837), .ZN(n15131) );
  OR2_X1 U13308 ( .A1(n14655), .A2(n10796), .ZN(n14734) );
  INV_X1 U13309 ( .A(n16595), .ZN(n10610) );
  INV_X1 U13310 ( .A(n16554), .ZN(n10580) );
  INV_X1 U13311 ( .A(n19826), .ZN(n16242) );
  NAND2_X1 U13312 ( .A1(n14644), .A2(n14643), .ZN(n14642) );
  INV_X1 U13313 ( .A(n18573), .ZN(n18673) );
  INV_X1 U13314 ( .A(n16970), .ZN(n17185) );
  AND2_X1 U13315 ( .A1(n11865), .A2(n11864), .ZN(n16970) );
  AND3_X1 U13316 ( .A1(n16047), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n13641), .ZN(n9876) );
  AND2_X1 U13317 ( .A1(n10845), .A2(n10844), .ZN(n9877) );
  NAND2_X1 U13318 ( .A1(n14379), .A2(n12909), .ZN(n14464) );
  NOR2_X1 U13319 ( .A1(n14747), .A2(n14775), .ZN(n9878) );
  OR2_X1 U13320 ( .A1(n17151), .A2(n17152), .ZN(n14617) );
  AND2_X1 U13321 ( .A1(n16574), .A2(n16573), .ZN(n9879) );
  INV_X1 U13322 ( .A(n16567), .ZN(n10584) );
  INV_X1 U13323 ( .A(n13775), .ZN(n10607) );
  INV_X1 U13324 ( .A(n13880), .ZN(n15621) );
  INV_X1 U13325 ( .A(n11488), .ZN(n10904) );
  INV_X1 U13326 ( .A(n11496), .ZN(n10507) );
  NOR2_X1 U13327 ( .A1(n13706), .A2(n10731), .ZN(n13710) );
  AND2_X1 U13328 ( .A1(n14173), .A2(n14297), .ZN(n13871) );
  INV_X1 U13329 ( .A(n16528), .ZN(n10519) );
  NAND2_X1 U13330 ( .A1(n12695), .A2(n12694), .ZN(n14505) );
  INV_X1 U13331 ( .A(n10948), .ZN(n10783) );
  INV_X1 U13332 ( .A(n17142), .ZN(n18291) );
  AOI21_X1 U13333 ( .B1(n17140), .B2(n17139), .A(n19573), .ZN(n17142) );
  NAND2_X1 U13334 ( .A1(n11446), .A2(n11445), .ZN(n11448) );
  AND2_X1 U13335 ( .A1(n15621), .A2(n15697), .ZN(n9880) );
  NAND2_X1 U13336 ( .A1(n14457), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14230) );
  AND2_X1 U13337 ( .A1(n18055), .A2(n10698), .ZN(n9881) );
  AND2_X1 U13338 ( .A1(n9759), .A2(n13558), .ZN(n9882) );
  OR2_X1 U13339 ( .A1(n18673), .A2(n18418), .ZN(n9883) );
  OR2_X1 U13340 ( .A1(n19771), .A2(n11507), .ZN(n13554) );
  NAND2_X1 U13341 ( .A1(n16568), .A2(n16567), .ZN(n9884) );
  NAND2_X1 U13342 ( .A1(n13689), .A2(n10721), .ZN(n10724) );
  AND2_X1 U13343 ( .A1(n19879), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n9885) );
  INV_X1 U13344 ( .A(n16214), .ZN(n10129) );
  INV_X1 U13345 ( .A(n14198), .ZN(n10775) );
  AND2_X1 U13346 ( .A1(n18573), .A2(n17071), .ZN(n17072) );
  INV_X1 U13347 ( .A(n10055), .ZN(n15574) );
  NAND2_X1 U13348 ( .A1(n13885), .A2(n15585), .ZN(n10055) );
  INV_X1 U13349 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15257) );
  NAND2_X1 U13350 ( .A1(n11865), .A2(n20545), .ZN(n17193) );
  INV_X1 U13351 ( .A(n9762), .ZN(n10651) );
  NAND2_X1 U13352 ( .A1(n13049), .A2(n10436), .ZN(n10439) );
  INV_X1 U13353 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n14457) );
  INV_X1 U13354 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12510) );
  OR2_X1 U13355 ( .A1(n18673), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9886) );
  AND2_X1 U13356 ( .A1(n9766), .A2(n15964), .ZN(n9887) );
  OR2_X1 U13357 ( .A1(n19730), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9888) );
  NOR2_X1 U13358 ( .A1(n13950), .A2(n13947), .ZN(n9889) );
  AND2_X1 U13359 ( .A1(n10316), .A2(n16944), .ZN(n9890) );
  AND2_X1 U13360 ( .A1(n12281), .A2(n16326), .ZN(n9891) );
  AND2_X1 U13361 ( .A1(n10802), .A2(n11878), .ZN(n9892) );
  AND2_X1 U13362 ( .A1(n10618), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n9893) );
  INV_X1 U13363 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13665) );
  INV_X1 U13364 ( .A(n11281), .ZN(n10171) );
  INV_X1 U13365 ( .A(n11931), .ZN(n17788) );
  INV_X1 U13366 ( .A(n17788), .ZN(n18089) );
  OR2_X2 U13367 ( .A1(n11923), .A2(n11921), .ZN(n18058) );
  INV_X1 U13368 ( .A(n12044), .ZN(n17817) );
  INV_X1 U13369 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10690) );
  INV_X1 U13370 ( .A(n19736), .ZN(n10538) );
  NOR2_X2 U13371 ( .A1(n19105), .A2(n18147), .ZN(n18148) );
  INV_X2 U13372 ( .A(n18148), .ZN(n18143) );
  NAND2_X1 U13373 ( .A1(n17386), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18451) );
  NOR2_X1 U13374 ( .A1(n14380), .A2(n14381), .ZN(n9894) );
  INV_X1 U13375 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10437) );
  INV_X1 U13376 ( .A(n10459), .ZN(n10458) );
  NOR2_X1 U13377 ( .A1(n12456), .A2(n12475), .ZN(n10459) );
  AND2_X1 U13378 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n9895)
         );
  AND2_X1 U13379 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n9896) );
  AND2_X1 U13380 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n9897)
         );
  AND2_X1 U13381 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n9898)
         );
  AND2_X1 U13382 ( .A1(n12292), .A2(n10860), .ZN(n9899) );
  INV_X1 U13383 ( .A(n15102), .ZN(n10777) );
  INV_X1 U13384 ( .A(n16623), .ZN(n10302) );
  NOR2_X1 U13385 ( .A1(n18900), .A2(n18889), .ZN(n17077) );
  INV_X1 U13386 ( .A(n11454), .ZN(n10893) );
  AND2_X1 U13387 ( .A1(n13099), .A2(n13098), .ZN(n9900) );
  NOR2_X1 U13388 ( .A1(n12158), .A2(n12183), .ZN(n17261) );
  AND2_X1 U13389 ( .A1(n13068), .A2(n13067), .ZN(n9901) );
  AND2_X1 U13390 ( .A1(n9899), .A2(n16306), .ZN(n9902) );
  AND2_X1 U13391 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n9903) );
  AND2_X1 U13392 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9904) );
  AND2_X1 U13393 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9905) );
  AND2_X1 U13394 ( .A1(n12630), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n9906) );
  INV_X1 U13395 ( .A(n9906), .ZN(n10387) );
  NAND2_X1 U13396 ( .A1(n10521), .A2(n10522), .ZN(n10525) );
  INV_X1 U13397 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15997) );
  AND2_X1 U13398 ( .A1(n10700), .A2(n10699), .ZN(n9907) );
  INV_X1 U13399 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9919) );
  INV_X1 U13400 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10759) );
  INV_X1 U13401 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14680) );
  NOR2_X1 U13402 ( .A1(n18619), .A2(n18905), .ZN(n18903) );
  INV_X1 U13403 ( .A(n18903), .ZN(n10766) );
  OR2_X1 U13404 ( .A1(n16719), .A2(n10927), .ZN(n9908) );
  INV_X1 U13405 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10438) );
  INV_X1 U13406 ( .A(n19820), .ZN(n19782) );
  OR2_X1 U13407 ( .A1(n16719), .A2(n13787), .ZN(n9909) );
  INV_X1 U13408 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10444) );
  INV_X1 U13409 ( .A(n10510), .ZN(n17015) );
  OR2_X1 U13410 ( .A1(n17012), .A2(n17013), .ZN(n10510) );
  INV_X1 U13411 ( .A(n10702), .ZN(n10701) );
  NAND2_X1 U13412 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .ZN(n10702) );
  INV_X1 U13413 ( .A(n13627), .ZN(n10553) );
  INV_X1 U13414 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10042) );
  AND2_X1 U13415 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n9910) );
  AND2_X1 U13416 ( .A1(n10939), .A2(n10322), .ZN(n9911) );
  INV_X1 U13417 ( .A(n10475), .ZN(n10474) );
  OR2_X1 U13418 ( .A1(n15017), .A2(n15452), .ZN(n9912) );
  INV_X1 U13419 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10555) );
  INV_X1 U13420 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n10683) );
  INV_X1 U13421 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U13422 ( .A1(n13972), .A2(n21273), .ZN(n15573) );
  AND2_X1 U13423 ( .A1(n10738), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9913) );
  INV_X1 U13424 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10746) );
  AND2_X1 U13425 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9914) );
  INV_X1 U13426 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10723) );
  INV_X1 U13427 ( .A(n10739), .ZN(n10738) );
  NAND2_X1 U13428 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10739) );
  INV_X1 U13429 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20393) );
  NAND2_X1 U13430 ( .A1(n19832), .A2(n14813), .ZN(n16354) );
  INV_X2 U13431 ( .A(n19832), .ZN(n16351) );
  OR2_X1 U13432 ( .A1(n19832), .A2(n11423), .ZN(n10010) );
  NAND2_X1 U13433 ( .A1(n19832), .A2(n12210), .ZN(n10009) );
  OAI21_X1 U13434 ( .B1(n16853), .B2(n16680), .A(n10284), .ZN(n10283) );
  NOR3_X2 U13435 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19576), .A3(
        n19219), .ZN(n19214) );
  NOR3_X2 U13436 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19576), .A3(
        n19196), .ZN(n19125) );
  NOR3_X2 U13437 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19576), .A3(
        n19289), .ZN(n19262) );
  AOI22_X2 U13438 ( .A1(DATAI_21_), .A2(n14553), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20829), .ZN(n21310) );
  NOR2_X2 U13439 ( .A1(n15573), .A2(n15405), .ZN(n20829) );
  NOR3_X2 U13440 ( .A1(n19576), .A2(n19553), .A3(n19196), .ZN(n19168) );
  OAI33_X1 U13441 ( .A1(n19418), .A2(n19364), .A3(n19221), .B1(n19220), .B2(
        n19130), .B3(n19073), .ZN(n9915) );
  OR2_X1 U13442 ( .A1(n19220), .A2(n19414), .ZN(n19221) );
  NAND2_X1 U13443 ( .A1(n17380), .A2(n19074), .ZN(n19220) );
  INV_X1 U13444 ( .A(n17182), .ZN(n16944) );
  NAND2_X2 U13445 ( .A1(n10086), .A2(n10084), .ZN(n10143) );
  NAND3_X1 U13446 ( .A1(n10287), .A2(n10291), .A3(n9916), .ZN(n10292) );
  NAND2_X1 U13447 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  NAND2_X1 U13448 ( .A1(n10190), .A2(n11195), .ZN(n10115) );
  INV_X2 U13449 ( .A(n11077), .ZN(n11628) );
  XNOR2_X2 U13450 ( .A(n12910), .B(n12798), .ZN(n15911) );
  NAND2_X2 U13451 ( .A1(n10425), .A2(n9921), .ZN(n18429) );
  NAND2_X1 U13452 ( .A1(n10926), .A2(n14927), .ZN(n9924) );
  NAND3_X1 U13453 ( .A1(n12043), .A2(n12045), .A3(n9926), .ZN(n9925) );
  NAND3_X1 U13454 ( .A1(n12041), .A2(n9930), .A3(n9929), .ZN(n9928) );
  AND2_X1 U13455 ( .A1(n12070), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9931) );
  NOR2_X1 U13456 ( .A1(n17817), .A2(n21495), .ZN(n9932) );
  OAI21_X1 U13457 ( .B1(n9933), .B2(n9935), .A(n12097), .ZN(n9934) );
  NAND3_X1 U13458 ( .A1(n12098), .A2(n18700), .A3(n12094), .ZN(n9936) );
  NAND2_X1 U13459 ( .A1(n9937), .A2(n12098), .ZN(n12099) );
  NAND2_X1 U13460 ( .A1(n9938), .A2(n9941), .ZN(n10227) );
  NAND2_X1 U13461 ( .A1(n9942), .A2(n18735), .ZN(n18734) );
  OAI211_X1 U13462 ( .C1(n9940), .C2(n9942), .A(n18723), .B(n9939), .ZN(n18721) );
  NAND2_X1 U13463 ( .A1(n9941), .A2(n19026), .ZN(n9939) );
  INV_X1 U13464 ( .A(n18735), .ZN(n9941) );
  NAND3_X1 U13465 ( .A1(n17271), .A2(n9944), .A3(n9861), .ZN(P3_U2834) );
  NOR2_X2 U13466 ( .A1(n10232), .A2(n18557), .ZN(n17069) );
  AND2_X2 U13467 ( .A1(n9947), .A2(n18476), .ZN(n18557) );
  INV_X2 U13468 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12163) );
  NAND2_X2 U13469 ( .A1(n15544), .A2(n15543), .ZN(n15507) );
  AND2_X2 U13470 ( .A1(n10625), .A2(n9867), .ZN(n18056) );
  NAND3_X1 U13471 ( .A1(n17769), .A2(n17768), .A3(n9888), .ZN(P3_U2671) );
  XNOR2_X2 U13472 ( .A(n9948), .B(n11139), .ZN(n11173) );
  NAND2_X1 U13473 ( .A1(n9952), .A2(n10665), .ZN(n9955) );
  NAND3_X1 U13474 ( .A1(n18762), .A2(n12118), .A3(n18287), .ZN(n9954) );
  NAND4_X1 U13475 ( .A1(n9956), .A2(n9960), .A3(n12074), .A4(n12076), .ZN(
        n9959) );
  NOR2_X1 U13476 ( .A1(n9829), .A2(n9957), .ZN(n9956) );
  INV_X2 U13477 ( .A(n11969), .ZN(n18073) );
  INV_X1 U13478 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n9962) );
  AND2_X2 U13479 ( .A1(n10657), .A2(n9855), .ZN(n12141) );
  OR2_X2 U13480 ( .A1(n18706), .A2(n18997), .ZN(n10657) );
  NOR2_X1 U13481 ( .A1(n12143), .A2(n10666), .ZN(n18682) );
  NAND3_X1 U13482 ( .A1(n11270), .A2(n11271), .A3(n11684), .ZN(n9964) );
  NAND2_X2 U13483 ( .A1(n10008), .A2(n10077), .ZN(n11271) );
  NOR2_X2 U13484 ( .A1(n18416), .A2(n17131), .ZN(n17236) );
  NAND2_X1 U13485 ( .A1(n9986), .A2(n9966), .ZN(P2_U3023) );
  OAI211_X1 U13486 ( .C1(n10545), .C2(n9839), .A(n9967), .B(n16993), .ZN(n9966) );
  NAND3_X1 U13487 ( .A1(n9968), .A2(n10139), .A3(n11867), .ZN(P2_U3026) );
  OAI21_X1 U13488 ( .B1(n10586), .B2(n10587), .A(n9736), .ZN(P3_U2799) );
  NAND2_X1 U13489 ( .A1(n10585), .A2(n18756), .ZN(n9969) );
  NAND4_X1 U13490 ( .A1(n9798), .A2(n10760), .A3(n18688), .A4(n18900), .ZN(
        n9976) );
  NAND2_X1 U13491 ( .A1(n12202), .A2(n10940), .ZN(n9977) );
  NAND2_X1 U13492 ( .A1(n18476), .A2(n9977), .ZN(n18468) );
  NAND3_X1 U13493 ( .A1(n10481), .A2(n10479), .A3(n10478), .ZN(n13988) );
  NAND2_X1 U13494 ( .A1(n14913), .A2(n10482), .ZN(n10478) );
  AND2_X1 U13495 ( .A1(n9752), .A2(n11173), .ZN(n10037) );
  NAND3_X1 U13496 ( .A1(n9991), .A2(n9990), .A3(n9989), .ZN(n9988) );
  INV_X1 U13497 ( .A(n10020), .ZN(n9989) );
  NAND2_X1 U13498 ( .A1(n10066), .A2(n11281), .ZN(n9990) );
  NAND2_X1 U13499 ( .A1(n10019), .A2(n10042), .ZN(n9991) );
  NAND2_X2 U13500 ( .A1(n11153), .A2(n11155), .ZN(n11140) );
  NAND2_X2 U13501 ( .A1(n11143), .A2(n11142), .ZN(n11155) );
  XNOR2_X2 U13502 ( .A(n10863), .B(n10862), .ZN(n11153) );
  NAND2_X1 U13503 ( .A1(n16594), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10271) );
  NAND3_X1 U13504 ( .A1(n10144), .A2(n9997), .A3(n9994), .ZN(n10200) );
  NAND2_X1 U13505 ( .A1(n11170), .A2(n9683), .ZN(n9999) );
  NAND2_X1 U13506 ( .A1(n11170), .A2(n9754), .ZN(n10003) );
  INV_X1 U13507 ( .A(n9999), .ZN(n20163) );
  OAI22_X1 U13508 ( .A1(n9999), .A2(n9998), .B1(n11205), .B2(n11296), .ZN(
        n11297) );
  NAND2_X1 U13509 ( .A1(n11170), .A2(n9755), .ZN(n10002) );
  NAND2_X1 U13510 ( .A1(n20163), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10123) );
  NAND2_X1 U13511 ( .A1(n20163), .A2(n20300), .ZN(n10001) );
  NAND3_X1 U13512 ( .A1(n10125), .A2(n10872), .A3(n10870), .ZN(n10004) );
  NAND4_X1 U13513 ( .A1(n10125), .A2(n10603), .A3(n10872), .A4(n10870), .ZN(
        n10006) );
  NAND3_X1 U13514 ( .A1(n10077), .A2(n11282), .A3(n10008), .ZN(n10022) );
  OAI21_X1 U13515 ( .B1(n16774), .B2(n16712), .A(n16530), .ZN(P2_U2992) );
  OAI21_X1 U13516 ( .B1(n16774), .B2(n17193), .A(n16773), .ZN(P2_U3024) );
  NAND2_X1 U13517 ( .A1(n9691), .A2(n11062), .ZN(n10013) );
  NAND2_X1 U13518 ( .A1(n10017), .A2(n10021), .ZN(n16685) );
  INV_X1 U13519 ( .A(n10172), .ZN(n10018) );
  INV_X1 U13520 ( .A(n10019), .ZN(n10021) );
  NAND2_X1 U13521 ( .A1(n10382), .A2(n10022), .ZN(n10019) );
  NAND2_X1 U13522 ( .A1(n10023), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11123) );
  OAI22_X1 U13523 ( .A1(n10023), .A2(n11117), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12503), .ZN(n10736) );
  AOI21_X1 U13524 ( .B1(n10023), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n9893), .ZN(n11138) );
  NAND2_X1 U13525 ( .A1(n10025), .A2(n10024), .ZN(n14550) );
  INV_X1 U13526 ( .A(n14549), .ZN(n10024) );
  NAND2_X1 U13527 ( .A1(n16281), .A2(n10026), .ZN(n10029) );
  INV_X1 U13528 ( .A(n12424), .ZN(n10027) );
  INV_X1 U13529 ( .A(n12425), .ZN(n10028) );
  XNOR2_X2 U13530 ( .A(n16305), .B(n12347), .ZN(n16299) );
  AND2_X2 U13531 ( .A1(n14653), .A2(n10247), .ZN(n12293) );
  NAND2_X1 U13532 ( .A1(n10126), .A2(n11147), .ZN(n11134) );
  NAND2_X2 U13533 ( .A1(n9793), .A2(n10033), .ZN(n10863) );
  NAND2_X1 U13534 ( .A1(n11104), .A2(n11115), .ZN(n10034) );
  NAND2_X1 U13535 ( .A1(n10037), .A2(n9703), .ZN(n11283) );
  NAND2_X1 U13536 ( .A1(n10288), .A2(n10037), .ZN(n10287) );
  INV_X1 U13537 ( .A(n10043), .ZN(n10060) );
  NAND2_X1 U13538 ( .A1(n10043), .A2(n20231), .ZN(n20237) );
  OAI22_X1 U13539 ( .A1(n10043), .A2(n11204), .B1(n19997), .B2(n11203), .ZN(
        n11209) );
  OAI22_X1 U13540 ( .A1(n20391), .A2(n11151), .B1(n10043), .B2(n11152), .ZN(
        n11163) );
  NAND3_X1 U13541 ( .A1(n11146), .A2(n10126), .A3(n11147), .ZN(n10045) );
  NAND2_X1 U13542 ( .A1(n10047), .A2(n11148), .ZN(n10046) );
  AND2_X2 U13543 ( .A1(n10049), .A2(n12515), .ZN(n12732) );
  AND2_X2 U13544 ( .A1(n10049), .A2(n12517), .ZN(n12733) );
  AND2_X2 U13545 ( .A1(n14489), .A2(n10049), .ZN(n12755) );
  AND2_X2 U13546 ( .A1(n14486), .A2(n10049), .ZN(n12739) );
  NAND2_X2 U13547 ( .A1(n15455), .A2(n15462), .ZN(n15456) );
  NAND2_X2 U13548 ( .A1(n9845), .A2(n13899), .ZN(n15455) );
  NAND3_X1 U13549 ( .A1(n16676), .A2(n10064), .A3(n16673), .ZN(n10063) );
  CLKBUF_X1 U13550 ( .A(n10066), .Z(n10065) );
  NAND2_X1 U13551 ( .A1(n10066), .A2(n16237), .ZN(n10087) );
  NOR2_X1 U13552 ( .A1(n11185), .A2(n10067), .ZN(n10088) );
  NAND3_X1 U13553 ( .A1(n10136), .A2(n10137), .A3(n10068), .ZN(n10266) );
  NAND2_X1 U13554 ( .A1(n10041), .A2(n10069), .ZN(n10068) );
  OAI21_X1 U13555 ( .B1(n20122), .B2(n20393), .A(n20300), .ZN(n10071) );
  NAND2_X1 U13556 ( .A1(n20264), .A2(n20300), .ZN(n10073) );
  NAND4_X1 U13557 ( .A1(n10117), .A2(n10265), .A3(n10118), .A4(n11329), .ZN(
        n10074) );
  NAND2_X1 U13558 ( .A1(n11342), .A2(n10075), .ZN(n10293) );
  NAND2_X1 U13559 ( .A1(n10085), .A2(n10075), .ZN(n10084) );
  NAND2_X2 U13560 ( .A1(n11344), .A2(n16646), .ZN(n10076) );
  NAND2_X1 U13561 ( .A1(n10076), .A2(n13600), .ZN(n10596) );
  NAND2_X1 U13562 ( .A1(n10076), .A2(n9680), .ZN(n10737) );
  NAND3_X1 U13563 ( .A1(n10076), .A2(n9680), .A3(n10474), .ZN(n10173) );
  NAND4_X1 U13564 ( .A1(n10079), .A2(n10268), .A3(n10078), .A4(n10081), .ZN(
        n10080) );
  AOI21_X1 U13565 ( .B1(n9715), .B2(n10601), .A(n9719), .ZN(n10079) );
  NAND2_X1 U13566 ( .A1(n10080), .A2(n14347), .ZN(n10190) );
  NAND2_X1 U13567 ( .A1(n9758), .A2(n11182), .ZN(n10081) );
  AOI21_X2 U13568 ( .B1(n16543), .B2(n16533), .A(n10083), .ZN(n16799) );
  NAND2_X2 U13569 ( .A1(n10176), .A2(n10179), .ZN(n16802) );
  NAND3_X1 U13570 ( .A1(n10093), .A2(n9866), .A3(n10089), .ZN(P2_U3015) );
  NAND2_X1 U13571 ( .A1(n10481), .A2(n10090), .ZN(n10089) );
  NOR2_X1 U13572 ( .A1(n10092), .A2(n10091), .ZN(n10090) );
  NAND3_X1 U13573 ( .A1(n10493), .A2(n10494), .A3(n10492), .ZN(n10093) );
  INV_X1 U13574 ( .A(n13745), .ZN(n10094) );
  AND2_X1 U13575 ( .A1(n10608), .A2(n13588), .ZN(n10096) );
  NAND2_X1 U13576 ( .A1(n9799), .A2(n10097), .ZN(n10099) );
  NAND2_X1 U13577 ( .A1(n10100), .A2(n10649), .ZN(n16621) );
  AOI21_X1 U13578 ( .B1(n11909), .B2(n16531), .A(n13549), .ZN(n11912) );
  NAND3_X1 U13579 ( .A1(n10109), .A2(n10111), .A3(n10108), .ZN(n16728) );
  NAND4_X1 U13580 ( .A1(n10109), .A2(n10111), .A3(n10108), .A4(n11531), .ZN(
        n10138) );
  INV_X1 U13581 ( .A(n16485), .ZN(n10110) );
  NAND2_X1 U13582 ( .A1(n10116), .A2(n11531), .ZN(n13803) );
  NAND2_X1 U13583 ( .A1(n10116), .A2(n16944), .ZN(n13796) );
  OAI211_X1 U13584 ( .C1(n14936), .C2(n17182), .A(n10799), .B(n10800), .ZN(
        P2_U3017) );
  NAND3_X1 U13585 ( .A1(n10275), .A2(n10123), .A3(n10277), .ZN(n10120) );
  AOI21_X1 U13586 ( .B1(n10125), .B2(n10872), .A(n13561), .ZN(n16525) );
  NAND2_X1 U13587 ( .A1(n10128), .A2(n10686), .ZN(n10184) );
  OAI21_X1 U13588 ( .B1(n10128), .B2(n10507), .A(n10505), .ZN(n16566) );
  OAI21_X1 U13589 ( .B1(n10128), .B2(n10507), .A(n10185), .ZN(n10188) );
  NAND2_X1 U13590 ( .A1(n16494), .A2(n10138), .ZN(P2_U2987) );
  NAND2_X1 U13591 ( .A1(n10143), .A2(n10140), .ZN(n10179) );
  NAND2_X1 U13592 ( .A1(n10141), .A2(n16697), .ZN(n10234) );
  NAND2_X1 U13593 ( .A1(n10141), .A2(n16993), .ZN(n10315) );
  INV_X1 U13594 ( .A(n10143), .ZN(n10381) );
  NAND2_X1 U13595 ( .A1(n10143), .A2(n13600), .ZN(n10594) );
  OAI21_X1 U13596 ( .B1(n16517), .B2(n10607), .A(n9756), .ZN(n10147) );
  NAND3_X1 U13597 ( .A1(n9843), .A2(n13381), .A3(n10148), .ZN(n13387) );
  OAI211_X1 U13598 ( .C1(n13382), .C2(n13359), .A(n10149), .B(n10559), .ZN(
        n10148) );
  AND2_X1 U13599 ( .A1(n13358), .A2(n13357), .ZN(n10149) );
  NAND2_X1 U13600 ( .A1(n10157), .A2(n11378), .ZN(n10165) );
  NAND2_X1 U13601 ( .A1(n10157), .A2(n16711), .ZN(n10169) );
  XNOR2_X1 U13602 ( .A(n10157), .B(n16711), .ZN(n16983) );
  NAND3_X1 U13604 ( .A1(n10163), .A2(n10207), .A3(n10206), .ZN(P2_U2991) );
  NAND2_X1 U13605 ( .A1(n10169), .A2(n11281), .ZN(n16687) );
  OR2_X1 U13606 ( .A1(n16711), .A2(n10171), .ZN(n10170) );
  NAND2_X1 U13607 ( .A1(n11271), .A2(n11684), .ZN(n10172) );
  NAND3_X1 U13608 ( .A1(n11596), .A2(n11597), .A3(n11595), .ZN(P2_U2994) );
  AND2_X1 U13609 ( .A1(n10189), .A2(n9762), .ZN(n11483) );
  NAND2_X1 U13610 ( .A1(n10323), .A2(n10196), .ZN(n16894) );
  XNOR2_X2 U13611 ( .A(n10200), .B(n11453), .ZN(n16661) );
  NAND4_X1 U13612 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n10201) );
  OAI22_X1 U13613 ( .A1(n19965), .A2(n11287), .B1(n11286), .B2(n20087), .ZN(
        n10202) );
  NAND3_X1 U13614 ( .A1(n10335), .A2(n10430), .A3(n10337), .ZN(n10203) );
  NAND2_X1 U13615 ( .A1(n10205), .A2(n10337), .ZN(n10204) );
  NAND3_X1 U13616 ( .A1(n10267), .A2(n16491), .A3(n16697), .ZN(n13800) );
  NAND3_X1 U13617 ( .A1(n10267), .A2(n16491), .A3(n16993), .ZN(n13793) );
  NAND2_X1 U13618 ( .A1(n10787), .A2(n11314), .ZN(n11315) );
  NAND3_X1 U13619 ( .A1(n10476), .A2(n10213), .A3(n10212), .ZN(P2_U2999) );
  OR2_X1 U13620 ( .A1(n16834), .A2(n16712), .ZN(n10212) );
  NAND3_X1 U13621 ( .A1(n10864), .A2(n10215), .A3(n9757), .ZN(n10214) );
  INV_X1 U13622 ( .A(n10216), .ZN(n11175) );
  OAI211_X1 U13623 ( .C1(n20024), .C2(n10274), .A(n9750), .B(n10217), .ZN(
        n10216) );
  NAND2_X1 U13624 ( .A1(n13664), .A2(n11531), .ZN(n10375) );
  NAND2_X2 U13625 ( .A1(n10416), .A2(n10415), .ZN(n12118) );
  INV_X2 U13626 ( .A(n18016), .ZN(n18076) );
  OR2_X2 U13627 ( .A1(n17069), .A2(n18673), .ZN(n10747) );
  OAI211_X1 U13628 ( .C1(n10234), .C2(n10486), .A(n10233), .B(n11900), .ZN(
        P2_U2993) );
  NAND2_X1 U13629 ( .A1(n9823), .A2(n11531), .ZN(n10233) );
  NAND2_X2 U13630 ( .A1(n11082), .A2(n19869), .ZN(n11096) );
  NAND2_X1 U13631 ( .A1(n10239), .A2(n16506), .ZN(P2_U2989) );
  NOR2_X1 U13632 ( .A1(n16497), .A2(n10790), .ZN(n10242) );
  INV_X1 U13633 ( .A(n12403), .ZN(n10246) );
  NOR2_X1 U13634 ( .A1(n16294), .A2(n12387), .ZN(n12403) );
  NAND3_X1 U13635 ( .A1(n9783), .A2(n10461), .A3(n10847), .ZN(n16373) );
  NAND2_X1 U13636 ( .A1(n9850), .A2(n16326), .ZN(n16323) );
  NAND3_X1 U13638 ( .A1(n10653), .A2(n10652), .A3(n13591), .ZN(n10252) );
  NAND3_X1 U13639 ( .A1(n9837), .A2(n10256), .A3(n11188), .ZN(n11676) );
  NAND4_X1 U13640 ( .A1(n10261), .A2(n10260), .A3(n10259), .A4(n10258), .ZN(
        n10257) );
  AND2_X2 U13641 ( .A1(n14018), .A2(n9860), .ZN(n11518) );
  NAND2_X2 U13642 ( .A1(n11489), .A2(n13539), .ZN(n14018) );
  AND2_X2 U13643 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11186) );
  INV_X2 U13644 ( .A(n12315), .ZN(n11044) );
  NAND2_X1 U13645 ( .A1(n13553), .A2(n10344), .ZN(n10264) );
  OR2_X2 U13646 ( .A1(n16500), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10267) );
  NAND2_X1 U13647 ( .A1(n10271), .A2(n16595), .ZN(n16576) );
  NAND2_X1 U13648 ( .A1(n10290), .A2(n10289), .ZN(n10288) );
  NAND2_X1 U13649 ( .A1(n11174), .A2(n9744), .ZN(n10291) );
  NAND2_X1 U13650 ( .A1(n12841), .A2(n10298), .ZN(n13854) );
  XNOR2_X1 U13651 ( .A(n10298), .B(n10634), .ZN(n13872) );
  INV_X1 U13652 ( .A(n15604), .ZN(n10305) );
  NAND4_X1 U13653 ( .A1(n10305), .A2(n15601), .A3(n15600), .A4(n13884), .ZN(
        n15564) );
  NAND3_X1 U13654 ( .A1(n10494), .A2(n10493), .A3(n10310), .ZN(n13989) );
  AND2_X1 U13655 ( .A1(n10496), .A2(n11531), .ZN(n10310) );
  NAND3_X1 U13656 ( .A1(n10313), .A2(n9890), .A3(n10311), .ZN(n10314) );
  OAI211_X1 U13657 ( .C1(n10315), .C2(n10486), .A(n10314), .B(n11893), .ZN(
        P2_U3025) );
  AND2_X1 U13658 ( .A1(n13896), .A2(n13895), .ZN(n10322) );
  AND2_X1 U13659 ( .A1(n11344), .A2(n10381), .ZN(n16649) );
  NAND3_X1 U13660 ( .A1(n10621), .A2(n11270), .A3(n10484), .ZN(n10615) );
  NAND3_X1 U13661 ( .A1(n10325), .A2(n15551), .A3(n9794), .ZN(n10324) );
  NAND4_X1 U13662 ( .A1(n10330), .A2(n13879), .A3(n10329), .A4(n10642), .ZN(
        n10641) );
  NAND4_X1 U13663 ( .A1(n13843), .A2(n13842), .A3(n13852), .A4(n13862), .ZN(
        n10329) );
  NAND2_X1 U13664 ( .A1(n10331), .A2(n13862), .ZN(n10330) );
  OAI21_X1 U13665 ( .B1(n10715), .B2(n17145), .A(n13860), .ZN(n10331) );
  NAND3_X1 U13666 ( .A1(n11180), .A2(n10333), .A3(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11210) );
  NAND2_X1 U13667 ( .A1(n10430), .A2(n10336), .ZN(n10334) );
  NOR2_X1 U13668 ( .A1(n11173), .A2(n11168), .ZN(n10648) );
  INV_X1 U13669 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10343) );
  OAI21_X1 U13670 ( .B1(n16485), .B2(n14908), .A(n10654), .ZN(n10653) );
  AND2_X1 U13671 ( .A1(n10865), .A2(n13588), .ZN(n10344) );
  NAND3_X1 U13672 ( .A1(n12799), .A2(n12798), .A3(n10782), .ZN(n10347) );
  NAND2_X1 U13673 ( .A1(n10347), .A2(n10346), .ZN(n12841) );
  INV_X1 U13674 ( .A(n12840), .ZN(n10346) );
  NAND2_X1 U13675 ( .A1(n9748), .A2(n9689), .ZN(n10349) );
  OAI21_X2 U13676 ( .B1(n18820), .B2(n10351), .A(n10350), .ZN(n19564) );
  INV_X1 U13677 ( .A(n14853), .ZN(n10357) );
  OAI21_X2 U13678 ( .B1(n10353), .B2(n10357), .A(n12114), .ZN(n19546) );
  NOR3_X2 U13679 ( .A1(n10357), .A2(n12103), .A3(n10355), .ZN(n19520) );
  NAND4_X1 U13680 ( .A1(n10366), .A2(n10361), .A3(n11954), .A4(n11955), .ZN(
        n12195) );
  NAND3_X1 U13681 ( .A1(n11960), .A2(n11957), .A3(n10363), .ZN(n10362) );
  NAND3_X1 U13682 ( .A1(n11967), .A2(n11968), .A3(n10369), .ZN(n10368) );
  NAND3_X1 U13683 ( .A1(n10375), .A2(n10374), .A3(n10931), .ZN(P2_U2984) );
  AOI21_X1 U13684 ( .B1(n11315), .B2(n11282), .A(n16966), .ZN(n10376) );
  NAND2_X1 U13685 ( .A1(n16510), .A2(n10379), .ZN(n10926) );
  NAND2_X1 U13686 ( .A1(n10685), .A2(n11282), .ZN(n10382) );
  OAI21_X1 U13687 ( .B1(n13829), .B2(n12888), .A(n10385), .ZN(n14377) );
  XNOR2_X2 U13688 ( .A(n12884), .B(n12883), .ZN(n13829) );
  NAND2_X1 U13689 ( .A1(n15008), .A2(n10390), .ZN(n14984) );
  NAND2_X1 U13690 ( .A1(n15008), .A2(n15009), .ZN(n14997) );
  NAND3_X1 U13691 ( .A1(n14538), .A2(n10393), .A3(n12927), .ZN(n14723) );
  NAND2_X1 U13692 ( .A1(n13829), .A2(n13871), .ZN(n13836) );
  INV_X1 U13693 ( .A(n15911), .ZN(n10399) );
  MUX2_X1 U13694 ( .A(n15909), .B(n21270), .S(n13829), .Z(n14519) );
  AND2_X1 U13695 ( .A1(n10419), .A2(n10418), .ZN(n12045) );
  NAND2_X1 U13696 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10418) );
  NAND4_X1 U13697 ( .A1(n10422), .A2(n13658), .A3(n10420), .A4(n9856), .ZN(
        P2_U3016) );
  NOR2_X2 U13698 ( .A1(n18420), .A2(n18421), .ZN(n18419) );
  NAND3_X1 U13699 ( .A1(n10426), .A2(n10746), .A3(n9797), .ZN(n10425) );
  NAND2_X1 U13700 ( .A1(n16510), .A2(n10655), .ZN(n14914) );
  INV_X1 U13701 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10440) );
  NAND2_X2 U13702 ( .A1(n14885), .A2(n14884), .ZN(n20637) );
  NAND2_X1 U13703 ( .A1(n10445), .A2(n9863), .ZN(n12865) );
  NOR2_X1 U13704 ( .A1(n10446), .A2(n11922), .ZN(n12044) );
  XNOR2_X1 U13705 ( .A(n12138), .B(n12137), .ZN(n18706) );
  NOR2_X2 U13706 ( .A1(n18710), .A2(n12135), .ZN(n12138) );
  NOR2_X2 U13707 ( .A1(n18739), .A2(n18738), .ZN(n18737) );
  NAND2_X1 U13708 ( .A1(n10451), .A2(n10450), .ZN(n10449) );
  INV_X1 U13709 ( .A(n12232), .ZN(n10451) );
  NAND2_X1 U13710 ( .A1(n10847), .A2(n9783), .ZN(n16267) );
  NAND2_X1 U13711 ( .A1(n10457), .A2(n10452), .ZN(n16364) );
  NAND2_X1 U13712 ( .A1(n10454), .A2(n10453), .ZN(n10452) );
  NAND3_X1 U13713 ( .A1(n10847), .A2(n9783), .A3(n10455), .ZN(n10454) );
  NAND3_X1 U13714 ( .A1(n10847), .A2(n9783), .A3(n10456), .ZN(n10457) );
  INV_X2 U13715 ( .A(n15908), .ZN(n12798) );
  NAND2_X1 U13716 ( .A1(n12799), .A2(n10463), .ZN(n10462) );
  INV_X2 U13717 ( .A(n12910), .ZN(n12799) );
  INV_X1 U13718 ( .A(n16829), .ZN(n10471) );
  NAND2_X1 U13719 ( .A1(n10622), .A2(n10472), .ZN(P2_U3029) );
  NAND2_X1 U13720 ( .A1(n10473), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13721 ( .A1(n16826), .A2(n10935), .ZN(n10473) );
  NAND3_X1 U13722 ( .A1(n10489), .A2(n11346), .A3(n10485), .ZN(n10491) );
  NAND2_X1 U13723 ( .A1(n10641), .A2(n10639), .ZN(n15551) );
  NAND2_X1 U13724 ( .A1(n11485), .A2(n11484), .ZN(n11489) );
  INV_X1 U13725 ( .A(n10866), .ZN(n10611) );
  NOR2_X1 U13726 ( .A1(n13589), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16496) );
  INV_X1 U13727 ( .A(n14019), .ZN(n11485) );
  INV_X1 U13728 ( .A(n10867), .ZN(n10609) );
  NAND2_X1 U13729 ( .A1(n16062), .A2(n10515), .ZN(n10514) );
  AND2_X1 U13730 ( .A1(n16229), .A2(n10523), .ZN(n10521) );
  NAND2_X1 U13731 ( .A1(n10520), .A2(n10522), .ZN(n16193) );
  INV_X1 U13732 ( .A(n10525), .ZN(n16206) );
  OR2_X1 U13733 ( .A1(n13709), .A2(n19778), .ZN(n10530) );
  NAND2_X1 U13734 ( .A1(n13709), .A2(n10528), .ZN(n10527) );
  NAND2_X1 U13735 ( .A1(n13709), .A2(n13708), .ZN(n10531) );
  NAND4_X1 U13736 ( .A1(n11037), .A2(n11035), .A3(n11036), .A4(n11034), .ZN(
        n10535) );
  NAND2_X1 U13737 ( .A1(n10534), .A2(n11006), .ZN(n10537) );
  NAND4_X1 U13738 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11033), .ZN(
        n10534) );
  AND2_X2 U13739 ( .A1(n10539), .A2(n10538), .ZN(n11865) );
  AOI21_X1 U13740 ( .B1(n10554), .B2(n10548), .A(n9853), .ZN(n13770) );
  NOR2_X1 U13741 ( .A1(n16744), .A2(n10553), .ZN(n10552) );
  NOR2_X1 U13742 ( .A1(n16742), .A2(n16744), .ZN(n16729) );
  NAND3_X1 U13743 ( .A1(n13376), .A2(n10561), .A3(n13370), .ZN(n10558) );
  NAND2_X1 U13744 ( .A1(n10575), .A2(n16606), .ZN(n16607) );
  XNOR2_X1 U13745 ( .A(n16669), .B(n10575), .ZN(n16973) );
  INV_X1 U13746 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10592) );
  INV_X2 U13747 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19696) );
  NAND2_X1 U13748 ( .A1(n16629), .A2(n10598), .ZN(n10597) );
  NAND2_X1 U13749 ( .A1(n16629), .A2(n9777), .ZN(n16870) );
  NAND2_X1 U13750 ( .A1(n16629), .A2(n16885), .ZN(n16604) );
  NAND2_X1 U13751 ( .A1(n10597), .A2(n16561), .ZN(n16563) );
  AND3_X1 U13752 ( .A1(n10619), .A2(n11061), .A3(n10617), .ZN(n10620) );
  AOI21_X1 U13753 ( .B1(n11105), .B2(n11054), .A(n10618), .ZN(n10617) );
  NAND2_X1 U13754 ( .A1(n11837), .A2(n11054), .ZN(n10619) );
  NAND2_X1 U13755 ( .A1(n11110), .A2(n10620), .ZN(n11111) );
  AOI21_X1 U13756 ( .B1(n10624), .B2(n16944), .A(n10623), .ZN(n10622) );
  INV_X2 U13757 ( .A(n19546), .ZN(n18949) );
  NAND2_X1 U13758 ( .A1(n12901), .A2(n17176), .ZN(n10636) );
  NAND2_X1 U13759 ( .A1(n15497), .A2(n13898), .ZN(n15437) );
  NAND3_X1 U13760 ( .A1(n15497), .A2(n13898), .A3(n10637), .ZN(n10638) );
  NAND2_X1 U13761 ( .A1(n10736), .A2(n11121), .ZN(n11143) );
  AND4_X2 U13762 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n9821), .ZN(
        n10862) );
  NAND3_X1 U13763 ( .A1(n10661), .A2(n10659), .A3(n10658), .ZN(n10664) );
  NAND2_X1 U13764 ( .A1(n18737), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10658) );
  NAND3_X1 U13765 ( .A1(n10661), .A2(n10662), .A3(n10658), .ZN(n18727) );
  NOR2_X1 U13766 ( .A1(n18737), .A2(n12127), .ZN(n12130) );
  INV_X1 U13767 ( .A(n10664), .ZN(n18725) );
  NAND2_X1 U13768 ( .A1(n20606), .A2(n10676), .ZN(n15188) );
  NAND3_X1 U13769 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .A3(n10683), .ZN(n10682) );
  INV_X2 U13770 ( .A(n17396), .ZN(n17696) );
  NOR2_X1 U13771 ( .A1(n17891), .A2(n18148), .ZN(n17894) );
  NAND2_X1 U13772 ( .A1(n17885), .A2(n10696), .ZN(P3_U2675) );
  NAND2_X1 U13773 ( .A1(n17935), .A2(n9907), .ZN(n17901) );
  NAND2_X1 U13774 ( .A1(n17935), .A2(n10701), .ZN(n17933) );
  INV_X1 U13775 ( .A(n10704), .ZN(n17910) );
  NAND3_X1 U13776 ( .A1(n17060), .A2(P3_EBX_REG_3__SCAN_IN), .A3(
        P3_EBX_REG_4__SCAN_IN), .ZN(n10705) );
  NOR2_X2 U13777 ( .A1(n18126), .A2(n18122), .ZN(n18120) );
  NAND2_X1 U13778 ( .A1(n10709), .A2(n10708), .ZN(n10707) );
  NOR2_X1 U13779 ( .A1(n16725), .A2(n16712), .ZN(n10711) );
  NAND2_X1 U13780 ( .A1(n13843), .A2(n13842), .ZN(n17144) );
  NAND2_X1 U13781 ( .A1(n13900), .A2(n10906), .ZN(n10905) );
  AND2_X2 U13782 ( .A1(n20942), .A2(n12711), .ZN(n14513) );
  NAND2_X1 U13783 ( .A1(n10718), .A2(n10717), .ZN(n20942) );
  INV_X1 U13784 ( .A(n20883), .ZN(n10718) );
  NAND2_X1 U13785 ( .A1(n16028), .A2(n10719), .ZN(n13705) );
  AND2_X1 U13786 ( .A1(n16519), .A2(n13704), .ZN(n10719) );
  INV_X1 U13787 ( .A(n10724), .ZN(n13692) );
  OAI21_X1 U13788 ( .B1(n10729), .B2(n19820), .A(n10725), .ZN(P2_U2826) );
  XNOR2_X1 U13789 ( .A(n15946), .B(n15947), .ZN(n10729) );
  INV_X1 U13790 ( .A(n10730), .ZN(n13687) );
  INV_X1 U13791 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10735) );
  OAI21_X1 U13792 ( .B1(n18701), .B2(n10740), .A(n18700), .ZN(n19001) );
  OR2_X1 U13793 ( .A1(n10741), .A2(n12083), .ZN(n18736) );
  NAND3_X1 U13794 ( .A1(n12199), .A2(n10742), .A3(n12201), .ZN(n10744) );
  NAND3_X1 U13795 ( .A1(n12199), .A2(n12201), .A3(n10943), .ZN(n18562) );
  NOR2_X1 U13796 ( .A1(n17072), .A2(n10746), .ZN(n10745) );
  NAND2_X1 U13797 ( .A1(n10748), .A2(n10751), .ZN(P3_U2831) );
  AND2_X1 U13798 ( .A1(n10755), .A2(n18962), .ZN(n10749) );
  NAND2_X1 U13799 ( .A1(n17217), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10758) );
  NOR2_X1 U13800 ( .A1(n17215), .A2(n10757), .ZN(n10756) );
  NOR2_X4 U13801 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14504) );
  AND2_X2 U13802 ( .A1(n14504), .A2(n14489), .ZN(n12748) );
  NAND3_X1 U13803 ( .A1(n10916), .A2(n12571), .A3(n12638), .ZN(n14056) );
  OAI211_X1 U13804 ( .C1(n15695), .C2(n15671), .A(n10781), .B(n10780), .ZN(
        P1_U2970) );
  NAND2_X1 U13805 ( .A1(n14868), .A2(n14984), .ZN(n14870) );
  NAND2_X1 U13806 ( .A1(n12799), .A2(n12798), .ZN(n12917) );
  AND2_X1 U13807 ( .A1(n10784), .A2(n11602), .ZN(n11071) );
  NAND3_X1 U13808 ( .A1(n11059), .A2(n11058), .A3(n10784), .ZN(n11077) );
  AND2_X2 U13809 ( .A1(n11015), .A2(n11063), .ZN(n10784) );
  NAND3_X1 U13810 ( .A1(n11643), .A2(n11060), .A3(n11607), .ZN(n11061) );
  NAND3_X1 U13811 ( .A1(n11134), .A2(n11533), .A3(n11146), .ZN(n16689) );
  AND2_X1 U13812 ( .A1(n12490), .A2(n9766), .ZN(n13788) );
  AND2_X2 U13813 ( .A1(n12490), .A2(n9887), .ZN(n13605) );
  INV_X1 U13814 ( .A(n14655), .ZN(n10795) );
  NAND2_X1 U13815 ( .A1(n10795), .A2(n9740), .ZN(n14740) );
  NAND2_X1 U13816 ( .A1(n10798), .A2(n9865), .ZN(n16329) );
  INV_X1 U13817 ( .A(n14923), .ZN(n15945) );
  AOI21_X1 U13818 ( .B1(n14923), .B2(n16970), .A(n10801), .ZN(n10800) );
  NAND2_X1 U13819 ( .A1(n11901), .A2(n9892), .ZN(n12482) );
  NAND3_X1 U13820 ( .A1(n11671), .A2(n11654), .A3(n10803), .ZN(n14269) );
  NAND2_X1 U13821 ( .A1(n11652), .A2(n11653), .ZN(n10803) );
  NAND3_X1 U13822 ( .A1(n11656), .A2(P2_REIP_REG_0__SCAN_IN), .A3(n11663), 
        .ZN(n10804) );
  NAND2_X1 U13823 ( .A1(n14268), .A2(n14269), .ZN(n11666) );
  NAND2_X1 U13824 ( .A1(n14747), .A2(n11692), .ZN(n10805) );
  NAND2_X1 U13825 ( .A1(n10805), .A2(n10806), .ZN(n14287) );
  AND2_X1 U13826 ( .A1(n13781), .A2(n10818), .ZN(n13622) );
  NAND2_X1 U13827 ( .A1(n13781), .A2(n13782), .ZN(n13780) );
  NOR2_X2 U13828 ( .A1(n14254), .A2(n10820), .ZN(n14439) );
  NOR2_X2 U13829 ( .A1(n14472), .A2(n10824), .ZN(n14809) );
  NAND2_X1 U13830 ( .A1(n10836), .A2(n10834), .ZN(n15118) );
  NAND2_X1 U13831 ( .A1(n12210), .A2(n10853), .ZN(n10850) );
  OAI211_X1 U13832 ( .C1(n12210), .C2(n10852), .A(n10851), .B(n10850), .ZN(
        n14522) );
  INV_X1 U13833 ( .A(n10863), .ZN(n10861) );
  AND2_X1 U13834 ( .A1(n10867), .A2(n16584), .ZN(n10865) );
  AND2_X2 U13835 ( .A1(n10868), .A2(n10932), .ZN(n10866) );
  NAND3_X1 U13836 ( .A1(n10892), .A2(n11457), .A3(n10895), .ZN(n11431) );
  INV_X2 U13837 ( .A(n11461), .ZN(n10895) );
  NOR2_X2 U13838 ( .A1(n15998), .A2(n11378), .ZN(n13589) );
  NAND2_X1 U13839 ( .A1(n11518), .A2(n10900), .ZN(n10899) );
  NAND2_X1 U13840 ( .A1(n11518), .A2(n11517), .ZN(n11869) );
  NAND2_X2 U13841 ( .A1(n10899), .A2(n10897), .ZN(n13570) );
  NOR2_X1 U13842 ( .A1(n15621), .A2(n15690), .ZN(n10913) );
  AND2_X2 U13843 ( .A1(n12467), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11355) );
  NAND2_X1 U13844 ( .A1(n14466), .A2(n14542), .ZN(n17151) );
  XNOR2_X1 U13845 ( .A(n11912), .B(n11911), .ZN(n16775) );
  NOR2_X1 U13846 ( .A1(n19696), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12168) );
  NOR2_X1 U13847 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  NAND2_X1 U13848 ( .A1(n17213), .A2(n18573), .ZN(n17217) );
  OAI21_X1 U13849 ( .B1(n13622), .B2(n13623), .A(n13648), .ZN(n16376) );
  NAND2_X1 U13850 ( .A1(n15081), .A2(n15080), .ZN(n15067) );
  AND2_X1 U13851 ( .A1(n14444), .A2(n14443), .ZN(n19814) );
  INV_X1 U13852 ( .A(n9809), .ZN(n13620) );
  INV_X1 U13854 ( .A(n13581), .ZN(n13584) );
  CLKBUF_X1 U13855 ( .A(n14823), .Z(n16144) );
  NAND2_X1 U13856 ( .A1(n14823), .A2(n11570), .ZN(n14822) );
  NOR2_X2 U13857 ( .A1(n14023), .A2(n16143), .ZN(n14823) );
  NAND2_X1 U13858 ( .A1(n11561), .A2(n11560), .ZN(n14023) );
  NAND2_X1 U13859 ( .A1(n11888), .A2(n11887), .ZN(n16043) );
  INV_X1 U13860 ( .A(n11884), .ZN(n11888) );
  NAND2_X1 U13861 ( .A1(n13488), .A2(n13487), .ZN(n15152) );
  CLKBUF_X1 U13862 ( .A(n14022), .Z(n14844) );
  INV_X1 U13863 ( .A(n14022), .ZN(n11561) );
  AND3_X1 U13864 ( .A1(n12670), .A2(n14587), .A3(n12645), .ZN(n12646) );
  NOR2_X2 U13865 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10955) );
  INV_X1 U13866 ( .A(n14377), .ZN(n12908) );
  AND2_X1 U13867 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  NOR2_X1 U13868 ( .A1(n12210), .A2(n11154), .ZN(n11170) );
  NOR2_X1 U13869 ( .A1(n12210), .A2(n11158), .ZN(n11166) );
  INV_X1 U13870 ( .A(n15185), .ZN(n13488) );
  AOI22_X1 U13871 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10963) );
  NAND2_X1 U13872 ( .A1(n16704), .A2(n11145), .ZN(n11150) );
  INV_X1 U13873 ( .A(n11055), .ZN(n11081) );
  XNOR2_X1 U13874 ( .A(n12731), .B(n12730), .ZN(n12901) );
  CLKBUF_X1 U13875 ( .A(n12463), .Z(n12457) );
  AOI22_X1 U13876 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11041) );
  NAND2_X1 U13877 ( .A1(n11065), .A2(n11063), .ZN(n14811) );
  AOI22_X1 U13878 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12740), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12519) );
  BUF_X1 U13879 ( .A(n12881), .Z(n12884) );
  NAND2_X1 U13880 ( .A1(n16265), .A2(n16715), .ZN(n13986) );
  NAND2_X1 U13881 ( .A1(n16265), .A2(n16970), .ZN(n13761) );
  INV_X1 U13882 ( .A(n14279), .ZN(n11712) );
  NAND2_X1 U13883 ( .A1(n14876), .A2(n14875), .ZN(n14879) );
  AOI21_X1 U13884 ( .B1(n14876), .B2(n20715), .A(n13979), .ZN(n13980) );
  NAND2_X1 U13885 ( .A1(n15907), .A2(n15911), .ZN(n21126) );
  NOR2_X1 U13886 ( .A1(n18197), .A2(n18191), .ZN(n18186) );
  INV_X1 U13887 ( .A(n15418), .ZN(n15407) );
  INV_X1 U13888 ( .A(n20641), .ZN(n20610) );
  NOR2_X1 U13889 ( .A1(n13429), .A2(n13428), .ZN(n10929) );
  OR2_X1 U13890 ( .A1(n16830), .A2(n16808), .ZN(n10930) );
  AND2_X1 U13891 ( .A1(n13663), .A2(n13662), .ZN(n10931) );
  AND4_X1 U13892 ( .A1(n13552), .A2(n13551), .A3(n13550), .A4(n11525), .ZN(
        n10932) );
  INV_X1 U13893 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19598) );
  OR2_X1 U13894 ( .A1(n18945), .A2(n18845), .ZN(n10933) );
  AND2_X1 U13895 ( .A1(n16351), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10934) );
  OR2_X1 U13896 ( .A1(n16810), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10935) );
  AND2_X1 U13897 ( .A1(n19040), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n10936) );
  NAND2_X2 U13898 ( .A1(n15418), .A2(n14588), .ZN(n15421) );
  AND2_X1 U13899 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10937) );
  INV_X1 U13900 ( .A(n12315), .ZN(n14662) );
  INV_X1 U13901 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n21624) );
  INV_X1 U13902 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11591) );
  AND2_X1 U13903 ( .A1(n13894), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10938) );
  INV_X1 U13904 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20783) );
  AND2_X1 U13905 ( .A1(n15509), .A2(n15508), .ZN(n10939) );
  OR3_X1 U13906 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n18501), .ZN(n10940) );
  INV_X1 U13907 ( .A(n13619), .ZN(n11808) );
  INV_X1 U13908 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19734) );
  AND2_X1 U13909 ( .A1(n14812), .A2(n17038), .ZN(n16464) );
  AND2_X1 U13910 ( .A1(n13730), .A2(n19832), .ZN(n10941) );
  AND2_X1 U13911 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .ZN(n10942) );
  INV_X2 U13912 ( .A(n18399), .ZN(n18403) );
  INV_X1 U13913 ( .A(n16712), .ZN(n16697) );
  NAND2_X1 U13914 ( .A1(n19738), .A2(n11590), .ZN(n16672) );
  AND2_X1 U13915 ( .A1(n16672), .A2(n14452), .ZN(n16715) );
  INV_X1 U13916 ( .A(n16715), .ZN(n16695) );
  INV_X1 U13917 ( .A(n21380), .ZN(n21392) );
  AND2_X1 U13918 ( .A1(n10618), .A2(n20528), .ZN(n19788) );
  OR2_X1 U13919 ( .A1(n18673), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10943) );
  OR2_X1 U13920 ( .A1(n19738), .A2(n11650), .ZN(n16680) );
  INV_X1 U13921 ( .A(n16680), .ZN(n11531) );
  INV_X1 U13922 ( .A(n13582), .ZN(n15984) );
  INV_X1 U13923 ( .A(n13549), .ZN(n11525) );
  INV_X1 U13924 ( .A(n12885), .ZN(n13339) );
  AND3_X1 U13925 ( .A1(n11015), .A2(n11075), .A3(n11064), .ZN(n10945) );
  INV_X1 U13926 ( .A(n15336), .ZN(n20651) );
  INV_X1 U13927 ( .A(n14429), .ZN(n15430) );
  INV_X1 U13928 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12666) );
  AND4_X1 U13929 ( .A1(n12566), .A2(n12565), .A3(n12564), .A4(n12563), .ZN(
        n10947) );
  INV_X1 U13930 ( .A(n12718), .ZN(n12697) );
  NAND2_X1 U13931 ( .A1(n12811), .A2(n12810), .ZN(n10948) );
  BUF_X4 U13932 ( .A(n13454), .Z(n13528) );
  NAND2_X1 U13933 ( .A1(n13912), .A2(n12637), .ZN(n12670) );
  INV_X1 U13934 ( .A(n13912), .ZN(n12633) );
  AND4_X1 U13935 ( .A1(n12514), .A2(n12513), .A3(n12512), .A4(n12511), .ZN(
        n10950) );
  INV_X1 U13936 ( .A(n11126), .ZN(n12506) );
  AND2_X1 U13937 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11087) );
  INV_X1 U13938 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13362) );
  NAND2_X1 U13939 ( .A1(n11064), .A2(n11065), .ZN(n11028) );
  AOI22_X1 U13940 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12713), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12511) );
  OR2_X1 U13941 ( .A1(n11369), .A2(n11368), .ZN(n11371) );
  OR2_X1 U13942 ( .A1(n12707), .A2(n12706), .ZN(n12708) );
  OR2_X1 U13943 ( .A1(n12821), .A2(n12820), .ZN(n13865) );
  OR2_X1 U13944 ( .A1(n12809), .A2(n12808), .ZN(n13845) );
  INV_X1 U13945 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11445) );
  INV_X1 U13946 ( .A(n11398), .ZN(n11397) );
  AOI22_X1 U13947 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11036) );
  BUF_X1 U13948 ( .A(n11077), .Z(n11643) );
  AOI22_X1 U13949 ( .A1(n11614), .A2(n11613), .B1(n11612), .B2(n11611), .ZN(
        n11620) );
  INV_X1 U13950 ( .A(n13047), .ZN(n13048) );
  INV_X1 U13951 ( .A(n12708), .ZN(n13830) );
  OR2_X1 U13952 ( .A1(n13867), .A2(n13866), .ZN(n13875) );
  NAND2_X1 U13953 ( .A1(n13839), .A2(n20733), .ZN(n13840) );
  AND2_X1 U13954 ( .A1(n12731), .A2(n12729), .ZN(n12712) );
  INV_X1 U13955 ( .A(n13710), .ZN(n13712) );
  OAI21_X2 U13956 ( .B1(n11425), .B2(n19879), .A(n11424), .ZN(n11462) );
  INV_X1 U13957 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11484) );
  INV_X1 U13958 ( .A(n11532), .ZN(n11533) );
  NAND2_X1 U13959 ( .A1(n11020), .A2(n11006), .ZN(n11027) );
  INV_X1 U13960 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n21487) );
  NOR2_X1 U13961 ( .A1(n11922), .A2(n17750), .ZN(n11931) );
  OR2_X1 U13962 ( .A1(n14566), .A2(n17176), .ZN(n12784) );
  INV_X1 U13963 ( .A(n13375), .ZN(n13391) );
  MUX2_X1 U13964 ( .A(n13521), .B(n13522), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13436) );
  AND2_X1 U13965 ( .A1(n14891), .A2(n14893), .ZN(n12927) );
  NOR2_X1 U13966 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12885) );
  INV_X1 U13967 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12864) );
  NAND2_X1 U13968 ( .A1(n20745), .A2(n13838), .ZN(n14625) );
  INV_X1 U13969 ( .A(n13570), .ZN(n13572) );
  INV_X1 U13970 ( .A(n11432), .ZN(n11429) );
  OR2_X1 U13971 ( .A1(n11405), .A2(n11404), .ZN(n11407) );
  INV_X1 U13972 ( .A(n11879), .ZN(n11878) );
  INV_X1 U13973 ( .A(n14025), .ZN(n11560) );
  NOR2_X1 U13974 ( .A1(n11378), .A2(n13787), .ZN(n13583) );
  INV_X1 U13975 ( .A(n13547), .ZN(n11524) );
  AND2_X1 U13976 ( .A1(n13641), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11435) );
  INV_X1 U13977 ( .A(n11623), .ZN(n11624) );
  INV_X1 U13978 ( .A(n11385), .ZN(n11602) );
  INV_X1 U13979 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n21568) );
  NOR2_X1 U13980 ( .A1(n12164), .A2(n12163), .ZN(n12172) );
  INV_X1 U13981 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n21691) );
  INV_X1 U13982 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21639) );
  INV_X1 U13983 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21702) );
  OR2_X1 U13984 ( .A1(n18887), .A2(n18942), .ZN(n18816) );
  INV_X1 U13985 ( .A(n12070), .ZN(n11976) );
  NAND2_X1 U13986 ( .A1(n12085), .A2(n12084), .ZN(n12088) );
  INV_X1 U13987 ( .A(n20622), .ZN(n20607) );
  OR2_X1 U13988 ( .A1(n14060), .A2(n21341), .ZN(n14196) );
  NAND2_X1 U13989 ( .A1(n12636), .A2(n14566), .ZN(n12677) );
  NAND2_X1 U13990 ( .A1(n12976), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13047) );
  INV_X1 U13991 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U13992 ( .A1(n13898), .A2(n9689), .ZN(n15470) );
  NAND2_X1 U13993 ( .A1(n21031), .A2(n17176), .ZN(n12797) );
  INV_X1 U13994 ( .A(n14739), .ZN(n11548) );
  NAND2_X1 U13995 ( .A1(n11407), .A2(n11406), .ZN(n11623) );
  INV_X1 U13996 ( .A(n12460), .ZN(n12469) );
  INV_X1 U13997 ( .A(n12406), .ZN(n16282) );
  INV_X1 U13998 ( .A(n16320), .ZN(n12292) );
  AND2_X1 U13999 ( .A1(n11813), .A2(n11812), .ZN(n16106) );
  INV_X1 U14000 ( .A(n14471), .ZN(n11779) );
  AND2_X1 U14001 ( .A1(n14677), .A2(n11842), .ZN(n14701) );
  INV_X1 U14002 ( .A(n13587), .ZN(n13588) );
  OR2_X1 U14003 ( .A1(n11523), .A2(n16779), .ZN(n11910) );
  INV_X1 U14004 ( .A(n11147), .ZN(n11148) );
  NAND2_X1 U14005 ( .A1(n11607), .A2(n11624), .ZN(n11625) );
  INV_X1 U14006 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U14007 ( .A1(n20403), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19891) );
  NAND2_X1 U14008 ( .A1(n18572), .A2(n18806), .ZN(n12202) );
  INV_X1 U14009 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U14010 ( .A1(n13402), .A2(n13394), .ZN(n13395) );
  AND2_X1 U14011 ( .A1(n13903), .A2(n17110), .ZN(n13425) );
  OR2_X1 U14012 ( .A1(n14175), .A2(n14196), .ZN(n14584) );
  INV_X1 U14013 ( .A(n13339), .ZN(n13332) );
  INV_X1 U14014 ( .A(n14376), .ZN(n12907) );
  OR3_X1 U14015 ( .A1(n15735), .A2(n15716), .A3(n13966), .ZN(n15707) );
  AND2_X1 U14016 ( .A1(n13501), .A2(n13500), .ZN(n15105) );
  OR3_X1 U14017 ( .A1(n20737), .A2(n17149), .A3(n14622), .ZN(n15891) );
  INV_X1 U14018 ( .A(n20756), .ZN(n20722) );
  AND2_X1 U14019 ( .A1(n14517), .A2(n21273), .ZN(n21270) );
  NOR2_X1 U14020 ( .A1(n21154), .A2(n20824), .ZN(n21096) );
  INV_X1 U14021 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21156) );
  AND2_X1 U14022 ( .A1(n21034), .A2(n20919), .ZN(n21236) );
  INV_X1 U14023 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n12628) );
  NAND2_X1 U14024 ( .A1(n13725), .A2(n19809), .ZN(n13726) );
  AND2_X1 U14025 ( .A1(n13615), .A2(n13614), .ZN(n15989) );
  NOR2_X2 U14026 ( .A1(n12482), .A2(n16037), .ZN(n16021) );
  INV_X1 U14027 ( .A(n19812), .ZN(n19789) );
  OR2_X1 U14028 ( .A1(n15942), .A2(n13732), .ZN(n19812) );
  AND3_X1 U14029 ( .A1(n11752), .A2(n11751), .A3(n11750), .ZN(n14016) );
  INV_X1 U14030 ( .A(n13753), .ZN(n12507) );
  OR2_X1 U14031 ( .A1(n16033), .A2(n13586), .ZN(n13775) );
  OR2_X1 U14032 ( .A1(n16154), .A2(n11495), .ZN(n16584) );
  INV_X1 U14033 ( .A(n14523), .ZN(n14524) );
  NAND2_X1 U14034 ( .A1(n17022), .A2(n14456), .ZN(n14458) );
  INV_X1 U14035 ( .A(n20528), .ZN(n20343) );
  OR2_X1 U14036 ( .A1(n20537), .A2(n20524), .ZN(n19909) );
  OR2_X1 U14037 ( .A1(n20537), .A2(n19998), .ZN(n19961) );
  OR2_X1 U14038 ( .A1(n19891), .A2(n11650), .ZN(n20352) );
  OR2_X1 U14039 ( .A1(n19891), .A2(n11082), .ZN(n20362) );
  INV_X1 U14040 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11127) );
  INV_X1 U14041 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20454) );
  NAND2_X1 U14042 ( .A1(n17709), .A2(n18302), .ZN(n17385) );
  AND2_X1 U14043 ( .A1(n18153), .A2(n10942), .ZN(n18154) );
  INV_X1 U14044 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21610) );
  INV_X1 U14045 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18602) );
  INV_X1 U14046 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18545) );
  INV_X1 U14047 ( .A(n18858), .ZN(n18945) );
  INV_X1 U14048 ( .A(n12098), .ZN(n12097) );
  NAND2_X1 U14049 ( .A1(n19557), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19340) );
  INV_X1 U14050 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19519) );
  INV_X1 U14051 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21398) );
  AND2_X1 U14052 ( .A1(n20638), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14884) );
  INV_X1 U14053 ( .A(n20655), .ZN(n15319) );
  OR2_X1 U14054 ( .A1(n15407), .A2(n14590), .ZN(n14877) );
  INV_X1 U14055 ( .A(n15399), .ZN(n15392) );
  AND2_X1 U14056 ( .A1(n14590), .A2(n14589), .ZN(n14588) );
  AND2_X1 U14057 ( .A1(n15673), .A2(n14210), .ZN(n15517) );
  INV_X1 U14058 ( .A(n15671), .ZN(n20716) );
  AND2_X1 U14059 ( .A1(n15833), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15810) );
  INV_X1 U14060 ( .A(n20781), .ZN(n20727) );
  INV_X1 U14061 ( .A(n20774), .ZN(n20736) );
  AND2_X1 U14062 ( .A1(n13944), .A2(n14180), .ZN(n20756) );
  INV_X1 U14063 ( .A(n21273), .ZN(n21266) );
  OAI211_X1 U14064 ( .C1(n20828), .C2(n21091), .A(n21096), .B(n20796), .ZN(
        n20830) );
  INV_X1 U14065 ( .A(n20785), .ZN(n20848) );
  OAI22_X1 U14066 ( .A1(n20859), .A2(n20858), .B1(n21034), .B2(n20974), .ZN(
        n20877) );
  INV_X1 U14067 ( .A(n20912), .ZN(n20904) );
  OAI21_X1 U14068 ( .B1(n20937), .B2(n20920), .A(n21236), .ZN(n20939) );
  INV_X1 U14069 ( .A(n20972), .ZN(n20996) );
  INV_X1 U14070 ( .A(n21029), .ZN(n21021) );
  INV_X1 U14071 ( .A(n21069), .ZN(n21080) );
  INV_X1 U14072 ( .A(n21084), .ZN(n21111) );
  INV_X1 U14073 ( .A(n21133), .ZN(n21144) );
  INV_X1 U14074 ( .A(n21149), .ZN(n21193) );
  OR2_X1 U14075 ( .A1(n9707), .A2(n20784), .ZN(n21148) );
  OR2_X1 U14076 ( .A1(n9707), .A2(n13816), .ZN(n21206) );
  INV_X1 U14077 ( .A(n20797), .ZN(n21275) );
  INV_X1 U14078 ( .A(n20808), .ZN(n21295) );
  AND2_X1 U14079 ( .A1(n20919), .A2(n20816), .ZN(n21306) );
  NAND2_X1 U14080 ( .A1(n9707), .A2(n20784), .ZN(n21125) );
  INV_X1 U14081 ( .A(n21409), .ZN(n21341) );
  INV_X1 U14082 ( .A(n21385), .ZN(n21387) );
  AND2_X1 U14084 ( .A1(n13734), .A2(n13724), .ZN(n19809) );
  OR2_X1 U14085 ( .A1(n14941), .A2(n13735), .ZN(n19807) );
  AND2_X1 U14086 ( .A1(n16036), .A2(n11881), .ZN(n16310) );
  OR2_X1 U14087 ( .A1(n14801), .A2(n14800), .ZN(n16344) );
  OR2_X1 U14088 ( .A1(n11707), .A2(n11706), .ZN(n14768) );
  INV_X1 U14089 ( .A(n19834), .ZN(n14785) );
  INV_X2 U14090 ( .A(n11650), .ZN(n14347) );
  INV_X1 U14091 ( .A(n14067), .ZN(n14143) );
  NAND3_X1 U14092 ( .A1(n11628), .A2(n14705), .A3(n13720), .ZN(n14046) );
  AND2_X1 U14093 ( .A1(n14834), .A2(n14825), .ZN(n16852) );
  INV_X1 U14094 ( .A(n16348), .ZN(n16880) );
  INV_X1 U14095 ( .A(n17180), .ZN(n16989) );
  INV_X1 U14096 ( .A(n17193), .ZN(n16993) );
  NAND2_X1 U14097 ( .A1(n11865), .A2(n11825), .ZN(n17180) );
  AND2_X1 U14098 ( .A1(n14709), .A2(n11633), .ZN(n20545) );
  INV_X1 U14099 ( .A(n14715), .ZN(n14344) );
  INV_X1 U14100 ( .A(n19929), .ZN(n19896) );
  NAND2_X1 U14101 ( .A1(n14458), .A2(n14457), .ZN(n19930) );
  OAI21_X1 U14102 ( .B1(n19969), .B2(n19968), .A(n19967), .ZN(n19990) );
  OAI21_X1 U14103 ( .B1(n20343), .B2(n19999), .A(n19996), .ZN(n20018) );
  AND2_X1 U14104 ( .A1(n20057), .A2(n20306), .ZN(n20051) );
  INV_X1 U14105 ( .A(n20154), .ZN(n20117) );
  OAI21_X1 U14106 ( .B1(n20125), .B2(n20124), .A(n20123), .ZN(n20150) );
  INV_X1 U14107 ( .A(n20023), .ZN(n20095) );
  NAND2_X1 U14108 ( .A1(n20165), .A2(n20164), .ZN(n20190) );
  OAI21_X1 U14109 ( .B1(n20203), .B2(n20219), .A(n20403), .ZN(n20221) );
  INV_X1 U14110 ( .A(n20263), .ZN(n20253) );
  NOR2_X2 U14111 ( .A1(n20270), .A2(n20269), .ZN(n20332) );
  OAI21_X1 U14112 ( .B1(n20349), .B2(n20348), .A(n20347), .ZN(n20385) );
  NOR2_X1 U14113 ( .A1(n20155), .A2(n17033), .ZN(n20307) );
  INV_X1 U14114 ( .A(n20363), .ZN(n20417) );
  INV_X1 U14115 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20464) );
  NOR2_X1 U14116 ( .A1(n19532), .A2(n17381), .ZN(n19510) );
  OR2_X1 U14117 ( .A1(n17414), .A2(n17413), .ZN(n17415) );
  NOR2_X1 U14118 ( .A1(n17757), .A2(n17399), .ZN(n17438) );
  NOR2_X1 U14119 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17491), .ZN(n17463) );
  NOR2_X1 U14120 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17533), .ZN(n17520) );
  NOR2_X1 U14121 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17555), .ZN(n17541) );
  NOR2_X1 U14122 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17603), .ZN(n17585) );
  NOR2_X1 U14123 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17624), .ZN(n17610) );
  NOR2_X1 U14124 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17700), .ZN(n17684) );
  INV_X1 U14125 ( .A(n17767), .ZN(n17751) );
  INV_X1 U14126 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18125) );
  INV_X1 U14127 ( .A(n18233), .ZN(n18222) );
  INV_X1 U14128 ( .A(n18263), .ZN(n18286) );
  INV_X1 U14129 ( .A(n18300), .ZN(n18341) );
  INV_X1 U14130 ( .A(n18943), .ZN(n18645) );
  OAI21_X1 U14131 ( .B1(n18444), .B2(n18970), .A(n12206), .ZN(n12207) );
  NOR2_X1 U14132 ( .A1(n18859), .A2(n12203), .ZN(n18806) );
  INV_X1 U14133 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21613) );
  INV_X1 U14134 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18905) );
  INV_X1 U14135 ( .A(n18920), .ZN(n18948) );
  AOI21_X2 U14136 ( .B1(n12198), .B2(n12197), .A(n19573), .ZN(n19039) );
  NAND2_X1 U14137 ( .A1(n19676), .A2(n19666), .ZN(n19726) );
  INV_X1 U14138 ( .A(n19167), .ZN(n19169) );
  NOR2_X1 U14139 ( .A1(n19553), .A2(n19072), .ZN(n19246) );
  CLKBUF_X1 U14140 ( .A(n19350), .Z(n19355) );
  INV_X1 U14141 ( .A(n19477), .ZN(n19430) );
  INV_X1 U14142 ( .A(n19716), .ZN(n19586) );
  INV_X1 U14143 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21543) );
  NAND2_X1 U14144 ( .A1(n14011), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n17040)
         );
  INV_X1 U14145 ( .A(U212), .ZN(n17313) );
  INV_X1 U14146 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21232) );
  NAND2_X1 U14147 ( .A1(n13534), .A2(n20627), .ZN(n13535) );
  INV_X1 U14148 ( .A(n20627), .ZN(n20648) );
  INV_X1 U14149 ( .A(n20650), .ZN(n15334) );
  OAI21_X1 U14150 ( .B1(n9900), .B2(n9786), .A(n15130), .ZN(n15545) );
  INV_X1 U14151 ( .A(n15629), .ZN(n15414) );
  AND2_X1 U14152 ( .A1(n14406), .A2(n14405), .ZN(n20825) );
  NOR2_X2 U14153 ( .A1(n15397), .A2(n14591), .ZN(n15419) );
  NAND2_X1 U14154 ( .A1(n20671), .A2(n14566), .ZN(n14325) );
  NAND2_X1 U14155 ( .A1(n20686), .A2(n20680), .ZN(n20678) );
  INV_X1 U14156 ( .A(n20671), .ZN(n20686) );
  NOR2_X1 U14157 ( .A1(n14384), .A2(n14383), .ZN(n15429) );
  INV_X2 U14158 ( .A(n15517), .ZN(n20720) );
  NAND2_X1 U14159 ( .A1(n13944), .A2(n13929), .ZN(n20774) );
  INV_X1 U14160 ( .A(n20757), .ZN(n20775) );
  NAND2_X1 U14161 ( .A1(n14512), .A2(n20824), .ZN(n20782) );
  AOI22_X1 U14162 ( .A1(n20795), .A2(n20793), .B1(n21089), .B2(n20789), .ZN(
        n20833) );
  OR2_X1 U14163 ( .A1(n20881), .A2(n21206), .ZN(n20866) );
  OR2_X1 U14164 ( .A1(n20881), .A2(n21231), .ZN(n20912) );
  OR2_X1 U14165 ( .A1(n20881), .A2(n21125), .ZN(n20927) );
  NAND2_X1 U14166 ( .A1(n21008), .A2(n20948), .ZN(n20972) );
  AOI22_X1 U14167 ( .A1(n20979), .A2(n20976), .B1(n21154), .B2(n20975), .ZN(
        n21001) );
  NAND2_X1 U14168 ( .A1(n21008), .A2(n20971), .ZN(n21029) );
  NAND2_X1 U14169 ( .A1(n21008), .A2(n21007), .ZN(n21044) );
  OR2_X1 U14170 ( .A1(n21126), .A2(n21148), .ZN(n21069) );
  AOI22_X1 U14171 ( .A1(n21094), .A2(n21090), .B1(n21089), .B2(n21088), .ZN(
        n21116) );
  OR2_X1 U14172 ( .A1(n21126), .A2(n21125), .ZN(n21149) );
  INV_X1 U14173 ( .A(n21294), .ZN(n21178) );
  OR2_X1 U14174 ( .A1(n21265), .A2(n21148), .ZN(n21213) );
  OR2_X1 U14175 ( .A1(n21265), .A2(n21206), .ZN(n21244) );
  OR2_X1 U14176 ( .A1(n21265), .A2(n21231), .ZN(n21291) );
  INV_X1 U14177 ( .A(n21397), .ZN(n21331) );
  NOR2_X1 U14178 ( .A1(n21392), .A2(n20566), .ZN(n21397) );
  INV_X1 U14179 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21353) );
  INV_X1 U14180 ( .A(n21381), .ZN(n21385) );
  INV_X1 U14181 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20198) );
  INV_X1 U14182 ( .A(n13739), .ZN(n13740) );
  INV_X1 U14183 ( .A(n19787), .ZN(n19815) );
  OR2_X1 U14184 ( .A1(n14841), .A2(n14840), .ZN(n16865) );
  INV_X1 U14185 ( .A(n19819), .ZN(n16238) );
  AND2_X1 U14186 ( .A1(n12478), .A2(n10538), .ZN(n19832) );
  AND2_X1 U14187 ( .A1(n14262), .A2(n10538), .ZN(n19840) );
  NAND2_X1 U14188 ( .A1(n14263), .A2(n19840), .ZN(n16475) );
  NAND2_X1 U14189 ( .A1(n14231), .A2(n11607), .ZN(n14360) );
  OR2_X1 U14190 ( .A1(n14230), .A2(n11127), .ZN(n15940) );
  OR2_X1 U14191 ( .A1(n14046), .A2(n14045), .ZN(n14067) );
  OR2_X1 U14192 ( .A1(n19738), .A2(n14347), .ZN(n16712) );
  NAND2_X1 U14193 ( .A1(n11865), .A2(n20546), .ZN(n17182) );
  INV_X1 U14194 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14714) );
  INV_X1 U14195 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17056) );
  NAND2_X1 U14196 ( .A1(n20160), .A2(n20057), .ZN(n19929) );
  AOI211_X2 U14197 ( .C1(n19932), .C2(n20528), .A(n19931), .B(n19930), .ZN(
        n19959) );
  INV_X1 U14198 ( .A(n19989), .ZN(n19987) );
  INV_X1 U14199 ( .A(n20019), .ZN(n20010) );
  INV_X1 U14200 ( .A(n20051), .ZN(n20049) );
  INV_X1 U14201 ( .A(n20108), .ZN(n20115) );
  NAND2_X1 U14202 ( .A1(n20307), .A2(n20160), .ZN(n20224) );
  AND2_X1 U14203 ( .A1(n20234), .A2(n20233), .ZN(n20252) );
  NAND2_X1 U14204 ( .A1(n20307), .A2(n20522), .ZN(n20295) );
  INV_X1 U14205 ( .A(n20435), .ZN(n20328) );
  NAND2_X1 U14206 ( .A1(n20307), .A2(n20306), .ZN(n20389) );
  NAND3_X1 U14207 ( .A1(n11127), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19736) );
  INV_X1 U14208 ( .A(n20520), .ZN(n20445) );
  NAND2_X1 U14209 ( .A1(n19734), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20557) );
  INV_X1 U14210 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19714) );
  AOI211_X1 U14211 ( .C1(n17417), .C2(n17771), .A(n17404), .B(n17403), .ZN(
        n17405) );
  INV_X1 U14212 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18072) );
  INV_X1 U14213 ( .A(n17715), .ZN(n17753) );
  AND2_X1 U14214 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18247), .ZN(n18250) );
  NOR2_X1 U14215 ( .A1(n12068), .A2(n12067), .ZN(n18278) );
  NAND2_X1 U14216 ( .A1(n18333), .A2(n18302), .ZN(n18318) );
  NAND2_X1 U14217 ( .A1(n18300), .A2(n18299), .ZN(n18340) );
  AOI211_X1 U14218 ( .C1(n18343), .C2(n19586), .A(n18342), .B(n18341), .ZN(
        n18388) );
  INV_X1 U14219 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21474) );
  AOI21_X1 U14220 ( .B1(n12208), .B2(n19039), .A(n12207), .ZN(n12209) );
  INV_X1 U14221 ( .A(n19055), .ZN(n18963) );
  INV_X1 U14222 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18900) );
  INV_X1 U14223 ( .A(n19047), .ZN(n19053) );
  AND2_X1 U14224 ( .A1(n19726), .A2(n17360), .ZN(n19710) );
  INV_X1 U14225 ( .A(n19215), .ZN(n19211) );
  INV_X1 U14226 ( .A(n19263), .ZN(n19261) );
  INV_X1 U14227 ( .A(n19311), .ZN(n19309) );
  INV_X1 U14228 ( .A(n19383), .ZN(n19376) );
  INV_X1 U14229 ( .A(n19401), .ZN(n19412) );
  INV_X1 U14230 ( .A(n19473), .ZN(n19433) );
  INV_X1 U14231 ( .A(n19303), .ZN(n19489) );
  INV_X1 U14232 ( .A(n17745), .ZN(n19581) );
  INV_X1 U14233 ( .A(n19663), .ZN(n19585) );
  OAI211_X1 U14234 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(P3_STATE_REG_1__SCAN_IN), .A(n19648), .B(n19598), .ZN(n19713) );
  INV_X1 U14235 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19606) );
  NAND2_X1 U14236 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n19723), .ZN(n19655) );
  NOR2_X1 U14237 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14014), .ZN(n17338)
         );
  INV_X1 U14238 ( .A(n17318), .ZN(n17316) );
  INV_X1 U14239 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20510) );
  OR4_X1 U14240 ( .A1(n14031), .A2(n14030), .A3(n14029), .A4(n14028), .ZN(
        P2_U2844) );
  INV_X1 U14241 ( .A(n12209), .ZN(P3_U2836) );
  NAND4_X1 U14242 ( .A1(n15350), .A2(n21430), .A3(n14001), .A4(n14000), .ZN(
        U214) );
  INV_X1 U14243 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11152) );
  NOR2_X4 U14244 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14676) );
  AND2_X4 U14245 ( .A1(n14676), .A2(n14599), .ZN(n12463) );
  AOI22_X1 U14246 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14247 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10958) );
  AND3_X4 U14248 ( .A1(n10952), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U14249 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10957) );
  AND3_X4 U14250 ( .A1(n10954), .A2(n10953), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12467) );
  AND2_X4 U14251 ( .A1(n10955), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12319) );
  AOI22_X1 U14252 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U14253 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10960) );
  NAND2_X1 U14254 ( .A1(n10960), .A2(n11006), .ZN(n10967) );
  AOI22_X1 U14255 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U14256 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U14257 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10961) );
  NAND4_X1 U14258 ( .A1(n10964), .A2(n10963), .A3(n10962), .A4(n10961), .ZN(
        n10965) );
  NAND2_X1 U14259 ( .A1(n10965), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10966) );
  AOI22_X1 U14260 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U14261 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U14262 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U14263 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10968) );
  NAND4_X1 U14264 ( .A1(n10971), .A2(n10970), .A3(n10969), .A4(n10968), .ZN(
        n10977) );
  AOI22_X1 U14265 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U14266 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14267 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10972) );
  NAND4_X1 U14268 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10976) );
  AOI22_X1 U14269 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U14270 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U14271 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10978) );
  NAND4_X1 U14272 ( .A1(n10981), .A2(n10980), .A3(n10979), .A4(n10978), .ZN(
        n10982) );
  NAND2_X1 U14273 ( .A1(n10982), .A2(n11006), .ZN(n10989) );
  AOI22_X1 U14274 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U14275 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14276 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U14277 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10983) );
  NAND4_X1 U14278 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n10987) );
  NAND2_X1 U14279 ( .A1(n10987), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10988) );
  AOI22_X1 U14280 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U14281 ( .A1(n9699), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9708), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U14282 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14283 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10990) );
  NAND4_X1 U14284 ( .A1(n10993), .A2(n10992), .A3(n10991), .A4(n10990), .ZN(
        n10994) );
  NAND2_X1 U14285 ( .A1(n10994), .A2(n11006), .ZN(n11001) );
  AOI22_X1 U14286 ( .A1(n9700), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14287 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U14288 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10996) );
  NAND4_X1 U14289 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n10999) );
  NAND2_X1 U14290 ( .A1(n10999), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11000) );
  NAND2_X2 U14291 ( .A1(n11081), .A2(n11064), .ZN(n11099) );
  AOI22_X1 U14292 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14293 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14294 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14295 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11002) );
  NAND4_X1 U14296 ( .A1(n11005), .A2(n11004), .A3(n11003), .A4(n11002), .ZN(
        n11007) );
  NAND2_X1 U14297 ( .A1(n11007), .A2(n11006), .ZN(n11014) );
  AOI22_X1 U14298 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12463), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U14299 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14300 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14301 ( .A1(n11044), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11008) );
  NAND4_X1 U14302 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11012) );
  NAND2_X1 U14303 ( .A1(n11012), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11013) );
  INV_X1 U14304 ( .A(n11062), .ZN(n11015) );
  AOI22_X1 U14305 ( .A1(n9699), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9709), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14306 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14307 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14308 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11016) );
  NAND4_X1 U14309 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11020) );
  AOI22_X1 U14310 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n9700), .ZN(n11024) );
  AOI22_X1 U14311 ( .A1(n9705), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14312 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14313 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11021) );
  NAND4_X1 U14314 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11025) );
  NAND2_X1 U14315 ( .A1(n11025), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11026) );
  AND2_X1 U14316 ( .A1(n11836), .A2(n11064), .ZN(n11070) );
  NAND2_X1 U14317 ( .A1(n11028), .A2(n19869), .ZN(n11029) );
  AOI22_X1 U14318 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9705), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14319 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14320 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U14321 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14322 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14323 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14324 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14325 ( .A1(n9706), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14326 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14327 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U14328 ( .A1(n12463), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U14329 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U14330 ( .A1(n11046), .A2(n11045), .ZN(n11050) );
  AOI22_X1 U14331 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14332 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U14333 ( .A1(n11048), .A2(n11047), .ZN(n11049) );
  NOR2_X1 U14334 ( .A1(n11050), .A2(n11049), .ZN(n11051) );
  NAND2_X1 U14335 ( .A1(n11051), .A2(n11006), .ZN(n11052) );
  AND2_X4 U14336 ( .A1(n11053), .A2(n11052), .ZN(n11385) );
  NOR2_X1 U14337 ( .A1(n11385), .A2(n14457), .ZN(n11054) );
  INV_X1 U14338 ( .A(n14811), .ZN(n11056) );
  NAND2_X1 U14339 ( .A1(n11056), .A2(n10945), .ZN(n11409) );
  NAND2_X1 U14340 ( .A1(n11409), .A2(n11057), .ZN(n11060) );
  NOR2_X1 U14341 ( .A1(n11836), .A2(n11064), .ZN(n11058) );
  AND2_X2 U14342 ( .A1(n11385), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11607) );
  NAND2_X1 U14343 ( .A1(n11099), .A2(n11635), .ZN(n11630) );
  AND2_X1 U14344 ( .A1(n11630), .A2(n14813), .ZN(n11067) );
  INV_X1 U14345 ( .A(n11632), .ZN(n11066) );
  NAND2_X1 U14346 ( .A1(n11067), .A2(n11639), .ZN(n11826) );
  NAND2_X1 U14347 ( .A1(n11826), .A2(n11075), .ZN(n11069) );
  INV_X1 U14348 ( .A(n11075), .ZN(n11082) );
  NAND2_X1 U14349 ( .A1(n11069), .A2(n11068), .ZN(n11104) );
  NAND2_X1 U14350 ( .A1(n14457), .A2(n11127), .ZN(n11118) );
  NOR2_X1 U14351 ( .A1(n14811), .A2(n11064), .ZN(n11076) );
  AND2_X4 U14352 ( .A1(n11079), .A2(n11115), .ZN(n12503) );
  AND2_X1 U14353 ( .A1(n14813), .A2(n11635), .ZN(n11097) );
  NAND2_X1 U14354 ( .A1(n15939), .A2(n11097), .ZN(n11821) );
  INV_X1 U14355 ( .A(n11821), .ZN(n11085) );
  NAND3_X1 U14356 ( .A1(n9698), .A2(n11602), .A3(n12213), .ZN(n11100) );
  NAND3_X1 U14357 ( .A1(n11082), .A2(n19869), .A3(n11087), .ZN(n11083) );
  NOR2_X1 U14358 ( .A1(n11100), .A2(n11083), .ZN(n11084) );
  AOI22_X1 U14359 ( .A1(n12503), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n11085), .B2(
        n11084), .ZN(n11095) );
  INV_X1 U14360 ( .A(n11629), .ZN(n11086) );
  NAND2_X1 U14361 ( .A1(n11086), .A2(n11087), .ZN(n11090) );
  INV_X1 U14362 ( .A(n11860), .ZN(n11088) );
  AOI22_X1 U14363 ( .A1(n11088), .A2(n11087), .B1(P2_STATE2_REG_1__SCAN_IN), 
        .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11089) );
  AND2_X1 U14364 ( .A1(n11090), .A2(n11089), .ZN(n11094) );
  INV_X1 U14365 ( .A(n11091), .ZN(n11092) );
  NAND2_X1 U14366 ( .A1(n11092), .A2(n11650), .ZN(n11103) );
  NAND2_X1 U14367 ( .A1(n13754), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11093) );
  INV_X1 U14368 ( .A(n11096), .ZN(n11098) );
  NAND3_X1 U14369 ( .A1(n11098), .A2(n11097), .A3(n15939), .ZN(n11101) );
  NAND2_X1 U14370 ( .A1(n11862), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11120) );
  NAND3_X1 U14371 ( .A1(n11120), .A2(n11103), .A3(n11102), .ZN(n11125) );
  INV_X1 U14372 ( .A(n11104), .ZN(n11107) );
  NAND2_X1 U14373 ( .A1(n11105), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11106) );
  NOR2_X1 U14374 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  AOI22_X1 U14375 ( .A1(n12503), .A2(P2_EBX_REG_0__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11109) );
  INV_X1 U14376 ( .A(n11109), .ZN(n11112) );
  NAND2_X1 U14377 ( .A1(n13754), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11110) );
  NOR2_X1 U14378 ( .A1(n11112), .A2(n11111), .ZN(n11113) );
  INV_X1 U14379 ( .A(n11115), .ZN(n11116) );
  NOR2_X1 U14380 ( .A1(n11116), .A2(n11096), .ZN(n11117) );
  NAND2_X1 U14381 ( .A1(n10618), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14382 ( .A1(n14457), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11122) );
  INV_X1 U14383 ( .A(n11133), .ZN(n11124) );
  INV_X1 U14384 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U14385 ( .A1(n12503), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U14386 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11128) );
  AOI21_X2 U14387 ( .B1(n11126), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11131), .ZN(n11147) );
  INV_X1 U14388 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n16705) );
  NAND2_X1 U14389 ( .A1(n12503), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14390 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11135) );
  OAI211_X1 U14391 ( .C1(n11876), .C2(n16705), .A(n11136), .B(n11135), .ZN(
        n11137) );
  XNOR2_X1 U14392 ( .A(n11532), .B(n11138), .ZN(n11139) );
  INV_X1 U14393 ( .A(n11173), .ZN(n16704) );
  BUF_X1 U14394 ( .A(n11140), .Z(n11141) );
  INV_X1 U14395 ( .A(n11157), .ZN(n11144) );
  OR2_X1 U14396 ( .A1(n11141), .A2(n11144), .ZN(n11179) );
  INV_X1 U14397 ( .A(n11179), .ZN(n11145) );
  BUF_X4 U14398 ( .A(n11149), .Z(n12210) );
  INV_X1 U14399 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11151) );
  BUF_X1 U14400 ( .A(n11153), .Z(n11154) );
  INV_X1 U14401 ( .A(n11155), .ZN(n11156) );
  INV_X1 U14402 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11161) );
  NAND3_X1 U14403 ( .A1(n11159), .A2(n12210), .A3(n11158), .ZN(n19997) );
  INV_X1 U14404 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11160) );
  OAI22_X1 U14405 ( .A1(n11323), .A2(n11161), .B1(n19997), .B2(n11160), .ZN(
        n11162) );
  NOR2_X1 U14406 ( .A1(n11163), .A2(n11162), .ZN(n11177) );
  INV_X1 U14407 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11167) );
  INV_X1 U14408 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11165) );
  INV_X1 U14409 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11171) );
  INV_X1 U14410 ( .A(n17184), .ZN(n11168) );
  NOR2_X1 U14411 ( .A1(n17184), .A2(n11154), .ZN(n11172) );
  NAND2_X1 U14412 ( .A1(n11173), .A2(n11172), .ZN(n11181) );
  INV_X1 U14413 ( .A(n11181), .ZN(n11182) );
  NOR2_X1 U14414 ( .A1(n9703), .A2(n11154), .ZN(n11184) );
  AOI22_X1 U14415 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11244), .B1(
        n11238), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U14416 ( .A1(n11186), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14601) );
  INV_X1 U14417 ( .A(n14601), .ZN(n11190) );
  AOI22_X1 U14418 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11187) );
  AND2_X2 U14419 ( .A1(n12466), .A2(n11006), .ZN(n11251) );
  AOI22_X1 U14420 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n11251), .ZN(n11194) );
  NAND2_X1 U14421 ( .A1(n11189), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11411) );
  AND2_X1 U14422 ( .A1(n12319), .A2(n11006), .ZN(n11713) );
  AOI22_X1 U14423 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n11713), .ZN(n11193) );
  AOI22_X1 U14424 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12330), .B1(
        n11358), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14425 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11355), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U14426 ( .A1(n11676), .A2(n11650), .ZN(n11195) );
  INV_X1 U14427 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17050) );
  INV_X1 U14428 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11196) );
  INV_X1 U14429 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11199) );
  INV_X1 U14430 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11198) );
  OAI22_X1 U14431 ( .A1(n11199), .A2(n20024), .B1(n19902), .B2(n11198), .ZN(
        n11202) );
  INV_X1 U14432 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11200) );
  NOR2_X1 U14433 ( .A1(n11202), .A2(n11201), .ZN(n11215) );
  INV_X1 U14434 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11204) );
  INV_X1 U14435 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11203) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11207) );
  INV_X1 U14437 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11206) );
  OAI22_X1 U14438 ( .A1(n11207), .A2(n20391), .B1(n11205), .B2(n11206), .ZN(
        n11208) );
  NOR2_X1 U14439 ( .A1(n11209), .A2(n11208), .ZN(n11214) );
  INV_X1 U14440 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11211) );
  OAI211_X1 U14441 ( .C1(n11289), .C2(n11211), .A(n14347), .B(n11210), .ZN(
        n11212) );
  AOI22_X1 U14442 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11217), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14443 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14444 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11713), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14445 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14446 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14447 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14448 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14449 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11223) );
  AND2_X1 U14450 ( .A1(n11653), .A2(n11650), .ZN(n14350) );
  AOI22_X1 U14451 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11250), .B1(
        n11217), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14452 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11358), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14453 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12330), .B1(
        n11713), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14454 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11251), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14455 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11237) );
  AOI22_X1 U14456 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11306), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14457 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11245), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14458 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14459 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11232) );
  NAND4_X1 U14460 ( .A1(n11235), .A2(n11234), .A3(n11233), .A4(n11232), .ZN(
        n11236) );
  NAND2_X1 U14461 ( .A1(n14350), .A2(n11662), .ZN(n11276) );
  INV_X1 U14462 ( .A(n11306), .ZN(n11242) );
  INV_X1 U14463 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11241) );
  INV_X1 U14464 ( .A(n11238), .ZN(n11240) );
  INV_X1 U14465 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11239) );
  OAI22_X1 U14466 ( .A1(n11242), .A2(n11241), .B1(n11240), .B2(n11239), .ZN(
        n11243) );
  INV_X1 U14467 ( .A(n11243), .ZN(n11249) );
  AOI22_X1 U14468 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11248) );
  INV_X2 U14469 ( .A(n14596), .ZN(n12337) );
  AOI22_X1 U14470 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14471 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11358), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11246) );
  NAND4_X1 U14472 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11257) );
  AOI22_X1 U14473 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11251), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14474 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14475 ( .A1(n12294), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14476 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11252) );
  NAND4_X1 U14477 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n11256) );
  OR2_X2 U14478 ( .A1(n11257), .A2(n11256), .ZN(n11386) );
  INV_X1 U14479 ( .A(n11386), .ZN(n11275) );
  NAND2_X1 U14480 ( .A1(n11276), .A2(n11275), .ZN(n11258) );
  AOI22_X1 U14481 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11217), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14482 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11238), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14483 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14484 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11259) );
  NAND4_X1 U14485 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(
        n11268) );
  AOI22_X1 U14486 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14487 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14488 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14489 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11263) );
  NAND4_X1 U14490 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(
        n11267) );
  INV_X1 U14491 ( .A(n11684), .ZN(n11282) );
  INV_X1 U14492 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17189) );
  NOR2_X1 U14493 ( .A1(n14350), .A2(n17189), .ZN(n11273) );
  INV_X1 U14494 ( .A(n11273), .ZN(n14352) );
  XNOR2_X1 U14495 ( .A(n11653), .B(n11662), .ZN(n11272) );
  OR2_X1 U14496 ( .A1(n14352), .A2(n11272), .ZN(n11274) );
  XNOR2_X1 U14497 ( .A(n11273), .B(n11272), .ZN(n14218) );
  NAND2_X1 U14498 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14218), .ZN(
        n14219) );
  NAND2_X1 U14499 ( .A1(n11274), .A2(n14219), .ZN(n11277) );
  XOR2_X1 U14500 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11277), .Z(
        n14951) );
  XNOR2_X1 U14501 ( .A(n11276), .B(n11275), .ZN(n14950) );
  NAND2_X1 U14502 ( .A1(n14951), .A2(n14950), .ZN(n11279) );
  NAND2_X1 U14503 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11277), .ZN(
        n11278) );
  NAND2_X1 U14504 ( .A1(n11279), .A2(n11278), .ZN(n11280) );
  INV_X1 U14505 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16985) );
  XNOR2_X1 U14506 ( .A(n11280), .B(n16985), .ZN(n16711) );
  NAND2_X1 U14507 ( .A1(n11280), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11281) );
  INV_X1 U14508 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11285) );
  INV_X1 U14509 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11284) );
  OAI22_X1 U14510 ( .A1(n11285), .A2(n11283), .B1(n19902), .B2(n11284), .ZN(
        n11288) );
  INV_X1 U14511 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11287) );
  INV_X1 U14512 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11286) );
  INV_X1 U14513 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11291) );
  INV_X1 U14514 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11290) );
  OAI22_X1 U14515 ( .A1(n11291), .A2(n20202), .B1(n11289), .B2(n11290), .ZN(
        n11292) );
  INV_X1 U14516 ( .A(n11292), .ZN(n11294) );
  NAND2_X1 U14517 ( .A1(n20122), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11293) );
  INV_X1 U14518 ( .A(n20024), .ZN(n20027) );
  INV_X1 U14519 ( .A(n11323), .ZN(n20059) );
  AOI22_X1 U14520 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20027), .B1(
        n20059), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11301) );
  INV_X1 U14521 ( .A(n20391), .ZN(n11295) );
  INV_X1 U14522 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11296) );
  INV_X1 U14523 ( .A(n11297), .ZN(n11300) );
  INV_X1 U14524 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14732) );
  INV_X1 U14525 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14526 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11217), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14527 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14528 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11713), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14529 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11302) );
  NAND4_X1 U14530 ( .A1(n11305), .A2(n11304), .A3(n11303), .A4(n11302), .ZN(
        n11312) );
  AOI22_X1 U14531 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14532 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14533 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14534 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U14535 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11311) );
  INV_X1 U14536 ( .A(n11688), .ZN(n11313) );
  NAND2_X1 U14537 ( .A1(n11313), .A2(n11650), .ZN(n11314) );
  INV_X1 U14538 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16966) );
  INV_X1 U14539 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n21603) );
  INV_X1 U14540 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11317) );
  INV_X1 U14541 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11316) );
  INV_X1 U14542 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11320) );
  INV_X1 U14543 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11319) );
  OAI22_X1 U14544 ( .A1(n11320), .A2(n11283), .B1(n20024), .B2(n11319), .ZN(
        n11325) );
  INV_X1 U14545 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11322) );
  INV_X1 U14546 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11321) );
  OAI22_X1 U14547 ( .A1(n11323), .A2(n11322), .B1(n19997), .B2(n11321), .ZN(
        n11324) );
  NOR2_X1 U14548 ( .A1(n11325), .A2(n11324), .ZN(n11329) );
  INV_X1 U14549 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11327) );
  INV_X1 U14550 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11326) );
  INV_X1 U14551 ( .A(n11289), .ZN(n20346) );
  AOI22_X1 U14552 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11217), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14553 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14554 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14555 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11330) );
  NAND4_X1 U14556 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11339) );
  AOI22_X1 U14557 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14558 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14559 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14560 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U14561 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  NAND2_X1 U14562 ( .A1(n11428), .A2(n11650), .ZN(n11340) );
  NAND2_X1 U14563 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U14564 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U14565 ( .A1(n9712), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14566 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11347) );
  NAND2_X1 U14567 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11354) );
  NAND2_X1 U14568 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11353) );
  NAND2_X1 U14569 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14570 ( .A1(n12337), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14571 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11366) );
  INV_X1 U14572 ( .A(n11355), .ZN(n11357) );
  INV_X1 U14573 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11356) );
  OR2_X1 U14574 ( .A1(n11357), .A2(n11356), .ZN(n11365) );
  INV_X1 U14575 ( .A(n11358), .ZN(n11360) );
  INV_X1 U14576 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11359) );
  OR2_X1 U14577 ( .A1(n11360), .A2(n11359), .ZN(n11364) );
  INV_X1 U14578 ( .A(n11713), .ZN(n11362) );
  INV_X1 U14579 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11361) );
  OR2_X1 U14580 ( .A1(n11362), .A2(n11361), .ZN(n11363) );
  NAND2_X1 U14581 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14582 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11372) );
  INV_X1 U14583 ( .A(n11367), .ZN(n11369) );
  INV_X1 U14584 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U14585 ( .A1(n12336), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11370) );
  AND4_X2 U14586 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n9808), .ZN(
        n11378) );
  INV_X1 U14587 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16937) );
  NAND4_X1 U14588 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11379) );
  NAND2_X1 U14589 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16839) );
  NOR2_X1 U14590 ( .A1(n11379), .A2(n16839), .ZN(n16811) );
  INV_X1 U14591 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16828) );
  INV_X1 U14592 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16825) );
  INV_X1 U14593 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16779) );
  NAND2_X1 U14594 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16812) );
  INV_X1 U14595 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11381) );
  NOR2_X1 U14596 ( .A1(n16812), .A2(n11381), .ZN(n11382) );
  NAND2_X1 U14597 ( .A1(n16811), .A2(n11382), .ZN(n16790) );
  INV_X1 U14598 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16533) );
  OR2_X1 U14599 ( .A1(n16790), .A2(n16533), .ZN(n11855) );
  NAND2_X1 U14600 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11383) );
  NOR2_X1 U14601 ( .A1(n11855), .A2(n11383), .ZN(n13599) );
  INV_X1 U14602 ( .A(n11387), .ZN(n11413) );
  NAND2_X1 U14603 ( .A1(n10954), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14604 ( .A1(n11413), .A2(n11384), .ZN(n11605) );
  INV_X1 U14605 ( .A(n11605), .ZN(n11600) );
  MUX2_X1 U14606 ( .A(n11653), .B(n11600), .S(n11402), .Z(n11463) );
  NAND2_X1 U14607 ( .A1(n11463), .A2(n11604), .ZN(n11392) );
  NAND2_X1 U14608 ( .A1(n11617), .A2(n11386), .ZN(n11391) );
  NAND2_X1 U14609 ( .A1(n11604), .A2(n11387), .ZN(n11389) );
  NAND2_X1 U14610 ( .A1(n14690), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14611 ( .A1(n11389), .A2(n11388), .ZN(n11394) );
  INV_X1 U14612 ( .A(n11393), .ZN(n11390) );
  XNOR2_X1 U14613 ( .A(n11394), .B(n11390), .ZN(n11598) );
  NAND2_X1 U14614 ( .A1(n11402), .A2(n11598), .ZN(n11611) );
  NAND2_X1 U14615 ( .A1(n11392), .A2(n11425), .ZN(n11403) );
  NAND2_X1 U14616 ( .A1(n11394), .A2(n11393), .ZN(n11396) );
  NAND2_X1 U14617 ( .A1(n20542), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11395) );
  NAND2_X1 U14618 ( .A1(n11399), .A2(n11398), .ZN(n11401) );
  NAND2_X1 U14619 ( .A1(n20533), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11400) );
  NAND2_X1 U14620 ( .A1(n11401), .A2(n11400), .ZN(n11405) );
  MUX2_X1 U14621 ( .A(n11684), .B(n11615), .S(n11402), .Z(n11618) );
  NAND3_X1 U14622 ( .A1(n11403), .A2(n11422), .A3(n11618), .ZN(n11408) );
  NOR2_X1 U14623 ( .A1(n14714), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14624 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14714), .ZN(
        n11406) );
  AND2_X1 U14625 ( .A1(n11408), .A2(n11623), .ZN(n20550) );
  INV_X1 U14626 ( .A(n11409), .ZN(n11410) );
  AND2_X1 U14627 ( .A1(n11410), .A2(n19869), .ZN(n14709) );
  AND2_X1 U14628 ( .A1(n11650), .A2(n11385), .ZN(n11633) );
  NAND2_X1 U14629 ( .A1(n20550), .A2(n20545), .ZN(n11648) );
  AND2_X1 U14630 ( .A1(n14601), .A2(n14714), .ZN(n14346) );
  NAND2_X1 U14631 ( .A1(n11411), .A2(n14346), .ZN(n11412) );
  INV_X1 U14632 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n14459) );
  NAND2_X1 U14633 ( .A1(n11412), .A2(n14459), .ZN(n17000) );
  XNOR2_X1 U14634 ( .A(n11604), .B(n11413), .ZN(n11599) );
  NAND2_X1 U14635 ( .A1(n11415), .A2(n11599), .ZN(n11414) );
  NAND2_X1 U14636 ( .A1(n11414), .A2(n11623), .ZN(n14702) );
  INV_X1 U14637 ( .A(n11415), .ZN(n11416) );
  NOR2_X1 U14638 ( .A1(n11416), .A2(n11605), .ZN(n11417) );
  NOR2_X1 U14639 ( .A1(n14702), .A2(n11417), .ZN(n11418) );
  MUX2_X1 U14640 ( .A(n17000), .B(n11418), .S(n11127), .Z(n20547) );
  AND2_X1 U14641 ( .A1(n14709), .A2(n11617), .ZN(n20546) );
  NAND2_X1 U14642 ( .A1(n20547), .A2(n20546), .ZN(n11419) );
  NAND2_X1 U14643 ( .A1(n11648), .A2(n11419), .ZN(n11420) );
  INV_X1 U14644 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11421) );
  MUX2_X1 U14645 ( .A(n11422), .B(n11421), .S(n19879), .Z(n11457) );
  INV_X1 U14646 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11423) );
  NOR2_X1 U14647 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11426) );
  MUX2_X1 U14648 ( .A(n11662), .B(n11426), .S(n19879), .Z(n11466) );
  NAND2_X1 U14649 ( .A1(n11462), .A2(n11466), .ZN(n11461) );
  INV_X1 U14650 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11427) );
  MUX2_X1 U14651 ( .A(n11688), .B(n11427), .S(n19879), .Z(n11454) );
  MUX2_X1 U14652 ( .A(n11428), .B(P2_EBX_REG_6__SCAN_IN), .S(n19879), .Z(
        n11432) );
  NAND2_X1 U14653 ( .A1(n11456), .A2(n11432), .ZN(n11433) );
  NAND2_X1 U14654 ( .A1(n11437), .A2(n11433), .ZN(n16214) );
  INV_X1 U14655 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11434) );
  MUX2_X1 U14656 ( .A(n11434), .B(n13641), .S(n13593), .Z(n11436) );
  NAND2_X1 U14657 ( .A1(n19879), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11439) );
  XNOR2_X1 U14658 ( .A(n11438), .B(n11439), .ZN(n16181) );
  NAND2_X1 U14659 ( .A1(n16181), .A2(n11435), .ZN(n16638) );
  XNOR2_X1 U14660 ( .A(n11437), .B(n11436), .ZN(n11443) );
  NAND2_X1 U14661 ( .A1(n11443), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16650) );
  AND2_X1 U14662 ( .A1(n16638), .A2(n16650), .ZN(n16623) );
  NAND2_X1 U14663 ( .A1(n19879), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11440) );
  XNOR2_X1 U14664 ( .A(n11444), .B(n11440), .ZN(n16172) );
  NAND2_X1 U14665 ( .A1(n16172), .A2(n13750), .ZN(n11441) );
  INV_X1 U14666 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16913) );
  NAND2_X1 U14667 ( .A1(n11441), .A2(n16913), .ZN(n16626) );
  NAND2_X1 U14668 ( .A1(n16181), .A2(n13750), .ZN(n11442) );
  INV_X1 U14669 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16926) );
  NAND2_X1 U14670 ( .A1(n11442), .A2(n16926), .ZN(n16639) );
  INV_X1 U14671 ( .A(n11443), .ZN(n16202) );
  NAND2_X1 U14672 ( .A1(n16202), .A2(n16937), .ZN(n16651) );
  AND2_X1 U14673 ( .A1(n16639), .A2(n16651), .ZN(n16624) );
  AND2_X1 U14674 ( .A1(n16626), .A2(n16624), .ZN(n16609) );
  NOR2_X1 U14675 ( .A1(n13593), .A2(n16166), .ZN(n11447) );
  NOR2_X4 U14676 ( .A1(n11438), .A2(n19879), .ZN(n13576) );
  AOI21_X1 U14677 ( .B1(n11448), .B2(n11447), .A(n13576), .ZN(n11449) );
  NAND2_X1 U14678 ( .A1(n11449), .A2(n14019), .ZN(n16167) );
  OR2_X1 U14679 ( .A1(n16167), .A2(n11378), .ZN(n11450) );
  INV_X1 U14680 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16602) );
  NAND2_X1 U14681 ( .A1(n11450), .A2(n16602), .ZN(n16613) );
  NAND2_X1 U14682 ( .A1(n13750), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11451) );
  OR2_X1 U14683 ( .A1(n16167), .A2(n11451), .ZN(n16612) );
  AND2_X1 U14684 ( .A1(n13641), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11452) );
  NAND2_X1 U14685 ( .A1(n16172), .A2(n11452), .ZN(n16625) );
  INV_X1 U14686 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14687 ( .A1(n9874), .A2(n10893), .ZN(n11455) );
  NAND2_X1 U14688 ( .A1(n11456), .A2(n11455), .ZN(n16224) );
  INV_X1 U14689 ( .A(n11457), .ZN(n11458) );
  NAND2_X1 U14690 ( .A1(n11458), .A2(n11461), .ZN(n11460) );
  NAND2_X1 U14691 ( .A1(n11460), .A2(n11459), .ZN(n16237) );
  OAI21_X1 U14692 ( .B1(n11462), .B2(n11466), .A(n11461), .ZN(n11469) );
  XNOR2_X1 U14693 ( .A(n11469), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14954) );
  MUX2_X1 U14694 ( .A(n11463), .B(P2_EBX_REG_0__SCAN_IN), .S(n19879), .Z(
        n16257) );
  NAND2_X1 U14695 ( .A1(n16257), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14354) );
  INV_X1 U14696 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14293) );
  NAND2_X1 U14697 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n11464) );
  NOR2_X1 U14698 ( .A1(n13593), .A2(n11464), .ZN(n11465) );
  NOR2_X1 U14699 ( .A1(n11466), .A2(n11465), .ZN(n19808) );
  NAND2_X1 U14700 ( .A1(n19808), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11468) );
  INV_X1 U14701 ( .A(n19808), .ZN(n11467) );
  AOI22_X1 U14702 ( .A1(n14354), .A2(n11468), .B1(n17017), .B2(n11467), .ZN(
        n14953) );
  NAND2_X1 U14703 ( .A1(n14954), .A2(n14953), .ZN(n14952) );
  INV_X1 U14704 ( .A(n11469), .ZN(n16247) );
  NAND2_X1 U14705 ( .A1(n16247), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11470) );
  NAND2_X1 U14706 ( .A1(n14952), .A2(n11470), .ZN(n16681) );
  NAND2_X1 U14707 ( .A1(n11459), .A2(n11471), .ZN(n11472) );
  NAND2_X1 U14708 ( .A1(n9874), .A2(n11472), .ZN(n19792) );
  NAND2_X1 U14709 ( .A1(n19792), .A2(n10042), .ZN(n11475) );
  OAI21_X1 U14710 ( .B1(n16681), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11475), .ZN(n11473) );
  INV_X1 U14711 ( .A(n11473), .ZN(n11474) );
  NAND3_X1 U14712 ( .A1(n16681), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n11475), .ZN(n11478) );
  INV_X1 U14713 ( .A(n19792), .ZN(n11476) );
  NAND2_X1 U14714 ( .A1(n11476), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11477) );
  AND2_X1 U14715 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  NAND2_X1 U14716 ( .A1(n16224), .A2(n16966), .ZN(n16606) );
  AND2_X1 U14717 ( .A1(n11481), .A2(n16606), .ZN(n11482) );
  OR2_X1 U14718 ( .A1(n14018), .A2(n11378), .ZN(n16595) );
  NAND2_X1 U14719 ( .A1(n19879), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11488) );
  INV_X1 U14720 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14721 ( .A1(n11491), .A2(n11486), .ZN(n11487) );
  NAND2_X1 U14722 ( .A1(n11500), .A2(n11487), .ZN(n11493) );
  INV_X1 U14723 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16857) );
  OAI21_X1 U14724 ( .B1(n11493), .B2(n11378), .A(n16857), .ZN(n16574) );
  NAND2_X1 U14725 ( .A1(n11489), .A2(n10904), .ZN(n11490) );
  NAND2_X1 U14726 ( .A1(n11491), .A2(n11490), .ZN(n16154) );
  OR2_X1 U14727 ( .A1(n16154), .A2(n11378), .ZN(n11492) );
  INV_X1 U14728 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16875) );
  NAND2_X1 U14729 ( .A1(n11492), .A2(n16875), .ZN(n16586) );
  AND2_X1 U14730 ( .A1(n16574), .A2(n16586), .ZN(n13544) );
  INV_X1 U14731 ( .A(n11493), .ZN(n16141) );
  AND2_X1 U14732 ( .A1(n13641), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U14733 ( .A1(n16141), .A2(n11494), .ZN(n16573) );
  NAND2_X1 U14734 ( .A1(n13750), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11495) );
  AND2_X1 U14735 ( .A1(n16573), .A2(n16584), .ZN(n11496) );
  NAND2_X1 U14736 ( .A1(n19879), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11499) );
  XNOR2_X1 U14737 ( .A(n11500), .B(n11499), .ZN(n16129) );
  NAND2_X1 U14738 ( .A1(n16129), .A2(n13750), .ZN(n11497) );
  INV_X1 U14739 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16561) );
  NAND2_X1 U14740 ( .A1(n11497), .A2(n16561), .ZN(n16568) );
  AND2_X1 U14741 ( .A1(n13641), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U14742 ( .A1(n16129), .A2(n11498), .ZN(n16567) );
  NAND2_X1 U14743 ( .A1(n19879), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11501) );
  INV_X1 U14744 ( .A(n11501), .ZN(n11502) );
  NAND2_X1 U14745 ( .A1(n9841), .A2(n11502), .ZN(n11503) );
  NAND2_X1 U14746 ( .A1(n11512), .A2(n11503), .ZN(n16116) );
  INV_X1 U14747 ( .A(n16553), .ZN(n11505) );
  OR2_X1 U14748 ( .A1(n16116), .A2(n11378), .ZN(n11504) );
  NAND2_X1 U14749 ( .A1(n11504), .A2(n16828), .ZN(n16554) );
  OR2_X1 U14750 ( .A1(n11512), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11510) );
  NAND3_X1 U14751 ( .A1(n11512), .A2(n19879), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n11506) );
  NAND3_X1 U14752 ( .A1(n11510), .A2(n13539), .A3(n11506), .ZN(n19771) );
  OAI21_X1 U14753 ( .B1(n19771), .B2(n11378), .A(n16825), .ZN(n11508) );
  NAND2_X1 U14754 ( .A1(n13750), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14755 ( .A1(n11508), .A2(n13554), .ZN(n13543) );
  INV_X1 U14756 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n21689) );
  NOR2_X1 U14757 ( .A1(n13593), .A2(n21689), .ZN(n11509) );
  NOR2_X1 U14758 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n11511) );
  AOI21_X1 U14759 ( .B1(n19760), .B2(n13750), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11515) );
  INV_X1 U14760 ( .A(n19760), .ZN(n11514) );
  NAND2_X1 U14761 ( .A1(n13750), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11513) );
  NOR2_X1 U14762 ( .A1(n11514), .A2(n11513), .ZN(n13557) );
  OR2_X1 U14763 ( .A1(n11515), .A2(n13557), .ZN(n16540) );
  INV_X1 U14764 ( .A(n11515), .ZN(n13546) );
  INV_X1 U14765 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U14766 ( .A1(n11516), .A2(n16098), .ZN(n11520) );
  NAND3_X1 U14767 ( .A1(n11520), .A2(n19879), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n11519) );
  OAI21_X1 U14768 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n19879), .ZN(n11517) );
  NAND2_X1 U14769 ( .A1(n11519), .A2(n11869), .ZN(n16090) );
  AND2_X1 U14770 ( .A1(n13641), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11522) );
  NAND2_X1 U14771 ( .A1(n16104), .A2(n11522), .ZN(n16531) );
  AOI21_X1 U14772 ( .B1(n16104), .B2(n13750), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13549) );
  NAND2_X1 U14773 ( .A1(n19879), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11526) );
  XNOR2_X1 U14774 ( .A(n11869), .B(n11526), .ZN(n16069) );
  AND2_X1 U14775 ( .A1(n13641), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11527) );
  AOI21_X1 U14776 ( .B1(n16069), .B2(n13750), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11868) );
  INV_X1 U14777 ( .A(n11868), .ZN(n13550) );
  INV_X1 U14778 ( .A(n11528), .ZN(n13558) );
  NAND2_X1 U14779 ( .A1(n13550), .A2(n13558), .ZN(n11529) );
  INV_X1 U14780 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n16691) );
  NAND2_X1 U14781 ( .A1(n12503), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14782 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11534) );
  OAI211_X1 U14783 ( .C1(n11876), .C2(n16691), .A(n11535), .B(n11534), .ZN(
        n11536) );
  AOI21_X1 U14784 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11536), .ZN(n16688) );
  INV_X1 U14785 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16223) );
  NAND2_X1 U14786 ( .A1(n12503), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11540) );
  NAND2_X1 U14787 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11539) );
  OAI211_X1 U14788 ( .C1(n11876), .C2(n16223), .A(n11540), .B(n11539), .ZN(
        n11541) );
  AOI21_X1 U14789 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11541), .ZN(n14656) );
  INV_X1 U14790 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n16211) );
  NAND2_X1 U14791 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11543) );
  AOI22_X1 U14792 ( .A1(n9694), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11542) );
  OAI211_X1 U14793 ( .C1(n13758), .C2(n16211), .A(n11543), .B(n11542), .ZN(
        n14735) );
  INV_X1 U14794 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n16654) );
  NAND2_X1 U14795 ( .A1(n12503), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11546) );
  NAND2_X1 U14796 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11545) );
  OAI211_X1 U14797 ( .C1(n11876), .C2(n16654), .A(n11546), .B(n11545), .ZN(
        n11547) );
  AOI21_X1 U14798 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11547), .ZN(n14739) );
  INV_X1 U14799 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20474) );
  NAND2_X1 U14800 ( .A1(n12503), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14801 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11549) );
  OAI211_X1 U14802 ( .C1(n11876), .C2(n20474), .A(n11550), .B(n11549), .ZN(
        n11551) );
  AOI21_X1 U14803 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11551), .ZN(n14765) );
  NAND2_X1 U14804 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11553) );
  AOI22_X1 U14805 ( .A1(n9694), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11552) );
  OAI211_X1 U14806 ( .C1(n11445), .C2(n13758), .A(n11553), .B(n11552), .ZN(
        n14790) );
  NAND2_X1 U14807 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11555) );
  AOI22_X1 U14808 ( .A1(n9694), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11554) );
  OAI211_X1 U14809 ( .C1(n16166), .C2(n13758), .A(n11555), .B(n11554), .ZN(
        n14845) );
  NAND2_X1 U14810 ( .A1(n14789), .A2(n14845), .ZN(n14022) );
  INV_X1 U14811 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14812 ( .A1(n12503), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U14813 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11556) );
  OAI211_X1 U14814 ( .C1(n11876), .C2(n11558), .A(n11557), .B(n11556), .ZN(
        n11559) );
  AOI21_X1 U14815 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11559), .ZN(n14025) );
  INV_X1 U14816 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20481) );
  NAND2_X1 U14817 ( .A1(n12503), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14818 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14819 ( .C1(n11876), .C2(n20481), .A(n11563), .B(n11562), .ZN(
        n11564) );
  AOI21_X1 U14820 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11564), .ZN(n16143) );
  INV_X1 U14821 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n16127) );
  NAND2_X1 U14822 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11566) );
  AOI22_X1 U14823 ( .A1(n9694), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11565) );
  OAI211_X1 U14824 ( .C1(n13758), .C2(n16127), .A(n11566), .B(n11565), .ZN(
        n14824) );
  NAND2_X1 U14825 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11568) );
  AOI22_X1 U14826 ( .A1(n9694), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11567) );
  OAI211_X1 U14827 ( .C1(n13758), .C2(n11569), .A(n11568), .B(n11567), .ZN(
        n14839) );
  AND2_X1 U14828 ( .A1(n14824), .A2(n14839), .ZN(n11570) );
  INV_X1 U14829 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20485) );
  NAND2_X1 U14830 ( .A1(n12503), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14831 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11571) );
  OAI211_X1 U14832 ( .C1(n11876), .C2(n20485), .A(n11572), .B(n11571), .ZN(
        n11573) );
  AOI21_X1 U14833 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11573), .ZN(n14833) );
  INV_X1 U14834 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20487) );
  NAND2_X1 U14835 ( .A1(n12503), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11576) );
  NAND2_X1 U14836 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11575) );
  OAI211_X1 U14837 ( .C1(n11876), .C2(n20487), .A(n11576), .B(n11575), .ZN(
        n11577) );
  AOI21_X1 U14838 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11577), .ZN(n16338) );
  INV_X1 U14839 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20488) );
  NAND2_X1 U14840 ( .A1(n12503), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14841 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11579) );
  OAI211_X1 U14842 ( .C1(n11876), .C2(n20488), .A(n11580), .B(n11579), .ZN(
        n11581) );
  AOI21_X1 U14843 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11581), .ZN(n16330) );
  NOR2_X2 U14844 ( .A1(n16329), .A2(n16330), .ZN(n16095) );
  NAND2_X1 U14845 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11583) );
  AOI22_X1 U14846 ( .A1(n9694), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11582) );
  OAI211_X1 U14847 ( .C1(n13758), .C2(n16098), .A(n11583), .B(n11582), .ZN(
        n16094) );
  AND2_X2 U14848 ( .A1(n16095), .A2(n16094), .ZN(n11901) );
  INV_X1 U14849 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11586) );
  NAND2_X1 U14850 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11585) );
  AOI22_X1 U14851 ( .A1(n9694), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11584) );
  OAI211_X1 U14852 ( .C1(n13758), .C2(n11586), .A(n11585), .B(n11584), .ZN(
        n11904) );
  INV_X1 U14853 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16067) );
  NAND2_X1 U14854 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11588) );
  AOI22_X1 U14855 ( .A1(n9694), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11587) );
  OAI211_X1 U14856 ( .C1(n13758), .C2(n16067), .A(n11588), .B(n11587), .ZN(
        n11589) );
  OAI21_X1 U14857 ( .B1(n11902), .B2(n11589), .A(n11880), .ZN(n16322) );
  INV_X1 U14858 ( .A(n16322), .ZN(n16073) );
  NOR2_X1 U14859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17019) );
  OR2_X1 U14860 ( .A1(n20528), .A2(n17019), .ZN(n20525) );
  NAND2_X1 U14861 ( .A1(n20525), .A2(n14457), .ZN(n11590) );
  AND2_X1 U14862 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14452) );
  INV_X1 U14863 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11592) );
  AND2_X2 U14864 ( .A1(n13681), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13683) );
  NOR2_X2 U14865 ( .A1(n13686), .A2(n21703), .ZN(n13689) );
  NAND2_X1 U14866 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11905), .ZN(
        n11894) );
  OAI21_X1 U14867 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11905), .A(
        n11894), .ZN(n16063) );
  NAND2_X1 U14868 ( .A1(n20198), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U14869 ( .A1(n14230), .A2(n13716), .ZN(n14355) );
  INV_X2 U14870 ( .A(n19788), .ZN(n16706) );
  INV_X1 U14871 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20493) );
  NOR2_X1 U14872 ( .A1(n16706), .A2(n20493), .ZN(n11857) );
  AOI21_X1 U14873 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n11857), .ZN(n11593) );
  OAI21_X1 U14874 ( .B1(n16063), .B2(n16710), .A(n11593), .ZN(n11594) );
  AOI21_X1 U14875 ( .B1(n16073), .B2(n16715), .A(n11594), .ZN(n11595) );
  NAND2_X1 U14876 ( .A1(n20454), .A2(n20464), .ZN(n20459) );
  OAI211_X1 U14877 ( .C1(n20454), .C2(n20464), .A(n19734), .B(n20459), .ZN(
        n15934) );
  NAND2_X1 U14878 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n17196) );
  AND2_X1 U14879 ( .A1(n20450), .A2(n17196), .ZN(n14335) );
  NAND2_X1 U14880 ( .A1(n11836), .A2(n14335), .ZN(n11627) );
  INV_X1 U14881 ( .A(n11598), .ZN(n11609) );
  OAI21_X1 U14882 ( .B1(n14347), .B2(n11600), .A(n11599), .ZN(n11601) );
  OAI21_X1 U14883 ( .B1(n11609), .B2(n14347), .A(n11601), .ZN(n11603) );
  NAND2_X1 U14884 ( .A1(n11603), .A2(n11602), .ZN(n11614) );
  INV_X1 U14885 ( .A(n11604), .ZN(n11606) );
  OAI21_X1 U14886 ( .B1(n11606), .B2(n11605), .A(n11617), .ZN(n11613) );
  INV_X1 U14887 ( .A(n11607), .ZN(n11608) );
  NAND2_X1 U14888 ( .A1(n11608), .A2(n14347), .ZN(n11610) );
  NAND2_X1 U14889 ( .A1(n11610), .A2(n11609), .ZN(n11612) );
  INV_X1 U14890 ( .A(n11620), .ZN(n11616) );
  NAND3_X1 U14891 ( .A1(n11620), .A2(n11619), .A3(n11618), .ZN(n11621) );
  NAND2_X1 U14892 ( .A1(n11626), .A2(n11602), .ZN(n11622) );
  NAND2_X1 U14893 ( .A1(n14699), .A2(n14347), .ZN(n14227) );
  NAND2_X1 U14894 ( .A1(n14705), .A2(n17196), .ZN(n14258) );
  NAND2_X1 U14895 ( .A1(n11628), .A2(n20450), .ZN(n11642) );
  NAND2_X1 U14896 ( .A1(n11630), .A2(n19869), .ZN(n11631) );
  NAND2_X1 U14897 ( .A1(n14345), .A2(n11631), .ZN(n11641) );
  NAND2_X1 U14898 ( .A1(n11632), .A2(n14813), .ZN(n11634) );
  NAND2_X1 U14899 ( .A1(n11634), .A2(n11633), .ZN(n11827) );
  NAND3_X1 U14900 ( .A1(n11650), .A2(n14813), .A3(n11635), .ZN(n11637) );
  NAND2_X1 U14901 ( .A1(n11385), .A2(n14813), .ZN(n11636) );
  NAND3_X1 U14902 ( .A1(n11637), .A2(n19869), .A3(n11636), .ZN(n11638) );
  AND4_X1 U14903 ( .A1(n11639), .A2(n11827), .A3(n11096), .A4(n11638), .ZN(
        n11640) );
  OAI211_X1 U14904 ( .C1(n14258), .C2(n11642), .A(n11641), .B(n11640), .ZN(
        n14337) );
  MUX2_X1 U14905 ( .A(n11643), .B(n19869), .S(n11650), .Z(n11644) );
  NOR2_X1 U14906 ( .A1(n11644), .A2(n14258), .ZN(n11645) );
  NOR2_X1 U14907 ( .A1(n14337), .A2(n11645), .ZN(n11647) );
  NAND3_X1 U14908 ( .A1(n20547), .A2(n14709), .A3(n14347), .ZN(n11646) );
  INV_X1 U14909 ( .A(n14264), .ZN(n14263) );
  NAND2_X1 U14910 ( .A1(n14263), .A2(n11808), .ZN(n11671) );
  AND2_X1 U14911 ( .A1(n11064), .A2(n20300), .ZN(n11651) );
  NAND2_X1 U14912 ( .A1(n14813), .A2(n20300), .ZN(n11655) );
  NAND2_X1 U14913 ( .A1(n20338), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16998) );
  NAND2_X1 U14914 ( .A1(n11655), .A2(n16998), .ZN(n11654) );
  INV_X1 U14915 ( .A(n11655), .ZN(n11663) );
  NOR2_X1 U14916 ( .A1(n11074), .A2(n11064), .ZN(n11656) );
  NAND2_X1 U14917 ( .A1(n9691), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11657) );
  OAI211_X1 U14918 ( .C1(n13619), .C2(n17189), .A(n20300), .B(n11657), .ZN(
        n11658) );
  INV_X1 U14919 ( .A(n11658), .ZN(n11659) );
  AOI22_X1 U14920 ( .A1(n11672), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11808), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U14921 ( .A1(n9809), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14922 ( .A1(n11661), .A2(n11660), .ZN(n11667) );
  XNOR2_X1 U14923 ( .A(n11666), .B(n11667), .ZN(n14442) );
  NAND2_X1 U14924 ( .A1(n11652), .A2(n11662), .ZN(n11665) );
  AOI22_X1 U14925 ( .A1(n14264), .A2(n11663), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11664) );
  AND2_X1 U14926 ( .A1(n11665), .A2(n11664), .ZN(n14441) );
  INV_X1 U14927 ( .A(n11667), .ZN(n11668) );
  NAND2_X1 U14928 ( .A1(n11666), .A2(n11668), .ZN(n11669) );
  NAND2_X1 U14929 ( .A1(n14444), .A2(n11669), .ZN(n11681) );
  NAND2_X1 U14930 ( .A1(n11652), .A2(n11386), .ZN(n11670) );
  OAI211_X1 U14931 ( .C1(n20300), .C2(n20542), .A(n11671), .B(n11670), .ZN(
        n11679) );
  XNOR2_X1 U14932 ( .A(n11681), .B(n11679), .ZN(n14644) );
  AOI22_X1 U14933 ( .A1(n9687), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14934 ( .A1(n13763), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11673) );
  AND2_X1 U14935 ( .A1(n11674), .A2(n11673), .ZN(n14643) );
  OAI22_X1 U14936 ( .A1(n13619), .A2(n16985), .B1(n20533), .B2(n20300), .ZN(
        n11675) );
  AOI21_X1 U14937 ( .B1(n13763), .B2(P2_REIP_REG_3__SCAN_IN), .A(n11675), .ZN(
        n11678) );
  AOI22_X1 U14938 ( .A1(n11652), .A2(n11676), .B1(n9687), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n11677) );
  AND2_X1 U14939 ( .A1(n11678), .A2(n11677), .ZN(n14749) );
  INV_X1 U14940 ( .A(n14749), .ZN(n11682) );
  INV_X1 U14941 ( .A(n11679), .ZN(n11680) );
  NAND2_X1 U14942 ( .A1(n11681), .A2(n11680), .ZN(n14748) );
  AND2_X1 U14943 ( .A1(n11682), .A2(n14748), .ZN(n11683) );
  NAND2_X1 U14944 ( .A1(n14642), .A2(n11683), .ZN(n14747) );
  AOI22_X1 U14945 ( .A1(n9687), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11687) );
  INV_X4 U14946 ( .A(n13620), .ZN(n13763) );
  NAND2_X1 U14947 ( .A1(n13763), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11686) );
  NAND2_X1 U14948 ( .A1(n11652), .A2(n11684), .ZN(n11685) );
  AND3_X1 U14949 ( .A1(n11687), .A2(n11686), .A3(n11685), .ZN(n14775) );
  AOI22_X1 U14950 ( .A1(n9687), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11690) );
  NAND2_X1 U14951 ( .A1(n11652), .A2(n11688), .ZN(n11689) );
  OAI211_X1 U14952 ( .C1(n13620), .C2(n16223), .A(n11690), .B(n11689), .ZN(
        n14772) );
  NAND2_X1 U14953 ( .A1(n11652), .A2(n11691), .ZN(n11692) );
  AOI22_X1 U14954 ( .A1(n9687), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U14955 ( .A1(n13763), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U14956 ( .A1(n11694), .A2(n11693), .ZN(n14288) );
  NAND2_X1 U14957 ( .A1(n11652), .A2(n13750), .ZN(n11695) );
  NAND2_X1 U14958 ( .A1(n14287), .A2(n11695), .ZN(n14274) );
  AOI22_X1 U14959 ( .A1(n9687), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U14960 ( .A1(n13763), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14961 ( .A1(n11697), .A2(n11696), .ZN(n14273) );
  NAND2_X1 U14962 ( .A1(n14274), .A2(n14273), .ZN(n14279) );
  AOI22_X1 U14963 ( .A1(n9687), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14964 ( .A1(n13763), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14965 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14966 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14967 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11238), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14968 ( .A1(n12336), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11698) );
  NAND4_X1 U14969 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n11707) );
  AOI22_X1 U14970 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12330), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14971 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14972 ( .A1(n12294), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11251), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14973 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U14974 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NAND2_X1 U14975 ( .A1(n11652), .A2(n14768), .ZN(n11708) );
  NAND2_X1 U14976 ( .A1(n11712), .A2(n11711), .ZN(n14254) );
  AOI22_X1 U14977 ( .A1(n9687), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U14978 ( .A1(n13763), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14979 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14980 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11358), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14981 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12330), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14982 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11251), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14983 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11723) );
  AOI22_X1 U14984 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11306), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14985 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11245), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14986 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14987 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11718) );
  NAND4_X1 U14988 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11722) );
  NAND2_X1 U14989 ( .A1(n11652), .A2(n14788), .ZN(n11724) );
  AOI22_X1 U14990 ( .A1(n9687), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11739) );
  NAND2_X1 U14991 ( .A1(n13763), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14992 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14993 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11238), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14994 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14995 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11727) );
  NAND4_X1 U14996 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11736) );
  AOI22_X1 U14997 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11251), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14998 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14999 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U15000 ( .A1(n12294), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11731) );
  NAND4_X1 U15001 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11735) );
  NAND2_X1 U15002 ( .A1(n11652), .A2(n14848), .ZN(n11737) );
  AOI22_X1 U15003 ( .A1(n9687), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U15004 ( .A1(n13763), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U15005 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U15006 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U15007 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U15008 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U15009 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11749) );
  AOI22_X1 U15010 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11306), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U15011 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11245), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U15012 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U15013 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11744) );
  NAND4_X1 U15014 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11748) );
  OR2_X1 U15015 ( .A1(n11749), .A2(n11748), .ZN(n16342) );
  NAND2_X1 U15016 ( .A1(n11652), .A2(n16342), .ZN(n11750) );
  AOI22_X1 U15017 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U15018 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U15019 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11238), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U15020 ( .A1(n12336), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11753) );
  NAND4_X1 U15021 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11762) );
  AOI22_X1 U15022 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11251), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U15023 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11245), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U15024 ( .A1(n11355), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U15025 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11757) );
  NAND4_X1 U15026 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11761) );
  NOR2_X1 U15027 ( .A1(n11762), .A2(n11761), .ZN(n16343) );
  AOI22_X1 U15028 ( .A1(n9687), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U15029 ( .A1(n13763), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11763) );
  OAI211_X1 U15030 ( .C1(n16343), .C2(n11765), .A(n11764), .B(n11763), .ZN(
        n14438) );
  NAND2_X1 U15031 ( .A1(n14439), .A2(n14438), .ZN(n14472) );
  AOI22_X1 U15032 ( .A1(n9687), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U15033 ( .A1(n13763), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U15034 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U15035 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U15036 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U15037 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11766) );
  NAND4_X1 U15038 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11775) );
  AOI22_X1 U15039 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U15040 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U15041 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U15042 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11770) );
  NAND4_X1 U15043 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11774) );
  OR2_X1 U15044 ( .A1(n11775), .A2(n11774), .ZN(n14802) );
  NAND2_X1 U15045 ( .A1(n11652), .A2(n14802), .ZN(n11776) );
  AOI22_X1 U15046 ( .A1(n9687), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U15047 ( .A1(n13763), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U15048 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U15049 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11238), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U15050 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U15051 ( .A1(n11244), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11780) );
  NAND4_X1 U15052 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11789) );
  AOI22_X1 U15053 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11245), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U15054 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U15055 ( .A1(n12294), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U15056 ( .A1(n11367), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11251), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U15057 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11788) );
  NAND2_X1 U15058 ( .A1(n11652), .A2(n14826), .ZN(n11790) );
  AOI22_X1 U15059 ( .A1(n9687), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U15060 ( .A1(n13763), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U15061 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U15062 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U15063 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U15064 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11793) );
  NAND4_X1 U15065 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11802) );
  AOI22_X1 U15066 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U15067 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U15068 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U15069 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11797) );
  NAND4_X1 U15070 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(
        n11801) );
  OR2_X1 U15071 ( .A1(n11802), .A2(n11801), .ZN(n14803) );
  NAND2_X1 U15072 ( .A1(n11652), .A2(n14803), .ZN(n11803) );
  AOI22_X1 U15073 ( .A1(n9687), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11807) );
  NAND2_X1 U15074 ( .A1(n13763), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U15075 ( .A1(n11807), .A2(n11806), .ZN(n14808) );
  NAND2_X1 U15076 ( .A1(n14809), .A2(n14808), .ZN(n14807) );
  AOI22_X1 U15077 ( .A1(n9687), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U15078 ( .A1(n13763), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11809) );
  INV_X1 U15079 ( .A(n16463), .ZN(n11811) );
  AOI22_X1 U15080 ( .A1(n9687), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U15081 ( .A1(n13763), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15082 ( .A1(n9687), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U15083 ( .A1(n13763), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11814) );
  NAND2_X1 U15084 ( .A1(n11815), .A2(n11814), .ZN(n16075) );
  AOI22_X1 U15085 ( .A1(n9687), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U15086 ( .A1(n13763), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11816) );
  NAND2_X1 U15087 ( .A1(n11817), .A2(n11816), .ZN(n11819) );
  NAND2_X1 U15088 ( .A1(n11818), .A2(n11819), .ZN(n11884) );
  OR2_X1 U15089 ( .A1(n11818), .A2(n11819), .ZN(n11820) );
  NAND2_X1 U15090 ( .A1(n11884), .A2(n11820), .ZN(n16442) );
  NAND2_X1 U15091 ( .A1(n14677), .A2(n11822), .ZN(n14597) );
  NAND2_X1 U15092 ( .A1(n11628), .A2(n11385), .ZN(n11823) );
  NAND2_X1 U15093 ( .A1(n14345), .A2(n11823), .ZN(n14708) );
  NAND2_X1 U15094 ( .A1(n14708), .A2(n14347), .ZN(n11824) );
  NAND2_X1 U15095 ( .A1(n14597), .A2(n11824), .ZN(n11825) );
  NAND2_X1 U15096 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n11843) );
  INV_X1 U15097 ( .A(n11843), .ZN(n14959) );
  AND2_X1 U15098 ( .A1(n14959), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14955) );
  NAND2_X1 U15099 ( .A1(n11826), .A2(n14347), .ZN(n14678) );
  AOI21_X1 U15100 ( .B1(n14678), .B2(n11827), .A(n11082), .ZN(n11835) );
  INV_X1 U15101 ( .A(n11840), .ZN(n12477) );
  NAND2_X1 U15102 ( .A1(n11828), .A2(n12477), .ZN(n14261) );
  INV_X1 U15103 ( .A(n11829), .ZN(n11830) );
  NAND2_X1 U15104 ( .A1(n11830), .A2(n11840), .ZN(n11831) );
  NAND2_X1 U15105 ( .A1(n11831), .A2(n15939), .ZN(n11832) );
  NAND2_X1 U15106 ( .A1(n11832), .A2(n11098), .ZN(n11833) );
  OAI211_X1 U15107 ( .C1(n19875), .C2(n15939), .A(n14261), .B(n11833), .ZN(
        n11834) );
  MUX2_X1 U15108 ( .A(n11837), .B(n11836), .S(n11385), .Z(n11838) );
  NAND2_X1 U15109 ( .A1(n14661), .A2(n11840), .ZN(n11841) );
  NAND2_X1 U15110 ( .A1(n11865), .A2(n11841), .ZN(n16806) );
  AND3_X1 U15111 ( .A1(n19869), .A2(n11650), .A3(n13593), .ZN(n11842) );
  INV_X1 U15112 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14958) );
  AND2_X1 U15113 ( .A1(n14958), .A2(n11843), .ZN(n11849) );
  NAND2_X1 U15114 ( .A1(n14956), .A2(n11849), .ZN(n14966) );
  INV_X1 U15115 ( .A(n11865), .ZN(n11844) );
  NAND2_X1 U15116 ( .A1(n11844), .A2(n16706), .ZN(n17183) );
  OAI211_X1 U15117 ( .C1(n14955), .C2(n16806), .A(n14966), .B(n17183), .ZN(
        n16984) );
  NAND2_X2 U15118 ( .A1(n16803), .A2(n16806), .ZN(n17188) );
  AND2_X1 U15119 ( .A1(n17188), .A2(n16985), .ZN(n11845) );
  AND2_X1 U15120 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16948) );
  NAND2_X1 U15121 ( .A1(n16948), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11852) );
  AND2_X1 U15122 ( .A1(n17188), .A2(n11852), .ZN(n11846) );
  NOR2_X1 U15123 ( .A1(n16937), .A2(n16926), .ZN(n11853) );
  INV_X1 U15124 ( .A(n11853), .ZN(n16922) );
  NAND2_X1 U15125 ( .A1(n17188), .A2(n16922), .ZN(n11847) );
  AND2_X1 U15126 ( .A1(n17188), .A2(n11855), .ZN(n11848) );
  NOR2_X1 U15127 ( .A1(n16844), .A2(n11848), .ZN(n16780) );
  INV_X1 U15128 ( .A(n14955), .ZN(n11850) );
  AOI21_X1 U15129 ( .B1(n16803), .B2(n11850), .A(n11849), .ZN(n11851) );
  NAND2_X1 U15130 ( .A1(n11851), .A2(n17188), .ZN(n16986) );
  NOR2_X2 U15131 ( .A1(n16974), .A2(n11852), .ZN(n16935) );
  AND2_X2 U15132 ( .A1(n16935), .A2(n11853), .ZN(n16910) );
  NOR2_X1 U15133 ( .A1(n11855), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U15134 ( .A1(n16910), .A2(n11854), .ZN(n16777) );
  NAND2_X1 U15135 ( .A1(n16780), .A2(n16777), .ZN(n11858) );
  INV_X1 U15136 ( .A(n16910), .ZN(n16884) );
  NOR4_X1 U15137 ( .A1(n16884), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16779), .A4(n11855), .ZN(n11856) );
  AOI211_X1 U15138 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n11858), .A(
        n11857), .B(n11856), .ZN(n11859) );
  OAI21_X1 U15139 ( .B1(n16442), .B2(n17180), .A(n11859), .ZN(n11866) );
  INV_X1 U15140 ( .A(n14708), .ZN(n11861) );
  NAND2_X1 U15141 ( .A1(n11861), .A2(n11860), .ZN(n14684) );
  NAND2_X1 U15142 ( .A1(n14684), .A2(n11650), .ZN(n11863) );
  INV_X1 U15143 ( .A(n11862), .ZN(n14594) );
  NAND2_X1 U15144 ( .A1(n11863), .A2(n14594), .ZN(n11864) );
  NOR2_X1 U15145 ( .A1(n11866), .A2(n9813), .ZN(n11867) );
  INV_X1 U15146 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n16316) );
  NOR2_X1 U15147 ( .A1(n13593), .A2(n16316), .ZN(n11870) );
  AOI21_X1 U15148 ( .B1(n9859), .B2(n11870), .A(n13576), .ZN(n11871) );
  AND2_X1 U15149 ( .A1(n13562), .A2(n11871), .ZN(n16055) );
  AND2_X1 U15150 ( .A1(n16055), .A2(n13641), .ZN(n11872) );
  NAND2_X1 U15151 ( .A1(n11872), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13560) );
  INV_X1 U15152 ( .A(n11872), .ZN(n11873) );
  INV_X1 U15153 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21546) );
  NAND2_X1 U15154 ( .A1(n11873), .A2(n21546), .ZN(n13551) );
  INV_X1 U15155 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20495) );
  NAND2_X1 U15156 ( .A1(n12503), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U15157 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11874) );
  OAI211_X1 U15158 ( .C1(n11876), .C2(n20495), .A(n11875), .B(n11874), .ZN(
        n11877) );
  AOI21_X1 U15159 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11877), .ZN(n11879) );
  NAND2_X1 U15160 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  INV_X1 U15161 ( .A(n13599), .ZN(n11882) );
  OR2_X1 U15162 ( .A1(n11882), .A2(n21546), .ZN(n13624) );
  AOI21_X1 U15163 ( .B1(n16910), .B2(n13599), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U15164 ( .A1(n19788), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11897) );
  OAI21_X1 U15165 ( .B1(n16754), .B2(n11883), .A(n11897), .ZN(n11892) );
  AOI22_X1 U15166 ( .A1(n9687), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11886) );
  NAND2_X1 U15167 ( .A1(n13763), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11885) );
  AND2_X1 U15168 ( .A1(n11886), .A2(n11885), .ZN(n11889) );
  INV_X1 U15169 ( .A(n11889), .ZN(n11887) );
  NAND2_X1 U15170 ( .A1(n11884), .A2(n11889), .ZN(n11890) );
  NAND2_X1 U15171 ( .A1(n16043), .A2(n11890), .ZN(n16429) );
  NOR2_X1 U15172 ( .A1(n16429), .A2(n17180), .ZN(n11891) );
  AOI211_X1 U15173 ( .C1(n16310), .C2(n16970), .A(n11892), .B(n11891), .ZN(
        n11893) );
  INV_X1 U15174 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16049) );
  NAND2_X1 U15175 ( .A1(n16049), .A2(n11894), .ZN(n11896) );
  AND2_X1 U15176 ( .A1(n11896), .A2(n13696), .ZN(n16053) );
  NAND2_X1 U15177 ( .A1(n16692), .A2(n16053), .ZN(n11898) );
  OAI211_X1 U15178 ( .C1(n16049), .C2(n16672), .A(n11898), .B(n11897), .ZN(
        n11899) );
  AOI21_X1 U15179 ( .B1(n16310), .B2(n16715), .A(n11899), .ZN(n11900) );
  INV_X1 U15180 ( .A(n11902), .ZN(n11903) );
  OAI21_X1 U15181 ( .B1(n11901), .B2(n11904), .A(n11903), .ZN(n16784) );
  AOI21_X1 U15182 ( .B1(n13693), .B2(n16082), .A(n11905), .ZN(n16085) );
  INV_X1 U15183 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n16079) );
  NOR2_X1 U15184 ( .A1(n16706), .A2(n16079), .ZN(n16776) );
  NOR2_X1 U15185 ( .A1(n16672), .A2(n16082), .ZN(n11906) );
  AOI211_X1 U15186 ( .C1(n16085), .C2(n16692), .A(n16776), .B(n11906), .ZN(
        n11907) );
  OAI21_X1 U15187 ( .B1(n16784), .B2(n16695), .A(n11907), .ZN(n11908) );
  AOI21_X1 U15188 ( .B1(n16786), .B2(n16697), .A(n11908), .ZN(n11914) );
  NAND2_X1 U15189 ( .A1(n11524), .A2(n11910), .ZN(n11911) );
  NAND2_X1 U15190 ( .A1(n16775), .A2(n11531), .ZN(n11913) );
  NAND2_X1 U15191 ( .A1(n11914), .A2(n11913), .ZN(P2_U2995) );
  INV_X2 U15192 ( .A(n11976), .ZN(n18094) );
  AOI22_X1 U15193 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12075), .ZN(n11919) );
  AOI22_X1 U15194 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11918) );
  INV_X2 U15195 ( .A(n17817), .ZN(n18095) );
  NOR2_X2 U15196 ( .A1(n11920), .A2(n11921), .ZN(n17806) );
  AOI22_X1 U15197 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U15198 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12071), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U15199 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11930) );
  AOI22_X1 U15200 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11928) );
  NOR2_X2 U15201 ( .A1(n17750), .A2(n11920), .ZN(n11998) );
  AOI22_X1 U15202 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11998), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11927) );
  INV_X2 U15203 ( .A(n9778), .ZN(n18006) );
  AOI22_X1 U15204 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15205 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11925) );
  NAND4_X1 U15206 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11929) );
  AOI22_X1 U15207 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9692), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15208 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15209 ( .A1(n17852), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11932) );
  OAI21_X1 U15210 ( .B1(n11969), .B2(n21639), .A(n11932), .ZN(n11938) );
  AOI22_X1 U15211 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11936) );
  INV_X2 U15212 ( .A(n17817), .ZN(n17807) );
  AOI22_X1 U15213 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15214 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15215 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11933) );
  NAND4_X1 U15216 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(
        n11937) );
  NOR2_X1 U15217 ( .A1(n19715), .A2(n9681), .ZN(n12179) );
  INV_X2 U15218 ( .A(n11999), .ZN(n18075) );
  AOI22_X1 U15219 ( .A1(n9702), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15220 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15221 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15222 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U15223 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11952) );
  AOI22_X1 U15224 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9693), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15225 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15226 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15227 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15228 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NAND2_X1 U15229 ( .A1(n12179), .A2(n18156), .ZN(n12158) );
  AOI22_X1 U15230 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11960) );
  INV_X2 U15231 ( .A(n11969), .ZN(n17911) );
  AOI22_X1 U15232 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15233 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11953) );
  OAI21_X1 U15234 ( .B1(n11974), .B2(n21691), .A(n11953), .ZN(n11958) );
  AOI22_X1 U15235 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15236 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11956) );
  INV_X2 U15237 ( .A(n11976), .ZN(n17852) );
  AOI22_X1 U15238 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15239 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15240 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9702), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U15241 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15242 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11961) );
  OAI21_X1 U15243 ( .B1(n9778), .B2(n21487), .A(n11961), .ZN(n11966) );
  AOI22_X1 U15244 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15245 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15246 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15247 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15248 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15249 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15250 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12040), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15251 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15252 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15253 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15254 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11975) );
  OAI21_X1 U15255 ( .B1(n11999), .B2(n21702), .A(n11975), .ZN(n11982) );
  AOI22_X1 U15256 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15257 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15258 ( .A1(n11931), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15259 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11977) );
  NAND4_X1 U15260 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(
        n11981) );
  AOI211_X1 U15261 ( .C1(n9696), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11982), .B(n11981), .ZN(n11983) );
  NAND3_X1 U15262 ( .A1(n11985), .A2(n11984), .A3(n11983), .ZN(n12113) );
  NOR2_X2 U15263 ( .A1(n19105), .A2(n19087), .ZN(n12148) );
  NOR2_X1 U15264 ( .A1(n19099), .A2(n12100), .ZN(n12101) );
  AOI22_X1 U15265 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15266 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15267 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15268 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U15269 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11995) );
  AOI22_X1 U15270 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15271 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15272 ( .A1(n9702), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15273 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U15274 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11994) );
  OR2_X1 U15275 ( .A1(n9681), .A2(n12147), .ZN(n12106) );
  NOR2_X1 U15276 ( .A1(n12101), .A2(n12106), .ZN(n11996) );
  OAI211_X1 U15277 ( .C1(n19091), .C2(n19547), .A(n12148), .B(n11996), .ZN(
        n12183) );
  AOI22_X1 U15278 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15279 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15280 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11997) );
  OAI21_X1 U15281 ( .B1(n17788), .B2(n21618), .A(n11997), .ZN(n12005) );
  AOI22_X1 U15282 ( .A1(n9693), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15283 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15284 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15285 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U15286 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12004) );
  NAND2_X1 U15287 ( .A1(n17261), .A2(n18267), .ZN(n18942) );
  INV_X1 U15288 ( .A(n18942), .ZN(n18803) );
  NAND2_X1 U15289 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18859) );
  NOR2_X1 U15290 ( .A1(n21613), .A2(n18545), .ZN(n18838) );
  AND3_X1 U15291 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18838), .ZN(n12115) );
  NAND2_X1 U15292 ( .A1(n12115), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18474) );
  NOR2_X1 U15293 ( .A1(n18805), .A2(n18474), .ZN(n12150) );
  INV_X1 U15294 ( .A(n12150), .ZN(n12203) );
  INV_X1 U15295 ( .A(n18806), .ZN(n12009) );
  NAND3_X1 U15296 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17230) );
  NOR2_X1 U15297 ( .A1(n12009), .A2(n17230), .ZN(n18780) );
  AOI22_X1 U15298 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15299 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9692), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15300 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15301 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12010) );
  NAND4_X1 U15302 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12019) );
  AOI22_X1 U15303 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15304 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15305 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12015) );
  INV_X2 U15306 ( .A(n18016), .ZN(n18043) );
  AOI22_X1 U15307 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U15308 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  AOI22_X1 U15309 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15310 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12028) );
  INV_X1 U15311 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21643) );
  AOI22_X1 U15312 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12020) );
  OAI21_X1 U15313 ( .B1(n17788), .B2(n21643), .A(n12020), .ZN(n12026) );
  AOI22_X1 U15314 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15315 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15316 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15317 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U15318 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12025) );
  AOI211_X1 U15319 ( .C1(n18105), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n12026), .B(n12025), .ZN(n12027) );
  NAND3_X1 U15320 ( .A1(n12029), .A2(n12028), .A3(n12027), .ZN(n12131) );
  AOI22_X1 U15321 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15322 ( .A1(n17773), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15323 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17806), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15324 ( .A1(n12040), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12030) );
  NAND4_X1 U15325 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12039) );
  AOI22_X1 U15326 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15327 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15328 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15329 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12070), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12034) );
  NAND4_X1 U15330 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n12038) );
  AOI22_X1 U15331 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15332 ( .A1(n17773), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11998), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15333 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18113), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n18107), .ZN(n12043) );
  AOI22_X1 U15334 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12040), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17806), .ZN(n12042) );
  AOI22_X1 U15335 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18112), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12071), .ZN(n12041) );
  INV_X1 U15336 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21495) );
  AOI22_X1 U15337 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15338 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15339 ( .A1(n12070), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12048) );
  OAI21_X1 U15340 ( .B1(n10946), .B2(n21702), .A(n12048), .ZN(n12054) );
  AOI22_X1 U15341 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15342 ( .A1(n17773), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15343 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15344 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17806), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12049) );
  NAND4_X1 U15345 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12053) );
  AOI211_X1 U15346 ( .C1(n18076), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n12054), .B(n12053), .ZN(n12055) );
  NAND3_X1 U15347 ( .A1(n12057), .A2(n12056), .A3(n12055), .ZN(n18282) );
  AOI22_X1 U15348 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15349 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18105), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15350 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15351 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U15352 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12068) );
  AOI22_X1 U15353 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15354 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15355 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15356 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15357 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12067) );
  INV_X1 U15358 ( .A(n18278), .ZN(n12084) );
  XOR2_X1 U15359 ( .A(n12095), .B(n12096), .Z(n12093) );
  XOR2_X1 U15360 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12093), .Z(
        n18701) );
  INV_X1 U15361 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19026) );
  XOR2_X1 U15362 ( .A(n18282), .B(n12069), .Z(n18735) );
  NAND2_X1 U15363 ( .A1(n18298), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12080) );
  XNOR2_X1 U15364 ( .A(n12118), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18765) );
  AOI22_X1 U15365 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15366 ( .A1(n11998), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12070), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15367 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17806), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15368 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12072) );
  INV_X1 U15369 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21634) );
  AOI22_X1 U15370 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15371 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12077) );
  INV_X1 U15372 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19693) );
  NOR2_X1 U15373 ( .A1(n9952), .A2(n19693), .ZN(n18771) );
  NAND2_X1 U15374 ( .A1(n18765), .A2(n18771), .ZN(n18764) );
  NAND2_X1 U15375 ( .A1(n12080), .A2(n18764), .ZN(n18753) );
  INV_X1 U15376 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19036) );
  NAND2_X1 U15377 ( .A1(n18753), .A2(n18754), .ZN(n18752) );
  OR2_X1 U15378 ( .A1(n19036), .A2(n12081), .ZN(n12082) );
  NAND2_X1 U15379 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12086), .ZN(
        n12087) );
  XNOR2_X1 U15380 ( .A(n12131), .B(n12088), .ZN(n12091) );
  NAND2_X1 U15381 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NAND2_X1 U15382 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12093), .ZN(
        n12094) );
  AOI21_X1 U15383 ( .B1(n18267), .B2(n17267), .A(n9684), .ZN(n12098) );
  NOR2_X1 U15384 ( .A1(n21474), .A2(n18966), .ZN(n18946) );
  NAND2_X1 U15385 ( .A1(n18946), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18920) );
  NAND2_X1 U15386 ( .A1(n18948), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18619) );
  NAND2_X1 U15387 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18903), .ZN(
        n18889) );
  NAND2_X1 U15388 ( .A1(n18780), .A2(n18887), .ZN(n18415) );
  NOR3_X2 U15389 ( .A1(n9681), .A2(n18156), .A3(n12195), .ZN(n12108) );
  NAND2_X1 U15390 ( .A1(n9728), .A2(n9681), .ZN(n12181) );
  NAND2_X1 U15391 ( .A1(n18342), .A2(n12181), .ZN(n17363) );
  NAND2_X1 U15392 ( .A1(n12147), .A2(n17363), .ZN(n14853) );
  NAND2_X1 U15393 ( .A1(n19524), .A2(n12101), .ZN(n17059) );
  NOR2_X1 U15394 ( .A1(n12104), .A2(n17059), .ZN(n12102) );
  NOR2_X1 U15395 ( .A1(n19095), .A2(n9681), .ZN(n12180) );
  NOR2_X1 U15396 ( .A1(n19076), .A2(n18343), .ZN(n12146) );
  OAI21_X1 U15397 ( .B1(n19105), .B2(n19547), .A(n12146), .ZN(n12184) );
  OAI21_X1 U15398 ( .B1(n12180), .B2(n12108), .A(n12184), .ZN(n12112) );
  AOI22_X1 U15399 ( .A1(n19087), .A2(n12104), .B1(n19091), .B2(n19547), .ZN(
        n12111) );
  AOI21_X1 U15400 ( .B1(n18197), .B2(n12107), .A(n19091), .ZN(n12105) );
  AOI21_X1 U15401 ( .B1(n12107), .B2(n12106), .A(n12105), .ZN(n12110) );
  NOR2_X1 U15402 ( .A1(n9681), .A2(n12107), .ZN(n12196) );
  OAI21_X1 U15403 ( .B1(n12108), .B2(n12196), .A(n19076), .ZN(n12109) );
  NAND3_X1 U15404 ( .A1(n12111), .A2(n12110), .A3(n12109), .ZN(n12182) );
  AOI21_X1 U15405 ( .B1(n12113), .B2(n12112), .A(n12182), .ZN(n12114) );
  NAND2_X1 U15406 ( .A1(n19520), .A2(n19521), .ZN(n19049) );
  INV_X1 U15407 ( .A(n19030), .ZN(n12117) );
  INV_X1 U15408 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19674) );
  INV_X1 U15409 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18984) );
  INV_X1 U15410 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18712) );
  NOR2_X1 U15411 ( .A1(n12128), .A2(n18712), .ZN(n18998) );
  NAND2_X1 U15412 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18998), .ZN(
        n18986) );
  NOR2_X1 U15413 ( .A1(n18984), .A2(n18986), .ZN(n18978) );
  NAND2_X1 U15414 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18978), .ZN(
        n18863) );
  OR2_X1 U15415 ( .A1(n19026), .A2(n18863), .ZN(n12149) );
  NOR3_X1 U15416 ( .A1(n19036), .A2(n19674), .A3(n12149), .ZN(n18877) );
  NAND2_X1 U15417 ( .A1(n17077), .A2(n18877), .ZN(n12155) );
  INV_X1 U15418 ( .A(n12155), .ZN(n18857) );
  INV_X1 U15419 ( .A(n18859), .ZN(n18507) );
  NAND2_X1 U15420 ( .A1(n18507), .A2(n12115), .ZN(n18823) );
  INV_X1 U15421 ( .A(n18823), .ZN(n18821) );
  NAND3_X1 U15422 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18857), .A3(
        n18821), .ZN(n12116) );
  NAND2_X1 U15423 ( .A1(n19546), .A2(n19693), .ZN(n18975) );
  INV_X1 U15424 ( .A(n18975), .ZN(n19028) );
  AOI21_X1 U15425 ( .B1(n19030), .B2(n12116), .A(n19028), .ZN(n18801) );
  OAI221_X1 U15426 ( .B1(n12117), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), 
        .C1(n12117), .C2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n18801), .ZN(
        n18789) );
  INV_X1 U15427 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18910) );
  NAND2_X1 U15428 ( .A1(n12125), .A2(n18282), .ZN(n12129) );
  NOR2_X1 U15429 ( .A1(n18278), .A2(n12129), .ZN(n12132) );
  NAND2_X1 U15430 ( .A1(n12132), .A2(n12131), .ZN(n12136) );
  NOR2_X1 U15431 ( .A1(n18271), .A2(n12136), .ZN(n12139) );
  NAND2_X1 U15432 ( .A1(n12139), .A2(n17262), .ZN(n12140) );
  NOR2_X1 U15433 ( .A1(n18298), .A2(n19693), .ZN(n12121) );
  NAND3_X1 U15434 ( .A1(n9952), .A2(n18298), .A3(n19693), .ZN(n12120) );
  OAI221_X1 U15435 ( .B1(n12121), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n9952), .C2(n18298), .A(n12120), .ZN(n18751) );
  NOR2_X1 U15436 ( .A1(n12122), .A2(n19036), .ZN(n12123) );
  XNOR2_X1 U15437 ( .A(n12129), .B(n18278), .ZN(n18726) );
  XNOR2_X1 U15438 ( .A(n12132), .B(n12131), .ZN(n12133) );
  NOR2_X2 U15439 ( .A1(n18711), .A2(n18712), .ZN(n18710) );
  NOR2_X1 U15440 ( .A1(n12134), .A2(n12133), .ZN(n12135) );
  XNOR2_X1 U15441 ( .A(n12136), .B(n18271), .ZN(n12137) );
  INV_X1 U15442 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18997) );
  XOR2_X1 U15443 ( .A(n12139), .B(n18267), .Z(n12142) );
  INV_X1 U15444 ( .A(n12140), .ZN(n12145) );
  OR2_X1 U15445 ( .A1(n12142), .A2(n12141), .ZN(n18694) );
  OAI21_X1 U15446 ( .B1(n12145), .B2(n12144), .A(n18694), .ZN(n12143) );
  NOR2_X1 U15447 ( .A1(n12147), .A2(n12146), .ZN(n19727) );
  NOR2_X1 U15448 ( .A1(n18156), .A2(n19091), .ZN(n19525) );
  INV_X1 U15449 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18793) );
  INV_X1 U15450 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18445) );
  NOR2_X1 U15451 ( .A1(n18793), .A2(n18445), .ZN(n17070) );
  OAI22_X1 U15452 ( .A1(n19548), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18949), .B2(n17070), .ZN(n12151) );
  NAND2_X1 U15453 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12156) );
  AOI21_X1 U15454 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18974) );
  NOR2_X1 U15455 ( .A1(n18974), .A2(n12149), .ZN(n18876) );
  NAND2_X1 U15456 ( .A1(n17077), .A2(n18876), .ZN(n18818) );
  NOR2_X1 U15457 ( .A1(n18859), .A2(n18818), .ZN(n18862) );
  NAND2_X1 U15458 ( .A1(n12150), .A2(n18862), .ZN(n18804) );
  NOR2_X1 U15459 ( .A1(n12156), .A2(n18804), .ZN(n18785) );
  AOI21_X1 U15460 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18785), .A(
        n19027), .ZN(n17078) );
  AOI211_X1 U15461 ( .C1(n18416), .C2(n19509), .A(n12151), .B(n17078), .ZN(
        n12152) );
  INV_X1 U15462 ( .A(n12152), .ZN(n12153) );
  AOI211_X2 U15463 ( .C1(n18803), .C2(n18415), .A(n18789), .B(n12153), .ZN(
        n18778) );
  AOI22_X1 U15464 ( .A1(n19509), .A2(n12154), .B1(n18943), .B2(n18803), .ZN(
        n18864) );
  INV_X1 U15465 ( .A(n17077), .ZN(n18865) );
  AOI21_X1 U15466 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19546), .A(
        n19049), .ZN(n19031) );
  OAI22_X1 U15467 ( .A1(n19027), .A2(n18818), .B1(n12155), .B2(n19031), .ZN(
        n17084) );
  INV_X1 U15468 ( .A(n17084), .ZN(n18787) );
  OAI21_X2 U15469 ( .B1(n18864), .B2(n18865), .A(n18787), .ZN(n18829) );
  NAND2_X1 U15470 ( .A1(n18806), .A2(n18829), .ZN(n12157) );
  OR2_X1 U15471 ( .A1(n12156), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18450) );
  OAI22_X1 U15472 ( .A1(n18778), .A2(n18445), .B1(n12157), .B2(n18450), .ZN(
        n12208) );
  INV_X1 U15473 ( .A(n12158), .ZN(n12187) );
  AOI21_X1 U15474 ( .B1(n19696), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12168), .ZN(n12188) );
  INV_X1 U15475 ( .A(n12168), .ZN(n12159) );
  OAI22_X1 U15476 ( .A1(n12161), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19557), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12169) );
  NOR2_X1 U15477 ( .A1(n12170), .A2(n12169), .ZN(n12162) );
  AOI22_X1 U15478 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19519), .B1(
        n12164), .B2(n12163), .ZN(n12173) );
  OAI21_X1 U15479 ( .B1(n19560), .B2(n12172), .A(n12173), .ZN(n12165) );
  OAI21_X1 U15480 ( .B1(n19519), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n12165), .ZN(n12166) );
  INV_X1 U15481 ( .A(n12166), .ZN(n12174) );
  NAND2_X1 U15482 ( .A1(n12168), .A2(n12189), .ZN(n12167) );
  OAI211_X1 U15483 ( .C1(n12168), .C2(n12189), .A(n12174), .B(n12167), .ZN(
        n12176) );
  XNOR2_X1 U15484 ( .A(n12170), .B(n12169), .ZN(n12175) );
  NAND2_X1 U15485 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19519), .ZN(
        n12171) );
  OAI22_X1 U15486 ( .A1(n12173), .A2(n19560), .B1(n12172), .B2(n12171), .ZN(
        n12191) );
  OAI21_X1 U15487 ( .B1(n12188), .B2(n12176), .A(n12192), .ZN(n19514) );
  NAND2_X1 U15488 ( .A1(n12192), .A2(n12176), .ZN(n19511) );
  INV_X1 U15489 ( .A(n9681), .ZN(n19083) );
  OAI21_X1 U15490 ( .B1(n19083), .B2(n18343), .A(n19713), .ZN(n12178) );
  NAND2_X1 U15491 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19716) );
  OAI21_X1 U15492 ( .B1(n12179), .B2(n12178), .A(n19716), .ZN(n17362) );
  NOR3_X1 U15493 ( .A1(n12180), .A2(n17357), .A3(n17362), .ZN(n12186) );
  OAI21_X1 U15494 ( .B1(n12183), .B2(n12182), .A(n12181), .ZN(n12185) );
  NAND2_X1 U15495 ( .A1(n12185), .A2(n12184), .ZN(n14854) );
  INV_X1 U15496 ( .A(n12188), .ZN(n12190) );
  NOR2_X1 U15497 ( .A1(n12190), .A2(n12189), .ZN(n12194) );
  INV_X1 U15498 ( .A(n12191), .ZN(n12193) );
  OAI21_X1 U15499 ( .B1(n12196), .B2(n12195), .A(n19513), .ZN(n12197) );
  INV_X1 U15500 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18637) );
  NAND3_X1 U15501 ( .A1(n21474), .A2(n18966), .A3(n18637), .ZN(n18583) );
  NOR3_X1 U15502 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n18583), .ZN(n18607) );
  INV_X1 U15503 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18881) );
  INV_X1 U15504 ( .A(n18572), .ZN(n18502) );
  NOR2_X1 U15505 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18573), .ZN(
        n18555) );
  NAND2_X1 U15506 ( .A1(n18555), .A2(n18545), .ZN(n18532) );
  NOR2_X1 U15507 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18532), .ZN(
        n18514) );
  INV_X1 U15508 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18516) );
  NAND2_X1 U15509 ( .A1(n18514), .A2(n18516), .ZN(n18501) );
  NAND2_X1 U15510 ( .A1(n18673), .A2(n18455), .ZN(n12204) );
  AOI21_X1 U15511 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n12205), .A(
        n17073), .ZN(n18444) );
  NAND3_X1 U15512 ( .A1(n17262), .A2(n17261), .A3(n19039), .ZN(n18970) );
  INV_X2 U15513 ( .A(n19055), .ZN(n19040) );
  NOR2_X2 U15514 ( .A1(n19040), .A2(n19039), .ZN(n19047) );
  AOI21_X1 U15515 ( .B1(n19047), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10936), .ZN(n12206) );
  INV_X1 U15516 ( .A(n14230), .ZN(n12219) );
  NAND2_X1 U15517 ( .A1(n11055), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U15518 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20227) );
  XNOR2_X1 U15519 ( .A(n20227), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19994) );
  AND2_X1 U15520 ( .A1(n19994), .A2(n20528), .ZN(n20266) );
  AOI21_X1 U15521 ( .B1(n12228), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n20266), .ZN(n12212) );
  NAND2_X1 U15522 ( .A1(n12228), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12217) );
  NAND2_X1 U15523 ( .A1(n20338), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20195) );
  NAND2_X1 U15524 ( .A1(n14690), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20297) );
  NAND2_X1 U15525 ( .A1(n20195), .A2(n20297), .ZN(n20342) );
  NAND2_X1 U15526 ( .A1(n20342), .A2(n20528), .ZN(n20197) );
  NAND2_X1 U15527 ( .A1(n12217), .A2(n20197), .ZN(n12218) );
  NAND2_X1 U15528 ( .A1(n14292), .A2(n14291), .ZN(n12223) );
  INV_X1 U15529 ( .A(n12220), .ZN(n12221) );
  NAND2_X1 U15530 ( .A1(n12223), .A2(n12222), .ZN(n14523) );
  OAI21_X1 U15531 ( .B1(n20227), .B2(n20542), .A(n20533), .ZN(n12226) );
  NAND2_X1 U15532 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20296) );
  INV_X1 U15533 ( .A(n20296), .ZN(n20341) );
  NAND2_X1 U15534 ( .A1(n20392), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20400) );
  AND3_X1 U15535 ( .A1(n12226), .A2(n20400), .A3(n20528), .ZN(n12227) );
  AOI21_X1 U15536 ( .B1(n12228), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12227), .ZN(n12229) );
  NAND2_X1 U15537 ( .A1(n12232), .A2(n12230), .ZN(n14780) );
  NAND2_X1 U15538 ( .A1(n11055), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12231) );
  INV_X1 U15539 ( .A(n16343), .ZN(n12236) );
  AND2_X1 U15540 ( .A1(n14788), .A2(n14768), .ZN(n12235) );
  AND3_X1 U15541 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__5__SCAN_IN), 
        .ZN(n12234) );
  AND2_X1 U15542 ( .A1(n16342), .A2(n14848), .ZN(n12233) );
  NAND4_X1 U15543 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n14800) );
  AOI22_X1 U15544 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15545 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15546 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15547 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12237) );
  NAND4_X1 U15548 ( .A1(n12240), .A2(n12239), .A3(n12238), .A4(n12237), .ZN(
        n12246) );
  AOI22_X1 U15549 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15550 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15551 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15552 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12241) );
  NAND4_X1 U15553 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12241), .ZN(
        n12245) );
  OR2_X1 U15554 ( .A1(n12246), .A2(n12245), .ZN(n14805) );
  AND2_X1 U15555 ( .A1(n14805), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12247) );
  NAND4_X1 U15556 ( .A1(n12247), .A2(n14803), .A3(n14826), .A4(n14802), .ZN(
        n12248) );
  NOR3_X1 U15557 ( .A1(n14800), .A2(n14652), .A3(n12248), .ZN(n12249) );
  AOI22_X1 U15558 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15559 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11358), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15560 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12330), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15561 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11251), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15562 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12259) );
  AOI22_X1 U15563 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11306), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15564 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11245), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15565 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15566 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12254) );
  NAND4_X1 U15567 ( .A1(n12257), .A2(n12256), .A3(n12255), .A4(n12254), .ZN(
        n12258) );
  NOR2_X1 U15568 ( .A1(n12259), .A2(n12258), .ZN(n16331) );
  AOI22_X1 U15569 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15570 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15571 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15572 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12260) );
  NAND4_X1 U15573 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12269) );
  AOI22_X1 U15574 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15575 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15576 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15577 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15578 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12268) );
  OR2_X1 U15579 ( .A1(n12269), .A2(n12268), .ZN(n16326) );
  AOI22_X1 U15580 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15581 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15582 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15583 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11251), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U15584 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12280) );
  AOI22_X1 U15585 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11244), .B1(
        n11306), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15586 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15587 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15588 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12275) );
  NAND4_X1 U15589 ( .A1(n12278), .A2(n12277), .A3(n12276), .A4(n12275), .ZN(
        n12279) );
  NOR2_X1 U15590 ( .A1(n12280), .A2(n12279), .ZN(n16324) );
  INV_X1 U15591 ( .A(n16324), .ZN(n12281) );
  AOI22_X1 U15592 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15593 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15594 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15595 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12282) );
  NAND4_X1 U15596 ( .A1(n12285), .A2(n12284), .A3(n12283), .A4(n12282), .ZN(
        n12291) );
  AOI22_X1 U15597 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15598 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15599 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15600 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12286) );
  NAND4_X1 U15601 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n12286), .ZN(
        n12290) );
  NOR2_X1 U15602 ( .A1(n12291), .A2(n12290), .ZN(n16320) );
  AOI22_X1 U15603 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15604 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15605 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15606 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12295) );
  NAND4_X1 U15607 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12304) );
  AOI22_X1 U15608 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15609 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15610 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15611 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12299) );
  NAND4_X1 U15612 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n12303) );
  NOR2_X1 U15613 ( .A1(n12304), .A2(n12303), .ZN(n16311) );
  AOI22_X1 U15614 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11250), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15615 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11355), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15616 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15617 ( .A1(n11251), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U15618 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12314) );
  AOI22_X1 U15619 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15620 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15621 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15622 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12309) );
  NAND4_X1 U15623 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12313) );
  OR2_X1 U15624 ( .A1(n12314), .A2(n12313), .ZN(n16306) );
  AOI22_X1 U15625 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12318) );
  INV_X1 U15626 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U15627 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12317) );
  AND2_X1 U15628 ( .A1(n12318), .A2(n12317), .ZN(n12322) );
  AOI22_X1 U15629 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12321) );
  XNOR2_X1 U15630 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12460) );
  NAND4_X1 U15631 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12460), .ZN(
        n12329) );
  AOI22_X1 U15632 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12324) );
  INV_X1 U15633 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20241) );
  AOI22_X1 U15634 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12323) );
  AND2_X1 U15635 ( .A1(n12324), .A2(n12323), .ZN(n12327) );
  AOI22_X1 U15636 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12326) );
  INV_X1 U15637 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n20169) );
  NAND4_X1 U15638 ( .A1(n12327), .A2(n12469), .A3(n12326), .A4(n12325), .ZN(
        n12328) );
  AND2_X1 U15639 ( .A1(n12329), .A2(n12328), .ZN(n12350) );
  NAND2_X1 U15640 ( .A1(n12350), .A2(n14347), .ZN(n12345) );
  AOI22_X1 U15641 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12294), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15642 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11358), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15643 ( .A1(n11245), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11251), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15644 ( .A1(n11355), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12331) );
  NAND4_X1 U15645 ( .A1(n12334), .A2(n12333), .A3(n12332), .A4(n12331), .ZN(
        n12344) );
  AOI22_X1 U15646 ( .A1(n11306), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11244), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15647 ( .A1(n11250), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15648 ( .A1(n11222), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12336), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15649 ( .A1(n11238), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12337), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12339) );
  NAND4_X1 U15650 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12343) );
  OR2_X1 U15651 ( .A1(n12344), .A2(n12343), .ZN(n12351) );
  XNOR2_X1 U15652 ( .A(n12345), .B(n12351), .ZN(n12347) );
  INV_X1 U15653 ( .A(n12350), .ZN(n12346) );
  NOR2_X1 U15654 ( .A1(n14347), .A2(n12346), .ZN(n16301) );
  NAND2_X1 U15655 ( .A1(n16299), .A2(n16301), .ZN(n16300) );
  INV_X1 U15656 ( .A(n12347), .ZN(n12348) );
  NAND2_X1 U15657 ( .A1(n16300), .A2(n12349), .ZN(n16296) );
  NAND2_X1 U15658 ( .A1(n12351), .A2(n12350), .ZN(n12369) );
  AOI22_X1 U15659 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15660 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12352) );
  AND2_X1 U15661 ( .A1(n12353), .A2(n12352), .ZN(n12356) );
  AOI22_X1 U15662 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U15663 ( .A1(n12356), .A2(n12355), .A3(n12354), .A4(n12460), .ZN(
        n12363) );
  AOI22_X1 U15664 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15665 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12357) );
  AND2_X1 U15666 ( .A1(n12358), .A2(n12357), .ZN(n12361) );
  AOI22_X1 U15667 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12360) );
  NAND4_X1 U15668 ( .A1(n12361), .A2(n12469), .A3(n12360), .A4(n12359), .ZN(
        n12362) );
  AND2_X1 U15669 ( .A1(n12363), .A2(n12362), .ZN(n12367) );
  XNOR2_X1 U15670 ( .A(n12369), .B(n12367), .ZN(n12364) );
  NAND2_X1 U15671 ( .A1(n12364), .A2(n12386), .ZN(n12366) );
  NAND2_X1 U15672 ( .A1(n11650), .A2(n12367), .ZN(n12365) );
  NAND2_X1 U15673 ( .A1(n12366), .A2(n12365), .ZN(n16295) );
  NAND2_X2 U15674 ( .A1(n16296), .A2(n16295), .ZN(n16294) );
  INV_X1 U15675 ( .A(n12367), .ZN(n12368) );
  NOR2_X1 U15676 ( .A1(n12369), .A2(n12368), .ZN(n12382) );
  AOI22_X1 U15677 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12371) );
  INV_X1 U15678 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U15679 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12370) );
  AND2_X1 U15680 ( .A1(n12371), .A2(n12370), .ZN(n12374) );
  AOI22_X1 U15681 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15682 ( .A1(n12374), .A2(n12373), .A3(n12372), .A4(n12460), .ZN(
        n12381) );
  AOI22_X1 U15683 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15684 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12375) );
  AND2_X1 U15685 ( .A1(n12376), .A2(n12375), .ZN(n12379) );
  AOI22_X1 U15686 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U15687 ( .A1(n12379), .A2(n12469), .A3(n12378), .A4(n12377), .ZN(
        n12380) );
  AND2_X1 U15688 ( .A1(n12381), .A2(n12380), .ZN(n12383) );
  NAND2_X1 U15689 ( .A1(n12382), .A2(n12383), .ZN(n12400) );
  INV_X1 U15690 ( .A(n12382), .ZN(n12384) );
  INV_X1 U15691 ( .A(n12383), .ZN(n12405) );
  NAND2_X1 U15692 ( .A1(n12384), .A2(n12405), .ZN(n12385) );
  AND3_X1 U15693 ( .A1(n12400), .A2(n12386), .A3(n12385), .ZN(n12404) );
  INV_X1 U15694 ( .A(n12404), .ZN(n12387) );
  AOI22_X1 U15695 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15696 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12388) );
  AND2_X1 U15697 ( .A1(n12389), .A2(n12388), .ZN(n12392) );
  AOI22_X1 U15698 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12391) );
  NAND4_X1 U15699 ( .A1(n12392), .A2(n12391), .A3(n12390), .A4(n12460), .ZN(
        n12399) );
  AOI22_X1 U15700 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15701 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12393) );
  AND2_X1 U15702 ( .A1(n12394), .A2(n12393), .ZN(n12397) );
  AOI22_X1 U15703 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15704 ( .A1(n12397), .A2(n12469), .A3(n12396), .A4(n12395), .ZN(
        n12398) );
  AND2_X1 U15705 ( .A1(n12399), .A2(n12398), .ZN(n12406) );
  AOI21_X1 U15706 ( .B1(n12400), .B2(n16282), .A(n14652), .ZN(n12401) );
  OR2_X1 U15707 ( .A1(n12400), .A2(n16282), .ZN(n12422) );
  NAND2_X1 U15708 ( .A1(n12401), .A2(n12422), .ZN(n16284) );
  INV_X1 U15709 ( .A(n16284), .ZN(n12402) );
  NAND2_X1 U15710 ( .A1(n12403), .A2(n12402), .ZN(n12407) );
  NOR2_X1 U15711 ( .A1(n14347), .A2(n12405), .ZN(n16291) );
  INV_X1 U15712 ( .A(n12422), .ZN(n12420) );
  AOI22_X1 U15713 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15714 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12408) );
  AND2_X1 U15715 ( .A1(n12409), .A2(n12408), .ZN(n12412) );
  AOI22_X1 U15716 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12411) );
  NAND4_X1 U15717 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12460), .ZN(
        n12419) );
  AOI22_X1 U15718 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11043), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15719 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12413) );
  AND2_X1 U15720 ( .A1(n12414), .A2(n12413), .ZN(n12417) );
  AOI22_X1 U15721 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12416) );
  NAND4_X1 U15722 ( .A1(n12417), .A2(n12469), .A3(n12416), .A4(n12415), .ZN(
        n12418) );
  AND2_X1 U15723 ( .A1(n12419), .A2(n12418), .ZN(n12426) );
  NAND2_X1 U15724 ( .A1(n12420), .A2(n12426), .ZN(n16270) );
  INV_X1 U15725 ( .A(n12426), .ZN(n12421) );
  AOI21_X1 U15726 ( .B1(n12422), .B2(n12421), .A(n14652), .ZN(n12423) );
  AND2_X1 U15727 ( .A1(n16270), .A2(n12423), .ZN(n12424) );
  NAND2_X1 U15728 ( .A1(n11650), .A2(n12426), .ZN(n16277) );
  INV_X1 U15729 ( .A(n16271), .ZN(n12439) );
  AOI22_X1 U15730 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15731 ( .A1(n9711), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12427) );
  AND2_X1 U15732 ( .A1(n12428), .A2(n12427), .ZN(n12431) );
  AOI22_X1 U15733 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12430) );
  NAND4_X1 U15734 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12460), .ZN(
        n12438) );
  AOI22_X1 U15735 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15736 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12432) );
  AND2_X1 U15737 ( .A1(n12433), .A2(n12432), .ZN(n12436) );
  AOI22_X1 U15738 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15739 ( .A1(n12436), .A2(n12469), .A3(n12435), .A4(n12434), .ZN(
        n12437) );
  AND2_X1 U15740 ( .A1(n12438), .A2(n12437), .ZN(n16272) );
  INV_X1 U15741 ( .A(n16270), .ZN(n12441) );
  AND2_X1 U15742 ( .A1(n16272), .A2(n14347), .ZN(n12440) );
  AND2_X1 U15743 ( .A1(n12441), .A2(n12440), .ZN(n12455) );
  AOI22_X1 U15744 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15745 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12442) );
  AND2_X1 U15746 ( .A1(n12443), .A2(n12442), .ZN(n12446) );
  AOI22_X1 U15747 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12445) );
  NAND4_X1 U15748 ( .A1(n12446), .A2(n12445), .A3(n12444), .A4(n12460), .ZN(
        n12453) );
  AOI22_X1 U15749 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12448) );
  INV_X1 U15750 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n21627) );
  AOI22_X1 U15751 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9709), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12447) );
  AND2_X1 U15752 ( .A1(n12448), .A2(n12447), .ZN(n12451) );
  AOI22_X1 U15753 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12450) );
  NAND4_X1 U15754 ( .A1(n12451), .A2(n12469), .A3(n12450), .A4(n12449), .ZN(
        n12452) );
  AND2_X1 U15755 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  NAND2_X1 U15756 ( .A1(n12455), .A2(n12454), .ZN(n12456) );
  OAI21_X1 U15757 ( .B1(n12455), .B2(n12454), .A(n12456), .ZN(n16266) );
  AOI22_X1 U15758 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9708), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15759 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U15760 ( .A1(n12459), .A2(n12458), .ZN(n12474) );
  AOI22_X1 U15761 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12466), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12461) );
  NAND3_X1 U15762 ( .A1(n12462), .A2(n12461), .A3(n12460), .ZN(n12473) );
  AOI22_X1 U15763 ( .A1(n12457), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15764 ( .A1(n9710), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14662), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12464) );
  NAND2_X1 U15765 ( .A1(n12465), .A2(n12464), .ZN(n12472) );
  AOI22_X1 U15766 ( .A1(n12467), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12468) );
  NAND3_X1 U15767 ( .A1(n12470), .A2(n12469), .A3(n12468), .ZN(n12471) );
  OAI22_X1 U15768 ( .A1(n12474), .A2(n12473), .B1(n12472), .B2(n12471), .ZN(
        n12475) );
  INV_X1 U15769 ( .A(n14699), .ZN(n12476) );
  INV_X1 U15770 ( .A(n14597), .ZN(n14700) );
  NAND2_X1 U15771 ( .A1(n12476), .A2(n14700), .ZN(n14339) );
  NAND2_X1 U15772 ( .A1(n14661), .A2(n12477), .ZN(n14595) );
  NAND2_X1 U15773 ( .A1(n14339), .A2(n14595), .ZN(n12478) );
  NAND2_X1 U15774 ( .A1(n9694), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12480) );
  NAND2_X1 U15775 ( .A1(n12503), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12479) );
  OAI211_X1 U15776 ( .C1(n11127), .C2(n13695), .A(n12480), .B(n12479), .ZN(
        n12481) );
  AOI21_X1 U15777 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12481), .ZN(n16037) );
  INV_X1 U15778 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16027) );
  NAND2_X1 U15779 ( .A1(n11126), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12484) );
  AOI22_X1 U15780 ( .A1(n9694), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12483) );
  OAI211_X1 U15781 ( .C1(n16027), .C2(n13758), .A(n12484), .B(n12483), .ZN(
        n16023) );
  NAND2_X1 U15782 ( .A1(n16021), .A2(n16023), .ZN(n16004) );
  NAND2_X1 U15783 ( .A1(n9694), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12487) );
  NAND2_X1 U15784 ( .A1(n12503), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12486) );
  NAND2_X1 U15785 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12485) );
  NAND3_X1 U15786 ( .A1(n12487), .A2(n12486), .A3(n12485), .ZN(n12488) );
  AOI21_X1 U15787 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12488), .ZN(n16005) );
  NAND2_X1 U15788 ( .A1(n9694), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U15789 ( .A1(n12503), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12491) );
  OAI211_X1 U15790 ( .C1(n11127), .C2(n15997), .A(n12492), .B(n12491), .ZN(
        n12493) );
  AOI21_X1 U15791 ( .B1(n11544), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12493), .ZN(n15992) );
  INV_X1 U15792 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16288) );
  NAND2_X1 U15793 ( .A1(n11544), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12495) );
  AOI22_X1 U15794 ( .A1(n9694), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12494) );
  OAI211_X1 U15795 ( .C1(n16288), .C2(n13758), .A(n12495), .B(n12494), .ZN(
        n13790) );
  INV_X1 U15796 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12498) );
  NAND2_X1 U15797 ( .A1(n11126), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12497) );
  AOI22_X1 U15798 ( .A1(n9694), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12496) );
  OAI211_X1 U15799 ( .C1(n12498), .C2(n13758), .A(n12497), .B(n12496), .ZN(
        n15964) );
  INV_X1 U15800 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U15801 ( .A1(n9694), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12500) );
  NAND2_X1 U15802 ( .A1(n12503), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12499) );
  OAI211_X1 U15803 ( .C1(n12506), .C2(n14927), .A(n12500), .B(n12499), .ZN(
        n13607) );
  INV_X1 U15804 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15950) );
  AOI22_X1 U15805 ( .A1(n9694), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12501) );
  OAI21_X1 U15806 ( .B1(n13758), .B2(n15950), .A(n12501), .ZN(n12502) );
  AOI21_X1 U15807 ( .B1(n11126), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12502), .ZN(n14916) );
  AOI22_X1 U15808 ( .A1(n9694), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12505) );
  NAND2_X1 U15809 ( .A1(n12503), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12504) );
  OAI211_X1 U15810 ( .C1(n12506), .C2(n10555), .A(n12505), .B(n12504), .ZN(
        n13753) );
  OAI21_X1 U15811 ( .B1(n16364), .B2(n16354), .A(n12508), .ZN(P2_U2857) );
  INV_X1 U15812 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12509) );
  INV_X1 U15813 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15814 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12741), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15815 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12513) );
  AND2_X2 U15816 ( .A1(n14504), .A2(n12515), .ZN(n12617) );
  AOI22_X1 U15817 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15818 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12733), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12521) );
  AND2_X2 U15819 ( .A1(n12517), .A2(n14178), .ZN(n12619) );
  AOI22_X1 U15820 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12520) );
  AND2_X2 U15821 ( .A1(n14504), .A2(n12517), .ZN(n12618) );
  AOI22_X1 U15822 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12618), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12518) );
  NAND2_X1 U15823 ( .A1(n10950), .A2(n12522), .ZN(n12634) );
  INV_X2 U15824 ( .A(n12634), .ZN(n12630) );
  NAND2_X1 U15825 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12526) );
  NAND2_X1 U15826 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12525) );
  NAND2_X1 U15827 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12524) );
  NAND2_X1 U15828 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12523) );
  NAND2_X1 U15829 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12530) );
  NAND2_X1 U15830 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12529) );
  NAND2_X1 U15831 ( .A1(n12618), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12528) );
  NAND2_X1 U15832 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12527) );
  NAND2_X1 U15833 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12534) );
  NAND2_X1 U15834 ( .A1(n12740), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12533) );
  NAND2_X1 U15835 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12532) );
  NAND2_X1 U15836 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U15837 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12538) );
  NAND2_X1 U15838 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12537) );
  NAND2_X1 U15839 ( .A1(n12713), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12536) );
  NAND2_X1 U15840 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12535) );
  NAND2_X1 U15841 ( .A1(n12630), .A2(n20812), .ZN(n12645) );
  INV_X1 U15842 ( .A(n12645), .ZN(n12571) );
  AOI22_X1 U15843 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15844 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15845 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12713), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15846 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15847 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12740), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15848 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15849 ( .A1(n12618), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12547) );
  NAND2_X4 U15850 ( .A1(n12552), .A2(n12551), .ZN(n14173) );
  AOI22_X1 U15851 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15852 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15853 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12713), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15854 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15855 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12740), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15856 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15857 ( .A1(n12618), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12557) );
  NAND2_X2 U15858 ( .A1(n12562), .A2(n12561), .ZN(n12637) );
  AOI22_X1 U15859 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12607), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15860 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12713), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15861 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15862 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15863 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15864 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15865 ( .A1(n12740), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12618), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U15866 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U15867 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U15868 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12573) );
  NAND2_X1 U15869 ( .A1(n12713), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U15870 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12579) );
  NAND2_X1 U15871 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12578) );
  NAND2_X1 U15872 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12577) );
  NAND2_X1 U15873 ( .A1(n12740), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12576) );
  NAND2_X1 U15874 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12583) );
  NAND2_X1 U15875 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U15876 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12581) );
  NAND2_X1 U15877 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12580) );
  NAND2_X1 U15878 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12587) );
  NAND2_X1 U15879 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12586) );
  NAND2_X1 U15880 ( .A1(n12618), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12585) );
  NAND2_X1 U15881 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12584) );
  NAND4_X4 U15882 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        n14566) );
  INV_X1 U15883 ( .A(n14056), .ZN(n12602) );
  AOI22_X1 U15884 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12732), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15885 ( .A1(n12740), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12607), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15886 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12741), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15887 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12619), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15888 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12601) );
  AOI22_X1 U15889 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12757), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15890 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12713), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15891 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12618), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15892 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12596) );
  NAND4_X1 U15893 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  NAND2_X1 U15894 ( .A1(n12602), .A2(n14587), .ZN(n12662) );
  INV_X1 U15895 ( .A(n12662), .ZN(n12629) );
  NAND2_X1 U15896 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12606) );
  NAND2_X1 U15897 ( .A1(n12732), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12605) );
  NAND2_X1 U15898 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12604) );
  NAND2_X1 U15899 ( .A1(n12713), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12603) );
  NAND2_X1 U15900 ( .A1(n12607), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12611) );
  NAND2_X1 U15901 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12610) );
  NAND2_X1 U15902 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12609) );
  NAND2_X1 U15903 ( .A1(n12740), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12608) );
  NAND2_X1 U15904 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12616) );
  NAND2_X1 U15905 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12615) );
  NAND2_X1 U15906 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12614) );
  NAND2_X1 U15907 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12613) );
  NAND2_X1 U15908 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12623) );
  NAND2_X1 U15909 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12622) );
  NAND2_X1 U15910 ( .A1(n12618), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12621) );
  NAND2_X1 U15911 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12620) );
  NAND4_X4 U15912 ( .A1(n12627), .A2(n12626), .A3(n12625), .A4(n12624), .ZN(
        n13430) );
  NAND2_X1 U15913 ( .A1(n12629), .A2(n9817), .ZN(n12653) );
  NAND2_X2 U15914 ( .A1(n12630), .A2(n14173), .ZN(n13912) );
  NAND2_X1 U15915 ( .A1(n13912), .A2(n14566), .ZN(n12631) );
  AND2_X1 U15916 ( .A1(n12631), .A2(n12677), .ZN(n13919) );
  NAND2_X1 U15917 ( .A1(n13919), .A2(n13052), .ZN(n12635) );
  NAND2_X1 U15918 ( .A1(n12658), .A2(n12671), .ZN(n14162) );
  NAND2_X1 U15919 ( .A1(n14162), .A2(n14587), .ZN(n13911) );
  NAND2_X1 U15920 ( .A1(n12676), .A2(n13912), .ZN(n12668) );
  NAND2_X1 U15921 ( .A1(n12635), .A2(n12668), .ZN(n12652) );
  BUF_X4 U15922 ( .A(n13430), .Z(n14297) );
  NAND2_X2 U15923 ( .A1(n13916), .A2(n12636), .ZN(n14055) );
  NAND2_X1 U15924 ( .A1(n12648), .A2(n14566), .ZN(n13432) );
  NAND2_X2 U15925 ( .A1(n13432), .A2(n13454), .ZN(n14158) );
  INV_X1 U15926 ( .A(n12638), .ZN(n13915) );
  NAND2_X1 U15927 ( .A1(n14158), .A2(n13915), .ZN(n13931) );
  NAND2_X1 U15928 ( .A1(n14566), .A2(n14198), .ZN(n12640) );
  OAI211_X1 U15929 ( .C1(n14054), .C2(n14055), .A(n13931), .B(n14174), .ZN(
        n12641) );
  INV_X1 U15930 ( .A(n12641), .ZN(n12651) );
  NAND2_X1 U15931 ( .A1(n13912), .A2(n14173), .ZN(n12642) );
  NAND2_X1 U15932 ( .A1(n12642), .A2(n20804), .ZN(n12643) );
  NAND2_X1 U15933 ( .A1(n12644), .A2(n12643), .ZN(n12647) );
  NAND2_X1 U15934 ( .A1(n12647), .A2(n12646), .ZN(n12669) );
  NAND2_X1 U15935 ( .A1(n14179), .A2(n17112), .ZN(n12649) );
  OAI21_X1 U15936 ( .B1(n12669), .B2(n12649), .A(n13916), .ZN(n12650) );
  NAND4_X1 U15937 ( .A1(n12653), .A2(n12652), .A3(n12651), .A4(n12650), .ZN(
        n12654) );
  NAND2_X1 U15938 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12690) );
  OAI21_X1 U15939 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n12690), .ZN(n21087) );
  NAND2_X1 U15940 ( .A1(n21329), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12683) );
  OAI21_X1 U15941 ( .B1(n13973), .B2(n21087), .A(n12683), .ZN(n12656) );
  INV_X1 U15942 ( .A(n12656), .ZN(n12657) );
  INV_X1 U15943 ( .A(n13409), .ZN(n12660) );
  NAND2_X1 U15944 ( .A1(n13904), .A2(n12658), .ZN(n12659) );
  OR2_X1 U15945 ( .A1(n14054), .A2(n14566), .ZN(n12661) );
  NOR2_X1 U15946 ( .A1(n12669), .A2(n12661), .ZN(n13396) );
  NAND2_X1 U15947 ( .A1(n13396), .A2(n17112), .ZN(n14175) );
  INV_X1 U15948 ( .A(n12662), .ZN(n17113) );
  NAND2_X1 U15949 ( .A1(n17113), .A2(n14297), .ZN(n12663) );
  NAND2_X1 U15950 ( .A1(n14175), .A2(n12663), .ZN(n13925) );
  OAI21_X2 U15951 ( .B1(n12664), .B2(n13925), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12682) );
  INV_X1 U15952 ( .A(n21329), .ZN(n17119) );
  MUX2_X1 U15953 ( .A(n17119), .B(n13973), .S(n21199), .Z(n12667) );
  NAND3_X1 U15954 ( .A1(n12668), .A2(n14297), .A3(n15918), .ZN(n12681) );
  NAND2_X1 U15955 ( .A1(n12669), .A2(n15267), .ZN(n13935) );
  NAND2_X1 U15956 ( .A1(n14980), .A2(n12670), .ZN(n12673) );
  INV_X1 U15957 ( .A(n17163), .ZN(n15931) );
  NOR2_X1 U15958 ( .A1(n15931), .A2(n17176), .ZN(n12672) );
  NAND2_X1 U15959 ( .A1(n14484), .A2(n12630), .ZN(n13939) );
  NAND2_X1 U15960 ( .A1(n13916), .A2(n14297), .ZN(n14199) );
  NAND4_X1 U15961 ( .A1(n12673), .A2(n12672), .A3(n13939), .A4(n14199), .ZN(
        n12675) );
  INV_X1 U15962 ( .A(n14174), .ZN(n12674) );
  NOR2_X1 U15963 ( .A1(n12675), .A2(n12674), .ZN(n12680) );
  INV_X1 U15964 ( .A(n12676), .ZN(n12678) );
  NAND2_X1 U15965 ( .A1(n12678), .A2(n14052), .ZN(n12679) );
  NAND4_X1 U15966 ( .A1(n12681), .A2(n13935), .A3(n12680), .A4(n12679), .ZN(
        n12729) );
  INV_X1 U15967 ( .A(n12682), .ZN(n12685) );
  NAND2_X1 U15968 ( .A1(n12683), .A2(n12655), .ZN(n12684) );
  NAND2_X1 U15969 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  OR2_X1 U15971 ( .A1(n12688), .A2(n12510), .ZN(n12693) );
  INV_X1 U15972 ( .A(n13973), .ZN(n12781) );
  INV_X1 U15973 ( .A(n12690), .ZN(n12689) );
  NAND2_X1 U15974 ( .A1(n12689), .A2(n21157), .ZN(n21117) );
  NAND2_X1 U15975 ( .A1(n12690), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12691) );
  NAND2_X1 U15976 ( .A1(n21117), .A2(n12691), .ZN(n20787) );
  AOI22_X1 U15977 ( .A1(n12781), .A2(n20787), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21329), .ZN(n12692) );
  NAND2_X1 U15978 ( .A1(n12696), .A2(n14505), .ZN(n14171) );
  AOI22_X1 U15979 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15980 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15981 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15982 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12698) );
  NAND4_X1 U15983 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12707) );
  AOI22_X1 U15984 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15985 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15986 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15987 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U15988 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12706) );
  OAI22_X2 U15989 ( .A1(n14171), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13830), 
        .B2(n12785), .ZN(n12710) );
  INV_X1 U15990 ( .A(n12784), .ZN(n12771) );
  XNOR2_X1 U15991 ( .A(n12710), .B(n12709), .ZN(n12881) );
  AOI22_X1 U15992 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15993 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15994 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15995 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12714) );
  NAND4_X1 U15996 ( .A1(n12717), .A2(n12716), .A3(n12715), .A4(n12714), .ZN(
        n12726) );
  INV_X2 U15997 ( .A(n12697), .ZN(n13316) );
  AOI22_X1 U15998 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15999 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U16000 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U16001 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12721) );
  NAND4_X1 U16002 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12725) );
  INV_X1 U16003 ( .A(n13821), .ZN(n12727) );
  NOR2_X1 U16004 ( .A1(n12727), .A2(n12785), .ZN(n12728) );
  INV_X1 U16005 ( .A(n12729), .ZN(n12730) );
  AOI22_X1 U16006 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U16007 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U16008 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12736) );
  INV_X1 U16009 ( .A(n12734), .ZN(n12825) );
  INV_X2 U16010 ( .A(n12825), .ZN(n14483) );
  AOI22_X1 U16011 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12735) );
  NAND4_X1 U16012 ( .A1(n12738), .A2(n12737), .A3(n12736), .A4(n12735), .ZN(
        n12747) );
  AOI22_X1 U16013 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U16014 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12740), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U16015 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U16016 ( .A1(n12618), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12742) );
  NAND4_X1 U16017 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12746) );
  NOR2_X1 U16018 ( .A1(n12785), .A2(n13876), .ZN(n12770) );
  AOI22_X1 U16019 ( .A1(n12748), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U16020 ( .A1(n12733), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U16021 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16022 ( .A1(n12739), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12750) );
  NAND4_X1 U16023 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12763) );
  AOI22_X1 U16024 ( .A1(n13123), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U16025 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16026 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12618), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16027 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12758) );
  NAND4_X1 U16028 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12762) );
  MUX2_X1 U16029 ( .A(n12769), .B(n12770), .S(n13820), .Z(n12764) );
  INV_X1 U16030 ( .A(n12764), .ZN(n12765) );
  INV_X1 U16031 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12768) );
  AOI21_X1 U16032 ( .B1(n13916), .B2(n13820), .A(n17176), .ZN(n12767) );
  INV_X1 U16033 ( .A(n12770), .ZN(n12774) );
  NAND2_X1 U16034 ( .A1(n13383), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12773) );
  NAND2_X1 U16035 ( .A1(n12771), .A2(n13821), .ZN(n12772) );
  INV_X1 U16036 ( .A(n12775), .ZN(n12776) );
  AOI21_X1 U16037 ( .B1(n12890), .B2(n12891), .A(n12778), .ZN(n12882) );
  NAND2_X1 U16038 ( .A1(n12881), .A2(n12882), .ZN(n12910) );
  OR2_X1 U16039 ( .A1(n12688), .A2(n14500), .ZN(n12783) );
  NAND3_X1 U16040 ( .A1(n21156), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21004) );
  INV_X1 U16041 ( .A(n21004), .ZN(n12779) );
  NAND2_X1 U16042 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12779), .ZN(
        n21002) );
  NAND2_X1 U16043 ( .A1(n21156), .A2(n21002), .ZN(n12780) );
  NOR3_X1 U16044 ( .A1(n21156), .A2(n21157), .A3(n13362), .ZN(n21274) );
  NAND2_X1 U16045 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21274), .ZN(
        n21259) );
  AOI22_X1 U16046 ( .A1(n12781), .A2(n21032), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21329), .ZN(n12782) );
  XNOR2_X2 U16047 ( .A(n14505), .B(n20913), .ZN(n21031) );
  AOI22_X1 U16048 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U16049 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16050 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16051 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U16052 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12795) );
  AOI22_X1 U16053 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U16054 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U16055 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U16056 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12790) );
  NAND4_X1 U16057 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12794) );
  AOI22_X1 U16058 ( .A1(n13394), .A2(n13846), .B1(n13383), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16059 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16060 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12720), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12802) );
  INV_X1 U16061 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21715) );
  AOI22_X1 U16062 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16063 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12800) );
  NAND4_X1 U16064 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n12809) );
  AOI22_X1 U16065 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13177), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U16066 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U16067 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12756), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U16068 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12804) );
  NAND4_X1 U16069 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12808) );
  NAND2_X1 U16070 ( .A1(n13394), .A2(n13845), .ZN(n12811) );
  NAND2_X1 U16071 ( .A1(n13383), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12810) );
  AOI22_X1 U16072 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16073 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16074 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16075 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12812) );
  NAND4_X1 U16076 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12821) );
  AOI22_X1 U16077 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16078 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U16079 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16080 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U16081 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12820) );
  NAND2_X1 U16082 ( .A1(n13394), .A2(n13865), .ZN(n12823) );
  NAND2_X1 U16083 ( .A1(n13383), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12822) );
  AOI22_X1 U16084 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U16085 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U16086 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12829) );
  INV_X1 U16087 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12826) );
  INV_X1 U16088 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12824) );
  OAI22_X1 U16089 ( .A1(n12697), .A2(n12826), .B1(n12825), .B2(n12824), .ZN(
        n12827) );
  INV_X1 U16090 ( .A(n12827), .ZN(n12828) );
  NAND4_X1 U16091 ( .A1(n12831), .A2(n12830), .A3(n12829), .A4(n12828), .ZN(
        n12837) );
  AOI22_X1 U16092 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16093 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16094 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16095 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12832) );
  NAND4_X1 U16096 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12836) );
  NAND2_X1 U16097 ( .A1(n13394), .A2(n13864), .ZN(n12839) );
  NAND2_X1 U16098 ( .A1(n13383), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12838) );
  NAND2_X1 U16099 ( .A1(n12839), .A2(n12838), .ZN(n12840) );
  INV_X1 U16100 ( .A(n13854), .ZN(n12842) );
  NAND2_X1 U16101 ( .A1(n12842), .A2(n9906), .ZN(n12848) );
  INV_X2 U16102 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21201) );
  INV_X2 U16103 ( .A(n10928), .ZN(n13333) );
  INV_X1 U16104 ( .A(n13340), .ZN(n13029) );
  INV_X1 U16105 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21587) );
  NAND2_X1 U16106 ( .A1(n12874), .A2(n21587), .ZN(n12844) );
  NAND2_X1 U16107 ( .A1(n12865), .A2(n12844), .ZN(n20595) );
  NAND2_X1 U16108 ( .A1(n20595), .A2(n12885), .ZN(n12845) );
  OAI21_X1 U16109 ( .B1(n13029), .B2(n21587), .A(n12845), .ZN(n12846) );
  AOI21_X1 U16110 ( .B1(n13333), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12846), .ZN(
        n12847) );
  NAND2_X1 U16111 ( .A1(n12848), .A2(n12847), .ZN(n14891) );
  AOI22_X1 U16112 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U16113 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U16114 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U16115 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12849) );
  NAND4_X1 U16116 ( .A1(n12852), .A2(n12851), .A3(n12850), .A4(n12849), .ZN(
        n12858) );
  AOI22_X1 U16117 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U16118 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16119 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U16120 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12853) );
  NAND4_X1 U16121 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12857) );
  OAI21_X1 U16122 ( .B1(n12858), .B2(n12857), .A(n9906), .ZN(n12862) );
  NAND2_X1 U16123 ( .A1(n13333), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12861) );
  INV_X1 U16124 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14905) );
  XNOR2_X1 U16125 ( .A(n12938), .B(n14905), .ZN(n15653) );
  NAND2_X1 U16126 ( .A1(n15653), .A2(n13332), .ZN(n12860) );
  NAND2_X1 U16127 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12859) );
  NAND4_X1 U16128 ( .A1(n12862), .A2(n12861), .A3(n12860), .A4(n12859), .ZN(
        n14893) );
  AOI22_X1 U16129 ( .A1(n13394), .A2(n13876), .B1(n13383), .B2(
        P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12863) );
  NAND2_X1 U16130 ( .A1(n12865), .A2(n12864), .ZN(n12866) );
  NAND2_X1 U16131 ( .A1(n12938), .A2(n12866), .ZN(n20586) );
  NAND2_X1 U16132 ( .A1(n20586), .A2(n13332), .ZN(n12868) );
  NAND2_X1 U16133 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12867) );
  NAND2_X1 U16134 ( .A1(n12868), .A2(n12867), .ZN(n12869) );
  AOI21_X1 U16135 ( .B1(n13333), .B2(P1_EAX_REG_7__SCAN_IN), .A(n12869), .ZN(
        n12870) );
  INV_X1 U16136 ( .A(n12871), .ZN(n12872) );
  NAND2_X1 U16137 ( .A1(n13844), .A2(n9906), .ZN(n12880) );
  INV_X1 U16138 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20624) );
  INV_X1 U16139 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12873) );
  OAI21_X1 U16140 ( .B1(n12923), .B2(n20624), .A(n12873), .ZN(n12875) );
  NAND2_X1 U16141 ( .A1(n12875), .A2(n12874), .ZN(n20611) );
  NAND2_X1 U16142 ( .A1(n20611), .A2(n12885), .ZN(n12877) );
  NAND2_X1 U16143 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12876) );
  NAND2_X1 U16144 ( .A1(n12877), .A2(n12876), .ZN(n12878) );
  AOI21_X1 U16145 ( .B1(n13333), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12878), .ZN(
        n12879) );
  NAND2_X1 U16146 ( .A1(n12880), .A2(n12879), .ZN(n14572) );
  INV_X1 U16147 ( .A(n12882), .ZN(n12883) );
  NAND2_X1 U16148 ( .A1(n13904), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12921) );
  XNOR2_X1 U16149 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15282) );
  AOI21_X1 U16150 ( .B1(n12885), .B2(n15282), .A(n13340), .ZN(n12887) );
  NAND2_X1 U16151 ( .A1(n13333), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12886) );
  OAI211_X1 U16152 ( .C1(n12921), .C2(n12510), .A(n12887), .B(n12886), .ZN(
        n12888) );
  INV_X1 U16153 ( .A(n12888), .ZN(n12889) );
  NAND2_X1 U16154 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12909) );
  INV_X1 U16155 ( .A(n12890), .ZN(n13825) );
  NAND2_X1 U16156 ( .A1(n20852), .A2(n9906), .ZN(n12897) );
  AOI22_X1 U16157 ( .A1(n13333), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21201), .ZN(n12895) );
  INV_X1 U16158 ( .A(n12921), .ZN(n12893) );
  NAND2_X1 U16159 ( .A1(n12893), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12894) );
  AND2_X1 U16160 ( .A1(n12895), .A2(n12894), .ZN(n12896) );
  NAND2_X1 U16161 ( .A1(n12897), .A2(n12896), .ZN(n14328) );
  NAND2_X1 U16162 ( .A1(n13816), .A2(n12630), .ZN(n12900) );
  NAND2_X1 U16163 ( .A1(n12900), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U16164 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12903) );
  NAND2_X1 U16165 ( .A1(n13333), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12902) );
  OAI211_X1 U16166 ( .C1(n12921), .C2(n12666), .A(n12903), .B(n12902), .ZN(
        n12904) );
  AOI21_X1 U16167 ( .B1(n20882), .B2(n9906), .A(n12904), .ZN(n14166) );
  OR2_X1 U16168 ( .A1(n14167), .A2(n14166), .ZN(n14169) );
  INV_X1 U16169 ( .A(n14166), .ZN(n12905) );
  OR2_X1 U16170 ( .A1(n12905), .A2(n13339), .ZN(n12906) );
  NAND2_X1 U16171 ( .A1(n14169), .A2(n12906), .ZN(n14327) );
  NAND2_X1 U16172 ( .A1(n14328), .A2(n14327), .ZN(n14376) );
  NAND2_X1 U16173 ( .A1(n12908), .A2(n12907), .ZN(n14379) );
  NAND2_X1 U16174 ( .A1(n15911), .A2(n9906), .ZN(n12916) );
  OAI21_X1 U16175 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12911), .A(
        n12923), .ZN(n15275) );
  AOI22_X1 U16176 ( .A1(n12885), .A2(n15275), .B1(n13340), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U16177 ( .A1(n13333), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12912) );
  OAI211_X1 U16178 ( .C1(n12921), .C2(n14500), .A(n12913), .B(n12912), .ZN(
        n12914) );
  INV_X1 U16179 ( .A(n12914), .ZN(n12915) );
  NAND2_X1 U16180 ( .A1(n12916), .A2(n12915), .ZN(n14465) );
  XNOR2_X1 U16181 ( .A(n12917), .B(n10948), .ZN(n13810) );
  INV_X1 U16182 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U16183 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12919) );
  NAND2_X1 U16184 ( .A1(n13333), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12918) );
  OAI211_X1 U16185 ( .C1(n12921), .C2(n12920), .A(n12919), .B(n12918), .ZN(
        n12922) );
  NAND2_X1 U16186 ( .A1(n12922), .A2(n13339), .ZN(n12925) );
  XNOR2_X1 U16187 ( .A(n12923), .B(n20624), .ZN(n20719) );
  NAND2_X1 U16188 ( .A1(n20719), .A2(n12885), .ZN(n12924) );
  NAND2_X1 U16189 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  AOI21_X1 U16190 ( .B1(n13810), .B2(n9906), .A(n12926), .ZN(n14539) );
  AOI22_X1 U16191 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13315), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16192 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16193 ( .A1(n13123), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16194 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12928) );
  NAND4_X1 U16195 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n12928), .ZN(
        n12937) );
  AOI22_X1 U16196 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16197 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16198 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U16199 ( .A1(n13297), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12932) );
  NAND4_X1 U16200 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n12936) );
  OAI21_X1 U16201 ( .B1(n12937), .B2(n12936), .A(n9906), .ZN(n12943) );
  NAND2_X1 U16202 ( .A1(n13333), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12942) );
  XNOR2_X1 U16203 ( .A(n12954), .B(n15257), .ZN(n15643) );
  NAND2_X1 U16204 ( .A1(n15643), .A2(n12885), .ZN(n12941) );
  NAND2_X1 U16205 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12940) );
  AOI22_X1 U16206 ( .A1(n13123), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16207 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16208 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U16209 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12944) );
  NAND4_X1 U16210 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12953) );
  AOI22_X1 U16211 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13315), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16212 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16213 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16214 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12948) );
  NAND4_X1 U16215 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n12948), .ZN(
        n12952) );
  OAI21_X1 U16216 ( .B1(n12953), .B2(n12952), .A(n9906), .ZN(n12958) );
  NAND2_X1 U16217 ( .A1(n13333), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12957) );
  XNOR2_X1 U16218 ( .A(n12960), .B(n12959), .ZN(n15637) );
  NAND2_X1 U16219 ( .A1(n15637), .A2(n13332), .ZN(n12956) );
  NAND2_X1 U16220 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12955) );
  NAND4_X1 U16221 ( .A1(n12958), .A2(n12957), .A3(n12956), .A4(n12955), .ZN(
        n15242) );
  NAND2_X1 U16222 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12961) );
  INV_X1 U16223 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15173) );
  XNOR2_X1 U16224 ( .A(n13047), .B(n15173), .ZN(n15581) );
  AOI22_X1 U16225 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16226 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16227 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16228 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12962) );
  NAND4_X1 U16229 ( .A1(n12965), .A2(n12964), .A3(n12963), .A4(n12962), .ZN(
        n12971) );
  AOI22_X1 U16230 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16231 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16232 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16233 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16234 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12970) );
  OAI21_X1 U16235 ( .B1(n12971), .B2(n12970), .A(n9906), .ZN(n12974) );
  NAND2_X1 U16236 ( .A1(n13333), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12973) );
  NAND2_X1 U16237 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12972) );
  NAND3_X1 U16238 ( .A1(n12974), .A2(n12973), .A3(n12972), .ZN(n12975) );
  AOI21_X1 U16239 ( .B1(n15581), .B2(n13332), .A(n12975), .ZN(n15169) );
  INV_X1 U16240 ( .A(n12976), .ZN(n12978) );
  INV_X1 U16241 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12977) );
  XNOR2_X1 U16242 ( .A(n12978), .B(n12977), .ZN(n15594) );
  NAND2_X1 U16243 ( .A1(n15594), .A2(n12885), .ZN(n12993) );
  AOI22_X1 U16244 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U16245 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U16246 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16247 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12979) );
  NAND4_X1 U16248 ( .A1(n12982), .A2(n12981), .A3(n12980), .A4(n12979), .ZN(
        n12988) );
  AOI22_X1 U16249 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16250 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16251 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16252 ( .A1(n13317), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12983) );
  NAND4_X1 U16253 ( .A1(n12986), .A2(n12985), .A3(n12984), .A4(n12983), .ZN(
        n12987) );
  OAI21_X1 U16254 ( .B1(n12988), .B2(n12987), .A(n9906), .ZN(n12991) );
  NAND2_X1 U16255 ( .A1(n13333), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U16256 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12989) );
  AND3_X1 U16257 ( .A1(n12991), .A2(n12990), .A3(n12989), .ZN(n12992) );
  NAND2_X1 U16258 ( .A1(n12993), .A2(n12992), .ZN(n15182) );
  INV_X1 U16259 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13010) );
  NOR2_X1 U16260 ( .A1(n13028), .A2(n13010), .ZN(n12994) );
  XNOR2_X1 U16261 ( .A(n12994), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15606) );
  NAND2_X1 U16262 ( .A1(n15606), .A2(n13332), .ZN(n13009) );
  AOI22_X1 U16263 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16264 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16265 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U16266 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12995) );
  NAND4_X1 U16267 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n13004) );
  AOI22_X1 U16268 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16269 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16270 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16271 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12999) );
  NAND4_X1 U16272 ( .A1(n13002), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13003) );
  OAI21_X1 U16273 ( .B1(n13004), .B2(n13003), .A(n9906), .ZN(n13007) );
  NAND2_X1 U16274 ( .A1(n13333), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13006) );
  NAND2_X1 U16275 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13005) );
  AND3_X1 U16276 ( .A1(n13007), .A2(n13006), .A3(n13005), .ZN(n13008) );
  NAND2_X1 U16277 ( .A1(n13009), .A2(n13008), .ZN(n15196) );
  XNOR2_X1 U16278 ( .A(n13028), .B(n13010), .ZN(n15617) );
  NAND2_X1 U16279 ( .A1(n15617), .A2(n13332), .ZN(n13025) );
  AOI22_X1 U16280 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12754), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16281 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16282 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U16283 ( .A1(n13317), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13011) );
  NAND4_X1 U16284 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13020) );
  AOI22_X1 U16285 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13315), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U16286 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U16287 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13302), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U16288 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13015) );
  NAND4_X1 U16289 ( .A1(n13018), .A2(n13017), .A3(n13016), .A4(n13015), .ZN(
        n13019) );
  OAI21_X1 U16290 ( .B1(n13020), .B2(n13019), .A(n9906), .ZN(n13023) );
  NAND2_X1 U16291 ( .A1(n13333), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U16292 ( .A1(n13340), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13021) );
  AND3_X1 U16293 ( .A1(n13023), .A2(n13022), .A3(n13021), .ZN(n13024) );
  NAND2_X1 U16294 ( .A1(n13025), .A2(n13024), .ZN(n15216) );
  NAND2_X1 U16295 ( .A1(n13026), .A2(n15232), .ZN(n13027) );
  NAND2_X1 U16296 ( .A1(n13028), .A2(n13027), .ZN(n15627) );
  NAND2_X1 U16297 ( .A1(n15627), .A2(n13332), .ZN(n13032) );
  NOR2_X1 U16298 ( .A1(n13029), .A2(n15232), .ZN(n13030) );
  AOI21_X1 U16299 ( .B1(n13333), .B2(P1_EAX_REG_11__SCAN_IN), .A(n13030), .ZN(
        n13031) );
  AND2_X1 U16300 ( .A1(n13032), .A2(n13031), .ZN(n15166) );
  AOI22_X1 U16301 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16302 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U16303 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16304 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13033) );
  NAND4_X1 U16305 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n13042) );
  AOI22_X1 U16306 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16307 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16308 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U16309 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13037) );
  NAND4_X1 U16310 ( .A1(n13040), .A2(n13039), .A3(n13038), .A4(n13037), .ZN(
        n13041) );
  OR2_X1 U16311 ( .A1(n13042), .A2(n13041), .ZN(n13043) );
  NAND2_X1 U16312 ( .A1(n9906), .A2(n13043), .ZN(n15229) );
  NAND2_X1 U16313 ( .A1(n15166), .A2(n15229), .ZN(n13044) );
  NAND4_X1 U16314 ( .A1(n15182), .A2(n15196), .A3(n15216), .A4(n13044), .ZN(
        n13045) );
  NOR2_X1 U16315 ( .A1(n15169), .A2(n13045), .ZN(n13046) );
  INV_X1 U16316 ( .A(n13049), .ZN(n13050) );
  NAND2_X1 U16317 ( .A1(n13050), .A2(n10437), .ZN(n13051) );
  NAND2_X1 U16318 ( .A1(n13083), .A2(n13051), .ZN(n15568) );
  OR2_X1 U16319 ( .A1(n15568), .A2(n13339), .ZN(n13068) );
  AOI22_X1 U16320 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16321 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16322 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16323 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13053) );
  NAND4_X1 U16324 ( .A1(n13056), .A2(n13055), .A3(n13054), .A4(n13053), .ZN(
        n13062) );
  AOI22_X1 U16325 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16326 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16327 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16328 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13057) );
  NAND4_X1 U16329 ( .A1(n13060), .A2(n13059), .A3(n13058), .A4(n13057), .ZN(
        n13061) );
  NOR2_X1 U16330 ( .A1(n13062), .A2(n13061), .ZN(n13066) );
  NAND2_X1 U16331 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13063) );
  NAND2_X1 U16332 ( .A1(n13339), .A2(n13063), .ZN(n13064) );
  AOI21_X1 U16333 ( .B1(n13333), .B2(P1_EAX_REG_16__SCAN_IN), .A(n13064), .ZN(
        n13065) );
  OAI21_X1 U16334 ( .B1(n13336), .B2(n13066), .A(n13065), .ZN(n13067) );
  XNOR2_X1 U16335 ( .A(n13083), .B(n10440), .ZN(n15559) );
  AOI22_X1 U16336 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U16337 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16338 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U16339 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13069) );
  NAND4_X1 U16340 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        n13078) );
  AOI22_X1 U16341 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16342 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16343 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16344 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13073) );
  NAND4_X1 U16345 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13077) );
  NOR2_X1 U16346 ( .A1(n13078), .A2(n13077), .ZN(n13080) );
  AOI22_X1 U16347 ( .A1(n13333), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13340), .ZN(n13079) );
  OAI21_X1 U16348 ( .B1(n13336), .B2(n13080), .A(n13079), .ZN(n13081) );
  AOI21_X1 U16349 ( .B1(n15559), .B2(n13332), .A(n13081), .ZN(n15140) );
  INV_X1 U16350 ( .A(n15140), .ZN(n13082) );
  NAND2_X1 U16351 ( .A1(n10439), .A2(n10438), .ZN(n13084) );
  NAND2_X1 U16352 ( .A1(n13114), .A2(n13084), .ZN(n15547) );
  AOI22_X1 U16353 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16354 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16355 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16356 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13085) );
  NAND4_X1 U16357 ( .A1(n13088), .A2(n13087), .A3(n13086), .A4(n13085), .ZN(
        n13094) );
  AOI22_X1 U16358 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16359 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16360 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16361 ( .A1(n13317), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13089) );
  NAND4_X1 U16362 ( .A1(n13092), .A2(n13091), .A3(n13090), .A4(n13089), .ZN(
        n13093) );
  NOR2_X1 U16363 ( .A1(n13094), .A2(n13093), .ZN(n13097) );
  OAI21_X1 U16364 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21232), .A(
        n21201), .ZN(n13096) );
  NAND2_X1 U16365 ( .A1(n13333), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n13095) );
  OAI211_X1 U16366 ( .C1(n13336), .C2(n13097), .A(n13096), .B(n13095), .ZN(
        n13098) );
  XNOR2_X1 U16367 ( .A(n13114), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15537) );
  AOI22_X1 U16368 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U16369 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U16370 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16371 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13100) );
  NAND4_X1 U16372 ( .A1(n13103), .A2(n13102), .A3(n13101), .A4(n13100), .ZN(
        n13109) );
  AOI22_X1 U16373 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16374 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16375 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16376 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13104) );
  NAND4_X1 U16377 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13108) );
  OR2_X1 U16378 ( .A1(n13109), .A2(n13108), .ZN(n13112) );
  INV_X1 U16379 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15381) );
  NAND2_X1 U16380 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13110) );
  OAI211_X1 U16381 ( .C1(n10928), .C2(n15381), .A(n13339), .B(n13110), .ZN(
        n13111) );
  AOI21_X1 U16382 ( .B1(n13309), .B2(n13112), .A(n13111), .ZN(n13113) );
  AOI21_X1 U16383 ( .B1(n15537), .B2(n13332), .A(n13113), .ZN(n15113) );
  INV_X1 U16384 ( .A(n13116), .ZN(n13117) );
  NAND2_X1 U16385 ( .A1(n13117), .A2(n10444), .ZN(n13118) );
  NAND2_X1 U16386 ( .A1(n13154), .A2(n13118), .ZN(n15528) );
  AOI22_X1 U16387 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16388 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16389 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12720), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16390 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13119) );
  NAND4_X1 U16391 ( .A1(n13122), .A2(n13121), .A3(n13120), .A4(n13119), .ZN(
        n13130) );
  AOI22_X1 U16392 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16393 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13127) );
  AOI22_X1 U16394 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U16395 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13125) );
  NAND4_X1 U16396 ( .A1(n13128), .A2(n13127), .A3(n13126), .A4(n13125), .ZN(
        n13129) );
  NOR2_X1 U16397 ( .A1(n13130), .A2(n13129), .ZN(n13134) );
  NAND2_X1 U16398 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13131) );
  NAND2_X1 U16399 ( .A1(n13339), .A2(n13131), .ZN(n13132) );
  AOI21_X1 U16400 ( .B1(n13333), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13132), .ZN(
        n13133) );
  OAI21_X1 U16401 ( .B1(n13336), .B2(n13134), .A(n13133), .ZN(n13135) );
  NAND2_X1 U16402 ( .A1(n13136), .A2(n13135), .ZN(n15102) );
  INV_X1 U16403 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15514) );
  INV_X1 U16404 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13137) );
  OAI21_X1 U16405 ( .B1(n13154), .B2(n15514), .A(n13137), .ZN(n13139) );
  NAND2_X1 U16406 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13138) );
  AND2_X1 U16407 ( .A1(n13139), .A2(n13170), .ZN(n15084) );
  AOI22_X1 U16408 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13315), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U16409 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U16410 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U16411 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13140) );
  NAND4_X1 U16412 ( .A1(n13143), .A2(n13142), .A3(n13141), .A4(n13140), .ZN(
        n13149) );
  AOI22_X1 U16413 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16414 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13146) );
  AOI22_X1 U16415 ( .A1(n13123), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U16416 ( .A1(n13297), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13144) );
  NAND4_X1 U16417 ( .A1(n13147), .A2(n13146), .A3(n13145), .A4(n13144), .ZN(
        n13148) );
  OR2_X1 U16418 ( .A1(n13149), .A2(n13148), .ZN(n13152) );
  INV_X1 U16419 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15370) );
  NAND2_X1 U16420 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13150) );
  OAI211_X1 U16421 ( .C1(n10928), .C2(n15370), .A(n13339), .B(n13150), .ZN(
        n13151) );
  AOI21_X1 U16422 ( .B1(n13309), .B2(n13152), .A(n13151), .ZN(n13153) );
  AOI21_X1 U16423 ( .B1(n15084), .B2(n13332), .A(n13153), .ZN(n15075) );
  XNOR2_X1 U16424 ( .A(n13154), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15516) );
  AOI22_X1 U16425 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16426 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16427 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16428 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13155) );
  NAND4_X1 U16429 ( .A1(n13158), .A2(n13157), .A3(n13156), .A4(n13155), .ZN(
        n13164) );
  AOI22_X1 U16430 ( .A1(n13123), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U16431 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13161) );
  AOI22_X1 U16432 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U16433 ( .A1(n13317), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13159) );
  NAND4_X1 U16434 ( .A1(n13162), .A2(n13161), .A3(n13160), .A4(n13159), .ZN(
        n13163) );
  OR2_X1 U16435 ( .A1(n13164), .A2(n13163), .ZN(n13168) );
  INV_X1 U16436 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U16437 ( .A1(n21201), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13165) );
  OAI211_X1 U16438 ( .C1(n10928), .C2(n13166), .A(n13339), .B(n13165), .ZN(
        n13167) );
  AOI21_X1 U16439 ( .B1(n13309), .B2(n13168), .A(n13167), .ZN(n13169) );
  AOI21_X1 U16440 ( .B1(n15516), .B2(n13332), .A(n13169), .ZN(n15097) );
  INV_X1 U16441 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21672) );
  NAND2_X1 U16442 ( .A1(n13170), .A2(n21672), .ZN(n13171) );
  AND2_X1 U16443 ( .A1(n13198), .A2(n13171), .ZN(n15491) );
  NOR2_X1 U16444 ( .A1(n21672), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13172) );
  AOI211_X1 U16445 ( .C1(n13333), .C2(P1_EAX_REG_23__SCAN_IN), .A(n13332), .B(
        n13172), .ZN(n13196) );
  AOI22_X1 U16446 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U16447 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16448 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16449 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13173) );
  NAND4_X1 U16450 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13183) );
  AOI22_X1 U16451 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U16452 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16453 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U16454 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13178) );
  NAND4_X1 U16455 ( .A1(n13181), .A2(n13180), .A3(n13179), .A4(n13178), .ZN(
        n13182) );
  NOR2_X1 U16456 ( .A1(n13183), .A2(n13182), .ZN(n13200) );
  AOI22_X1 U16457 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U16458 ( .A1(n13123), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U16459 ( .A1(n12749), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U16460 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13184) );
  NAND4_X1 U16461 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13193) );
  AOI22_X1 U16462 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16463 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13177), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16464 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U16465 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13188) );
  NAND4_X1 U16466 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13192) );
  NOR2_X1 U16467 ( .A1(n13193), .A2(n13192), .ZN(n13201) );
  XOR2_X1 U16468 ( .A(n13200), .B(n13201), .Z(n13194) );
  NAND2_X1 U16469 ( .A1(n13309), .A2(n13194), .ZN(n13195) );
  AOI22_X1 U16470 ( .A1(n15491), .A2(n13332), .B1(n13196), .B2(n13195), .ZN(
        n15062) );
  INV_X1 U16471 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U16472 ( .A1(n13198), .A2(n13197), .ZN(n13199) );
  NAND2_X1 U16473 ( .A1(n13216), .A2(n13199), .ZN(n15485) );
  NOR2_X1 U16474 ( .A1(n13201), .A2(n13200), .ZN(n13220) );
  AOI22_X1 U16475 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16476 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U16477 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U16478 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13202) );
  NAND4_X1 U16479 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n13211) );
  INV_X1 U16480 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21558) );
  AOI22_X1 U16481 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U16482 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U16483 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U16484 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13206) );
  NAND4_X1 U16485 ( .A1(n13209), .A2(n13208), .A3(n13207), .A4(n13206), .ZN(
        n13210) );
  OR2_X1 U16486 ( .A1(n13211), .A2(n13210), .ZN(n13219) );
  XNOR2_X1 U16487 ( .A(n13220), .B(n13219), .ZN(n13214) );
  AOI21_X1 U16488 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n21201), .A(
        n13332), .ZN(n13213) );
  NAND2_X1 U16489 ( .A1(n13333), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n13212) );
  OAI211_X1 U16490 ( .C1(n13214), .C2(n13336), .A(n13213), .B(n13212), .ZN(
        n13215) );
  OAI21_X1 U16491 ( .B1(n15485), .B2(n13339), .A(n13215), .ZN(n15049) );
  NAND2_X1 U16492 ( .A1(n13216), .A2(n21575), .ZN(n13217) );
  AND2_X1 U16493 ( .A1(n13237), .A2(n13217), .ZN(n15474) );
  NOR2_X1 U16494 ( .A1(n21575), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13218) );
  AOI211_X1 U16495 ( .C1(n13333), .C2(P1_EAX_REG_25__SCAN_IN), .A(n13332), .B(
        n13218), .ZN(n13234) );
  NAND2_X1 U16496 ( .A1(n13220), .A2(n13219), .ZN(n13239) );
  AOI22_X1 U16497 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13315), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U16498 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U16499 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U16500 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13222) );
  NAND4_X1 U16501 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13231) );
  AOI22_X1 U16502 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13229) );
  AOI22_X1 U16503 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13228) );
  AOI22_X1 U16504 ( .A1(n13297), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12756), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16505 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13226) );
  NAND4_X1 U16506 ( .A1(n13229), .A2(n13228), .A3(n13227), .A4(n13226), .ZN(
        n13230) );
  NOR2_X1 U16507 ( .A1(n13231), .A2(n13230), .ZN(n13240) );
  XOR2_X1 U16508 ( .A(n13239), .B(n13240), .Z(n13232) );
  NAND2_X1 U16509 ( .A1(n13232), .A2(n13309), .ZN(n13233) );
  AOI22_X1 U16510 ( .A1(n15474), .A2(n13332), .B1(n13234), .B2(n13233), .ZN(
        n15036) );
  INV_X1 U16511 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U16512 ( .A1(n13237), .A2(n13236), .ZN(n13238) );
  NAND2_X1 U16513 ( .A1(n13256), .A2(n13238), .ZN(n15465) );
  NOR2_X1 U16514 ( .A1(n13240), .A2(n13239), .ZN(n13259) );
  AOI22_X1 U16515 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16516 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16517 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16518 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U16519 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13250) );
  AOI22_X1 U16520 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16521 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16522 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13246) );
  INV_X1 U16523 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n21517) );
  AOI22_X1 U16524 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13245) );
  NAND4_X1 U16525 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13249) );
  OR2_X1 U16526 ( .A1(n13250), .A2(n13249), .ZN(n13258) );
  XNOR2_X1 U16527 ( .A(n13259), .B(n13258), .ZN(n13253) );
  AOI21_X1 U16528 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21201), .A(
        n13332), .ZN(n13252) );
  NAND2_X1 U16529 ( .A1(n13333), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13251) );
  OAI211_X1 U16530 ( .C1(n13253), .C2(n13336), .A(n13252), .B(n13251), .ZN(
        n13254) );
  OAI21_X1 U16531 ( .B1(n15465), .B2(n13339), .A(n13254), .ZN(n15023) );
  INV_X1 U16532 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21419) );
  INV_X1 U16533 ( .A(n13256), .ZN(n13255) );
  AOI21_X1 U16534 ( .B1(n21419), .B2(n13256), .A(n13274), .ZN(n15454) );
  NOR2_X1 U16535 ( .A1(n21419), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13257) );
  AOI211_X1 U16536 ( .C1(n13333), .C2(P1_EAX_REG_27__SCAN_IN), .A(n13332), .B(
        n13257), .ZN(n13273) );
  NAND2_X1 U16537 ( .A1(n13259), .A2(n13258), .ZN(n13278) );
  AOI22_X1 U16538 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12720), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U16539 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U16540 ( .A1(n13297), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U16541 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13260) );
  NAND4_X1 U16542 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        n13270) );
  AOI22_X1 U16543 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13315), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U16544 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12749), .B1(
        n13316), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U16545 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12754), .B1(
        n13177), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U16546 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13124), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13265) );
  NAND4_X1 U16547 ( .A1(n13268), .A2(n13267), .A3(n13266), .A4(n13265), .ZN(
        n13269) );
  NOR2_X1 U16548 ( .A1(n13270), .A2(n13269), .ZN(n13279) );
  XOR2_X1 U16549 ( .A(n13278), .B(n13279), .Z(n13271) );
  NAND2_X1 U16550 ( .A1(n13271), .A2(n13309), .ZN(n13272) );
  AOI22_X1 U16551 ( .A1(n15454), .A2(n13332), .B1(n13273), .B2(n13272), .ZN(
        n15009) );
  INV_X1 U16552 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U16553 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  NAND2_X1 U16554 ( .A1(n13313), .A2(n13277), .ZN(n15448) );
  NOR2_X1 U16555 ( .A1(n13279), .A2(n13278), .ZN(n13296) );
  AOI22_X1 U16556 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U16557 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16558 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16559 ( .A1(n13124), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13280) );
  NAND4_X1 U16560 ( .A1(n13283), .A2(n13282), .A3(n13281), .A4(n13280), .ZN(
        n13289) );
  AOI22_X1 U16561 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U16562 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U16563 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U16564 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13284) );
  NAND4_X1 U16565 ( .A1(n13287), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n13288) );
  OR2_X1 U16566 ( .A1(n13289), .A2(n13288), .ZN(n13295) );
  XNOR2_X1 U16567 ( .A(n13296), .B(n13295), .ZN(n13292) );
  AOI21_X1 U16568 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21201), .A(
        n13332), .ZN(n13291) );
  NAND2_X1 U16569 ( .A1(n13333), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13290) );
  OAI211_X1 U16570 ( .C1(n13292), .C2(n13336), .A(n13291), .B(n13290), .ZN(
        n13293) );
  OAI21_X1 U16571 ( .B1(n15448), .B2(n13339), .A(n13293), .ZN(n14998) );
  XNOR2_X1 U16572 ( .A(n13313), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14888) );
  INV_X1 U16573 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14865) );
  NOR2_X1 U16574 ( .A1(n14865), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13294) );
  AOI211_X1 U16575 ( .C1(n13333), .C2(P1_EAX_REG_29__SCAN_IN), .A(n13332), .B(
        n13294), .ZN(n13312) );
  NAND2_X1 U16576 ( .A1(n13296), .A2(n13295), .ZN(n13328) );
  AOI22_X1 U16577 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U16578 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16579 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U16580 ( .A1(n13177), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13298) );
  NAND4_X1 U16581 ( .A1(n13301), .A2(n13300), .A3(n13299), .A4(n13298), .ZN(
        n13308) );
  AOI22_X1 U16582 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U16583 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16584 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16585 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13124), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13303) );
  NAND4_X1 U16586 ( .A1(n13306), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13307) );
  NOR2_X1 U16587 ( .A1(n13308), .A2(n13307), .ZN(n13329) );
  XOR2_X1 U16588 ( .A(n13328), .B(n13329), .Z(n13310) );
  NAND2_X1 U16589 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  AOI22_X1 U16590 ( .A1(n14888), .A2(n13332), .B1(n13312), .B2(n13311), .ZN(
        n14867) );
  INV_X1 U16591 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13342) );
  XNOR2_X1 U16592 ( .A(n13343), .B(n13342), .ZN(n15433) );
  AOI22_X1 U16593 ( .A1(n13315), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12749), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16594 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13320) );
  AOI22_X1 U16595 ( .A1(n13316), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14483), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U16596 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13317), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13318) );
  NAND4_X1 U16597 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n13327) );
  AOI22_X1 U16598 ( .A1(n13302), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13123), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U16599 ( .A1(n13221), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13297), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16600 ( .A1(n12757), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12618), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16601 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13264), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13322) );
  NAND4_X1 U16602 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13326) );
  NOR2_X1 U16603 ( .A1(n13327), .A2(n13326), .ZN(n13331) );
  NOR2_X1 U16604 ( .A1(n13329), .A2(n13328), .ZN(n13330) );
  XOR2_X1 U16605 ( .A(n13331), .B(n13330), .Z(n13337) );
  AOI21_X1 U16606 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21201), .A(
        n13332), .ZN(n13335) );
  NAND2_X1 U16607 ( .A1(n13333), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13334) );
  OAI211_X1 U16608 ( .C1(n13337), .C2(n13336), .A(n13335), .B(n13334), .ZN(
        n13338) );
  OAI21_X1 U16609 ( .B1(n15433), .B2(n13339), .A(n13338), .ZN(n14985) );
  AOI22_X1 U16610 ( .A1(n13333), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13340), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13341) );
  INV_X1 U16611 ( .A(n14876), .ZN(n13536) );
  INV_X1 U16612 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13344) );
  INV_X1 U16613 ( .A(n14885), .ZN(n13408) );
  NAND2_X1 U16614 ( .A1(n13394), .A2(n14297), .ZN(n13347) );
  NAND2_X1 U16615 ( .A1(n12658), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13346) );
  NAND2_X1 U16616 ( .A1(n13347), .A2(n13346), .ZN(n13356) );
  INV_X1 U16617 ( .A(n13356), .ZN(n13348) );
  NAND2_X1 U16618 ( .A1(n13348), .A2(n14297), .ZN(n13382) );
  MUX2_X1 U16619 ( .A(n13362), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13361) );
  NAND2_X1 U16620 ( .A1(n21199), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13350) );
  XNOR2_X1 U16621 ( .A(n13361), .B(n13360), .ZN(n13397) );
  INV_X1 U16622 ( .A(n13397), .ZN(n13359) );
  NAND2_X1 U16623 ( .A1(n12658), .A2(n14566), .ZN(n13349) );
  NAND2_X1 U16624 ( .A1(n13349), .A2(n17112), .ZN(n13367) );
  OAI21_X1 U16625 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21199), .A(
        n13350), .ZN(n13351) );
  INV_X1 U16626 ( .A(n13351), .ZN(n13352) );
  OAI211_X1 U16627 ( .C1(n14054), .C2(n13916), .A(n13367), .B(n13352), .ZN(
        n13355) );
  NAND2_X1 U16628 ( .A1(n13394), .A2(n13352), .ZN(n13353) );
  NAND2_X1 U16629 ( .A1(n13375), .A2(n13353), .ZN(n13354) );
  OAI211_X1 U16630 ( .C1(n13356), .C2(n13359), .A(n13355), .B(n13354), .ZN(
        n13358) );
  NAND2_X1 U16631 ( .A1(n13356), .A2(n13359), .ZN(n13357) );
  NAND2_X1 U16632 ( .A1(n13361), .A2(n13360), .ZN(n13364) );
  NAND2_X1 U16633 ( .A1(n13362), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13363) );
  NAND2_X1 U16634 ( .A1(n13364), .A2(n13363), .ZN(n13372) );
  XNOR2_X1 U16635 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13371) );
  XNOR2_X1 U16636 ( .A(n13372), .B(n13371), .ZN(n13399) );
  INV_X1 U16637 ( .A(n13399), .ZN(n13368) );
  NAND2_X1 U16638 ( .A1(n13394), .A2(n13368), .ZN(n13365) );
  OAI211_X1 U16639 ( .C1(n13368), .C2(n13380), .A(n13365), .B(n13367), .ZN(
        n13366) );
  INV_X1 U16640 ( .A(n13367), .ZN(n13369) );
  NAND3_X1 U16641 ( .A1(n13369), .A2(n13368), .A3(n13394), .ZN(n13370) );
  NAND2_X1 U16642 ( .A1(n13372), .A2(n13371), .ZN(n13374) );
  NAND2_X1 U16643 ( .A1(n21157), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13373) );
  XNOR2_X1 U16644 ( .A(n13379), .B(n13378), .ZN(n13398) );
  NAND2_X1 U16645 ( .A1(n13391), .A2(n13398), .ZN(n13376) );
  NOR2_X1 U16646 ( .A1(n14500), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13377) );
  AND2_X1 U16647 ( .A1(n13390), .A2(n13388), .ZN(n13400) );
  NAND2_X1 U16648 ( .A1(n13400), .A2(n13380), .ZN(n13381) );
  INV_X1 U16649 ( .A(n13382), .ZN(n13385) );
  AND2_X1 U16650 ( .A1(n13383), .A2(n13400), .ZN(n13384) );
  AOI22_X1 U16651 ( .A1(n13385), .A2(n13384), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17176), .ZN(n13386) );
  NAND2_X1 U16652 ( .A1(n13387), .A2(n13386), .ZN(n13393) );
  NAND2_X1 U16653 ( .A1(n20783), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13389) );
  NAND2_X1 U16654 ( .A1(n13391), .A2(n13402), .ZN(n13392) );
  NOR4_X1 U16655 ( .A1(n13400), .A2(n13399), .A3(n13398), .A4(n13397), .ZN(
        n13401) );
  OR2_X1 U16656 ( .A1(n13402), .A2(n13401), .ZN(n14060) );
  INV_X1 U16657 ( .A(n14060), .ZN(n13403) );
  NAND2_X1 U16658 ( .A1(n14061), .A2(n13403), .ZN(n14050) );
  AND2_X1 U16659 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n17176), .ZN(n13405) );
  INV_X1 U16660 ( .A(n17172), .ZN(n21413) );
  NAND2_X1 U16661 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21413), .ZN(n17120) );
  INV_X1 U16662 ( .A(n17120), .ZN(n13404) );
  AOI22_X1 U16663 ( .A1(n12885), .A2(n13405), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n13404), .ZN(n13406) );
  NAND2_X1 U16664 ( .A1(n20781), .A2(n13406), .ZN(n13407) );
  OR2_X2 U16665 ( .A1(n21407), .A2(n13407), .ZN(n20638) );
  NAND2_X1 U16666 ( .A1(n13409), .A2(n21332), .ZN(n14298) );
  NAND2_X1 U16667 ( .A1(n17112), .A2(n14298), .ZN(n13903) );
  AND2_X1 U16668 ( .A1(n21409), .A2(n21232), .ZN(n17110) );
  NAND3_X1 U16669 ( .A1(n15281), .A2(P1_REIP_REG_3__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20632) );
  AND2_X1 U16670 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n13410) );
  NAND2_X1 U16671 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .ZN(n13414) );
  AND2_X1 U16672 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n13415) );
  NAND2_X1 U16673 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n13416) );
  AND2_X1 U16674 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15159) );
  NAND2_X1 U16675 ( .A1(n15159), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n13411) );
  AND2_X1 U16676 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n13418) );
  NAND2_X1 U16677 ( .A1(n15127), .A2(n13418), .ZN(n15100) );
  NAND2_X1 U16678 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n13412) );
  INV_X1 U16679 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21373) );
  AND2_X1 U16680 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15032) );
  NAND2_X1 U16681 ( .A1(n15032), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15017) );
  INV_X1 U16682 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15452) );
  INV_X1 U16683 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21386) );
  INV_X1 U16684 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15431) );
  NAND2_X1 U16685 ( .A1(n20645), .A2(n20638), .ZN(n20585) );
  INV_X1 U16686 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21374) );
  INV_X1 U16687 ( .A(n20638), .ZN(n13413) );
  NAND2_X1 U16688 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n15270) );
  NOR4_X1 U16689 ( .A1(n13413), .A2(n21353), .A3(n21398), .A4(n15270), .ZN(
        n20615) );
  NAND3_X1 U16690 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20615), .ZN(n20584) );
  INV_X1 U16691 ( .A(n13416), .ZN(n15154) );
  AND3_X1 U16692 ( .A1(n15154), .A2(n15159), .A3(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n13417) );
  NAND2_X1 U16693 ( .A1(n13418), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n13419) );
  INV_X1 U16694 ( .A(n15091), .ZN(n13420) );
  AND2_X1 U16695 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n13421) );
  NAND2_X1 U16696 ( .A1(n15013), .A2(n13421), .ZN(n14886) );
  NOR2_X1 U16697 ( .A1(n21386), .A2(n14886), .ZN(n13422) );
  NAND2_X1 U16698 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n13422), .ZN(n13423) );
  NAND2_X1 U16699 ( .A1(n20585), .A2(n13423), .ZN(n14995) );
  NAND2_X1 U16700 ( .A1(n13430), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13531) );
  INV_X1 U16701 ( .A(n13531), .ZN(n13424) );
  NOR2_X1 U16702 ( .A1(n13425), .A2(n13424), .ZN(n13426) );
  AND2_X2 U16703 ( .A1(n13533), .A2(n13426), .ZN(n20641) );
  AOI22_X1 U16704 ( .A1(n20641), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20608), .ZN(n13427) );
  OAI21_X1 U16705 ( .B1(n14995), .B2(n10683), .A(n13427), .ZN(n13428) );
  AND2_X1 U16706 ( .A1(n13433), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13431) );
  AOI21_X1 U16707 ( .B1(n14158), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13431), .ZN(
        n14989) );
  NAND2_X2 U16708 ( .A1(n12639), .A2(n14163), .ZN(n13521) );
  OR2_X1 U16709 ( .A1(n14163), .A2(n13522), .ZN(n13460) );
  NAND2_X1 U16710 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13433), .ZN(
        n13434) );
  AND2_X1 U16711 ( .A1(n13460), .A2(n13434), .ZN(n13435) );
  NAND2_X1 U16712 ( .A1(n13436), .A2(n13435), .ZN(n13439) );
  NAND2_X1 U16713 ( .A1(n13522), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13438) );
  INV_X1 U16714 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14170) );
  NAND2_X1 U16715 ( .A1(n13454), .A2(n14170), .ZN(n13437) );
  NAND2_X1 U16716 ( .A1(n13438), .A2(n13437), .ZN(n14159) );
  XNOR2_X1 U16717 ( .A(n13439), .B(n14159), .ZN(n14330) );
  NAND2_X1 U16718 ( .A1(n14330), .A2(n14163), .ZN(n14332) );
  NAND2_X1 U16719 ( .A1(n14332), .A2(n13439), .ZN(n14380) );
  OR2_X1 U16720 ( .A1(n13521), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13444) );
  INV_X1 U16721 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20754) );
  NAND2_X1 U16722 ( .A1(n13522), .A2(n20754), .ZN(n13442) );
  INV_X1 U16723 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U16724 ( .A1(n14163), .A2(n13440), .ZN(n13441) );
  NAND3_X1 U16725 ( .A1(n13442), .A2(n13454), .A3(n13441), .ZN(n13443) );
  AND2_X1 U16726 ( .A1(n13444), .A2(n13443), .ZN(n14381) );
  INV_X1 U16727 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13445) );
  NAND2_X1 U16728 ( .A1(n13502), .A2(n13445), .ZN(n13448) );
  NAND2_X1 U16729 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13446) );
  OAI211_X1 U16730 ( .C1(n13433), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13518), .B(
        n13446), .ZN(n13447) );
  OR2_X1 U16731 ( .A1(n13521), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n13453) );
  INV_X1 U16732 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20733) );
  NAND2_X1 U16733 ( .A1(n13518), .A2(n20733), .ZN(n13451) );
  INV_X1 U16734 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U16735 ( .A1(n14163), .A2(n13449), .ZN(n13450) );
  NAND3_X1 U16736 ( .A1(n13451), .A2(n13528), .A3(n13450), .ZN(n13452) );
  NAND2_X1 U16737 ( .A1(n13453), .A2(n13452), .ZN(n14542) );
  NAND2_X1 U16738 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13455) );
  OAI211_X1 U16739 ( .C1(n13433), .C2(P1_EBX_REG_5__SCAN_IN), .A(n13518), .B(
        n13455), .ZN(n13456) );
  OAI21_X1 U16740 ( .B1(n13520), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13456), .ZN(
        n17152) );
  MUX2_X1 U16741 ( .A(n13520), .B(n13528), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13458) );
  OR2_X1 U16742 ( .A1(n14158), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13457) );
  NAND2_X1 U16743 ( .A1(n13458), .A2(n13457), .ZN(n15325) );
  INV_X1 U16744 ( .A(n15325), .ZN(n13463) );
  MUX2_X1 U16745 ( .A(n13521), .B(n13518), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13462) );
  NAND2_X1 U16746 ( .A1(n13433), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13459) );
  AND2_X1 U16747 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  NAND2_X1 U16748 ( .A1(n13462), .A2(n13461), .ZN(n14618) );
  OR2_X1 U16749 ( .A1(n13521), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13467) );
  INV_X1 U16750 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15884) );
  NAND2_X1 U16751 ( .A1(n13518), .A2(n15884), .ZN(n13465) );
  INV_X1 U16752 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U16753 ( .A1(n14163), .A2(n14898), .ZN(n13464) );
  NAND3_X1 U16754 ( .A1(n13465), .A2(n13528), .A3(n13464), .ZN(n13466) );
  MUX2_X1 U16755 ( .A(n13520), .B(n13528), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13469) );
  OR2_X1 U16756 ( .A1(n14158), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13468) );
  AND2_X2 U16757 ( .A1(n14894), .A2(n14730), .ZN(n15251) );
  OR2_X1 U16758 ( .A1(n13521), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13474) );
  INV_X1 U16759 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15633) );
  NAND2_X1 U16760 ( .A1(n13522), .A2(n15633), .ZN(n13472) );
  INV_X1 U16761 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13470) );
  NAND2_X1 U16762 ( .A1(n14163), .A2(n13470), .ZN(n13471) );
  NAND3_X1 U16763 ( .A1(n13472), .A2(n13528), .A3(n13471), .ZN(n13473) );
  NAND2_X1 U16764 ( .A1(n13474), .A2(n13473), .ZN(n15250) );
  MUX2_X1 U16765 ( .A(n13520), .B(n13528), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13475) );
  OAI21_X1 U16766 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14158), .A(
        n13475), .ZN(n15230) );
  MUX2_X1 U16767 ( .A(n13521), .B(n13518), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13477) );
  NAND2_X1 U16768 ( .A1(n13433), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13476) );
  NAND2_X1 U16769 ( .A1(n13477), .A2(n13476), .ZN(n15218) );
  INV_X1 U16770 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15316) );
  NAND2_X1 U16771 ( .A1(n13502), .A2(n15316), .ZN(n13480) );
  NAND2_X1 U16772 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13478) );
  OAI211_X1 U16773 ( .C1(n13433), .C2(P1_EBX_REG_13__SCAN_IN), .A(n13522), .B(
        n13478), .ZN(n13479) );
  NAND2_X1 U16774 ( .A1(n15218), .A2(n15200), .ZN(n13481) );
  OR2_X1 U16775 ( .A1(n13521), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n13484) );
  INV_X1 U16776 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21709) );
  NAND2_X1 U16777 ( .A1(n13518), .A2(n21709), .ZN(n13482) );
  OAI211_X1 U16778 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n13433), .A(n13482), .B(
        n13528), .ZN(n13483) );
  NAND2_X1 U16779 ( .A1(n13484), .A2(n13483), .ZN(n15183) );
  NAND2_X1 U16780 ( .A1(n15202), .A2(n15183), .ZN(n15185) );
  NAND2_X1 U16781 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13485) );
  OAI211_X1 U16782 ( .C1(n13433), .C2(P1_EBX_REG_15__SCAN_IN), .A(n13522), .B(
        n13485), .ZN(n13486) );
  OAI21_X1 U16783 ( .B1(n13520), .B2(P1_EBX_REG_15__SCAN_IN), .A(n13486), .ZN(
        n15170) );
  INV_X1 U16784 ( .A(n15170), .ZN(n13487) );
  OR2_X1 U16785 ( .A1(n13521), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n13491) );
  INV_X1 U16786 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15806) );
  NAND2_X1 U16787 ( .A1(n13518), .A2(n15806), .ZN(n13489) );
  OAI211_X1 U16788 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n13433), .A(n13489), .B(
        n13528), .ZN(n13490) );
  INV_X1 U16789 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21516) );
  NAND2_X1 U16790 ( .A1(n13502), .A2(n21516), .ZN(n13494) );
  NAND2_X1 U16791 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13492) );
  OAI211_X1 U16792 ( .C1(n13433), .C2(P1_EBX_REG_17__SCAN_IN), .A(n13518), .B(
        n13492), .ZN(n13493) );
  MUX2_X1 U16793 ( .A(n13521), .B(n13518), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13496) );
  NAND2_X1 U16794 ( .A1(n13433), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13495) );
  NAND2_X1 U16795 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13497) );
  OAI211_X1 U16796 ( .C1(n13433), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13518), .B(
        n13497), .ZN(n13498) );
  OAI21_X1 U16797 ( .B1(n13520), .B2(P1_EBX_REG_19__SCAN_IN), .A(n13498), .ZN(
        n15119) );
  OR2_X1 U16798 ( .A1(n13521), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n13501) );
  INV_X1 U16799 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15509) );
  NAND2_X1 U16800 ( .A1(n13518), .A2(n15509), .ZN(n13499) );
  OAI211_X1 U16801 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n13433), .A(n13499), .B(
        n13528), .ZN(n13500) );
  INV_X1 U16802 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15308) );
  NAND2_X1 U16803 ( .A1(n13502), .A2(n15308), .ZN(n13505) );
  NAND2_X1 U16804 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13503) );
  OAI211_X1 U16805 ( .C1(n13433), .C2(P1_EBX_REG_21__SCAN_IN), .A(n13522), .B(
        n13503), .ZN(n13504) );
  AND2_X1 U16806 ( .A1(n13505), .A2(n13504), .ZN(n15094) );
  OR2_X1 U16807 ( .A1(n13521), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13508) );
  INV_X1 U16808 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U16809 ( .A1(n13522), .A2(n15499), .ZN(n13506) );
  OAI211_X1 U16810 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n13433), .A(n13506), .B(
        n13528), .ZN(n13507) );
  NAND2_X1 U16811 ( .A1(n13508), .A2(n13507), .ZN(n15080) );
  NAND2_X1 U16812 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13509) );
  OAI211_X1 U16813 ( .C1(n13433), .C2(P1_EBX_REG_23__SCAN_IN), .A(n13518), .B(
        n13509), .ZN(n13510) );
  OAI21_X1 U16814 ( .B1(n13520), .B2(P1_EBX_REG_23__SCAN_IN), .A(n13510), .ZN(
        n15068) );
  NOR2_X2 U16815 ( .A1(n15067), .A2(n15068), .ZN(n15070) );
  MUX2_X1 U16816 ( .A(n13521), .B(n13522), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13512) );
  NAND2_X1 U16817 ( .A1(n13433), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13511) );
  NAND2_X1 U16818 ( .A1(n13512), .A2(n13511), .ZN(n15050) );
  NAND2_X1 U16819 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13513) );
  OAI211_X1 U16820 ( .C1(n13433), .C2(P1_EBX_REG_25__SCAN_IN), .A(n13518), .B(
        n13513), .ZN(n13514) );
  OAI21_X1 U16821 ( .B1(n13520), .B2(P1_EBX_REG_25__SCAN_IN), .A(n13514), .ZN(
        n15039) );
  MUX2_X1 U16822 ( .A(n13521), .B(n13518), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13516) );
  NAND2_X1 U16823 ( .A1(n13433), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13515) );
  AND2_X1 U16824 ( .A1(n13516), .A2(n13515), .ZN(n15026) );
  NAND2_X1 U16825 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13517) );
  OAI211_X1 U16826 ( .C1(n13433), .C2(P1_EBX_REG_27__SCAN_IN), .A(n13518), .B(
        n13517), .ZN(n13519) );
  OAI21_X1 U16827 ( .B1(n13520), .B2(P1_EBX_REG_27__SCAN_IN), .A(n13519), .ZN(
        n15010) );
  OR2_X1 U16828 ( .A1(n13521), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13525) );
  INV_X1 U16829 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U16830 ( .A1(n13522), .A2(n15444), .ZN(n13523) );
  OAI211_X1 U16831 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n13433), .A(n13523), .B(
        n13528), .ZN(n13524) );
  NAND2_X1 U16832 ( .A1(n13525), .A2(n13524), .ZN(n14999) );
  INV_X1 U16833 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14874) );
  NAND2_X1 U16834 ( .A1(n14163), .A2(n14874), .ZN(n13527) );
  OR2_X1 U16835 ( .A1(n14158), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13526) );
  NAND2_X1 U16836 ( .A1(n13526), .A2(n13527), .ZN(n14987) );
  MUX2_X1 U16837 ( .A(n13527), .B(n14987), .S(n13528), .Z(n14872) );
  OR2_X2 U16838 ( .A1(n14871), .A2(n14872), .ZN(n14986) );
  AOI22_X1 U16839 ( .A1(n14158), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13433), .ZN(n13529) );
  INV_X1 U16840 ( .A(n15300), .ZN(n13534) );
  NOR2_X1 U16841 ( .A1(n13531), .A2(n17110), .ZN(n13532) );
  OAI211_X1 U16842 ( .C1(n13536), .C2(n15269), .A(n10929), .B(n13535), .ZN(
        P1_U2809) );
  INV_X1 U16843 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n21506) );
  NOR2_X1 U16844 ( .A1(n13593), .A2(n21506), .ZN(n13563) );
  NOR2_X1 U16845 ( .A1(n13593), .A2(n16027), .ZN(n13571) );
  INV_X1 U16846 ( .A(n13571), .ZN(n13537) );
  NAND2_X2 U16847 ( .A1(n13570), .A2(n13537), .ZN(n13574) );
  NOR2_X2 U16848 ( .A1(n13574), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13565) );
  INV_X1 U16849 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16292) );
  NAND2_X1 U16850 ( .A1(n13565), .A2(n16292), .ZN(n13578) );
  INV_X1 U16851 ( .A(n13578), .ZN(n13538) );
  NAND2_X1 U16852 ( .A1(n13538), .A2(n16288), .ZN(n13580) );
  NAND2_X1 U16853 ( .A1(n19879), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13540) );
  INV_X1 U16854 ( .A(n13540), .ZN(n13541) );
  NAND2_X1 U16855 ( .A1(n13580), .A2(n13541), .ZN(n13542) );
  NAND2_X1 U16856 ( .A1(n13635), .A2(n13542), .ZN(n15974) );
  INV_X1 U16857 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16719) );
  INV_X1 U16858 ( .A(n13543), .ZN(n16547) );
  AND2_X1 U16859 ( .A1(n16554), .A2(n13544), .ZN(n13545) );
  NAND4_X1 U16860 ( .A1(n13546), .A2(n16547), .A3(n13545), .A4(n16568), .ZN(
        n13548) );
  NOR2_X1 U16861 ( .A1(n13548), .A2(n13547), .ZN(n13552) );
  INV_X1 U16862 ( .A(n13554), .ZN(n13556) );
  NAND3_X1 U16863 ( .A1(n16553), .A2(n16567), .A3(n16573), .ZN(n13555) );
  NOR3_X1 U16864 ( .A1(n13557), .A2(n13556), .A3(n13555), .ZN(n13559) );
  AOI21_X1 U16865 ( .B1(n13563), .B2(n13562), .A(n13570), .ZN(n16047) );
  AOI21_X1 U16866 ( .B1(n16047), .B2(n13750), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16523) );
  INV_X1 U16867 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16008) );
  NOR2_X1 U16868 ( .A1(n13593), .A2(n16008), .ZN(n13564) );
  AOI21_X1 U16869 ( .B1(n13574), .B2(n13564), .A(n13576), .ZN(n13566) );
  INV_X1 U16870 ( .A(n13565), .ZN(n13568) );
  AND2_X1 U16871 ( .A1(n13566), .A2(n13568), .ZN(n16019) );
  NAND2_X1 U16872 ( .A1(n16019), .A2(n13750), .ZN(n16507) );
  INV_X1 U16873 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16511) );
  NOR2_X1 U16874 ( .A1(n13593), .A2(n16292), .ZN(n13567) );
  AOI21_X1 U16875 ( .B1(n13568), .B2(n13567), .A(n13576), .ZN(n13569) );
  NAND2_X1 U16876 ( .A1(n13578), .A2(n13569), .ZN(n15998) );
  INV_X1 U16877 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16732) );
  NAND2_X1 U16878 ( .A1(n13572), .A2(n13571), .ZN(n13573) );
  NAND2_X1 U16879 ( .A1(n13574), .A2(n13573), .ZN(n16033) );
  OR2_X1 U16880 ( .A1(n16033), .A2(n11378), .ZN(n13575) );
  XNOR2_X1 U16881 ( .A(n13575), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16518) );
  NOR2_X1 U16882 ( .A1(n13593), .A2(n16288), .ZN(n13577) );
  AOI21_X1 U16883 ( .B1(n13578), .B2(n13577), .A(n13576), .ZN(n13579) );
  AND2_X1 U16884 ( .A1(n13580), .A2(n13579), .ZN(n13582) );
  AOI21_X1 U16885 ( .B1(n13582), .B2(n13750), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13581) );
  INV_X1 U16886 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13787) );
  NAND2_X1 U16887 ( .A1(n13750), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13586) );
  OAI21_X1 U16888 ( .B1(n16507), .B2(n16511), .A(n13775), .ZN(n13587) );
  NAND2_X1 U16889 ( .A1(n13589), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16495) );
  NAND2_X1 U16890 ( .A1(n16495), .A2(n13590), .ZN(n16484) );
  INV_X1 U16891 ( .A(n16484), .ZN(n13591) );
  NAND2_X1 U16892 ( .A1(n16486), .A2(n16719), .ZN(n13633) );
  INV_X1 U16893 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n13592) );
  NOR2_X1 U16894 ( .A1(n13593), .A2(n13592), .ZN(n13634) );
  INV_X1 U16895 ( .A(n13634), .ZN(n13594) );
  XOR2_X1 U16896 ( .A(n13594), .B(n13635), .Z(n15957) );
  INV_X1 U16897 ( .A(n15957), .ZN(n13595) );
  NAND2_X1 U16898 ( .A1(n13595), .A2(n13750), .ZN(n14909) );
  XNOR2_X1 U16899 ( .A(n14909), .B(n14927), .ZN(n13596) );
  AND3_X1 U16900 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13598) );
  AND2_X1 U16901 ( .A1(n13599), .A2(n13598), .ZN(n13602) );
  OAI21_X1 U16902 ( .B1(n15966), .B2(n13607), .A(n13606), .ZN(n16274) );
  INV_X1 U16903 ( .A(n16274), .ZN(n16481) );
  AOI22_X1 U16904 ( .A1(n9687), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13609) );
  NAND2_X1 U16905 ( .A1(n13763), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U16906 ( .A1(n9687), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13611) );
  NAND2_X1 U16907 ( .A1(n13763), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n13610) );
  NAND2_X1 U16908 ( .A1(n13611), .A2(n13610), .ZN(n16026) );
  NAND2_X1 U16909 ( .A1(n16024), .A2(n16026), .ZN(n16014) );
  AOI22_X1 U16910 ( .A1(n9687), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U16911 ( .A1(n13763), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13612) );
  NOR2_X2 U16912 ( .A1(n16014), .A2(n16015), .ZN(n15987) );
  AOI22_X1 U16913 ( .A1(n9687), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U16914 ( .A1(n13763), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n13614) );
  INV_X1 U16915 ( .A(n15989), .ZN(n13616) );
  AOI22_X1 U16916 ( .A1(n9687), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13618) );
  NAND2_X1 U16917 ( .A1(n13763), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U16918 ( .A1(n13618), .A2(n13617), .ZN(n13782) );
  AOI222_X1 U16919 ( .A1(n13763), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n9687), 
        .B2(P2_EAX_REG_27__SCAN_IN), .C1(n13649), .C2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15967) );
  INV_X1 U16920 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14233) );
  INV_X1 U16921 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20508) );
  OAI222_X1 U16922 ( .A1(n14233), .A2(n13621), .B1(n20508), .B2(n13620), .C1(
        n13619), .C2(n14927), .ZN(n13623) );
  INV_X1 U16923 ( .A(n13624), .ZN(n13625) );
  NAND2_X1 U16924 ( .A1(n16910), .A2(n13625), .ZN(n16764) );
  NAND2_X1 U16925 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16755) );
  NOR3_X1 U16926 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16755), .ZN(n16742) );
  NOR2_X1 U16927 ( .A1(n16959), .A2(n17188), .ZN(n13769) );
  INV_X1 U16928 ( .A(n16755), .ZN(n13626) );
  OAI21_X1 U16929 ( .B1(n13769), .B2(n13626), .A(n16754), .ZN(n16744) );
  AND2_X1 U16930 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13627) );
  INV_X1 U16931 ( .A(n13769), .ZN(n16899) );
  NAND2_X1 U16932 ( .A1(n13653), .A2(n16899), .ZN(n16720) );
  NOR2_X1 U16933 ( .A1(n13784), .A2(n10553), .ZN(n13772) );
  NAND2_X1 U16934 ( .A1(n13772), .A2(n16719), .ZN(n16718) );
  NAND2_X1 U16935 ( .A1(n16720), .A2(n16718), .ZN(n14930) );
  OR2_X1 U16936 ( .A1(n16706), .A2(n20508), .ZN(n16477) );
  INV_X1 U16937 ( .A(n16477), .ZN(n13629) );
  INV_X1 U16938 ( .A(n13772), .ZN(n14924) );
  NOR3_X1 U16939 ( .A1(n14924), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16719), .ZN(n13628) );
  AOI211_X1 U16940 ( .C1(n14930), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n13629), .B(n13628), .ZN(n13630) );
  OAI21_X1 U16941 ( .B1(n16376), .B2(n17180), .A(n13630), .ZN(n13631) );
  INV_X1 U16942 ( .A(n13631), .ZN(n13632) );
  INV_X1 U16943 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14926) );
  INV_X1 U16944 ( .A(n16486), .ZN(n13639) );
  AND2_X1 U16945 ( .A1(n13633), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14910) );
  NAND2_X1 U16946 ( .A1(n19879), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13636) );
  OAI21_X1 U16947 ( .B1(n13640), .B2(n11378), .A(n14926), .ZN(n14911) );
  NAND2_X1 U16948 ( .A1(n14927), .A2(n16719), .ZN(n14908) );
  AOI21_X1 U16949 ( .B1(n13750), .B2(n14908), .A(n16484), .ZN(n13642) );
  INV_X1 U16950 ( .A(n13640), .ZN(n15948) );
  NAND3_X1 U16951 ( .A1(n15948), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13641), .ZN(n14912) );
  OAI21_X1 U16952 ( .B1(n13642), .B2(n15957), .A(n14912), .ZN(n13643) );
  NAND2_X1 U16953 ( .A1(n19879), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U16954 ( .A1(n13725), .A2(n13750), .ZN(n13646) );
  NAND2_X1 U16955 ( .A1(n13646), .A2(n10555), .ZN(n13744) );
  NAND2_X1 U16956 ( .A1(n9733), .A2(n13744), .ZN(n13647) );
  AOI222_X1 U16957 ( .A1(n13763), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n9687), 
        .B2(P2_EAX_REG_29__SCAN_IN), .C1(n13649), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U16958 ( .A1(n9687), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13649), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13651) );
  NAND2_X1 U16959 ( .A1(n13763), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13650) );
  NAND2_X1 U16960 ( .A1(n13651), .A2(n13650), .ZN(n13762) );
  OR2_X1 U16961 ( .A1(n16360), .A2(n17180), .ZN(n13657) );
  NAND3_X1 U16962 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13766) );
  NOR2_X1 U16963 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13766), .ZN(
        n13655) );
  INV_X1 U16964 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13652) );
  NOR2_X1 U16965 ( .A1(n16706), .A2(n13652), .ZN(n13659) );
  NOR3_X1 U16966 ( .A1(n9811), .A2(n13769), .A3(n10555), .ZN(n13654) );
  AOI211_X1 U16967 ( .C1(n13772), .C2(n13655), .A(n13659), .B(n13654), .ZN(
        n13656) );
  NAND2_X1 U16968 ( .A1(n13730), .A2(n16970), .ZN(n13658) );
  NAND2_X1 U16969 ( .A1(n13730), .A2(n16715), .ZN(n13663) );
  INV_X1 U16970 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15970) );
  XNOR2_X1 U16971 ( .A(n13711), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13731) );
  AOI21_X1 U16972 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n13659), .ZN(n13660) );
  OAI21_X1 U16973 ( .B1(n13731), .B2(n16710), .A(n13660), .ZN(n13661) );
  INV_X1 U16974 ( .A(n13661), .ZN(n13662) );
  AOI21_X1 U16975 ( .B1(n13665), .B2(n13691), .A(n13694), .ZN(n13666) );
  INV_X1 U16976 ( .A(n13666), .ZN(n19765) );
  INV_X1 U16977 ( .A(n13688), .ZN(n13667) );
  OAI21_X1 U16978 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n13667), .A(
        n10724), .ZN(n16558) );
  INV_X1 U16979 ( .A(n16558), .ZN(n13690) );
  AOI21_X1 U16980 ( .B1(n21703), .B2(n13686), .A(n13689), .ZN(n16578) );
  NAND2_X1 U16981 ( .A1(n21718), .A2(n13684), .ZN(n13668) );
  AND2_X1 U16982 ( .A1(n13668), .A2(n10730), .ZN(n16597) );
  NOR2_X1 U16983 ( .A1(n13683), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13669) );
  NOR2_X1 U16984 ( .A1(n13685), .A2(n13669), .ZN(n16633) );
  NOR2_X1 U16985 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n13679), .ZN(
        n13670) );
  NOR2_X1 U16986 ( .A1(n13681), .A2(n13670), .ZN(n16655) );
  OAI21_X1 U16987 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13671), .ZN(n16244) );
  AND2_X1 U16988 ( .A1(n17015), .A2(n16244), .ZN(n16229) );
  INV_X1 U16989 ( .A(n13674), .ZN(n13673) );
  NAND2_X1 U16990 ( .A1(n11591), .A2(n13671), .ZN(n13672) );
  NAND2_X1 U16991 ( .A1(n13673), .A2(n13672), .ZN(n16709) );
  NOR2_X1 U16992 ( .A1(n13674), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13675) );
  NOR2_X1 U16993 ( .A1(n13677), .A2(n13675), .ZN(n19802) );
  NOR2_X1 U16994 ( .A1(n13677), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13678) );
  NOR2_X1 U16995 ( .A1(n13676), .A2(n13678), .ZN(n16670) );
  INV_X1 U16996 ( .A(n13679), .ZN(n13680) );
  OAI21_X1 U16997 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13676), .A(
        n13680), .ZN(n16663) );
  OR2_X1 U16998 ( .A1(n16655), .A2(n16193), .ZN(n16182) );
  NOR2_X1 U16999 ( .A1(n13681), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13682) );
  NOR2_X1 U17000 ( .A1(n13683), .A2(n13682), .ZN(n16641) );
  OAI21_X1 U17001 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13685), .A(
        n13684), .ZN(n16616) );
  OAI21_X1 U17002 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13687), .A(
        n13686), .ZN(n16590) );
  NAND2_X1 U17003 ( .A1(n16147), .A2(n16590), .ZN(n16134) );
  NOR2_X1 U17004 ( .A1(n16578), .A2(n16134), .ZN(n16121) );
  OAI21_X1 U17005 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13689), .A(
        n13688), .ZN(n16565) );
  NAND2_X1 U17006 ( .A1(n16121), .A2(n16565), .ZN(n16111) );
  NOR2_X1 U17007 ( .A1(n13690), .A2(n16111), .ZN(n19777) );
  OAI21_X1 U17008 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13692), .A(
        n13691), .ZN(n19779) );
  AND2_X1 U17009 ( .A1(n19777), .A2(n19779), .ZN(n19766) );
  NAND2_X1 U17010 ( .A1(n19765), .A2(n19766), .ZN(n19763) );
  INV_X1 U17011 ( .A(n19763), .ZN(n16096) );
  OAI21_X1 U17012 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13694), .A(
        n13693), .ZN(n16534) );
  NAND2_X1 U17013 ( .A1(n16096), .A2(n16534), .ZN(n16086) );
  NOR2_X1 U17014 ( .A1(n16085), .A2(n16086), .ZN(n16062) );
  AND2_X1 U17015 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  OR2_X1 U17016 ( .A1(n13697), .A2(n13700), .ZN(n16528) );
  NAND2_X1 U17017 ( .A1(n13711), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13699) );
  INV_X1 U17018 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13698) );
  INV_X1 U17019 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13768) );
  NOR2_X1 U17020 ( .A1(n13700), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13701) );
  OR2_X1 U17021 ( .A1(n13702), .A2(n13701), .ZN(n16519) );
  OR2_X1 U17022 ( .A1(n13702), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13703) );
  AND2_X1 U17023 ( .A1(n13703), .A2(n13706), .ZN(n16512) );
  INV_X1 U17024 ( .A(n16512), .ZN(n13704) );
  NAND2_X1 U17025 ( .A1(n13705), .A2(n9682), .ZN(n15995) );
  INV_X1 U17026 ( .A(n13706), .ZN(n13707) );
  OAI21_X1 U17027 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13707), .A(
        n9760), .ZN(n16502) );
  NAND2_X1 U17028 ( .A1(n15995), .A2(n16502), .ZN(n15977) );
  INV_X1 U17029 ( .A(n15977), .ZN(n13709) );
  INV_X1 U17030 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21655) );
  AOI21_X1 U17031 ( .B1(n21655), .B2(n9760), .A(n9873), .ZN(n15982) );
  INV_X1 U17032 ( .A(n15982), .ZN(n13708) );
  OAI21_X1 U17033 ( .B1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n9873), .A(
        n9761), .ZN(n16490) );
  AOI21_X1 U17034 ( .B1(n10735), .B2(n9761), .A(n13710), .ZN(n15961) );
  INV_X1 U17035 ( .A(n13711), .ZN(n13715) );
  INV_X1 U17036 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13713) );
  NAND2_X1 U17037 ( .A1(n13713), .A2(n13712), .ZN(n13714) );
  NAND2_X1 U17038 ( .A1(n13715), .A2(n13714), .ZN(n15947) );
  NAND2_X1 U17039 ( .A1(n15946), .A2(n15947), .ZN(n14945) );
  INV_X1 U17040 ( .A(n13716), .ZN(n13718) );
  NOR2_X1 U17041 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U17042 ( .A1(n13718), .A2(n13717), .ZN(n19820) );
  NOR2_X1 U17043 ( .A1(n14345), .A2(n19736), .ZN(n13719) );
  NAND2_X1 U17044 ( .A1(n13719), .A2(n14705), .ZN(n19796) );
  NOR2_X1 U17045 ( .A1(n11602), .A2(n19736), .ZN(n13720) );
  NAND2_X1 U17046 ( .A1(n19796), .A2(n14046), .ZN(n15942) );
  AND2_X1 U17047 ( .A1(n17196), .A2(n20198), .ZN(n13728) );
  INV_X1 U17048 ( .A(n13728), .ZN(n13721) );
  NOR2_X1 U17049 ( .A1(n15934), .A2(n13721), .ZN(n13733) );
  INV_X1 U17050 ( .A(n13733), .ZN(n13722) );
  NOR2_X1 U17051 ( .A1(n14347), .A2(n13722), .ZN(n13723) );
  AND2_X1 U17052 ( .A1(n11385), .A2(n13723), .ZN(n14721) );
  NOR2_X1 U17053 ( .A1(n14046), .A2(n13728), .ZN(n13734) );
  AND2_X1 U17054 ( .A1(n14347), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13724) );
  OAI21_X1 U17055 ( .B1(n16360), .B2(n19813), .A(n13726), .ZN(n13727) );
  INV_X1 U17056 ( .A(n14046), .ZN(n14036) );
  AND2_X1 U17057 ( .A1(n14347), .A2(n13728), .ZN(n13729) );
  NAND2_X1 U17058 ( .A1(n13730), .A2(n19819), .ZN(n13741) );
  NOR2_X2 U17059 ( .A1(n19778), .A2(n19820), .ZN(n19764) );
  NAND2_X1 U17060 ( .A1(n19764), .A2(n13731), .ZN(n14944) );
  NOR2_X1 U17061 ( .A1(n20300), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20298) );
  NAND3_X1 U17062 ( .A1(n11127), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20298), 
        .ZN(n17194) );
  NAND3_X1 U17063 ( .A1(n19820), .A2(n16706), .A3(n17194), .ZN(n13732) );
  NOR2_X1 U17064 ( .A1(n14154), .A2(n13733), .ZN(n14941) );
  INV_X1 U17065 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13757) );
  AND2_X1 U17066 ( .A1(n13734), .A2(n13757), .ZN(n13735) );
  AOI22_X1 U17067 ( .A1(n19789), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19807), .ZN(n13737) );
  NAND2_X1 U17068 ( .A1(n19787), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13736) );
  OAI211_X1 U17069 ( .C1(n13738), .C2(n14944), .A(n13737), .B(n13736), .ZN(
        n13739) );
  NAND4_X1 U17070 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        P2_U2825) );
  INV_X1 U17071 ( .A(n13746), .ZN(n13749) );
  NOR2_X1 U17072 ( .A1(n13747), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13748) );
  MUX2_X1 U17073 ( .A(n13749), .B(n13748), .S(n19879), .Z(n14947) );
  NAND2_X1 U17074 ( .A1(n14947), .A2(n13750), .ZN(n13751) );
  XOR2_X1 U17075 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13751), .Z(
        n13752) );
  NAND2_X1 U17076 ( .A1(n14915), .A2(n13753), .ZN(n13760) );
  NAND2_X1 U17077 ( .A1(n11126), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13756) );
  AOI22_X1 U17078 ( .A1(n9694), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13755) );
  OAI211_X1 U17079 ( .C1(n13758), .C2(n13757), .A(n13756), .B(n13755), .ZN(
        n13759) );
  XNOR2_X2 U17080 ( .A(n13760), .B(n13759), .ZN(n16265) );
  NAND2_X1 U17081 ( .A1(n14931), .A2(n13762), .ZN(n13765) );
  AOI222_X1 U17082 ( .A1(n13763), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n9687), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n13649), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13764) );
  NOR3_X1 U17083 ( .A1(n10555), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13766), .ZN(n13771) );
  INV_X1 U17084 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n13767) );
  NOR2_X1 U17085 ( .A1(n16706), .A2(n13767), .ZN(n13982) );
  AOI211_X1 U17086 ( .C1(n13772), .C2(n13771), .A(n13982), .B(n13770), .ZN(
        n13773) );
  INV_X1 U17087 ( .A(n16496), .ZN(n13776) );
  INV_X1 U17088 ( .A(n13777), .ZN(n13778) );
  OR2_X1 U17089 ( .A1(n13781), .A2(n13782), .ZN(n13783) );
  AND2_X1 U17090 ( .A1(n13780), .A2(n13783), .ZN(n16397) );
  NAND2_X1 U17091 ( .A1(n19788), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13797) );
  INV_X1 U17092 ( .A(n13784), .ZN(n16733) );
  XNOR2_X1 U17093 ( .A(n16732), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13785) );
  NAND2_X1 U17094 ( .A1(n16733), .A2(n13785), .ZN(n13786) );
  OAI211_X1 U17095 ( .C1(n16729), .C2(n13787), .A(n13797), .B(n13786), .ZN(
        n13792) );
  INV_X1 U17096 ( .A(n13788), .ZN(n13789) );
  OAI21_X1 U17097 ( .B1(n9835), .B2(n13790), .A(n13789), .ZN(n16287) );
  NOR2_X1 U17098 ( .A1(n16287), .A2(n17185), .ZN(n13791) );
  AOI211_X1 U17099 ( .C1(n16989), .C2(n16397), .A(n13792), .B(n13791), .ZN(
        n13794) );
  NAND2_X1 U17100 ( .A1(n13796), .A2(n13795), .ZN(P2_U3020) );
  OAI21_X1 U17101 ( .B1(n16672), .B2(n21655), .A(n13797), .ZN(n13799) );
  NOR2_X1 U17102 ( .A1(n16287), .A2(n16695), .ZN(n13798) );
  AOI211_X1 U17103 ( .C1(n16692), .C2(n15982), .A(n13799), .B(n13798), .ZN(
        n13801) );
  NAND2_X1 U17104 ( .A1(n13803), .A2(n13802), .ZN(P2_U2988) );
  INV_X1 U17105 ( .A(n13871), .ZN(n13853) );
  NOR2_X1 U17106 ( .A1(n9689), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13901) );
  NAND2_X1 U17107 ( .A1(n13821), .A2(n13820), .ZN(n13831) );
  NAND2_X1 U17108 ( .A1(n13831), .A2(n13830), .ZN(n13848) );
  INV_X1 U17109 ( .A(n13846), .ZN(n13806) );
  XNOR2_X1 U17110 ( .A(n13848), .B(n13806), .ZN(n13807) );
  NAND2_X1 U17111 ( .A1(n13807), .A2(n14052), .ZN(n13808) );
  NAND2_X1 U17112 ( .A1(n13809), .A2(n20733), .ZN(n13815) );
  NAND2_X1 U17113 ( .A1(n13810), .A2(n13871), .ZN(n13814) );
  NAND2_X1 U17114 ( .A1(n13848), .A2(n13846), .ZN(n13811) );
  XNOR2_X1 U17115 ( .A(n13811), .B(n13845), .ZN(n13812) );
  NAND2_X1 U17116 ( .A1(n13812), .A2(n14052), .ZN(n13813) );
  NAND2_X1 U17117 ( .A1(n13814), .A2(n13813), .ZN(n20711) );
  AND2_X1 U17118 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20725) );
  AOI22_X1 U17119 ( .A1(n13815), .A2(n20711), .B1(n20725), .B2(n14626), .ZN(
        n13843) );
  NAND2_X1 U17120 ( .A1(n20784), .A2(n13871), .ZN(n13819) );
  NAND2_X1 U17121 ( .A1(n13916), .A2(n12637), .ZN(n13832) );
  OAI21_X1 U17122 ( .B1(n21412), .B2(n13820), .A(n13832), .ZN(n13817) );
  INV_X1 U17123 ( .A(n13817), .ZN(n13818) );
  NAND2_X1 U17124 ( .A1(n13819), .A2(n13818), .ZN(n14208) );
  OAI21_X1 U17125 ( .B1(n13821), .B2(n13820), .A(n13831), .ZN(n13822) );
  OAI211_X1 U17126 ( .C1(n13822), .C2(n21412), .A(n20804), .B(n14173), .ZN(
        n13823) );
  INV_X1 U17127 ( .A(n13823), .ZN(n13824) );
  OAI21_X2 U17128 ( .B1(n13825), .B2(n17112), .A(n13824), .ZN(n13826) );
  XNOR2_X1 U17129 ( .A(n14207), .B(n13826), .ZN(n15672) );
  NAND2_X1 U17130 ( .A1(n15672), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20758) );
  INV_X1 U17131 ( .A(n13826), .ZN(n13827) );
  OR2_X1 U17132 ( .A1(n13827), .A2(n14207), .ZN(n13828) );
  XNOR2_X1 U17133 ( .A(n13837), .B(n20754), .ZN(n14478) );
  XNOR2_X1 U17134 ( .A(n13831), .B(n13830), .ZN(n13834) );
  INV_X1 U17135 ( .A(n13832), .ZN(n13833) );
  AOI21_X1 U17136 ( .B1(n13834), .B2(n14052), .A(n13833), .ZN(n13835) );
  NAND2_X1 U17137 ( .A1(n13836), .A2(n13835), .ZN(n14477) );
  NAND2_X1 U17138 ( .A1(n14478), .A2(n14477), .ZN(n20745) );
  NAND2_X1 U17139 ( .A1(n13837), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13838) );
  OR2_X1 U17140 ( .A1(n14626), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13841) );
  INV_X1 U17141 ( .A(n20711), .ZN(n13839) );
  NAND3_X1 U17142 ( .A1(n14625), .A2(n13841), .A3(n13840), .ZN(n13842) );
  AND2_X1 U17143 ( .A1(n13846), .A2(n13845), .ZN(n13847) );
  NAND2_X1 U17144 ( .A1(n13848), .A2(n13847), .ZN(n13867) );
  XNOR2_X1 U17145 ( .A(n13867), .B(n13865), .ZN(n13849) );
  NAND2_X1 U17146 ( .A1(n13849), .A2(n14052), .ZN(n13850) );
  INV_X1 U17147 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17149) );
  NAND2_X1 U17148 ( .A1(n13851), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13852) );
  OR2_X1 U17149 ( .A1(n13854), .A2(n13853), .ZN(n13859) );
  INV_X1 U17150 ( .A(n13867), .ZN(n13855) );
  NAND2_X1 U17151 ( .A1(n13855), .A2(n13865), .ZN(n13856) );
  XNOR2_X1 U17152 ( .A(n13856), .B(n13864), .ZN(n13857) );
  NAND2_X1 U17153 ( .A1(n13857), .A2(n14052), .ZN(n13858) );
  INV_X1 U17154 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15892) );
  NAND2_X1 U17155 ( .A1(n14610), .A2(n15892), .ZN(n13860) );
  INV_X1 U17156 ( .A(n14610), .ZN(n13861) );
  NAND2_X1 U17157 ( .A1(n13861), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13862) );
  NAND2_X1 U17158 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  INV_X1 U17159 ( .A(n13876), .ZN(n13868) );
  XNOR2_X1 U17160 ( .A(n13875), .B(n13868), .ZN(n13869) );
  NOR2_X1 U17161 ( .A1(n13869), .A2(n21412), .ZN(n13870) );
  AOI21_X1 U17162 ( .B1(n13872), .B2(n13871), .A(n13870), .ZN(n13873) );
  INV_X1 U17163 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15889) );
  NAND2_X1 U17164 ( .A1(n13873), .A2(n15889), .ZN(n15658) );
  INV_X1 U17165 ( .A(n13873), .ZN(n13874) );
  INV_X1 U17166 ( .A(n13875), .ZN(n13877) );
  NAND3_X1 U17167 ( .A1(n13877), .A2(n14052), .A3(n13876), .ZN(n13878) );
  NAND2_X1 U17168 ( .A1(n9697), .A2(n13878), .ZN(n15647) );
  OR2_X1 U17169 ( .A1(n15647), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13879) );
  INV_X1 U17170 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15850) );
  NAND2_X1 U17171 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13881) );
  NAND2_X1 U17172 ( .A1(n9697), .A2(n13881), .ZN(n15600) );
  INV_X1 U17173 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13882) );
  NAND2_X1 U17174 ( .A1(n13880), .A2(n13882), .ZN(n13883) );
  NAND2_X1 U17175 ( .A1(n13880), .A2(n21709), .ZN(n13884) );
  OR2_X1 U17176 ( .A1(n9697), .A2(n21709), .ZN(n13885) );
  INV_X1 U17177 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15816) );
  XNOR2_X1 U17178 ( .A(n13880), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15566) );
  NAND2_X1 U17179 ( .A1(n13880), .A2(n15816), .ZN(n15576) );
  NAND2_X1 U17180 ( .A1(n15566), .A2(n15576), .ZN(n13886) );
  NAND2_X1 U17181 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U17182 ( .A1(n9689), .A2(n13887), .ZN(n13888) );
  NOR2_X1 U17183 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13890) );
  OR2_X1 U17184 ( .A1(n13880), .A2(n15850), .ZN(n15602) );
  NOR2_X1 U17185 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13889) );
  OR2_X1 U17186 ( .A1(n13880), .A2(n13889), .ZN(n15598) );
  INV_X1 U17187 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15879) );
  OAI211_X1 U17188 ( .C1(n13890), .C2(n13880), .A(n15563), .B(n15552), .ZN(
        n13892) );
  XNOR2_X1 U17189 ( .A(n9697), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15543) );
  NAND2_X1 U17190 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15770) );
  INV_X1 U17191 ( .A(n15770), .ZN(n13894) );
  NAND2_X1 U17192 ( .A1(n15498), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13898) );
  INV_X1 U17193 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13896) );
  INV_X1 U17194 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13895) );
  INV_X1 U17195 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15508) );
  NAND2_X1 U17196 ( .A1(n13897), .A2(n15621), .ZN(n15497) );
  AND2_X1 U17197 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15724) );
  NAND2_X1 U17198 ( .A1(n15724), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15716) );
  NAND2_X1 U17199 ( .A1(n15437), .A2(n15716), .ZN(n13899) );
  INV_X1 U17200 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15748) );
  INV_X1 U17201 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15725) );
  INV_X1 U17202 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15738) );
  NAND3_X1 U17203 ( .A1(n15748), .A2(n15725), .A3(n15738), .ZN(n15439) );
  NOR2_X1 U17204 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15697) );
  AND2_X1 U17205 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15696) );
  INV_X1 U17206 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15690) );
  AND2_X1 U17207 ( .A1(n13903), .A2(n21409), .ZN(n13906) );
  NAND2_X1 U17208 ( .A1(n14590), .A2(n14566), .ZN(n13905) );
  AOI21_X1 U17209 ( .B1(n13902), .B2(n13906), .A(n13905), .ZN(n13907) );
  INV_X1 U17210 ( .A(n14196), .ZN(n13909) );
  NAND2_X1 U17211 ( .A1(n14297), .A2(n14298), .ZN(n13908) );
  NAND2_X1 U17212 ( .A1(n13909), .A2(n13908), .ZN(n13910) );
  NOR2_X1 U17213 ( .A1(n15918), .A2(n17112), .ZN(n13941) );
  INV_X1 U17214 ( .A(n13911), .ZN(n13914) );
  NAND2_X1 U17215 ( .A1(n12633), .A2(n20812), .ZN(n13913) );
  AOI21_X1 U17216 ( .B1(n15918), .B2(n13916), .A(n13915), .ZN(n13917) );
  INV_X1 U17217 ( .A(n17102), .ZN(n13918) );
  OR2_X1 U17218 ( .A1(n14061), .A2(n13918), .ZN(n13921) );
  INV_X1 U17219 ( .A(n13919), .ZN(n13920) );
  NAND2_X1 U17220 ( .A1(n12668), .A2(n13920), .ZN(n13934) );
  NAND2_X1 U17221 ( .A1(n13921), .A2(n13934), .ZN(n14195) );
  AOI21_X1 U17222 ( .B1(n14579), .B2(n13941), .A(n14195), .ZN(n13922) );
  INV_X1 U17223 ( .A(n13928), .ZN(n13923) );
  NAND2_X1 U17224 ( .A1(n13923), .A2(n12632), .ZN(n13924) );
  OAI211_X1 U17225 ( .C1(n17102), .C2(n14054), .A(n14576), .B(n13924), .ZN(
        n13926) );
  OR2_X1 U17226 ( .A1(n13926), .A2(n13925), .ZN(n13927) );
  OAI22_X1 U17227 ( .A1(n14051), .A2(n14297), .B1(n12632), .B2(n13928), .ZN(
        n13929) );
  INV_X1 U17228 ( .A(n13930), .ZN(n13933) );
  OAI21_X1 U17229 ( .B1(n14179), .B2(n14199), .A(n13931), .ZN(n13932) );
  AOI21_X1 U17230 ( .B1(n13933), .B2(n14297), .A(n13932), .ZN(n13936) );
  AND3_X1 U17231 ( .A1(n13936), .A2(n13935), .A3(n13934), .ZN(n14177) );
  INV_X1 U17232 ( .A(n14199), .ZN(n15271) );
  NAND2_X1 U17233 ( .A1(n15271), .A2(n14054), .ZN(n14172) );
  MUX2_X1 U17234 ( .A(n13937), .B(n20804), .S(n14566), .Z(n13938) );
  NAND4_X1 U17235 ( .A1(n14177), .A2(n13939), .A3(n14172), .A4(n13938), .ZN(
        n13940) );
  NAND2_X1 U17236 ( .A1(n13944), .A2(n13940), .ZN(n20769) );
  NAND2_X1 U17237 ( .A1(n13944), .A2(n14495), .ZN(n20771) );
  INV_X1 U17238 ( .A(n15893), .ZN(n20761) );
  NAND2_X1 U17239 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13964) );
  AND2_X1 U17240 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15869) );
  NAND3_X1 U17241 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15827) );
  INV_X1 U17242 ( .A(n15827), .ZN(n15864) );
  NAND2_X1 U17243 ( .A1(n15869), .A2(n15864), .ZN(n15842) );
  NAND4_X1 U17244 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(n20725), .ZN(n14616) );
  INV_X1 U17245 ( .A(n14616), .ZN(n13942) );
  NAND3_X1 U17246 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n13942), .ZN(n13943) );
  NOR2_X1 U17247 ( .A1(n15842), .A2(n13943), .ZN(n13957) );
  AOI21_X1 U17248 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13957), .A(
        n20723), .ZN(n13947) );
  OR2_X1 U17249 ( .A1(n20769), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13946) );
  OR2_X1 U17250 ( .A1(n13944), .A2(n20727), .ZN(n13945) );
  NAND3_X1 U17251 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15828) );
  INV_X1 U17252 ( .A(n15842), .ZN(n15851) );
  INV_X1 U17253 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20770) );
  INV_X1 U17254 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20768) );
  OAI21_X1 U17255 ( .B1(n20770), .B2(n20768), .A(n20754), .ZN(n20721) );
  AND2_X1 U17256 ( .A1(n20725), .A2(n20721), .ZN(n13948) );
  AND2_X1 U17257 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13948), .ZN(
        n14613) );
  NAND2_X1 U17258 ( .A1(n15851), .A2(n14613), .ZN(n13956) );
  OAI21_X1 U17259 ( .B1(n15828), .B2(n13956), .A(n20756), .ZN(n13949) );
  NAND2_X1 U17260 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15804) );
  NOR2_X1 U17261 ( .A1(n15804), .A2(n15806), .ZN(n15795) );
  NAND2_X1 U17262 ( .A1(n15795), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15786) );
  OR2_X1 U17263 ( .A1(n15786), .A2(n13895), .ZN(n13962) );
  NOR2_X1 U17264 ( .A1(n13951), .A2(n15863), .ZN(n15766) );
  AOI21_X1 U17265 ( .B1(n15893), .B2(n13964), .A(n15766), .ZN(n15749) );
  INV_X1 U17266 ( .A(n15749), .ZN(n13952) );
  NOR2_X1 U17267 ( .A1(n13952), .A2(n15893), .ZN(n13954) );
  INV_X1 U17268 ( .A(n13954), .ZN(n13953) );
  OAI21_X1 U17269 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20722), .A(
        n15749), .ZN(n15734) );
  INV_X1 U17270 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14186) );
  NOR2_X1 U17271 ( .A1(n13954), .A2(n14186), .ZN(n13968) );
  NAND2_X1 U17272 ( .A1(n13957), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13961) );
  NAND2_X1 U17273 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13955) );
  NOR2_X1 U17274 ( .A1(n13956), .A2(n13955), .ZN(n15832) );
  NAND2_X1 U17275 ( .A1(n20756), .A2(n15832), .ZN(n13960) );
  INV_X1 U17276 ( .A(n13957), .ZN(n13958) );
  OR2_X1 U17277 ( .A1(n20771), .A2(n13958), .ZN(n13959) );
  OAI211_X1 U17278 ( .C1(n20769), .C2(n13961), .A(n13960), .B(n13959), .ZN(
        n15833) );
  INV_X1 U17279 ( .A(n13962), .ZN(n13963) );
  NAND2_X1 U17280 ( .A1(n15810), .A2(n13963), .ZN(n15777) );
  NOR2_X1 U17281 ( .A1(n15777), .A2(n15770), .ZN(n15754) );
  INV_X1 U17282 ( .A(n13964), .ZN(n13965) );
  NAND2_X1 U17283 ( .A1(n15754), .A2(n13965), .ZN(n15735) );
  INV_X1 U17284 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13966) );
  INV_X1 U17285 ( .A(n15707), .ZN(n15687) );
  NAND3_X1 U17286 ( .A1(n15687), .A2(n15696), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15679) );
  INV_X1 U17287 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15680) );
  NOR3_X1 U17288 ( .A1(n15679), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15680), .ZN(n13967) );
  NOR2_X1 U17289 ( .A1(n20781), .A2(n10683), .ZN(n13977) );
  AOI211_X1 U17290 ( .C1(n15677), .C2(n13968), .A(n13967), .B(n13977), .ZN(
        n13969) );
  NAND2_X1 U17291 ( .A1(n13971), .A2(n20716), .ZN(n13981) );
  NAND3_X1 U17292 ( .A1(n17176), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17168) );
  INV_X1 U17293 ( .A(n17168), .ZN(n13972) );
  NAND2_X1 U17294 ( .A1(n21266), .A2(n13973), .ZN(n21408) );
  NAND2_X1 U17295 ( .A1(n21408), .A2(n17176), .ZN(n13974) );
  NAND2_X1 U17296 ( .A1(n17176), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17114) );
  NAND2_X1 U17297 ( .A1(n21232), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13975) );
  NAND2_X1 U17298 ( .A1(n17114), .A2(n13975), .ZN(n14210) );
  NOR2_X1 U17299 ( .A1(n14885), .A2(n20720), .ZN(n13976) );
  AOI211_X1 U17300 ( .C1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n20709), .A(
        n13977), .B(n13976), .ZN(n13978) );
  INV_X1 U17301 ( .A(n13978), .ZN(n13979) );
  NAND2_X1 U17302 ( .A1(n13981), .A2(n13980), .ZN(P1_U2968) );
  AOI21_X1 U17303 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13982), .ZN(n13983) );
  OAI21_X1 U17304 ( .B1(n16710), .B2(n13984), .A(n13983), .ZN(n13985) );
  INV_X1 U17305 ( .A(n13985), .ZN(n13987) );
  NAND2_X1 U17306 ( .A1(n9832), .A2(n13989), .ZN(P2_U2983) );
  NOR2_X1 U17307 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21427) );
  NOR3_X1 U17308 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13992) );
  NOR4_X1 U17309 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13991) );
  NOR4_X1 U17310 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_2__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13990) );
  AND4_X1 U17311 ( .A1(n21427), .A2(n13992), .A3(n13991), .A4(n13990), .ZN(
        n13998) );
  NOR4_X1 U17312 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13996) );
  NOR4_X1 U17313 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13995) );
  NOR4_X1 U17314 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13994) );
  NOR4_X1 U17315 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13993) );
  AND4_X1 U17316 ( .A1(n13996), .A2(n13995), .A3(n13994), .A4(n13993), .ZN(
        n13997) );
  NAND2_X1 U17317 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  NOR2_X1 U17318 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(n21543), .ZN(n21430) );
  INV_X1 U17319 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21406) );
  NOR2_X1 U17320 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(n21406), .ZN(n14001) );
  NOR4_X1 U17321 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n14000) );
  NOR4_X1 U17322 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n14005) );
  NOR4_X1 U17323 ( .A1(P2_ADDRESS_REG_5__SCAN_IN), .A2(
        P2_ADDRESS_REG_4__SCAN_IN), .A3(P2_ADDRESS_REG_3__SCAN_IN), .A4(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n14004) );
  NOR4_X1 U17324 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n14003) );
  NOR4_X1 U17325 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n14002) );
  AND4_X1 U17326 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14010) );
  NOR4_X1 U17327 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n14008) );
  NOR4_X1 U17328 ( .A1(P2_ADDRESS_REG_9__SCAN_IN), .A2(
        P2_ADDRESS_REG_8__SCAN_IN), .A3(P2_ADDRESS_REG_7__SCAN_IN), .A4(
        P2_ADDRESS_REG_6__SCAN_IN), .ZN(n14007) );
  NOR4_X1 U17329 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n14006) );
  AND4_X1 U17330 ( .A1(n14008), .A2(n14007), .A3(n14006), .A4(n20510), .ZN(
        n14009) );
  NAND2_X1 U17331 ( .A1(n14010), .A2(n14009), .ZN(n14011) );
  NOR2_X1 U17332 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n14013) );
  NOR4_X1 U17333 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14012) );
  NAND4_X1 U17334 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n14013), .A4(n14012), .ZN(n14014) );
  NOR2_X1 U17335 ( .A1(n17040), .A2(n14014), .ZN(n17274) );
  INV_X2 U17336 ( .A(n17349), .ZN(U215) );
  AOI211_X1 U17337 ( .C1(n16597), .C2(n14015), .A(n16147), .B(n16195), .ZN(
        n14031) );
  OAI22_X1 U17338 ( .A1(n19774), .A2(n11484), .B1(n21718), .B2(n19815), .ZN(
        n14030) );
  AND2_X1 U17339 ( .A1(n14285), .A2(n14016), .ZN(n14017) );
  OR2_X1 U17340 ( .A1(n14017), .A2(n14439), .ZN(n19837) );
  AOI211_X1 U17341 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n14019), .A(n19791), .B(
        n14018), .ZN(n14020) );
  AOI211_X1 U17342 ( .C1(n19789), .C2(P2_REIP_REG_11__SCAN_IN), .A(n19788), 
        .B(n14020), .ZN(n14021) );
  OAI21_X1 U17343 ( .B1(n19837), .B2(n19813), .A(n14021), .ZN(n14029) );
  INV_X1 U17344 ( .A(n14023), .ZN(n14024) );
  AOI21_X1 U17345 ( .B1(n14025), .B2(n14844), .A(n14024), .ZN(n16892) );
  INV_X1 U17346 ( .A(n16892), .ZN(n14027) );
  INV_X1 U17347 ( .A(n16597), .ZN(n14026) );
  OAI22_X1 U17348 ( .A1(n14027), .A2(n16238), .B1(n14026), .B2(n19826), .ZN(
        n14028) );
  INV_X1 U17349 ( .A(HOLD), .ZN(n21335) );
  INV_X1 U17350 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21637) );
  NAND2_X1 U17351 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21347) );
  OAI21_X1 U17352 ( .B1(n21335), .B2(n12628), .A(n21347), .ZN(n14032) );
  OAI21_X1 U17353 ( .B1(n21335), .B2(n21637), .A(n14032), .ZN(n14033) );
  OAI211_X1 U17354 ( .C1(n12628), .C2(n21409), .A(n14033), .B(n14298), .ZN(
        P1_U3195) );
  NAND2_X1 U17355 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17196), .ZN(n14757) );
  OAI21_X1 U17356 ( .B1(n20198), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14757), 
        .ZN(n14034) );
  AOI21_X1 U17357 ( .B1(n14034), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14035) );
  NAND2_X1 U17358 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n16997) );
  NOR2_X1 U17359 ( .A1(n16997), .A2(n14457), .ZN(n17203) );
  NOR2_X1 U17360 ( .A1(n14035), .A2(n17203), .ZN(P2_U3178) );
  AND2_X1 U17361 ( .A1(n20528), .A2(n11127), .ZN(n14039) );
  AOI211_X1 U17362 ( .C1(n19796), .C2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n14039), 
        .B(n14036), .ZN(n14037) );
  INV_X1 U17363 ( .A(n14037), .ZN(P2_U2814) );
  INV_X1 U17364 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n14038) );
  INV_X1 U17365 ( .A(n17019), .ZN(n20523) );
  NAND2_X1 U17366 ( .A1(n20393), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17195) );
  OAI22_X1 U17367 ( .A1(n15942), .A2(n14038), .B1(n20523), .B2(n17195), .ZN(
        P2_U2816) );
  INV_X1 U17368 ( .A(n15939), .ZN(n14042) );
  INV_X1 U17369 ( .A(n15942), .ZN(n14041) );
  OAI21_X1 U17370 ( .B1(n14039), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n14041), 
        .ZN(n14040) );
  OAI21_X1 U17371 ( .B1(n14042), .B2(n14041), .A(n14040), .ZN(P2_U3612) );
  NAND2_X1 U17372 ( .A1(n21273), .A2(n17174), .ZN(n20564) );
  INV_X1 U17373 ( .A(n20564), .ZN(n14979) );
  AOI21_X1 U17374 ( .B1(n14043), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14979), 
        .ZN(n14044) );
  NAND2_X1 U17375 ( .A1(n14384), .A2(n14044), .ZN(P1_U2801) );
  NAND2_X1 U17376 ( .A1(n14347), .A2(n17196), .ZN(n14045) );
  INV_X1 U17377 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14049) );
  INV_X1 U17378 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n14047) );
  INV_X1 U17379 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n15403) );
  INV_X2 U17380 ( .A(n17040), .ZN(n17038) );
  MUX2_X1 U17381 ( .A(n14047), .B(n15403), .S(n17038), .Z(n14635) );
  INV_X1 U17382 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n14048) );
  OAI222_X1 U17383 ( .A1(n14066), .A2(n14049), .B1(n14067), .B2(n14635), .C1(
        n14048), .C2(n14154), .ZN(P2_U2982) );
  AOI22_X1 U17384 ( .A1(n14579), .A2(n14055), .B1(n14051), .B2(n14050), .ZN(
        n20560) );
  OAI21_X1 U17385 ( .B1(n15271), .B2(n14052), .A(n14298), .ZN(n14053) );
  NAND2_X1 U17386 ( .A1(n14053), .A2(n21409), .ZN(n21410) );
  NAND2_X1 U17387 ( .A1(n20560), .A2(n21410), .ZN(n17104) );
  INV_X1 U17388 ( .A(n20561), .ZN(n14295) );
  NAND2_X1 U17389 ( .A1(n17104), .A2(n14295), .ZN(n20568) );
  INV_X1 U17390 ( .A(n20568), .ZN(n14065) );
  INV_X1 U17391 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n14064) );
  AND2_X1 U17392 ( .A1(n14055), .A2(n14054), .ZN(n14057) );
  OAI21_X1 U17393 ( .B1(n17102), .B2(n14057), .A(n14056), .ZN(n14058) );
  MUX2_X1 U17394 ( .A(n14180), .B(n14058), .S(n14579), .Z(n14059) );
  AOI21_X1 U17395 ( .B1(n14061), .B2(n14060), .A(n14059), .ZN(n14062) );
  INV_X1 U17396 ( .A(n14587), .ZN(n20826) );
  NOR2_X1 U17397 ( .A1(n14062), .A2(n20826), .ZN(n17106) );
  NAND2_X1 U17398 ( .A1(n17106), .A2(n14065), .ZN(n14063) );
  OAI21_X1 U17399 ( .B1(n14065), .B2(n14064), .A(n14063), .ZN(P1_U3484) );
  INV_X1 U17400 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14071) );
  NAND2_X1 U17401 ( .A1(n14151), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n14070) );
  INV_X1 U17402 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n14069) );
  NAND2_X1 U17403 ( .A1(n17038), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14068) );
  OAI21_X1 U17404 ( .B1(n17038), .B2(n14069), .A(n14068), .ZN(n16422) );
  NAND2_X1 U17405 ( .A1(n14143), .A2(n16422), .ZN(n14122) );
  OAI211_X1 U17406 ( .C1(n14154), .C2(n14071), .A(n14070), .B(n14122), .ZN(
        P2_U2958) );
  INV_X1 U17407 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14075) );
  NAND2_X1 U17408 ( .A1(n14151), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14074) );
  INV_X1 U17409 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n14073) );
  NAND2_X1 U17410 ( .A1(n17038), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14072) );
  OAI21_X1 U17411 ( .B1(n17038), .B2(n14073), .A(n14072), .ZN(n16400) );
  NAND2_X1 U17412 ( .A1(n14143), .A2(n16400), .ZN(n14129) );
  OAI211_X1 U17413 ( .C1(n14154), .C2(n14075), .A(n14074), .B(n14129), .ZN(
        P2_U2961) );
  INV_X1 U17414 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14079) );
  NAND2_X1 U17415 ( .A1(n14151), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14078) );
  INV_X1 U17416 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n14077) );
  NAND2_X1 U17417 ( .A1(n17038), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14076) );
  OAI21_X1 U17418 ( .B1(n17038), .B2(n14077), .A(n14076), .ZN(n16407) );
  NAND2_X1 U17419 ( .A1(n14143), .A2(n16407), .ZN(n14126) );
  OAI211_X1 U17420 ( .C1(n14154), .C2(n14079), .A(n14078), .B(n14126), .ZN(
        P2_U2960) );
  INV_X1 U17421 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n21685) );
  NAND2_X1 U17422 ( .A1(n14151), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14080) );
  MUX2_X1 U17423 ( .A(BUF2_REG_14__SCAN_IN), .B(BUF1_REG_14__SCAN_IN), .S(
        n17038), .Z(n16356) );
  NAND2_X1 U17424 ( .A1(n14143), .A2(n16356), .ZN(n14145) );
  OAI211_X1 U17425 ( .C1(n21685), .C2(n14154), .A(n14080), .B(n14145), .ZN(
        P2_U2966) );
  INV_X1 U17426 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U17427 ( .A1(n14151), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n14083) );
  INV_X1 U17428 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n14082) );
  NAND2_X1 U17429 ( .A1(n17038), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14081) );
  OAI21_X1 U17430 ( .B1(n17038), .B2(n14082), .A(n14081), .ZN(n19870) );
  NAND2_X1 U17431 ( .A1(n14143), .A2(n19870), .ZN(n14110) );
  OAI211_X1 U17432 ( .C1(n14154), .C2(n14253), .A(n14083), .B(n14110), .ZN(
        P2_U2954) );
  INV_X1 U17433 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17434 ( .A1(n14151), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14086) );
  INV_X1 U17435 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U17436 ( .A1(n17038), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14084) );
  OAI21_X1 U17437 ( .B1(n17038), .B2(n14085), .A(n14084), .ZN(n16392) );
  NAND2_X1 U17438 ( .A1(n14143), .A2(n16392), .ZN(n14134) );
  OAI211_X1 U17439 ( .C1(n14154), .C2(n14250), .A(n14086), .B(n14134), .ZN(
        P2_U2962) );
  INV_X1 U17440 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U17441 ( .A1(n14151), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n14089) );
  INV_X1 U17442 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n14088) );
  NAND2_X1 U17443 ( .A1(n17038), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14087) );
  OAI21_X1 U17444 ( .B1(n17038), .B2(n14088), .A(n14087), .ZN(n17046) );
  NAND2_X1 U17445 ( .A1(n14143), .A2(n17046), .ZN(n14094) );
  OAI211_X1 U17446 ( .C1(n14154), .C2(n14090), .A(n14089), .B(n14094), .ZN(
        P2_U2953) );
  NAND2_X1 U17447 ( .A1(n14151), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14093) );
  INV_X1 U17448 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n14092) );
  NAND2_X1 U17449 ( .A1(n17038), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14091) );
  OAI21_X1 U17450 ( .B1(n17038), .B2(n14092), .A(n14091), .ZN(n16377) );
  NAND2_X1 U17451 ( .A1(n14143), .A2(n16377), .ZN(n14139) );
  OAI211_X1 U17452 ( .C1(n14154), .C2(n14233), .A(n14093), .B(n14139), .ZN(
        P2_U2964) );
  INV_X1 U17453 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n14235) );
  NAND2_X1 U17454 ( .A1(n14151), .A2(P2_LWORD_REG_1__SCAN_IN), .ZN(n14095) );
  OAI211_X1 U17455 ( .C1(n14154), .C2(n14235), .A(n14095), .B(n14094), .ZN(
        P2_U2968) );
  INV_X1 U17456 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14099) );
  NAND2_X1 U17457 ( .A1(n14151), .A2(P2_UWORD_REG_3__SCAN_IN), .ZN(n14098) );
  INV_X1 U17458 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n14097) );
  NAND2_X1 U17459 ( .A1(n17038), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14096) );
  OAI21_X1 U17460 ( .B1(n17038), .B2(n14097), .A(n14096), .ZN(n16448) );
  NAND2_X1 U17461 ( .A1(n14143), .A2(n16448), .ZN(n14113) );
  OAI211_X1 U17462 ( .C1(n14154), .C2(n14099), .A(n14098), .B(n14113), .ZN(
        P2_U2955) );
  INV_X1 U17463 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n21552) );
  NAND2_X1 U17464 ( .A1(n14151), .A2(P2_UWORD_REG_5__SCAN_IN), .ZN(n14102) );
  INV_X1 U17465 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n14101) );
  NAND2_X1 U17466 ( .A1(n17038), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14100) );
  OAI21_X1 U17467 ( .B1(n17038), .B2(n14101), .A(n14100), .ZN(n19880) );
  NAND2_X1 U17468 ( .A1(n14143), .A2(n19880), .ZN(n14147) );
  OAI211_X1 U17469 ( .C1(n14154), .C2(n21552), .A(n14102), .B(n14147), .ZN(
        P2_U2957) );
  INV_X1 U17470 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U17471 ( .A1(n14151), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n14105) );
  INV_X1 U17472 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n14104) );
  NAND2_X1 U17473 ( .A1(n17038), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14103) );
  OAI21_X1 U17474 ( .B1(n17038), .B2(n14104), .A(n14103), .ZN(n16438) );
  NAND2_X1 U17475 ( .A1(n14143), .A2(n16438), .ZN(n14115) );
  OAI211_X1 U17476 ( .C1(n14154), .C2(n14248), .A(n14105), .B(n14115), .ZN(
        P2_U2956) );
  INV_X1 U17477 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14109) );
  NAND2_X1 U17478 ( .A1(n14151), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n14108) );
  INV_X1 U17479 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n14107) );
  NAND2_X1 U17480 ( .A1(n17038), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14106) );
  OAI21_X1 U17481 ( .B1(n17038), .B2(n14107), .A(n14106), .ZN(n16414) );
  NAND2_X1 U17482 ( .A1(n14143), .A2(n16414), .ZN(n14124) );
  OAI211_X1 U17483 ( .C1(n14154), .C2(n14109), .A(n14108), .B(n14124), .ZN(
        P2_U2959) );
  INV_X1 U17484 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n14112) );
  NAND2_X1 U17485 ( .A1(n14151), .A2(P2_LWORD_REG_2__SCAN_IN), .ZN(n14111) );
  OAI211_X1 U17486 ( .C1(n14154), .C2(n14112), .A(n14111), .B(n14110), .ZN(
        P2_U2969) );
  INV_X1 U17487 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19858) );
  NAND2_X1 U17488 ( .A1(n14151), .A2(P2_LWORD_REG_3__SCAN_IN), .ZN(n14114) );
  OAI211_X1 U17489 ( .C1(n14154), .C2(n19858), .A(n14114), .B(n14113), .ZN(
        P2_U2970) );
  INV_X1 U17490 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n14117) );
  NAND2_X1 U17491 ( .A1(n14151), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n14116) );
  OAI211_X1 U17492 ( .C1(n14154), .C2(n14117), .A(n14116), .B(n14115), .ZN(
        P2_U2971) );
  INV_X1 U17493 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14121) );
  NAND2_X1 U17494 ( .A1(n14151), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14120) );
  INV_X1 U17495 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U17496 ( .A1(n17038), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14118) );
  OAI21_X1 U17497 ( .B1(n17038), .B2(n14119), .A(n14118), .ZN(n14815) );
  NAND2_X1 U17498 ( .A1(n14143), .A2(n14815), .ZN(n14152) );
  OAI211_X1 U17499 ( .C1(n14154), .C2(n14121), .A(n14120), .B(n14152), .ZN(
        P2_U2952) );
  INV_X1 U17500 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n14290) );
  NAND2_X1 U17501 ( .A1(n14151), .A2(P2_LWORD_REG_6__SCAN_IN), .ZN(n14123) );
  OAI211_X1 U17502 ( .C1(n14154), .C2(n14290), .A(n14123), .B(n14122), .ZN(
        P2_U2973) );
  INV_X1 U17503 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n14276) );
  NAND2_X1 U17504 ( .A1(n14151), .A2(P2_LWORD_REG_7__SCAN_IN), .ZN(n14125) );
  OAI211_X1 U17505 ( .C1(n14154), .C2(n14276), .A(n14125), .B(n14124), .ZN(
        P2_U2974) );
  INV_X1 U17506 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n14128) );
  NAND2_X1 U17507 ( .A1(n14151), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n14127) );
  OAI211_X1 U17508 ( .C1(n14154), .C2(n14128), .A(n14127), .B(n14126), .ZN(
        P2_U2975) );
  INV_X1 U17509 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17510 ( .A1(n14151), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14130) );
  OAI211_X1 U17511 ( .C1(n14154), .C2(n14131), .A(n14130), .B(n14129), .ZN(
        P2_U2976) );
  INV_X1 U17512 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U17513 ( .A1(n14151), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14133) );
  INV_X1 U17514 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21476) );
  NAND2_X1 U17515 ( .A1(n17038), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14132) );
  OAI21_X1 U17516 ( .B1(n17038), .B2(n21476), .A(n14132), .ZN(n19833) );
  NAND2_X1 U17517 ( .A1(n14143), .A2(n19833), .ZN(n14137) );
  OAI211_X1 U17518 ( .C1(n14245), .C2(n14154), .A(n14133), .B(n14137), .ZN(
        P2_U2963) );
  INV_X1 U17519 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n14136) );
  NAND2_X1 U17520 ( .A1(n14151), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14135) );
  OAI211_X1 U17521 ( .C1(n14154), .C2(n14136), .A(n14135), .B(n14134), .ZN(
        P2_U2977) );
  INV_X1 U17522 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19850) );
  NAND2_X1 U17523 ( .A1(n14151), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14138) );
  OAI211_X1 U17524 ( .C1(n19850), .C2(n14154), .A(n14138), .B(n14137), .ZN(
        P2_U2978) );
  INV_X1 U17525 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n14141) );
  NAND2_X1 U17526 ( .A1(n14151), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14140) );
  OAI211_X1 U17527 ( .C1(n14154), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        P2_U2979) );
  INV_X1 U17528 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19847) );
  NAND2_X1 U17529 ( .A1(n14151), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n14144) );
  INV_X1 U17530 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18400) );
  NAND2_X1 U17531 ( .A1(n17038), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14142) );
  OAI21_X1 U17532 ( .B1(n17038), .B2(n18400), .A(n14142), .ZN(n16365) );
  NAND2_X1 U17533 ( .A1(n14143), .A2(n16365), .ZN(n14149) );
  OAI211_X1 U17534 ( .C1(n19847), .C2(n14154), .A(n14144), .B(n14149), .ZN(
        P2_U2980) );
  INV_X1 U17535 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19845) );
  NAND2_X1 U17536 ( .A1(n14151), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14146) );
  OAI211_X1 U17537 ( .C1(n19845), .C2(n14154), .A(n14146), .B(n14145), .ZN(
        P2_U2981) );
  INV_X1 U17538 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n14242) );
  NAND2_X1 U17539 ( .A1(n14151), .A2(P2_LWORD_REG_5__SCAN_IN), .ZN(n14148) );
  OAI211_X1 U17540 ( .C1(n14154), .C2(n14242), .A(n14148), .B(n14147), .ZN(
        P2_U2972) );
  INV_X1 U17541 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U17542 ( .A1(n14151), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14150) );
  OAI211_X1 U17543 ( .C1(n14240), .C2(n14154), .A(n14150), .B(n14149), .ZN(
        P2_U2965) );
  INV_X1 U17544 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U17545 ( .A1(n14151), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n14153) );
  OAI211_X1 U17546 ( .C1(n14154), .C2(n14251), .A(n14153), .B(n14152), .ZN(
        P2_U2967) );
  NAND2_X1 U17547 ( .A1(n14347), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14155) );
  INV_X1 U17548 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n16260) );
  MUX2_X1 U17549 ( .A(n16260), .B(n17184), .S(n19832), .Z(n14157) );
  OAI21_X1 U17550 ( .B1(n17033), .B2(n16354), .A(n14157), .ZN(P2_U2887) );
  OR2_X1 U17551 ( .A1(n14158), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14160) );
  NAND2_X1 U17552 ( .A1(n14160), .A2(n14159), .ZN(n20773) );
  NAND2_X1 U17553 ( .A1(n14579), .A2(n14180), .ZN(n14203) );
  NAND2_X1 U17554 ( .A1(n20826), .A2(n20812), .ZN(n14161) );
  NOR2_X1 U17555 ( .A1(n14162), .A2(n14161), .ZN(n14581) );
  NAND3_X1 U17556 ( .A1(n14581), .A2(n14484), .A3(n14163), .ZN(n14164) );
  NAND2_X1 U17557 ( .A1(n14203), .A2(n14164), .ZN(n14165) );
  NAND2_X1 U17558 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  NAND2_X1 U17559 ( .A1(n14169), .A2(n14168), .ZN(n15297) );
  NAND2_X2 U17560 ( .A1(n20655), .A2(n14587), .ZN(n15336) );
  OAI222_X1 U17561 ( .A1(n20773), .A2(n15334), .B1(n14170), .B2(n20655), .C1(
        n15297), .C2(n15336), .ZN(P1_U2872) );
  AND3_X1 U17562 ( .A1(n14174), .A2(n14173), .A3(n14172), .ZN(n14176) );
  AND3_X1 U17563 ( .A1(n14177), .A2(n14176), .A3(n14175), .ZN(n14485) );
  XNOR2_X1 U17564 ( .A(n14178), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14187) );
  NOR2_X1 U17565 ( .A1(n14179), .A2(n14187), .ZN(n14182) );
  INV_X1 U17566 ( .A(n14180), .ZN(n14181) );
  NAND2_X1 U17567 ( .A1(n14181), .A2(n14576), .ZN(n14493) );
  AOI22_X1 U17568 ( .A1(n14485), .A2(n14182), .B1(n14493), .B2(n14187), .ZN(
        n14185) );
  NAND2_X1 U17569 ( .A1(n14495), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14183) );
  NAND2_X1 U17570 ( .A1(n14495), .A2(n12655), .ZN(n15917) );
  MUX2_X1 U17571 ( .A(n14183), .B(n15917), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n14184) );
  OAI211_X1 U17572 ( .C1(n21152), .C2(n14485), .A(n14185), .B(n14184), .ZN(
        n14481) );
  OAI22_X1 U17573 ( .A1(n14186), .A2(n20768), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15922) );
  INV_X1 U17574 ( .A(n15922), .ZN(n14189) );
  NOR2_X1 U17575 ( .A1(n17174), .A2(n20770), .ZN(n15923) );
  INV_X1 U17576 ( .A(n14187), .ZN(n14188) );
  AOI222_X1 U17577 ( .A1(n14481), .A2(n17163), .B1(n14189), .B2(n15923), .C1(
        n17123), .C2(n14188), .ZN(n14206) );
  OR2_X1 U17578 ( .A1(n14495), .A2(n13902), .ZN(n14193) );
  AND2_X1 U17579 ( .A1(n14297), .A2(n21409), .ZN(n14190) );
  NAND2_X1 U17580 ( .A1(n17113), .A2(n14190), .ZN(n14577) );
  OAI21_X1 U17581 ( .B1(n21341), .B2(n14298), .A(n14577), .ZN(n14192) );
  INV_X1 U17582 ( .A(n14576), .ZN(n14191) );
  AOI21_X1 U17583 ( .B1(n14193), .B2(n14192), .A(n14191), .ZN(n14194) );
  OR2_X1 U17584 ( .A1(n14579), .A2(n14194), .ZN(n14202) );
  INV_X1 U17585 ( .A(n14195), .ZN(n14197) );
  OAI211_X1 U17586 ( .C1(n14199), .C2(n14198), .A(n14197), .B(n14584), .ZN(
        n14200) );
  INV_X1 U17587 ( .A(n14200), .ZN(n14201) );
  NOR2_X1 U17588 ( .A1(n17176), .A2(n17177), .ZN(n14511) );
  NAND2_X1 U17589 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n14511), .ZN(n14204) );
  OAI21_X1 U17590 ( .B1(n17090), .B2(n20561), .A(n14204), .ZN(n17162) );
  AOI21_X1 U17591 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n17176), .A(n17162), 
        .ZN(n15926) );
  NAND2_X1 U17592 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15926), .ZN(
        n14205) );
  OAI21_X1 U17593 ( .B1(n14206), .B2(n15926), .A(n14205), .ZN(P1_U3472) );
  OAI21_X1 U17594 ( .B1(n14208), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14207), .ZN(n20776) );
  INV_X1 U17595 ( .A(n15297), .ZN(n14209) );
  NAND2_X1 U17596 ( .A1(n14209), .A2(n20715), .ZN(n14213) );
  OR2_X1 U17597 ( .A1(n20709), .A2(n14210), .ZN(n14211) );
  AOI22_X1 U17598 ( .A1(n14211), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20727), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n14212) );
  OAI211_X1 U17599 ( .C1(n15671), .C2(n20776), .A(n14213), .B(n14212), .ZN(
        P1_U2999) );
  INV_X1 U17600 ( .A(n20882), .ZN(n14535) );
  OAI22_X1 U17601 ( .A1(n14535), .A2(n14485), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15918), .ZN(n17089) );
  OAI22_X1 U17602 ( .A1(n15929), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17174), .ZN(n14214) );
  AOI21_X1 U17603 ( .B1(n17089), .B2(n17163), .A(n14214), .ZN(n14217) );
  INV_X1 U17604 ( .A(n14495), .ZN(n14215) );
  NOR2_X1 U17605 ( .A1(n14215), .A2(n12666), .ZN(n17088) );
  AOI22_X1 U17606 ( .A1(n17088), .A2(n17163), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15926), .ZN(n14216) );
  OAI21_X1 U17607 ( .B1(n14217), .B2(n15926), .A(n14216), .ZN(P1_U3474) );
  INV_X1 U17608 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21708) );
  OR2_X1 U17609 ( .A1(n14218), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14220) );
  NAND2_X1 U17610 ( .A1(n14220), .A2(n14219), .ZN(n14448) );
  INV_X1 U17611 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20465) );
  OR2_X1 U17612 ( .A1(n16706), .A2(n20465), .ZN(n14446) );
  INV_X1 U17613 ( .A(n14446), .ZN(n14221) );
  AOI21_X1 U17614 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14221), .ZN(n14224) );
  XNOR2_X1 U17615 ( .A(n19808), .B(n17017), .ZN(n14222) );
  XNOR2_X1 U17616 ( .A(n14354), .B(n14222), .ZN(n14445) );
  NAND2_X1 U17617 ( .A1(n11531), .A2(n14445), .ZN(n14223) );
  OAI211_X1 U17618 ( .C1(n14448), .C2(n16712), .A(n14224), .B(n14223), .ZN(
        n14225) );
  AOI21_X1 U17619 ( .B1(n16692), .B2(n21708), .A(n14225), .ZN(n14226) );
  OAI21_X1 U17620 ( .B1(n11158), .B2(n16695), .A(n14226), .ZN(P2_U3013) );
  NAND2_X1 U17621 ( .A1(n14336), .A2(n10538), .ZN(n14228) );
  INV_X1 U17622 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17348) );
  INV_X1 U17623 ( .A(n19862), .ZN(n14231) );
  INV_X1 U17624 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n21619) );
  OAI222_X1 U17625 ( .A1(n19842), .A2(n17348), .B1(n14360), .B2(n21685), .C1(
        n15940), .C2(n21619), .ZN(P2_U2921) );
  INV_X1 U17626 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14234) );
  INV_X1 U17627 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n14232) );
  OAI222_X1 U17628 ( .A1(n14234), .A2(n19842), .B1(n14360), .B2(n14233), .C1(
        n15940), .C2(n14232), .ZN(P2_U2923) );
  INV_X1 U17629 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n14236) );
  INV_X1 U17630 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n21688) );
  OAI222_X1 U17631 ( .A1(n14236), .A2(n19842), .B1(n15940), .B2(n21688), .C1(
        n14235), .C2(n19862), .ZN(P2_U2950) );
  INV_X1 U17632 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n14238) );
  INV_X1 U17633 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14237) );
  OAI222_X1 U17634 ( .A1(n14238), .A2(n19842), .B1(n14360), .B2(n21552), .C1(
        n15940), .C2(n14237), .ZN(P2_U2930) );
  INV_X1 U17635 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14241) );
  INV_X1 U17636 ( .A(P2_UWORD_REG_13__SCAN_IN), .ZN(n14239) );
  OAI222_X1 U17637 ( .A1(n14241), .A2(n19842), .B1(n14360), .B2(n14240), .C1(
        n15940), .C2(n14239), .ZN(P2_U2922) );
  INV_X1 U17638 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n14243) );
  INV_X1 U17639 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n21504) );
  OAI222_X1 U17640 ( .A1(n14243), .A2(n19842), .B1(n15940), .B2(n21504), .C1(
        n14242), .C2(n19862), .ZN(P2_U2946) );
  INV_X1 U17641 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14246) );
  INV_X1 U17642 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n14244) );
  OAI222_X1 U17643 ( .A1(n14246), .A2(n19842), .B1(n14360), .B2(n14245), .C1(
        n15940), .C2(n14244), .ZN(P2_U2924) );
  INV_X1 U17644 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n21636) );
  INV_X1 U17645 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14247) );
  OAI222_X1 U17646 ( .A1(n14360), .A2(n14248), .B1(n19842), .B2(n21636), .C1(
        n15940), .C2(n14247), .ZN(P2_U2931) );
  INV_X1 U17647 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n21621) );
  INV_X1 U17648 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n14249) );
  OAI222_X1 U17649 ( .A1(n14360), .A2(n14250), .B1(n19842), .B2(n21621), .C1(
        n15940), .C2(n14249), .ZN(P2_U2925) );
  INV_X1 U17650 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17320) );
  INV_X1 U17651 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n21612) );
  OAI222_X1 U17652 ( .A1(n19862), .A2(n14251), .B1(n19842), .B2(n17320), .C1(
        n15940), .C2(n21612), .ZN(P2_U2951) );
  INV_X1 U17653 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n21559) );
  INV_X1 U17654 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14252) );
  OAI222_X1 U17655 ( .A1(n14360), .A2(n14253), .B1(n19842), .B2(n21559), .C1(
        n15940), .C2(n14252), .ZN(P2_U2933) );
  INV_X1 U17656 ( .A(n14255), .ZN(n14256) );
  AOI21_X1 U17657 ( .B1(n14257), .B2(n14254), .A(n14256), .ZN(n16918) );
  INV_X1 U17658 ( .A(n16918), .ZN(n14267) );
  INV_X1 U17659 ( .A(n14258), .ZN(n14259) );
  AND3_X1 U17660 ( .A1(n14708), .A2(n14259), .A3(n15939), .ZN(n14260) );
  AOI21_X1 U17661 ( .B1(n14699), .B2(n14701), .A(n14260), .ZN(n14340) );
  NAND2_X1 U17662 ( .A1(n14340), .A2(n14261), .ZN(n14262) );
  AND2_X1 U17663 ( .A1(n14264), .A2(n14813), .ZN(n14265) );
  AOI22_X1 U17664 ( .A1(n14785), .A2(n16400), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n16465), .ZN(n14266) );
  OAI21_X1 U17665 ( .B1(n14267), .B2(n19836), .A(n14266), .ZN(P2_U2910) );
  INV_X1 U17666 ( .A(n14815), .ZN(n19863) );
  OAI21_X1 U17667 ( .B1(n14269), .B2(n14268), .A(n11666), .ZN(n17179) );
  INV_X1 U17668 ( .A(n17179), .ZN(n16256) );
  NOR2_X1 U17669 ( .A1(n17033), .A2(n17179), .ZN(n14528) );
  INV_X1 U17670 ( .A(n14528), .ZN(n14270) );
  INV_X1 U17671 ( .A(n16475), .ZN(n16372) );
  OAI211_X1 U17672 ( .C1(n20116), .C2(n16256), .A(n14270), .B(n16372), .ZN(
        n14272) );
  AOI22_X1 U17673 ( .A1(n16472), .A2(n16256), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n16465), .ZN(n14271) );
  OAI211_X1 U17674 ( .C1(n19863), .C2(n19834), .A(n14272), .B(n14271), .ZN(
        P2_U2919) );
  INV_X1 U17675 ( .A(n16414), .ZN(n19893) );
  OR2_X1 U17676 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  AND2_X1 U17677 ( .A1(n14279), .A2(n14275), .ZN(n16940) );
  INV_X1 U17678 ( .A(n16940), .ZN(n14277) );
  OAI222_X1 U17679 ( .A1(n19834), .A2(n19893), .B1(n14277), .B2(n19836), .C1(
        n14276), .C2(n19840), .ZN(P2_U2912) );
  INV_X1 U17680 ( .A(n16407), .ZN(n14282) );
  INV_X1 U17681 ( .A(n14254), .ZN(n14278) );
  AOI21_X1 U17682 ( .B1(n14280), .B2(n14279), .A(n14278), .ZN(n16928) );
  INV_X1 U17683 ( .A(n16928), .ZN(n14281) );
  OAI222_X1 U17684 ( .A1(n19834), .A2(n14282), .B1(n14281), .B2(n19836), .C1(
        n14128), .C2(n19840), .ZN(P2_U2911) );
  INV_X1 U17685 ( .A(n16392), .ZN(n14286) );
  NAND2_X1 U17686 ( .A1(n14255), .A2(n14283), .ZN(n14284) );
  NAND2_X1 U17687 ( .A1(n14285), .A2(n14284), .ZN(n16903) );
  OAI222_X1 U17688 ( .A1(n19834), .A2(n14286), .B1(n16903), .B2(n19836), .C1(
        n14136), .C2(n19840), .ZN(P2_U2909) );
  INV_X1 U17689 ( .A(n16422), .ZN(n19884) );
  OAI21_X1 U17690 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n16205) );
  OAI222_X1 U17691 ( .A1(n19834), .A2(n19884), .B1(n16205), .B2(n19836), .C1(
        n14290), .C2(n19840), .ZN(P2_U2913) );
  MUX2_X1 U17692 ( .A(n14293), .B(n11158), .S(n19832), .Z(n14294) );
  OAI21_X1 U17693 ( .B1(n19998), .B2(n16354), .A(n14294), .ZN(P2_U2886) );
  INV_X1 U17694 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U17695 ( .A1(n14495), .A2(n14295), .ZN(n14296) );
  OAI22_X1 U17696 ( .A1(n14384), .A2(n14297), .B1(n14579), .B2(n14296), .ZN(
        n14299) );
  INV_X1 U17697 ( .A(n14298), .ZN(n17111) );
  INV_X1 U17698 ( .A(n17177), .ZN(n17170) );
  NAND2_X1 U17699 ( .A1(n17176), .A2(n17170), .ZN(n20680) );
  INV_X2 U17700 ( .A(n20680), .ZN(n20684) );
  AOI22_X1 U17701 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14300) );
  OAI21_X1 U17702 ( .B1(n14301), .B2(n14325), .A(n14300), .ZN(P1_U2920) );
  INV_X1 U17703 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17704 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14302) );
  OAI21_X1 U17705 ( .B1(n14303), .B2(n14325), .A(n14302), .ZN(P1_U2907) );
  INV_X1 U17706 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14305) );
  AOI22_X1 U17707 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14304) );
  OAI21_X1 U17708 ( .B1(n14305), .B2(n14325), .A(n14304), .ZN(P1_U2918) );
  AOI22_X1 U17709 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14306) );
  OAI21_X1 U17710 ( .B1(n15381), .B2(n14325), .A(n14306), .ZN(P1_U2917) );
  INV_X1 U17711 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14308) );
  AOI22_X1 U17712 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14307) );
  OAI21_X1 U17713 ( .B1(n14308), .B2(n14325), .A(n14307), .ZN(P1_U2913) );
  INV_X1 U17714 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U17715 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14309) );
  OAI21_X1 U17716 ( .B1(n14310), .B2(n14325), .A(n14309), .ZN(P1_U2912) );
  INV_X1 U17717 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17718 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14311) );
  OAI21_X1 U17719 ( .B1(n14312), .B2(n14325), .A(n14311), .ZN(P1_U2909) );
  INV_X1 U17720 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U17721 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14313) );
  OAI21_X1 U17722 ( .B1(n14314), .B2(n14325), .A(n14313), .ZN(P1_U2916) );
  INV_X1 U17723 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U17724 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U17725 ( .B1(n14316), .B2(n14325), .A(n14315), .ZN(P1_U2906) );
  AOI22_X1 U17726 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14317) );
  OAI21_X1 U17727 ( .B1(n15370), .B2(n14325), .A(n14317), .ZN(P1_U2914) );
  AOI22_X1 U17728 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14318) );
  OAI21_X1 U17729 ( .B1(n13166), .B2(n14325), .A(n14318), .ZN(P1_U2915) );
  INV_X1 U17730 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U17731 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14319) );
  OAI21_X1 U17732 ( .B1(n14320), .B2(n14325), .A(n14319), .ZN(P1_U2919) );
  INV_X1 U17733 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21622) );
  AOI22_X1 U17734 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14321) );
  OAI21_X1 U17735 ( .B1(n21622), .B2(n14325), .A(n14321), .ZN(P1_U2911) );
  INV_X1 U17736 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17737 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14322) );
  OAI21_X1 U17738 ( .B1(n14323), .B2(n14325), .A(n14322), .ZN(P1_U2910) );
  INV_X1 U17739 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14326) );
  AOI22_X1 U17740 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14324) );
  OAI21_X1 U17741 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(P1_U2908) );
  OR2_X1 U17742 ( .A1(n14328), .A2(n14327), .ZN(n14329) );
  AND2_X1 U17743 ( .A1(n14376), .A2(n14329), .ZN(n20634) );
  INV_X1 U17744 ( .A(n20634), .ZN(n14636) );
  INV_X1 U17745 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14334) );
  INV_X1 U17746 ( .A(n14330), .ZN(n14331) );
  NAND2_X1 U17747 ( .A1(n14331), .A2(n13433), .ZN(n14333) );
  AND2_X1 U17748 ( .A1(n14333), .A2(n14332), .ZN(n20763) );
  OAI222_X1 U17749 ( .A1(n15336), .A2(n14636), .B1(n20655), .B2(n14334), .C1(
        n15334), .C2(n20763), .ZN(P1_U2871) );
  NAND2_X1 U17750 ( .A1(n14336), .A2(n14335), .ZN(n14342) );
  INV_X1 U17751 ( .A(n14337), .ZN(n14338) );
  AND3_X1 U17752 ( .A1(n14340), .A2(n14339), .A3(n14338), .ZN(n14341) );
  AOI21_X1 U17753 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n14457), .A(n17203), 
        .ZN(n14722) );
  AND2_X1 U17754 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14459), .ZN(n14343) );
  OAI22_X1 U17755 ( .A1(n14344), .A2(n19736), .B1(n14722), .B2(n14343), .ZN(
        n17023) );
  INV_X1 U17756 ( .A(n17023), .ZN(n17030) );
  NOR2_X1 U17757 ( .A1(n17030), .A2(n20523), .ZN(n17027) );
  INV_X1 U17758 ( .A(n17027), .ZN(n14349) );
  NOR2_X1 U17759 ( .A1(n14347), .A2(n14346), .ZN(n14348) );
  NAND2_X1 U17760 ( .A1(n11086), .A2(n14348), .ZN(n14710) );
  OAI22_X1 U17761 ( .A1(n14349), .A2(n14710), .B1(n14714), .B2(n17023), .ZN(
        P2_U3595) );
  NAND2_X1 U17762 ( .A1(n14350), .A2(n17189), .ZN(n14351) );
  NAND2_X1 U17763 ( .A1(n14352), .A2(n14351), .ZN(n17192) );
  INV_X1 U17764 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n14353) );
  OR2_X1 U17765 ( .A1(n16706), .A2(n14353), .ZN(n17190) );
  OAI21_X1 U17766 ( .B1(n16712), .B2(n17192), .A(n17190), .ZN(n14358) );
  OAI21_X1 U17767 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16257), .A(
        n14354), .ZN(n17181) );
  OAI21_X1 U17768 ( .B1(n16707), .B2(n14355), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14356) );
  OAI21_X1 U17769 ( .B1(n17181), .B2(n16680), .A(n14356), .ZN(n14357) );
  AOI211_X1 U17770 ( .C1(n11168), .C2(n16715), .A(n14358), .B(n14357), .ZN(
        n14359) );
  INV_X1 U17771 ( .A(n14359), .ZN(P2_U3014) );
  INV_X1 U17772 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17773 ( .A1(n14373), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14361) );
  OAI21_X1 U17774 ( .B1(n19842), .B2(n14362), .A(n14361), .ZN(P2_U2935) );
  INV_X1 U17775 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n14364) );
  AOI22_X1 U17776 ( .A1(n14373), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n14363) );
  OAI21_X1 U17777 ( .B1(n19842), .B2(n14364), .A(n14363), .ZN(P2_U2928) );
  INV_X1 U17778 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U17779 ( .A1(n14373), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n14365) );
  OAI21_X1 U17780 ( .B1(n19842), .B2(n14366), .A(n14365), .ZN(P2_U2934) );
  INV_X1 U17781 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U17782 ( .A1(n14373), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n14367) );
  OAI21_X1 U17783 ( .B1(n19842), .B2(n14368), .A(n14367), .ZN(P2_U2929) );
  INV_X1 U17784 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U17785 ( .A1(n14373), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n14369) );
  OAI21_X1 U17786 ( .B1(n19842), .B2(n14370), .A(n14369), .ZN(P2_U2932) );
  INV_X1 U17787 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17788 ( .A1(n14373), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14371) );
  OAI21_X1 U17789 ( .B1(n19842), .B2(n14372), .A(n14371), .ZN(P2_U2927) );
  INV_X1 U17790 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U17791 ( .A1(n14373), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n19859), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14374) );
  OAI21_X1 U17792 ( .B1(n19842), .B2(n14375), .A(n14374), .ZN(P2_U2926) );
  NAND2_X1 U17793 ( .A1(n14377), .A2(n14376), .ZN(n14378) );
  NAND2_X1 U17794 ( .A1(n14379), .A2(n14378), .ZN(n15290) );
  AOI21_X1 U17795 ( .B1(n14381), .B2(n14380), .A(n9894), .ZN(n20747) );
  AOI22_X1 U17796 ( .A1(n20650), .A2(n20747), .B1(n15319), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14382) );
  OAI21_X1 U17797 ( .B1(n15290), .B2(n15336), .A(n14382), .ZN(P1_U2870) );
  NOR2_X2 U17798 ( .A1(n20706), .A2(n17112), .ZN(n20698) );
  NAND2_X1 U17799 ( .A1(n15405), .A2(DATAI_1_), .ZN(n14386) );
  NAND2_X1 U17800 ( .A1(n15350), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14385) );
  AND2_X1 U17801 ( .A1(n14386), .A2(n14385), .ZN(n15389) );
  INV_X1 U17802 ( .A(n15389), .ZN(n14554) );
  NAND2_X1 U17803 ( .A1(n20698), .A2(n14554), .ZN(n14437) );
  AND2_X2 U17804 ( .A1(n15429), .A2(n17112), .ZN(n14429) );
  AOI22_X1 U17805 ( .A1(n14429), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U17806 ( .A1(n14437), .A2(n14387), .ZN(P1_U2953) );
  NAND2_X1 U17807 ( .A1(n15405), .A2(DATAI_4_), .ZN(n14389) );
  NAND2_X1 U17808 ( .A1(n15350), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14388) );
  AND2_X1 U17809 ( .A1(n14389), .A2(n14388), .ZN(n15377) );
  INV_X1 U17810 ( .A(n15377), .ZN(n20811) );
  NAND2_X1 U17811 ( .A1(n20698), .A2(n20811), .ZN(n14418) );
  AOI22_X1 U17812 ( .A1(n14429), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U17813 ( .A1(n14418), .A2(n14390), .ZN(P1_U2956) );
  INV_X1 U17814 ( .A(DATAI_2_), .ZN(n14392) );
  NAND2_X1 U17815 ( .A1(n15350), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14391) );
  OAI21_X1 U17816 ( .B1(n15350), .B2(n14392), .A(n14391), .ZN(n20803) );
  NAND2_X1 U17817 ( .A1(n20698), .A2(n20803), .ZN(n14433) );
  AOI22_X1 U17818 ( .A1(n14429), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U17819 ( .A1(n14433), .A2(n14393), .ZN(P1_U2954) );
  NAND2_X1 U17820 ( .A1(n15405), .A2(DATAI_6_), .ZN(n14395) );
  NAND2_X1 U17821 ( .A1(n15350), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14394) );
  AND2_X1 U17822 ( .A1(n14395), .A2(n14394), .ZN(n15420) );
  INV_X1 U17823 ( .A(n15420), .ZN(n20820) );
  NAND2_X1 U17824 ( .A1(n20698), .A2(n20820), .ZN(n14404) );
  AOI22_X1 U17825 ( .A1(n14429), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U17826 ( .A1(n14404), .A2(n14396), .ZN(P1_U2943) );
  INV_X1 U17827 ( .A(DATAI_8_), .ZN(n14398) );
  NAND2_X1 U17828 ( .A1(n15350), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14397) );
  OAI21_X1 U17829 ( .B1(n15350), .B2(n14398), .A(n14397), .ZN(n15416) );
  NAND2_X1 U17830 ( .A1(n20698), .A2(n15416), .ZN(n14423) );
  AOI22_X1 U17831 ( .A1(n14429), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U17832 ( .A1(n14423), .A2(n14399), .ZN(P1_U2960) );
  INV_X1 U17833 ( .A(DATAI_5_), .ZN(n14401) );
  NAND2_X1 U17834 ( .A1(n15350), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14400) );
  OAI21_X1 U17835 ( .B1(n15350), .B2(n14401), .A(n14400), .ZN(n20816) );
  NAND2_X1 U17836 ( .A1(n20698), .A2(n20816), .ZN(n14416) );
  AOI22_X1 U17837 ( .A1(n14429), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n14402) );
  NAND2_X1 U17838 ( .A1(n14416), .A2(n14402), .ZN(P1_U2957) );
  AOI22_X1 U17839 ( .A1(n14429), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U17840 ( .A1(n14404), .A2(n14403), .ZN(P1_U2958) );
  NAND2_X1 U17841 ( .A1(n15405), .A2(DATAI_7_), .ZN(n14406) );
  NAND2_X1 U17842 ( .A1(n15350), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14405) );
  INV_X1 U17843 ( .A(n20825), .ZN(n14407) );
  NAND2_X1 U17844 ( .A1(n20698), .A2(n14407), .ZN(n14410) );
  AOI22_X1 U17845 ( .A1(n14429), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U17846 ( .A1(n14410), .A2(n14408), .ZN(P1_U2944) );
  AOI22_X1 U17847 ( .A1(n14429), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U17848 ( .A1(n14410), .A2(n14409), .ZN(P1_U2959) );
  NAND2_X1 U17849 ( .A1(n15405), .A2(DATAI_10_), .ZN(n14412) );
  NAND2_X1 U17850 ( .A1(n15350), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14411) );
  AND2_X1 U17851 ( .A1(n14412), .A2(n14411), .ZN(n15415) );
  INV_X1 U17852 ( .A(n15415), .ZN(n14413) );
  NAND2_X1 U17853 ( .A1(n20698), .A2(n14413), .ZN(n14428) );
  AOI22_X1 U17854 ( .A1(n14429), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20706), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14414) );
  NAND2_X1 U17855 ( .A1(n14428), .A2(n14414), .ZN(P1_U2962) );
  AOI22_X1 U17856 ( .A1(n14429), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14415) );
  NAND2_X1 U17857 ( .A1(n14416), .A2(n14415), .ZN(P1_U2942) );
  AOI22_X1 U17858 ( .A1(n14429), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14417) );
  NAND2_X1 U17859 ( .A1(n14418), .A2(n14417), .ZN(P1_U2941) );
  INV_X1 U17860 ( .A(DATAI_0_), .ZN(n14420) );
  NAND2_X1 U17861 ( .A1(n15350), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14419) );
  OAI21_X1 U17862 ( .B1(n15350), .B2(n14420), .A(n14419), .ZN(n15396) );
  NAND2_X1 U17863 ( .A1(n20698), .A2(n15396), .ZN(n14435) );
  AOI22_X1 U17864 ( .A1(n14429), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n14421) );
  NAND2_X1 U17865 ( .A1(n14435), .A2(n14421), .ZN(P1_U2952) );
  AOI22_X1 U17866 ( .A1(n14429), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14422) );
  NAND2_X1 U17867 ( .A1(n14423), .A2(n14422), .ZN(P1_U2945) );
  NAND2_X1 U17868 ( .A1(n15405), .A2(DATAI_3_), .ZN(n14425) );
  NAND2_X1 U17869 ( .A1(n15350), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14424) );
  AND2_X1 U17870 ( .A1(n14425), .A2(n14424), .ZN(n15382) );
  INV_X1 U17871 ( .A(n15382), .ZN(n20807) );
  NAND2_X1 U17872 ( .A1(n20698), .A2(n20807), .ZN(n14431) );
  AOI22_X1 U17873 ( .A1(n14429), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20706), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n14426) );
  NAND2_X1 U17874 ( .A1(n14431), .A2(n14426), .ZN(P1_U2955) );
  AOI22_X1 U17875 ( .A1(n14429), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14427) );
  NAND2_X1 U17876 ( .A1(n14428), .A2(n14427), .ZN(P1_U2947) );
  AOI22_X1 U17877 ( .A1(n14429), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U17878 ( .A1(n14431), .A2(n14430), .ZN(P1_U2940) );
  AOI22_X1 U17879 ( .A1(n14429), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14432) );
  NAND2_X1 U17880 ( .A1(n14433), .A2(n14432), .ZN(P1_U2939) );
  AOI22_X1 U17881 ( .A1(n14429), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14434) );
  NAND2_X1 U17882 ( .A1(n14435), .A2(n14434), .ZN(P1_U2937) );
  AOI22_X1 U17883 ( .A1(n14429), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U17884 ( .A1(n14437), .A2(n14436), .ZN(P1_U2938) );
  XNOR2_X1 U17885 ( .A(n14439), .B(n14438), .ZN(n16878) );
  AOI22_X1 U17886 ( .A1(n14785), .A2(n16377), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n16465), .ZN(n14440) );
  OAI21_X1 U17887 ( .B1(n16878), .B2(n19836), .A(n14440), .ZN(P2_U2907) );
  INV_X1 U17888 ( .A(n17188), .ZN(n16810) );
  AOI211_X1 U17889 ( .C1(n17189), .C2(n17017), .A(n14959), .B(n16810), .ZN(
        n14451) );
  OR2_X1 U17890 ( .A1(n14442), .A2(n14441), .ZN(n14443) );
  AOI22_X1 U17891 ( .A1(n16944), .A2(n14445), .B1(n16970), .B2(n19818), .ZN(
        n14447) );
  OAI211_X1 U17892 ( .C1(n19814), .C2(n17180), .A(n14447), .B(n14446), .ZN(
        n14450) );
  OAI22_X1 U17893 ( .A1(n17183), .A2(n17017), .B1(n17193), .B2(n14448), .ZN(
        n14449) );
  OR3_X1 U17894 ( .A1(n14451), .A2(n14450), .A3(n14449), .ZN(P2_U3045) );
  NOR2_X1 U17895 ( .A1(n19814), .A2(n20300), .ZN(n14454) );
  INV_X1 U17896 ( .A(n20525), .ZN(n17002) );
  NOR3_X1 U17897 ( .A1(n19998), .A2(n17002), .A3(n14452), .ZN(n14453) );
  AOI211_X1 U17898 ( .C1(n20521), .C2(n19998), .A(n14454), .B(n14453), .ZN(
        n14463) );
  NAND2_X1 U17899 ( .A1(n11127), .A2(n20393), .ZN(n14455) );
  NAND2_X1 U17900 ( .A1(n20547), .A2(n14459), .ZN(n14460) );
  NAND2_X1 U17901 ( .A1(n14460), .A2(n17203), .ZN(n14461) );
  NAND2_X1 U17902 ( .A1(n19930), .A2(n14461), .ZN(n20540) );
  INV_X1 U17903 ( .A(n20540), .ZN(n20543) );
  NAND2_X1 U17904 ( .A1(n20543), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14462) );
  OAI21_X1 U17905 ( .B1(n14463), .B2(n20543), .A(n14462), .ZN(P2_U3604) );
  XNOR2_X1 U17906 ( .A(n14464), .B(n14465), .ZN(n15280) );
  INV_X1 U17907 ( .A(n14466), .ZN(n14467) );
  OAI21_X1 U17908 ( .B1(n9894), .B2(n14468), .A(n14467), .ZN(n15274) );
  INV_X1 U17909 ( .A(n15274), .ZN(n20735) );
  AOI22_X1 U17910 ( .A1(n20650), .A2(n20735), .B1(n15319), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14469) );
  OAI21_X1 U17911 ( .B1(n15280), .B2(n15336), .A(n14469), .ZN(P1_U2869) );
  NAND2_X1 U17912 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  NAND2_X1 U17913 ( .A1(n14470), .A2(n14473), .ZN(n16859) );
  AOI22_X1 U17914 ( .A1(n14785), .A2(n16365), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n16465), .ZN(n14474) );
  OAI21_X1 U17915 ( .B1(n16859), .B2(n19836), .A(n14474), .ZN(P2_U2906) );
  AOI22_X1 U17916 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20727), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14475) );
  OAI21_X1 U17917 ( .B1(n20720), .B2(n15282), .A(n14475), .ZN(n14476) );
  INV_X1 U17918 ( .A(n14476), .ZN(n14480) );
  OR2_X1 U17919 ( .A1(n14478), .A2(n14477), .ZN(n20746) );
  NAND3_X1 U17920 ( .A1(n20746), .A2(n20745), .A3(n20716), .ZN(n14479) );
  OAI211_X1 U17921 ( .C1(n15290), .C2(n15573), .A(n14480), .B(n14479), .ZN(
        P1_U2997) );
  NOR2_X1 U17922 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n17174), .ZN(n14509) );
  MUX2_X1 U17923 ( .A(n14481), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17090), .Z(n17096) );
  AOI22_X1 U17924 ( .A1(n14509), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17096), .B2(n17174), .ZN(n14503) );
  INV_X1 U17925 ( .A(n14485), .ZN(n15920) );
  AOI21_X1 U17926 ( .B1(n14178), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14482) );
  NOR2_X1 U17927 ( .A1(n14483), .A2(n14482), .ZN(n15928) );
  NAND3_X1 U17928 ( .A1(n14485), .A2(n14484), .A3(n15928), .ZN(n14497) );
  INV_X1 U17929 ( .A(n14486), .ZN(n14488) );
  NAND2_X1 U17930 ( .A1(n14489), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14487) );
  NAND2_X1 U17931 ( .A1(n14488), .A2(n14487), .ZN(n14494) );
  MUX2_X1 U17932 ( .A(n14488), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14178), .Z(n14491) );
  INV_X1 U17933 ( .A(n14489), .ZN(n14490) );
  NAND2_X1 U17934 ( .A1(n14491), .A2(n14490), .ZN(n14492) );
  AOI22_X1 U17935 ( .A1(n14495), .A2(n14494), .B1(n14493), .B2(n14492), .ZN(
        n14496) );
  OAI211_X1 U17936 ( .C1(n14500), .C2(n15917), .A(n14497), .B(n14496), .ZN(
        n14498) );
  AOI21_X1 U17937 ( .B1(n21031), .B2(n15920), .A(n14498), .ZN(n15932) );
  INV_X1 U17938 ( .A(n17090), .ZN(n14499) );
  MUX2_X1 U17939 ( .A(n14500), .B(n15932), .S(n14499), .Z(n17098) );
  INV_X1 U17940 ( .A(n17098), .ZN(n14501) );
  AOI22_X1 U17941 ( .A1(n14509), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n17174), .B2(n14501), .ZN(n14502) );
  NOR2_X1 U17942 ( .A1(n14503), .A2(n14502), .ZN(n17099) );
  INV_X1 U17943 ( .A(n17099), .ZN(n14510) );
  INV_X1 U17944 ( .A(n20913), .ZN(n21151) );
  NOR2_X1 U17945 ( .A1(n14505), .A2(n21151), .ZN(n14506) );
  XNOR2_X1 U17946 ( .A(n14506), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20621) );
  NOR2_X1 U17947 ( .A1(n20621), .A2(n14175), .ZN(n17164) );
  OAI21_X1 U17948 ( .B1(n17164), .B2(n17090), .A(n17174), .ZN(n14507) );
  AOI21_X1 U17949 ( .B1(n17090), .B2(n12920), .A(n14507), .ZN(n14508) );
  AOI21_X1 U17950 ( .B1(n14509), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n14508), .ZN(n17108) );
  OAI21_X1 U17951 ( .B1(n14510), .B2(n14504), .A(n17108), .ZN(n14533) );
  OAI21_X1 U17952 ( .B1(n14533), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14511), .ZN(
        n14512) );
  NAND2_X1 U17953 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21091), .ZN(n15910) );
  INV_X1 U17954 ( .A(n15910), .ZN(n14534) );
  NAND2_X1 U17955 ( .A1(n9707), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14517) );
  OAI21_X1 U17956 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9707), .A(n21270), 
        .ZN(n14514) );
  OAI21_X1 U17957 ( .B1(n14534), .B2(n21153), .A(n14514), .ZN(n14515) );
  NAND2_X1 U17958 ( .A1(n20782), .A2(n14515), .ZN(n14516) );
  OAI21_X1 U17959 ( .B1(n20782), .B2(n13362), .A(n14516), .ZN(P1_U3477) );
  NOR2_X1 U17960 ( .A1(n21152), .A2(n14534), .ZN(n14520) );
  INV_X1 U17961 ( .A(n14517), .ZN(n14518) );
  AND2_X1 U17962 ( .A1(n14518), .A2(n21273), .ZN(n15909) );
  OAI21_X1 U17963 ( .B1(n14520), .B2(n14519), .A(n20782), .ZN(n14521) );
  OAI21_X1 U17964 ( .B1(n20782), .B2(n21157), .A(n14521), .ZN(P1_U3476) );
  AOI21_X1 U17965 ( .B1(n20537), .B2(n19828), .A(n14525), .ZN(n14526) );
  INV_X1 U17966 ( .A(n14526), .ZN(P2_U2885) );
  NAND2_X1 U17967 ( .A1(n19998), .A2(n19814), .ZN(n14639) );
  OAI21_X1 U17968 ( .B1(n19998), .B2(n19814), .A(n14639), .ZN(n14527) );
  NOR2_X1 U17969 ( .A1(n14527), .A2(n14528), .ZN(n14641) );
  AOI21_X1 U17970 ( .B1(n14528), .B2(n14527), .A(n14641), .ZN(n14532) );
  INV_X1 U17971 ( .A(n19814), .ZN(n14529) );
  AOI22_X1 U17972 ( .A1(n16472), .A2(n14529), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n16465), .ZN(n14531) );
  NAND2_X1 U17973 ( .A1(n14785), .A2(n17046), .ZN(n14530) );
  OAI211_X1 U17974 ( .C1(n14532), .C2(n16475), .A(n14531), .B(n14530), .ZN(
        P2_U2918) );
  NOR2_X1 U17975 ( .A1(n14533), .A2(n17177), .ZN(n17117) );
  OAI22_X1 U17976 ( .A1(n13816), .A2(n21266), .B1(n14535), .B2(n14534), .ZN(
        n14536) );
  OAI21_X1 U17977 ( .B1(n17117), .B2(n14536), .A(n20782), .ZN(n14537) );
  OAI21_X1 U17978 ( .B1(n20782), .B2(n21199), .A(n14537), .ZN(P1_U3478) );
  AND2_X1 U17979 ( .A1(n14540), .A2(n14539), .ZN(n14541) );
  OR2_X1 U17980 ( .A1(n14538), .A2(n14541), .ZN(n20620) );
  OR2_X1 U17981 ( .A1(n14466), .A2(n14542), .ZN(n14543) );
  NAND2_X1 U17982 ( .A1(n17151), .A2(n14543), .ZN(n20729) );
  INV_X1 U17983 ( .A(n20729), .ZN(n20628) );
  AOI22_X1 U17984 ( .A1(n20650), .A2(n20628), .B1(n15319), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n14544) );
  OAI21_X1 U17985 ( .B1(n20620), .B2(n15336), .A(n14544), .ZN(P1_U2868) );
  NAND2_X1 U17986 ( .A1(n14470), .A2(n14545), .ZN(n14546) );
  NAND2_X1 U17987 ( .A1(n14632), .A2(n14546), .ZN(n16850) );
  AOI22_X1 U17988 ( .A1(n14785), .A2(n16356), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n16465), .ZN(n14547) );
  OAI21_X1 U17989 ( .B1(n16850), .B2(n19836), .A(n14547), .ZN(P2_U2905) );
  NOR2_X1 U17990 ( .A1(n11180), .A2(n16351), .ZN(n14551) );
  AOI21_X1 U17991 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16351), .A(n14551), .ZN(
        n14552) );
  OAI21_X1 U17992 ( .B1(n20155), .B2(n16354), .A(n14552), .ZN(P2_U2884) );
  AOI22_X1 U17993 ( .A1(DATAI_17_), .A2(n14553), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20829), .ZN(n20894) );
  AOI22_X1 U17994 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20829), .B1(DATAI_25_), 
        .B2(n14553), .ZN(n21284) );
  INV_X1 U17995 ( .A(n21284), .ZN(n21167) );
  INV_X1 U17996 ( .A(n21280), .ZN(n21170) );
  INV_X1 U17997 ( .A(n21152), .ZN(n14555) );
  OR2_X1 U17998 ( .A1(n21031), .A2(n14555), .ZN(n20854) );
  NAND3_X1 U17999 ( .A1(n21156), .A2(n21157), .A3(n13362), .ZN(n20791) );
  NOR2_X1 U18000 ( .A1(n21199), .A2(n20791), .ZN(n20847) );
  INV_X1 U18001 ( .A(n20847), .ZN(n14568) );
  OAI21_X1 U18002 ( .B1(n20854), .B2(n20942), .A(n14568), .ZN(n14558) );
  INV_X1 U18003 ( .A(n20791), .ZN(n14560) );
  AOI22_X1 U18004 ( .A1(n14558), .A2(n21273), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14560), .ZN(n20834) );
  INV_X1 U18005 ( .A(n20827), .ZN(n14567) );
  NAND2_X1 U18006 ( .A1(n14567), .A2(n13430), .ZN(n20800) );
  OAI22_X1 U18007 ( .A1(n21170), .A2(n20834), .B1(n20800), .B2(n14568), .ZN(
        n14557) );
  AOI21_X1 U18008 ( .B1(n20848), .B2(n21167), .A(n14557), .ZN(n14565) );
  NOR2_X1 U18009 ( .A1(n14558), .A2(n21266), .ZN(n14559) );
  OAI21_X1 U18010 ( .B1(n20881), .B2(n21232), .A(n14559), .ZN(n14563) );
  OAI21_X1 U18011 ( .B1(n21273), .B2(n14560), .A(n21272), .ZN(n14561) );
  INV_X1 U18012 ( .A(n14561), .ZN(n14562) );
  NAND2_X1 U18013 ( .A1(n20849), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14564) );
  OAI211_X1 U18014 ( .C1(n20894), .C2(n20866), .A(n14565), .B(n14564), .ZN(
        P1_U3042) );
  AOI22_X1 U18015 ( .A1(DATAI_16_), .A2(n14553), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20829), .ZN(n20797) );
  AOI22_X1 U18016 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20829), .B1(DATAI_24_), 
        .B2(n14553), .ZN(n21278) );
  INV_X1 U18017 ( .A(n21278), .ZN(n21163) );
  INV_X1 U18018 ( .A(n21264), .ZN(n21166) );
  NAND2_X1 U18019 ( .A1(n14567), .A2(n14566), .ZN(n20790) );
  OAI22_X1 U18020 ( .A1(n21166), .A2(n20834), .B1(n20790), .B2(n14568), .ZN(
        n14569) );
  AOI21_X1 U18021 ( .B1(n20848), .B2(n21163), .A(n14569), .ZN(n14571) );
  NAND2_X1 U18022 ( .A1(n20849), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14570) );
  OAI211_X1 U18023 ( .C1(n20797), .C2(n20866), .A(n14571), .B(n14570), .ZN(
        P1_U3041) );
  INV_X1 U18024 ( .A(n14572), .ZN(n14575) );
  INV_X1 U18025 ( .A(n14538), .ZN(n14574) );
  NAND2_X1 U18026 ( .A1(n14538), .A2(n14572), .ZN(n15332) );
  INV_X1 U18027 ( .A(n15332), .ZN(n14573) );
  AOI21_X1 U18028 ( .B1(n14575), .B2(n14574), .A(n14573), .ZN(n20652) );
  INV_X1 U18029 ( .A(n20652), .ZN(n14593) );
  INV_X1 U18030 ( .A(n14580), .ZN(n14582) );
  NAND2_X1 U18031 ( .A1(n14582), .A2(n14581), .ZN(n14583) );
  AOI21_X4 U18032 ( .B1(n14586), .B2(n14585), .A(n20561), .ZN(n15418) );
  NAND2_X1 U18033 ( .A1(n12658), .A2(n14587), .ZN(n14589) );
  INV_X1 U18034 ( .A(n15419), .ZN(n15408) );
  AOI22_X1 U18035 ( .A1(n15408), .A2(n20816), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n15407), .ZN(n14592) );
  OAI21_X1 U18036 ( .B1(n14593), .B2(n15421), .A(n14592), .ZN(P1_U2899) );
  INV_X1 U18037 ( .A(n20155), .ZN(n20530) );
  INV_X1 U18038 ( .A(n17022), .ZN(n17200) );
  NAND3_X1 U18039 ( .A1(n20530), .A2(n17200), .A3(n17023), .ZN(n14609) );
  OR2_X1 U18040 ( .A1(n11180), .A2(n14661), .ZN(n14607) );
  NAND2_X1 U18041 ( .A1(n14595), .A2(n14594), .ZN(n14671) );
  OAI21_X1 U18042 ( .B1(n14662), .B2(n11006), .A(n14596), .ZN(n14605) );
  INV_X1 U18043 ( .A(n14701), .ZN(n14598) );
  NAND2_X1 U18044 ( .A1(n14598), .A2(n14597), .ZN(n14665) );
  NAND2_X1 U18045 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14674) );
  INV_X1 U18046 ( .A(n14599), .ZN(n21424) );
  INV_X1 U18047 ( .A(n21424), .ZN(n21674) );
  NAND2_X1 U18048 ( .A1(n14674), .A2(n21674), .ZN(n14663) );
  XNOR2_X1 U18049 ( .A(n14663), .B(n11006), .ZN(n14600) );
  NAND2_X1 U18050 ( .A1(n14665), .A2(n14600), .ZN(n14603) );
  OAI211_X1 U18051 ( .C1(n11186), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14684), .B(n14601), .ZN(n14602) );
  NAND2_X1 U18052 ( .A1(n14603), .A2(n14602), .ZN(n14604) );
  AOI21_X1 U18053 ( .B1(n14671), .B2(n14605), .A(n14604), .ZN(n14606) );
  AND2_X1 U18054 ( .A1(n14607), .A2(n14606), .ZN(n14692) );
  INV_X1 U18055 ( .A(n14692), .ZN(n14694) );
  AOI22_X1 U18056 ( .A1(n14694), .A2(n17027), .B1(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17030), .ZN(n14608) );
  NAND2_X1 U18057 ( .A1(n14609), .A2(n14608), .ZN(P2_U3596) );
  XNOR2_X1 U18058 ( .A(n14610), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14611) );
  XNOR2_X1 U18059 ( .A(n14612), .B(n14611), .ZN(n15670) );
  INV_X1 U18060 ( .A(n20723), .ZN(n20724) );
  INV_X1 U18061 ( .A(n14613), .ZN(n14614) );
  NAND2_X1 U18062 ( .A1(n20756), .A2(n14614), .ZN(n14615) );
  NAND2_X1 U18063 ( .A1(n20772), .A2(n14615), .ZN(n17156) );
  AOI21_X1 U18064 ( .B1(n14616), .B2(n20724), .A(n17156), .ZN(n15865) );
  INV_X1 U18065 ( .A(n15865), .ZN(n15895) );
  INV_X1 U18066 ( .A(n14618), .ZN(n15326) );
  XNOR2_X1 U18067 ( .A(n14617), .B(n15326), .ZN(n20598) );
  NAND2_X1 U18068 ( .A1(n20727), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n15667) );
  OAI21_X1 U18069 ( .B1(n20774), .B2(n20598), .A(n15667), .ZN(n14619) );
  AOI21_X1 U18070 ( .B1(n15895), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14619), .ZN(n14624) );
  AND2_X1 U18071 ( .A1(n20771), .A2(n20770), .ZN(n20760) );
  NAND2_X1 U18072 ( .A1(n15845), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20755) );
  NAND2_X1 U18073 ( .A1(n14620), .A2(n20722), .ZN(n14621) );
  NAND2_X1 U18074 ( .A1(n14621), .A2(n20721), .ZN(n20737) );
  INV_X1 U18075 ( .A(n20725), .ZN(n14622) );
  INV_X1 U18076 ( .A(n15891), .ZN(n15885) );
  NAND2_X1 U18077 ( .A1(n15885), .A2(n15892), .ZN(n14623) );
  OAI211_X1 U18078 ( .C1(n15670), .C2(n20775), .A(n14624), .B(n14623), .ZN(
        P1_U3025) );
  XNOR2_X1 U18079 ( .A(n14625), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14628) );
  INV_X1 U18080 ( .A(n14626), .ZN(n14627) );
  NOR2_X1 U18081 ( .A1(n14628), .A2(n14627), .ZN(n20710) );
  AOI21_X1 U18082 ( .B1(n14628), .B2(n14627), .A(n20710), .ZN(n20739) );
  NAND2_X1 U18083 ( .A1(n20739), .A2(n20716), .ZN(n14631) );
  AND2_X1 U18084 ( .A1(n20727), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20734) );
  NOR2_X1 U18085 ( .A1(n20720), .A2(n15275), .ZN(n14629) );
  AOI211_X1 U18086 ( .C1(n20709), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20734), .B(n14629), .ZN(n14630) );
  OAI211_X1 U18087 ( .C1(n15573), .C2(n15280), .A(n14631), .B(n14630), .ZN(
        P1_U2996) );
  AOI21_X1 U18088 ( .B1(n14633), .B2(n14632), .A(n14809), .ZN(n14634) );
  INV_X1 U18089 ( .A(n14634), .ZN(n16833) );
  OAI222_X1 U18090 ( .A1(n19834), .A2(n14635), .B1(n16833), .B2(n19836), .C1(
        n14048), .C2(n19840), .ZN(P2_U2904) );
  INV_X1 U18091 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20682) );
  OAI222_X1 U18092 ( .A1(n15421), .A2(n14636), .B1(n15419), .B2(n15389), .C1(
        n15418), .C2(n20682), .ZN(P1_U2903) );
  INV_X1 U18093 ( .A(n20803), .ZN(n14637) );
  INV_X1 U18094 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20679) );
  OAI222_X1 U18095 ( .A1(n15421), .A2(n15290), .B1(n15419), .B2(n14637), .C1(
        n15418), .C2(n20679), .ZN(P1_U2902) );
  INV_X1 U18096 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20676) );
  OAI222_X1 U18097 ( .A1(n15421), .A2(n15280), .B1(n15419), .B2(n15382), .C1(
        n15418), .C2(n20676), .ZN(P1_U2901) );
  INV_X1 U18098 ( .A(n15396), .ZN(n14638) );
  INV_X1 U18099 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20687) );
  OAI222_X1 U18100 ( .A1(n15421), .A2(n15297), .B1(n15419), .B2(n14638), .C1(
        n15418), .C2(n20687), .ZN(P1_U2904) );
  INV_X1 U18101 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20674) );
  OAI222_X1 U18102 ( .A1(n15421), .A2(n20620), .B1(n15377), .B2(n15419), .C1(
        n15418), .C2(n20674), .ZN(P1_U2900) );
  INV_X1 U18103 ( .A(n14639), .ZN(n14640) );
  NOR2_X1 U18104 ( .A1(n14641), .A2(n14640), .ZN(n14647) );
  INV_X1 U18105 ( .A(n20537), .ZN(n16255) );
  OR2_X1 U18106 ( .A1(n14644), .A2(n14643), .ZN(n14645) );
  AND2_X1 U18107 ( .A1(n14642), .A2(n14645), .ZN(n16252) );
  NAND2_X1 U18108 ( .A1(n16255), .A2(n16252), .ZN(n14744) );
  OAI21_X1 U18109 ( .B1(n16255), .B2(n16252), .A(n14744), .ZN(n14646) );
  NOR2_X1 U18110 ( .A1(n14647), .A2(n14646), .ZN(n14746) );
  AOI21_X1 U18111 ( .B1(n14647), .B2(n14646), .A(n14746), .ZN(n14650) );
  INV_X1 U18112 ( .A(n16252), .ZN(n20535) );
  AOI22_X1 U18113 ( .A1(n16472), .A2(n20535), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n16465), .ZN(n14649) );
  NAND2_X1 U18114 ( .A1(n14785), .A2(n19870), .ZN(n14648) );
  OAI211_X1 U18115 ( .C1(n14650), .C2(n16475), .A(n14649), .B(n14648), .ZN(
        P2_U2917) );
  INV_X1 U18116 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14651) );
  NOR2_X1 U18117 ( .A1(n14652), .A2(n14651), .ZN(n14781) );
  NAND2_X1 U18118 ( .A1(n14653), .A2(n14781), .ZN(n14801) );
  XNOR2_X1 U18119 ( .A(n14784), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14660) );
  AND2_X1 U18120 ( .A1(n14655), .A2(n14656), .ZN(n14657) );
  NOR2_X1 U18121 ( .A1(n14654), .A2(n14657), .ZN(n16971) );
  NOR2_X1 U18122 ( .A1(n19832), .A2(n11427), .ZN(n14658) );
  AOI21_X1 U18123 ( .B1(n16971), .B2(n19832), .A(n14658), .ZN(n14659) );
  OAI21_X1 U18124 ( .B1(n14660), .B2(n16354), .A(n14659), .ZN(P2_U2882) );
  INV_X1 U18125 ( .A(n14661), .ZN(n14687) );
  NAND2_X1 U18126 ( .A1(n12315), .A2(n14663), .ZN(n14664) );
  INV_X1 U18127 ( .A(n14664), .ZN(n14670) );
  NAND2_X1 U18128 ( .A1(n14665), .A2(n14664), .ZN(n14668) );
  XNOR2_X1 U18129 ( .A(n21674), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14666) );
  NAND2_X1 U18130 ( .A1(n14684), .A2(n14666), .ZN(n14667) );
  NAND2_X1 U18131 ( .A1(n14668), .A2(n14667), .ZN(n14669) );
  AOI21_X1 U18132 ( .B1(n14671), .B2(n14670), .A(n14669), .ZN(n14672) );
  NAND2_X1 U18133 ( .A1(n14673), .A2(n14672), .ZN(n17028) );
  MUX2_X1 U18134 ( .A(n21424), .B(n17028), .S(n14715), .Z(n14717) );
  NAND2_X1 U18135 ( .A1(n19818), .A2(n14687), .ZN(n14683) );
  INV_X1 U18136 ( .A(n14674), .ZN(n14675) );
  NOR2_X1 U18137 ( .A1(n14676), .A2(n14675), .ZN(n14681) );
  INV_X1 U18138 ( .A(n14677), .ZN(n14679) );
  NAND2_X1 U18139 ( .A1(n14679), .A2(n14678), .ZN(n14685) );
  AOI22_X1 U18140 ( .A1(n14681), .A2(n14685), .B1(n14684), .B2(n14680), .ZN(
        n14682) );
  NAND2_X1 U18141 ( .A1(n14683), .A2(n14682), .ZN(n17020) );
  OAI21_X1 U18142 ( .B1(n17020), .B2(n20338), .A(n20227), .ZN(n14688) );
  MUX2_X1 U18143 ( .A(n14685), .B(n14684), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14686) );
  AOI21_X1 U18144 ( .B1(n11168), .B2(n14687), .A(n14686), .ZN(n17004) );
  NAND2_X1 U18145 ( .A1(n14688), .A2(n17004), .ZN(n14689) );
  OAI211_X1 U18146 ( .C1(n14690), .C2(n17020), .A(n14689), .B(n14715), .ZN(
        n14691) );
  AOI21_X1 U18147 ( .B1(n14692), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n14691), .ZN(n14693) );
  OAI21_X1 U18148 ( .B1(n14717), .B2(n20542), .A(n14693), .ZN(n14697) );
  NAND2_X1 U18149 ( .A1(n20542), .A2(n20533), .ZN(n19960) );
  INV_X1 U18150 ( .A(n19960), .ZN(n19962) );
  NAND2_X1 U18151 ( .A1(n14717), .A2(n19962), .ZN(n14696) );
  MUX2_X1 U18152 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14694), .S(
        n14715), .Z(n14718) );
  NAND2_X1 U18153 ( .A1(n14718), .A2(n20533), .ZN(n14695) );
  NAND3_X1 U18154 ( .A1(n14697), .A2(n14696), .A3(n14695), .ZN(n14698) );
  NAND2_X1 U18155 ( .A1(n14698), .A2(n17137), .ZN(n14720) );
  MUX2_X1 U18156 ( .A(n14701), .B(n14700), .S(n14699), .Z(n14704) );
  AND2_X1 U18157 ( .A1(n14708), .A2(n14702), .ZN(n14703) );
  NOR2_X1 U18158 ( .A1(n14704), .A2(n14703), .ZN(n20553) );
  OAI21_X1 U18159 ( .B1(n15939), .B2(n20450), .A(n17196), .ZN(n14706) );
  AND2_X1 U18160 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  AND2_X1 U18161 ( .A1(n14708), .A2(n14707), .ZN(n19737) );
  OAI21_X1 U18162 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19737), .ZN(n14712) );
  NAND2_X1 U18163 ( .A1(n14709), .A2(n11385), .ZN(n14711) );
  AND3_X1 U18164 ( .A1(n14712), .A2(n14711), .A3(n14710), .ZN(n14713) );
  OAI211_X1 U18165 ( .C1(n14715), .C2(n14714), .A(n20553), .B(n14713), .ZN(
        n14716) );
  AOI21_X1 U18166 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(n14719) );
  AND2_X1 U18167 ( .A1(n14720), .A2(n14719), .ZN(n17206) );
  AOI21_X1 U18168 ( .B1(n11628), .B2(n14721), .A(n19736), .ZN(n17198) );
  AOI21_X1 U18169 ( .B1(n17206), .B2(n17198), .A(n19859), .ZN(n14761) );
  OAI21_X1 U18170 ( .B1(n14761), .B2(n20300), .A(n14722), .ZN(P2_U3593) );
  AND2_X1 U18171 ( .A1(n14723), .A2(n14724), .ZN(n14726) );
  OR2_X1 U18172 ( .A1(n14726), .A2(n14725), .ZN(n15263) );
  INV_X1 U18173 ( .A(DATAI_9_), .ZN(n14728) );
  NAND2_X1 U18174 ( .A1(n15350), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14727) );
  OAI21_X1 U18175 ( .B1(n15350), .B2(n14728), .A(n14727), .ZN(n15423) );
  AOI22_X1 U18176 ( .A1(n15408), .A2(n15423), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15407), .ZN(n14729) );
  OAI21_X1 U18177 ( .B1(n15263), .B2(n15421), .A(n14729), .ZN(P1_U2895) );
  INV_X1 U18178 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21508) );
  NOR2_X1 U18179 ( .A1(n14894), .A2(n14730), .ZN(n14731) );
  OR2_X1 U18180 ( .A1(n15251), .A2(n14731), .ZN(n15877) );
  OAI222_X1 U18181 ( .A1(n15263), .A2(n15336), .B1(n20655), .B2(n21508), .C1(
        n15877), .C2(n15334), .ZN(P1_U2863) );
  NOR2_X1 U18182 ( .A1(n14801), .A2(n14732), .ZN(n14733) );
  NAND3_X1 U18183 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14767) );
  OAI211_X1 U18184 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14733), .A(
        n14767), .B(n19828), .ZN(n14738) );
  OR2_X1 U18185 ( .A1(n14654), .A2(n14735), .ZN(n14736) );
  AND2_X1 U18186 ( .A1(n14734), .A2(n14736), .ZN(n16956) );
  INV_X1 U18187 ( .A(n16956), .ZN(n16217) );
  MUX2_X1 U18188 ( .A(n16217), .B(n16211), .S(n16351), .Z(n14737) );
  NAND2_X1 U18189 ( .A1(n14738), .A2(n14737), .ZN(P2_U2881) );
  XOR2_X1 U18190 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14767), .Z(n14743)
         );
  INV_X1 U18191 ( .A(n14734), .ZN(n14741) );
  OAI21_X1 U18192 ( .B1(n14741), .B2(n11548), .A(n14764), .ZN(n16942) );
  MUX2_X1 U18193 ( .A(n16942), .B(n11434), .S(n16351), .Z(n14742) );
  OAI21_X1 U18194 ( .B1(n14743), .B2(n16354), .A(n14742), .ZN(P2_U2880) );
  INV_X1 U18195 ( .A(n14744), .ZN(n14745) );
  NOR2_X1 U18196 ( .A1(n14746), .A2(n14745), .ZN(n14753) );
  NAND2_X1 U18197 ( .A1(n14642), .A2(n14748), .ZN(n14750) );
  NAND2_X1 U18198 ( .A1(n14750), .A2(n14749), .ZN(n14751) );
  AND2_X1 U18199 ( .A1(n14747), .A2(n14751), .ZN(n20529) );
  XOR2_X1 U18200 ( .A(n20529), .B(n20155), .Z(n14752) );
  NOR2_X1 U18201 ( .A1(n14753), .A2(n14752), .ZN(n14778) );
  AOI21_X1 U18202 ( .B1(n14753), .B2(n14752), .A(n14778), .ZN(n14756) );
  INV_X1 U18203 ( .A(n16448), .ZN(n17053) );
  OAI22_X1 U18204 ( .A1(n19834), .A2(n17053), .B1(n19840), .B2(n19858), .ZN(
        n14754) );
  AOI21_X1 U18205 ( .B1(n16472), .B2(n20529), .A(n14754), .ZN(n14755) );
  OAI21_X1 U18206 ( .B1(n14756), .B2(n16475), .A(n14755), .ZN(P2_U2916) );
  OAI21_X1 U18207 ( .B1(n20523), .B2(n14757), .A(n19736), .ZN(n14760) );
  INV_X1 U18208 ( .A(n17196), .ZN(n20456) );
  NAND2_X1 U18209 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n20456), .ZN(n14758) );
  AOI21_X1 U18210 ( .B1(n14761), .B2(n17195), .A(n14758), .ZN(n14759) );
  AOI211_X1 U18211 ( .C1(n14761), .C2(n14760), .A(n19782), .B(n14759), .ZN(
        n14762) );
  INV_X1 U18212 ( .A(n14762), .ZN(P2_U3177) );
  AOI21_X1 U18213 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14766) );
  INV_X1 U18214 ( .A(n14766), .ZN(n16930) );
  INV_X1 U18215 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n21653) );
  NOR2_X1 U18216 ( .A1(n14767), .A2(n21653), .ZN(n14769) );
  NAND2_X1 U18217 ( .A1(n14769), .A2(n14768), .ZN(n14847) );
  OAI211_X1 U18218 ( .C1(n14769), .C2(n14768), .A(n14847), .B(n19828), .ZN(
        n14771) );
  NAND2_X1 U18219 ( .A1(n16351), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14770) );
  OAI211_X1 U18220 ( .C1(n16930), .C2(n16351), .A(n14771), .B(n14770), .ZN(
        P2_U2879) );
  OR2_X1 U18221 ( .A1(n9878), .A2(n14772), .ZN(n14773) );
  NAND2_X1 U18222 ( .A1(n14774), .A2(n14773), .ZN(n16961) );
  NOR2_X1 U18223 ( .A1(n20530), .A2(n20529), .ZN(n14777) );
  AND2_X1 U18224 ( .A1(n14747), .A2(n14775), .ZN(n14776) );
  OR2_X1 U18225 ( .A1(n9878), .A2(n14776), .ZN(n14796) );
  OAI21_X1 U18226 ( .B1(n14778), .B2(n14777), .A(n14796), .ZN(n14795) );
  INV_X1 U18227 ( .A(n14780), .ZN(n14782) );
  NOR3_X1 U18228 ( .A1(n14779), .A2(n14782), .A3(n14781), .ZN(n14783) );
  NOR2_X1 U18229 ( .A1(n14784), .A2(n14783), .ZN(n19829) );
  NAND3_X1 U18230 ( .A1(n14795), .A2(n16372), .A3(n19829), .ZN(n14787) );
  AOI22_X1 U18231 ( .A1(n14785), .A2(n19880), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n16465), .ZN(n14786) );
  OAI211_X1 U18232 ( .C1(n19836), .C2(n16961), .A(n14787), .B(n14786), .ZN(
        P2_U2914) );
  INV_X1 U18233 ( .A(n14788), .ZN(n14846) );
  XNOR2_X1 U18234 ( .A(n14847), .B(n14846), .ZN(n14794) );
  NOR2_X1 U18235 ( .A1(n14763), .A2(n14790), .ZN(n14791) );
  OR2_X1 U18236 ( .A1(n14789), .A2(n14791), .ZN(n16915) );
  NOR2_X1 U18237 ( .A1(n16915), .A2(n16351), .ZN(n14792) );
  AOI21_X1 U18238 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n16351), .A(n14792), .ZN(
        n14793) );
  OAI21_X1 U18239 ( .B1(n14794), .B2(n16354), .A(n14793), .ZN(P2_U2878) );
  XNOR2_X1 U18240 ( .A(n14795), .B(n19829), .ZN(n14799) );
  INV_X1 U18241 ( .A(n14796), .ZN(n19795) );
  INV_X1 U18242 ( .A(n16438), .ZN(n19876) );
  OAI22_X1 U18243 ( .A1(n19834), .A2(n19876), .B1(n19840), .B2(n14117), .ZN(
        n14797) );
  AOI21_X1 U18244 ( .B1(n19795), .B2(n16472), .A(n14797), .ZN(n14798) );
  OAI21_X1 U18245 ( .B1(n14799), .B2(n16475), .A(n14798), .ZN(P2_U2915) );
  INV_X1 U18246 ( .A(n14802), .ZN(n14838) );
  NOR2_X1 U18247 ( .A1(n16344), .A2(n14838), .ZN(n14827) );
  NAND2_X1 U18248 ( .A1(n14827), .A2(n14826), .ZN(n14832) );
  INV_X1 U18249 ( .A(n14803), .ZN(n14831) );
  NOR2_X1 U18250 ( .A1(n14832), .A2(n14831), .ZN(n14806) );
  OAI21_X1 U18251 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n16341) );
  OR2_X1 U18252 ( .A1(n14809), .A2(n14808), .ZN(n14810) );
  NAND2_X1 U18253 ( .A1(n14807), .A2(n14810), .ZN(n16819) );
  INV_X1 U18254 ( .A(n16819), .ZN(n19783) );
  NAND2_X1 U18255 ( .A1(n19840), .A2(n11056), .ZN(n14816) );
  INV_X1 U18256 ( .A(n14816), .ZN(n14812) );
  INV_X1 U18257 ( .A(n16464), .ZN(n14819) );
  INV_X1 U18258 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n19865) );
  AND2_X1 U18259 ( .A1(n19879), .A2(n14813), .ZN(n14814) );
  AOI22_X1 U18260 ( .A1(n16466), .A2(n14815), .B1(n16465), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14818) );
  INV_X1 U18261 ( .A(n16470), .ZN(n14938) );
  NAND2_X1 U18262 ( .A1(n14938), .A2(BUF2_REG_16__SCAN_IN), .ZN(n14817) );
  OAI211_X1 U18263 ( .C1(n14819), .C2(n19865), .A(n14818), .B(n14817), .ZN(
        n14820) );
  AOI21_X1 U18264 ( .B1(n19783), .B2(n16472), .A(n14820), .ZN(n14821) );
  OAI21_X1 U18265 ( .B1(n16475), .B2(n16341), .A(n14821), .ZN(P2_U2903) );
  AND2_X1 U18266 ( .A1(n16144), .A2(n14839), .ZN(n14841) );
  OR2_X1 U18267 ( .A1(n14841), .A2(n14824), .ZN(n14825) );
  INV_X1 U18268 ( .A(n16852), .ZN(n14830) );
  OAI211_X1 U18269 ( .C1(n14827), .C2(n14826), .A(n14832), .B(n19828), .ZN(
        n14829) );
  NAND2_X1 U18270 ( .A1(n16351), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14828) );
  OAI211_X1 U18271 ( .C1(n14830), .C2(n16351), .A(n14829), .B(n14828), .ZN(
        P2_U2873) );
  XNOR2_X1 U18272 ( .A(n14832), .B(n14831), .ZN(n14837) );
  XOR2_X1 U18273 ( .A(n14834), .B(n14833), .Z(n16836) );
  NAND2_X1 U18274 ( .A1(n16836), .A2(n19832), .ZN(n14836) );
  NAND2_X1 U18275 ( .A1(n16351), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14835) );
  OAI211_X1 U18276 ( .C1(n14837), .C2(n16354), .A(n14836), .B(n14835), .ZN(
        P2_U2872) );
  XNOR2_X1 U18277 ( .A(n16344), .B(n14838), .ZN(n14843) );
  NOR2_X1 U18278 ( .A1(n16144), .A2(n14839), .ZN(n14840) );
  MUX2_X1 U18279 ( .A(n16865), .B(n11569), .S(n16351), .Z(n14842) );
  OAI21_X1 U18280 ( .B1(n14843), .B2(n16354), .A(n14842), .ZN(P2_U2874) );
  OAI21_X1 U18281 ( .B1(n14789), .B2(n14845), .A(n14844), .ZN(n16896) );
  NOR2_X1 U18282 ( .A1(n14847), .A2(n14846), .ZN(n14849) );
  NAND2_X1 U18283 ( .A1(n14849), .A2(n14848), .ZN(n16350) );
  OAI211_X1 U18284 ( .C1(n14849), .C2(n14848), .A(n16350), .B(n19828), .ZN(
        n14851) );
  NAND2_X1 U18285 ( .A1(n16351), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14850) );
  OAI211_X1 U18286 ( .C1(n16896), .C2(n16351), .A(n14851), .B(n14850), .ZN(
        P2_U2877) );
  OAI21_X1 U18287 ( .B1(n19533), .B2(n12163), .A(n19519), .ZN(n14852) );
  NAND2_X1 U18288 ( .A1(n19532), .A2(n14852), .ZN(n19518) );
  NOR2_X1 U18289 ( .A1(n19726), .A2(n19518), .ZN(n14859) );
  NOR2_X1 U18290 ( .A1(n17357), .A2(n19586), .ZN(n14856) );
  NAND2_X1 U18291 ( .A1(n19715), .A2(n10355), .ZN(n19567) );
  AOI21_X1 U18292 ( .B1(n14853), .B2(n19567), .A(n19713), .ZN(n18299) );
  AOI21_X1 U18293 ( .B1(n14856), .B2(n18299), .A(n14854), .ZN(n14857) );
  NAND2_X1 U18294 ( .A1(n19513), .A2(n14855), .ZN(n17057) );
  NAND3_X1 U18295 ( .A1(n14857), .A2(n17057), .A3(n17140), .ZN(n19545) );
  NOR2_X1 U18296 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19666), .ZN(n19075) );
  INV_X1 U18297 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19065) );
  NAND3_X1 U18298 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19664)
         );
  NOR2_X1 U18299 ( .A1(n19065), .A2(n19664), .ZN(n14858) );
  MUX2_X1 U18300 ( .A(n14859), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19697), .Z(P3_U3284) );
  OAI211_X1 U18301 ( .C1(n19533), .C2(n12163), .A(n17817), .B(n19519), .ZN(
        n19064) );
  NOR2_X1 U18302 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n19064), .ZN(n14860) );
  INV_X1 U18303 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n17380) );
  NAND2_X1 U18304 ( .A1(n19519), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19678) );
  OAI21_X1 U18305 ( .B1(n14860), .B2(n19664), .A(n19220), .ZN(n19071) );
  INV_X1 U18306 ( .A(n19071), .ZN(n14861) );
  NOR2_X1 U18307 ( .A1(n19072), .A2(n19666), .ZN(n19073) );
  NAND2_X1 U18308 ( .A1(n19575), .A2(n19666), .ZN(n17360) );
  NOR2_X1 U18309 ( .A1(n19676), .A2(n19714), .ZN(n18741) );
  NOR2_X1 U18310 ( .A1(n19710), .A2(n18741), .ZN(n17066) );
  NOR2_X1 U18311 ( .A1(n19073), .A2(n17066), .ZN(n17067) );
  NOR2_X1 U18312 ( .A1(n14861), .A2(n17067), .ZN(n14863) );
  NAND3_X1 U18313 ( .A1(n19575), .A2(n19666), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19414) );
  INV_X1 U18314 ( .A(n19414), .ZN(n19067) );
  NOR2_X1 U18315 ( .A1(n19666), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19110) );
  OR2_X1 U18316 ( .A1(n19110), .A2(n14861), .ZN(n17065) );
  OR2_X1 U18317 ( .A1(n19067), .A2(n17065), .ZN(n14862) );
  MUX2_X1 U18318 ( .A(n14863), .B(n14862), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XNOR2_X1 U18319 ( .A(n14864), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15695) );
  NAND2_X1 U18320 ( .A1(n20727), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15689) );
  OAI21_X1 U18321 ( .B1(n15673), .B2(n14865), .A(n15689), .ZN(n14869) );
  NAND2_X1 U18322 ( .A1(n14871), .A2(n14872), .ZN(n14873) );
  NAND2_X1 U18323 ( .A1(n14986), .A2(n14873), .ZN(n15686) );
  OAI222_X1 U18324 ( .A1(n15336), .A2(n14870), .B1(n14874), .B2(n20655), .C1(
        n15686), .C2(n15334), .ZN(P1_U2843) );
  INV_X1 U18325 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19890) );
  AND2_X1 U18326 ( .A1(n15418), .A2(n20826), .ZN(n14875) );
  AOI22_X1 U18327 ( .A1(n15401), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15407), .ZN(n14878) );
  OAI211_X1 U18328 ( .C1(n15399), .C2(n19890), .A(n14879), .B(n14878), .ZN(
        P1_U2873) );
  INV_X1 U18329 ( .A(n15397), .ZN(n15390) );
  INV_X1 U18330 ( .A(DATAI_13_), .ZN(n14880) );
  INV_X1 U18331 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n17301) );
  MUX2_X1 U18332 ( .A(n14880), .B(n17301), .S(n15350), .Z(n20694) );
  OAI22_X1 U18333 ( .A1(n15390), .A2(n20694), .B1(n15418), .B2(n14303), .ZN(
        n14881) );
  AOI21_X1 U18334 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n15392), .A(n14881), .ZN(
        n14883) );
  NAND2_X1 U18335 ( .A1(n15401), .A2(DATAI_29_), .ZN(n14882) );
  OAI211_X1 U18336 ( .C1(n14870), .C2(n15421), .A(n14883), .B(n14882), .ZN(
        P1_U2875) );
  AOI22_X1 U18337 ( .A1(n20641), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20608), .ZN(n14887) );
  AOI21_X1 U18338 ( .B1(n9725), .B2(n21386), .A(n14889), .ZN(n14890) );
  OAI21_X1 U18339 ( .B1(n14870), .B2(n15269), .A(n14890), .ZN(P1_U2811) );
  INV_X1 U18340 ( .A(n14891), .ZN(n15333) );
  INV_X1 U18341 ( .A(n14892), .ZN(n15322) );
  NOR2_X1 U18342 ( .A1(n15330), .A2(n15322), .ZN(n15323) );
  OAI21_X1 U18343 ( .B1(n15323), .B2(n14893), .A(n14723), .ZN(n15650) );
  INV_X1 U18344 ( .A(n14894), .ZN(n14897) );
  NAND2_X1 U18345 ( .A1(n15327), .A2(n14895), .ZN(n14896) );
  NAND2_X1 U18346 ( .A1(n14897), .A2(n14896), .ZN(n15883) );
  OAI22_X1 U18347 ( .A1(n15883), .A2(n15334), .B1(n14898), .B2(n20655), .ZN(
        n14899) );
  INV_X1 U18348 ( .A(n14899), .ZN(n14900) );
  OAI21_X1 U18349 ( .B1(n15650), .B2(n15336), .A(n14900), .ZN(P1_U2864) );
  INV_X1 U18350 ( .A(n20585), .ZN(n20614) );
  NOR2_X1 U18351 ( .A1(n20614), .A2(n14901), .ZN(n15262) );
  NOR2_X1 U18352 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20594), .ZN(n14903) );
  NAND2_X1 U18353 ( .A1(n20638), .A2(n14979), .ZN(n20622) );
  AOI211_X1 U18354 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n14903), .A(n14902), .B(
        n20607), .ZN(n14904) );
  OAI21_X1 U18355 ( .B1(n14905), .B2(n20636), .A(n14904), .ZN(n14906) );
  AOI21_X1 U18356 ( .B1(n15262), .B2(P1_REIP_REG_8__SCAN_IN), .A(n14906), .ZN(
        n14907) );
  OAI21_X1 U18357 ( .B1(n15650), .B2(n15269), .A(n14907), .ZN(P1_U2832) );
  AOI21_X1 U18358 ( .B1(n14916), .B2(n13606), .A(n14915), .ZN(n14923) );
  NAND2_X1 U18359 ( .A1(n14923), .A2(n16715), .ZN(n14920) );
  OR2_X1 U18360 ( .A1(n15947), .A2(n16710), .ZN(n14918) );
  INV_X1 U18361 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n15949) );
  NOR2_X1 U18362 ( .A1(n16706), .A2(n15949), .ZN(n14929) );
  AOI21_X1 U18363 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14929), .ZN(n14917) );
  AND2_X1 U18364 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  AOI21_X1 U18365 ( .B1(n16697), .B2(n14935), .A(n14921), .ZN(n14922) );
  OAI21_X1 U18366 ( .B1(n14936), .B2(n16680), .A(n14922), .ZN(P2_U2985) );
  AOI21_X1 U18367 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14926), .A(
        n14927), .ZN(n14925) );
  AOI211_X1 U18368 ( .C1(n14927), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        n14928) );
  AOI211_X1 U18369 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14930), .A(
        n14929), .B(n14928), .ZN(n14934) );
  AOI21_X1 U18370 ( .B1(n13648), .B2(n14932), .A(n14931), .ZN(n16370) );
  NAND2_X1 U18371 ( .A1(n16370), .A2(n16989), .ZN(n14933) );
  AOI22_X1 U18372 ( .A1(n16464), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n16465), .ZN(n14940) );
  NAND2_X1 U18373 ( .A1(n14938), .A2(BUF2_REG_31__SCAN_IN), .ZN(n14939) );
  OAI211_X1 U18374 ( .C1(n14937), .C2(n16441), .A(n14940), .B(n14939), .ZN(
        P2_U2888) );
  NAND2_X1 U18375 ( .A1(n16265), .A2(n19819), .ZN(n14949) );
  AOI22_X1 U18376 ( .A1(n19789), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n14941), .ZN(n14943) );
  NAND2_X1 U18377 ( .A1(n19787), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14942) );
  OAI211_X1 U18378 ( .C1(n14945), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14946) );
  AOI21_X1 U18379 ( .B1(n14947), .B2(n19809), .A(n14946), .ZN(n14948) );
  OAI211_X1 U18380 ( .C1(n14937), .C2(n19813), .A(n14949), .B(n14948), .ZN(
        P2_U2824) );
  OAI21_X1 U18381 ( .B1(n14959), .B2(n16806), .A(n17183), .ZN(n14969) );
  XNOR2_X1 U18382 ( .A(n14951), .B(n14950), .ZN(n14974) );
  OAI21_X1 U18383 ( .B1(n14954), .B2(n14953), .A(n14952), .ZN(n14973) );
  INV_X1 U18384 ( .A(n14973), .ZN(n14957) );
  AOI22_X1 U18385 ( .A1(n16944), .A2(n14957), .B1(n14956), .B2(n14955), .ZN(
        n14965) );
  NAND2_X1 U18386 ( .A1(n14959), .A2(n14958), .ZN(n14960) );
  OR2_X1 U18387 ( .A1(n16806), .A2(n14960), .ZN(n14962) );
  NOR2_X1 U18388 ( .A1(n16706), .A2(n11130), .ZN(n14971) );
  INV_X1 U18389 ( .A(n14971), .ZN(n14961) );
  OAI211_X1 U18390 ( .C1(n16252), .C2(n17180), .A(n14962), .B(n14961), .ZN(
        n14963) );
  INV_X1 U18391 ( .A(n14963), .ZN(n14964) );
  OAI211_X1 U18392 ( .C1(n17193), .C2(n14974), .A(n14965), .B(n14964), .ZN(
        n14968) );
  INV_X1 U18393 ( .A(n14966), .ZN(n14967) );
  AOI211_X1 U18394 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n14969), .A(
        n14968), .B(n14967), .ZN(n14970) );
  OAI21_X1 U18395 ( .B1(n9703), .B2(n17185), .A(n14970), .ZN(P2_U3044) );
  INV_X1 U18396 ( .A(n16244), .ZN(n14977) );
  AOI21_X1 U18397 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14971), .ZN(n14972) );
  OAI21_X1 U18398 ( .B1(n16680), .B2(n14973), .A(n14972), .ZN(n14976) );
  NOR2_X1 U18399 ( .A1(n14974), .A2(n16712), .ZN(n14975) );
  AOI211_X1 U18400 ( .C1(n16692), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n14978) );
  OAI21_X1 U18401 ( .B1(n10864), .B2(n16695), .A(n14978), .ZN(P2_U3012) );
  OR2_X1 U18402 ( .A1(n14979), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14982) );
  INV_X1 U18403 ( .A(n14980), .ZN(n14981) );
  MUX2_X1 U18404 ( .A(n14982), .B(n14981), .S(n21407), .Z(P1_U3487) );
  AOI21_X1 U18405 ( .B1(n9725), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14996) );
  AOI21_X1 U18406 ( .B1(n14985), .B2(n14984), .A(n14983), .ZN(n15435) );
  NAND2_X1 U18407 ( .A1(n15435), .A2(n20601), .ZN(n14994) );
  INV_X1 U18408 ( .A(n14986), .ZN(n14988) );
  OAI22_X1 U18409 ( .A1(n14988), .A2(n13528), .B1(n14871), .B2(n14987), .ZN(
        n14990) );
  XNOR2_X1 U18410 ( .A(n14990), .B(n14989), .ZN(n15683) );
  AOI22_X1 U18411 ( .A1(n20641), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20608), .ZN(n14991) );
  OAI21_X1 U18412 ( .B1(n20637), .B2(n15433), .A(n14991), .ZN(n14992) );
  AOI21_X1 U18413 ( .B1(n15683), .B2(n20627), .A(n14992), .ZN(n14993) );
  OAI211_X1 U18414 ( .C1(n14996), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        P1_U2810) );
  AOI21_X1 U18415 ( .B1(n14998), .B2(n14997), .A(n14866), .ZN(n15450) );
  INV_X1 U18416 ( .A(n15450), .ZN(n15349) );
  INV_X1 U18417 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15446) );
  OAI21_X1 U18418 ( .B1(n15012), .B2(n14999), .A(n14871), .ZN(n15700) );
  NOR2_X1 U18419 ( .A1(n15700), .A2(n20648), .ZN(n15005) );
  AOI22_X1 U18420 ( .A1(n20641), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20608), .ZN(n15003) );
  INV_X1 U18421 ( .A(n15000), .ZN(n15001) );
  NAND2_X1 U18422 ( .A1(n15001), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15002) );
  OAI211_X1 U18423 ( .C1(n20637), .C2(n15448), .A(n15003), .B(n15002), .ZN(
        n15004) );
  OAI21_X1 U18424 ( .B1(n15349), .B2(n15269), .A(n15007), .ZN(P1_U2812) );
  OAI21_X1 U18425 ( .B1(n15008), .B2(n15009), .A(n14997), .ZN(n15460) );
  AND2_X1 U18426 ( .A1(n15024), .A2(n15010), .ZN(n15011) );
  NOR2_X1 U18427 ( .A1(n15012), .A2(n15011), .ZN(n15705) );
  INV_X1 U18428 ( .A(n15013), .ZN(n15014) );
  NAND2_X1 U18429 ( .A1(n20585), .A2(n15014), .ZN(n15028) );
  NAND2_X1 U18430 ( .A1(n15294), .A2(n15454), .ZN(n15016) );
  AOI22_X1 U18431 ( .A1(n20641), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20608), .ZN(n15015) );
  OAI211_X1 U18432 ( .C1(n15452), .C2(n15028), .A(n15016), .B(n15015), .ZN(
        n15019) );
  INV_X1 U18433 ( .A(n15059), .ZN(n15038) );
  NOR3_X1 U18434 ( .A1(n15038), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15017), 
        .ZN(n15018) );
  AOI211_X1 U18435 ( .C1(n20627), .C2(n15705), .A(n15019), .B(n15018), .ZN(
        n15020) );
  OAI21_X1 U18436 ( .B1(n15460), .B2(n15269), .A(n15020), .ZN(P1_U2813) );
  AOI21_X1 U18437 ( .B1(n15023), .B2(n15022), .A(n15008), .ZN(n15467) );
  INV_X1 U18438 ( .A(n15467), .ZN(n15358) );
  INV_X1 U18439 ( .A(n15024), .ZN(n15025) );
  AOI21_X1 U18440 ( .B1(n15026), .B2(n15041), .A(n15025), .ZN(n15719) );
  NOR2_X1 U18441 ( .A1(n20637), .A2(n15465), .ZN(n15030) );
  INV_X1 U18442 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U18443 ( .A1(n20641), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20608), .ZN(n15027) );
  OAI21_X1 U18444 ( .B1(n15028), .B2(n15031), .A(n15027), .ZN(n15029) );
  AOI211_X1 U18445 ( .C1(n15719), .C2(n20627), .A(n15030), .B(n15029), .ZN(
        n15034) );
  NAND3_X1 U18446 ( .A1(n15059), .A2(n15032), .A3(n15031), .ZN(n15033) );
  OAI211_X1 U18447 ( .C1(n15358), .C2(n15269), .A(n15034), .B(n15033), .ZN(
        P1_U2814) );
  OAI21_X1 U18448 ( .B1(n15035), .B2(n15036), .A(n15022), .ZN(n15477) );
  XNOR2_X1 U18449 ( .A(P1_REIP_REG_24__SCAN_IN), .B(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15037) );
  NOR2_X1 U18450 ( .A1(n15038), .A2(n15037), .ZN(n15047) );
  NAND2_X1 U18451 ( .A1(n15052), .A2(n15039), .ZN(n15040) );
  NAND2_X1 U18452 ( .A1(n15041), .A2(n15040), .ZN(n15732) );
  NAND2_X1 U18453 ( .A1(n20585), .A2(n15042), .ZN(n15064) );
  INV_X1 U18454 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21659) );
  AOI22_X1 U18455 ( .A1(n20641), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20608), .ZN(n15043) );
  OAI21_X1 U18456 ( .B1(n15064), .B2(n21659), .A(n15043), .ZN(n15044) );
  AOI21_X1 U18457 ( .B1(n15294), .B2(n15474), .A(n15044), .ZN(n15045) );
  OAI21_X1 U18458 ( .B1(n15732), .B2(n20648), .A(n15045), .ZN(n15046) );
  NOR2_X1 U18459 ( .A1(n15047), .A2(n15046), .ZN(n15048) );
  OAI21_X1 U18460 ( .B1(n15477), .B2(n15269), .A(n15048), .ZN(P1_U2815) );
  AOI21_X1 U18461 ( .B1(n15049), .B2(n9716), .A(n15035), .ZN(n15487) );
  INV_X1 U18462 ( .A(n15487), .ZN(n15366) );
  INV_X1 U18463 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15058) );
  OR2_X1 U18464 ( .A1(n15070), .A2(n15050), .ZN(n15051) );
  NAND2_X1 U18465 ( .A1(n15052), .A2(n15051), .ZN(n15733) );
  INV_X1 U18466 ( .A(n15485), .ZN(n15055) );
  AOI22_X1 U18467 ( .A1(n20641), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20608), .ZN(n15053) );
  OAI21_X1 U18468 ( .B1(n15064), .B2(n15058), .A(n15053), .ZN(n15054) );
  AOI21_X1 U18469 ( .B1(n15294), .B2(n15055), .A(n15054), .ZN(n15056) );
  OAI21_X1 U18470 ( .B1(n15733), .B2(n20648), .A(n15056), .ZN(n15057) );
  AOI21_X1 U18471 ( .B1(n15059), .B2(n15058), .A(n15057), .ZN(n15060) );
  OAI21_X1 U18472 ( .B1(n15366), .B2(n15269), .A(n15060), .ZN(P1_U2816) );
  OAI21_X1 U18473 ( .B1(n15061), .B2(n15062), .A(n9716), .ZN(n15490) );
  INV_X1 U18474 ( .A(n15063), .ZN(n15066) );
  INV_X1 U18475 ( .A(n15064), .ZN(n15065) );
  OAI21_X1 U18476 ( .B1(n15066), .B2(P1_REIP_REG_23__SCAN_IN), .A(n15065), 
        .ZN(n15074) );
  INV_X1 U18477 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21540) );
  OAI22_X1 U18478 ( .A1(n20610), .A2(n21540), .B1(n21672), .B2(n20636), .ZN(
        n15072) );
  AND2_X1 U18479 ( .A1(n15067), .A2(n15068), .ZN(n15069) );
  OR2_X1 U18480 ( .A1(n15070), .A2(n15069), .ZN(n15744) );
  NOR2_X1 U18481 ( .A1(n15744), .A2(n20648), .ZN(n15071) );
  AOI211_X1 U18482 ( .C1(n15294), .C2(n15491), .A(n15072), .B(n15071), .ZN(
        n15073) );
  OAI211_X1 U18483 ( .C1(n15490), .C2(n15269), .A(n15074), .B(n15073), .ZN(
        P1_U2817) );
  INV_X1 U18484 ( .A(n15097), .ZN(n15077) );
  INV_X1 U18485 ( .A(n15075), .ZN(n15076) );
  OAI21_X1 U18486 ( .B1(n9787), .B2(n15077), .A(n15076), .ZN(n15078) );
  INV_X1 U18487 ( .A(n15078), .ZN(n15079) );
  OR2_X1 U18488 ( .A1(n15079), .A2(n15061), .ZN(n15501) );
  INV_X1 U18489 ( .A(n15080), .ZN(n15083) );
  INV_X1 U18490 ( .A(n15081), .ZN(n15093) );
  INV_X1 U18491 ( .A(n15067), .ZN(n15082) );
  AOI21_X1 U18492 ( .B1(n15083), .B2(n15093), .A(n15082), .ZN(n15758) );
  INV_X1 U18493 ( .A(n15084), .ZN(n15503) );
  AOI22_X1 U18494 ( .A1(n20641), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20608), .ZN(n15087) );
  NAND3_X1 U18495 ( .A1(n20585), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n15085), 
        .ZN(n15086) );
  OAI211_X1 U18496 ( .C1(n20637), .C2(n15503), .A(n15087), .B(n15086), .ZN(
        n15089) );
  INV_X1 U18497 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15513) );
  NOR3_X1 U18498 ( .A1(n15100), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n15513), 
        .ZN(n15088) );
  AOI211_X1 U18499 ( .C1(n15758), .C2(n20627), .A(n15089), .B(n15088), .ZN(
        n15090) );
  OAI21_X1 U18500 ( .B1(n15269), .B2(n15501), .A(n15090), .ZN(P1_U2818) );
  NAND2_X1 U18501 ( .A1(n20585), .A2(n15091), .ZN(n15107) );
  AOI22_X1 U18502 ( .A1(n20641), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20608), .ZN(n15092) );
  OAI21_X1 U18503 ( .B1(n15107), .B2(n15513), .A(n15092), .ZN(n15096) );
  OAI21_X1 U18504 ( .B1(n15094), .B2(n15104), .A(n15093), .ZN(n15769) );
  NOR2_X1 U18505 ( .A1(n15769), .A2(n20648), .ZN(n15095) );
  AOI211_X1 U18506 ( .C1(n15294), .C2(n15516), .A(n15096), .B(n15095), .ZN(
        n15099) );
  XNOR2_X1 U18507 ( .A(n9787), .B(n15097), .ZN(n15307) );
  NAND2_X1 U18508 ( .A1(n15307), .A2(n20601), .ZN(n15098) );
  OAI211_X1 U18509 ( .C1(n15100), .C2(P1_REIP_REG_21__SCAN_IN), .A(n15099), 
        .B(n15098), .ZN(P1_U2819) );
  INV_X1 U18510 ( .A(n15101), .ZN(n15103) );
  OAI21_X1 U18511 ( .B1(n15103), .B2(n10777), .A(n9787), .ZN(n15525) );
  AOI21_X1 U18512 ( .B1(n15105), .B2(n15120), .A(n15104), .ZN(n15773) );
  AOI22_X1 U18513 ( .A1(n20641), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20608), .ZN(n15106) );
  OAI21_X1 U18514 ( .B1(n20637), .B2(n15528), .A(n15106), .ZN(n15110) );
  NAND3_X1 U18515 ( .A1(n15115), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n15108) );
  INV_X1 U18516 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15526) );
  AOI21_X1 U18517 ( .B1(n15108), .B2(n15526), .A(n15107), .ZN(n15109) );
  AOI211_X1 U18518 ( .C1(n15773), .C2(n20627), .A(n15110), .B(n15109), .ZN(
        n15111) );
  OAI21_X1 U18519 ( .B1(n15269), .B2(n15525), .A(n15111), .ZN(P1_U2820) );
  OR2_X1 U18520 ( .A1(n15112), .A2(n15113), .ZN(n15114) );
  NAND2_X1 U18521 ( .A1(n15101), .A2(n15114), .ZN(n15536) );
  INV_X1 U18522 ( .A(n15115), .ZN(n15116) );
  NOR2_X1 U18523 ( .A1(n15116), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15137) );
  AND2_X1 U18524 ( .A1(n20585), .A2(n15117), .ZN(n15142) );
  OAI21_X1 U18525 ( .B1(n15137), .B2(n15142), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15129) );
  INV_X1 U18526 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21571) );
  INV_X1 U18527 ( .A(n15118), .ZN(n15132) );
  INV_X1 U18528 ( .A(n15119), .ZN(n15121) );
  OAI21_X1 U18529 ( .B1(n15132), .B2(n15121), .A(n15120), .ZN(n15781) );
  INV_X1 U18530 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15123) );
  NAND2_X1 U18531 ( .A1(n20641), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n15122) );
  OAI211_X1 U18532 ( .C1(n20636), .C2(n15123), .A(n15122), .B(n20622), .ZN(
        n15124) );
  AOI21_X1 U18533 ( .B1(n15294), .B2(n15537), .A(n15124), .ZN(n15125) );
  OAI21_X1 U18534 ( .B1(n15781), .B2(n20648), .A(n15125), .ZN(n15126) );
  AOI21_X1 U18535 ( .B1(n15127), .B2(n21571), .A(n15126), .ZN(n15128) );
  OAI211_X1 U18536 ( .C1(n15536), .C2(n15269), .A(n15129), .B(n15128), .ZN(
        P1_U2821) );
  INV_X1 U18537 ( .A(n15112), .ZN(n15130) );
  AOI21_X1 U18538 ( .B1(n15133), .B2(n15131), .A(n15132), .ZN(n15791) );
  NAND2_X1 U18539 ( .A1(n20641), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n15134) );
  OAI211_X1 U18540 ( .C1(n20636), .C2(n10438), .A(n15134), .B(n20622), .ZN(
        n15135) );
  AOI21_X1 U18541 ( .B1(n15142), .B2(P1_REIP_REG_18__SCAN_IN), .A(n15135), 
        .ZN(n15136) );
  OAI21_X1 U18542 ( .B1(n20637), .B2(n15547), .A(n15136), .ZN(n15138) );
  AOI211_X1 U18543 ( .C1(n15791), .C2(n20627), .A(n15138), .B(n15137), .ZN(
        n15139) );
  OAI21_X1 U18544 ( .B1(n15269), .B2(n15545), .A(n15139), .ZN(P1_U2822) );
  AOI21_X1 U18545 ( .B1(n15140), .B2(n9724), .A(n9786), .ZN(n15561) );
  INV_X1 U18546 ( .A(n15561), .ZN(n15395) );
  INV_X1 U18547 ( .A(n15159), .ZN(n15141) );
  NOR2_X1 U18548 ( .A1(n15177), .A2(n15141), .ZN(n15143) );
  OAI21_X1 U18549 ( .B1(n15143), .B2(P1_REIP_REG_17__SCAN_IN), .A(n15142), 
        .ZN(n15151) );
  OR2_X1 U18550 ( .A1(n15145), .A2(n15144), .ZN(n15146) );
  AND2_X1 U18551 ( .A1(n15131), .A2(n15146), .ZN(n15800) );
  NOR2_X1 U18552 ( .A1(n20610), .A2(n21516), .ZN(n15147) );
  AOI211_X1 U18553 ( .C1(n20608), .C2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20607), .B(n15147), .ZN(n15148) );
  OAI21_X1 U18554 ( .B1(n20637), .B2(n15559), .A(n15148), .ZN(n15149) );
  AOI21_X1 U18555 ( .B1(n15800), .B2(n20627), .A(n15149), .ZN(n15150) );
  OAI211_X1 U18556 ( .C1(n15395), .C2(n15269), .A(n15151), .B(n15150), .ZN(
        P1_U2823) );
  OAI21_X1 U18557 ( .B1(n9784), .B2(n9901), .A(n9724), .ZN(n15572) );
  XNOR2_X1 U18558 ( .A(n15152), .B(n15153), .ZN(n15813) );
  INV_X1 U18559 ( .A(n15813), .ZN(n15163) );
  NAND2_X1 U18560 ( .A1(n15204), .A2(n15154), .ZN(n15155) );
  NAND2_X1 U18561 ( .A1(n20585), .A2(n15155), .ZN(n15189) );
  INV_X1 U18562 ( .A(n15189), .ZN(n15175) );
  NAND2_X1 U18563 ( .A1(n20641), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15156) );
  OAI211_X1 U18564 ( .C1(n20636), .C2(n10437), .A(n15156), .B(n20622), .ZN(
        n15157) );
  AOI21_X1 U18565 ( .B1(n15175), .B2(P1_REIP_REG_16__SCAN_IN), .A(n15157), 
        .ZN(n15158) );
  OAI21_X1 U18566 ( .B1(n20637), .B2(n15568), .A(n15158), .ZN(n15162) );
  INV_X1 U18567 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21367) );
  INV_X1 U18568 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15160) );
  AOI211_X1 U18569 ( .C1(n21367), .C2(n15160), .A(n15159), .B(n15177), .ZN(
        n15161) );
  AOI211_X1 U18570 ( .C1(n20627), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15164) );
  OAI21_X1 U18571 ( .B1(n15269), .B2(n15572), .A(n15164), .ZN(P1_U2824) );
  INV_X1 U18572 ( .A(n15165), .ZN(n15167) );
  INV_X1 U18573 ( .A(n15166), .ZN(n15194) );
  NAND2_X1 U18574 ( .A1(n15165), .A2(n15194), .ZN(n15195) );
  OAI21_X1 U18575 ( .B1(n15167), .B2(n15229), .A(n15195), .ZN(n15168) );
  NAND2_X1 U18576 ( .A1(n15197), .A2(n15182), .ZN(n15181) );
  AOI21_X1 U18577 ( .B1(n15181), .B2(n15169), .A(n9784), .ZN(n15583) );
  INV_X1 U18578 ( .A(n15583), .ZN(n15406) );
  NAND2_X1 U18579 ( .A1(n15185), .A2(n15170), .ZN(n15171) );
  AND2_X1 U18580 ( .A1(n15152), .A2(n15171), .ZN(n15819) );
  NAND2_X1 U18581 ( .A1(n20641), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15172) );
  OAI211_X1 U18582 ( .C1(n20636), .C2(n15173), .A(n15172), .B(n20622), .ZN(
        n15174) );
  AOI21_X1 U18583 ( .B1(n15175), .B2(P1_REIP_REG_15__SCAN_IN), .A(n15174), 
        .ZN(n15176) );
  OAI21_X1 U18584 ( .B1(n20637), .B2(n15581), .A(n15176), .ZN(n15179) );
  NOR2_X1 U18585 ( .A1(n15177), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15178) );
  AOI211_X1 U18586 ( .C1(n15819), .C2(n20627), .A(n15179), .B(n15178), .ZN(
        n15180) );
  OAI21_X1 U18587 ( .B1(n15269), .B2(n15406), .A(n15180), .ZN(P1_U2825) );
  OAI21_X1 U18588 ( .B1(n15197), .B2(n15182), .A(n15181), .ZN(n15591) );
  OR2_X1 U18589 ( .A1(n15202), .A2(n15183), .ZN(n15184) );
  AND2_X1 U18590 ( .A1(n15185), .A2(n15184), .ZN(n15826) );
  AOI21_X1 U18591 ( .B1(n20608), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20607), .ZN(n15187) );
  NAND2_X1 U18592 ( .A1(n20641), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n15186) );
  OAI211_X1 U18593 ( .C1(n20637), .C2(n15594), .A(n15187), .B(n15186), .ZN(
        n15192) );
  INV_X1 U18594 ( .A(n15188), .ZN(n15213) );
  AOI21_X1 U18595 ( .B1(n15213), .B2(P1_REIP_REG_13__SCAN_IN), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15190) );
  NOR2_X1 U18596 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  AOI211_X1 U18597 ( .C1(n15826), .C2(n20627), .A(n15192), .B(n15191), .ZN(
        n15193) );
  OAI21_X1 U18598 ( .B1(n15269), .B2(n15591), .A(n15193), .ZN(P1_U2826) );
  OAI21_X1 U18599 ( .B1(n15165), .B2(n15194), .A(n15195), .ZN(n15228) );
  OAI21_X1 U18600 ( .B1(n15228), .B2(n15229), .A(n15195), .ZN(n15217) );
  NAND2_X1 U18601 ( .A1(n15217), .A2(n15216), .ZN(n15215) );
  INV_X1 U18602 ( .A(n15196), .ZN(n15198) );
  AOI21_X1 U18603 ( .B1(n15215), .B2(n15198), .A(n15197), .ZN(n15608) );
  INV_X1 U18604 ( .A(n15608), .ZN(n15411) );
  INV_X1 U18605 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15212) );
  INV_X1 U18606 ( .A(n15199), .ZN(n15201) );
  AOI21_X1 U18607 ( .B1(n15201), .B2(n15218), .A(n15200), .ZN(n15203) );
  OR2_X1 U18608 ( .A1(n15203), .A2(n15202), .ZN(n15836) );
  NOR2_X1 U18609 ( .A1(n15836), .A2(n20648), .ZN(n15211) );
  INV_X1 U18610 ( .A(n15204), .ZN(n15205) );
  AND2_X1 U18611 ( .A1(n20585), .A2(n15205), .ZN(n15222) );
  INV_X1 U18612 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15207) );
  NAND2_X1 U18613 ( .A1(n20641), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n15206) );
  OAI211_X1 U18614 ( .C1(n20636), .C2(n15207), .A(n15206), .B(n20622), .ZN(
        n15208) );
  AOI21_X1 U18615 ( .B1(n15222), .B2(P1_REIP_REG_13__SCAN_IN), .A(n15208), 
        .ZN(n15209) );
  OAI21_X1 U18616 ( .B1(n20637), .B2(n15606), .A(n15209), .ZN(n15210) );
  AOI211_X1 U18617 ( .C1(n15213), .C2(n15212), .A(n15211), .B(n15210), .ZN(
        n15214) );
  OAI21_X1 U18618 ( .B1(n15411), .B2(n15269), .A(n15214), .ZN(P1_U2827) );
  OAI21_X1 U18619 ( .B1(n15217), .B2(n15216), .A(n15215), .ZN(n15614) );
  XNOR2_X1 U18620 ( .A(n15199), .B(n15218), .ZN(n15849) );
  NAND2_X1 U18621 ( .A1(n20608), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15219) );
  NAND2_X1 U18622 ( .A1(n15219), .A2(n20622), .ZN(n15220) );
  AOI21_X1 U18623 ( .B1(n20641), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15220), .ZN(
        n15221) );
  OAI21_X1 U18624 ( .B1(n20637), .B2(n15617), .A(n15221), .ZN(n15226) );
  AOI21_X1 U18625 ( .B1(n9872), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15224) );
  INV_X1 U18626 ( .A(n15222), .ZN(n15223) );
  NOR2_X1 U18627 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  AOI211_X1 U18628 ( .C1(n20627), .C2(n15849), .A(n15226), .B(n15225), .ZN(
        n15227) );
  OAI21_X1 U18629 ( .B1(n15269), .B2(n15614), .A(n15227), .ZN(P1_U2828) );
  XOR2_X1 U18630 ( .A(n15229), .B(n15228), .Z(n15629) );
  INV_X1 U18631 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15240) );
  NOR2_X1 U18632 ( .A1(n20637), .A2(n15627), .ZN(n15239) );
  NAND2_X1 U18633 ( .A1(n15249), .A2(n15230), .ZN(n15231) );
  NAND2_X1 U18634 ( .A1(n15199), .A2(n15231), .ZN(n15856) );
  OAI21_X1 U18635 ( .B1(n20636), .B2(n15232), .A(n20622), .ZN(n15236) );
  INV_X1 U18636 ( .A(n15233), .ZN(n15234) );
  NAND2_X1 U18637 ( .A1(n20585), .A2(n15234), .ZN(n15245) );
  NOR2_X1 U18638 ( .A1(n15245), .A2(n15240), .ZN(n15235) );
  AOI211_X1 U18639 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n20641), .A(n15236), .B(
        n15235), .ZN(n15237) );
  OAI21_X1 U18640 ( .B1(n20648), .B2(n15856), .A(n15237), .ZN(n15238) );
  AOI211_X1 U18641 ( .C1(n9872), .C2(n15240), .A(n15239), .B(n15238), .ZN(
        n15241) );
  OAI21_X1 U18642 ( .B1(n15414), .B2(n15269), .A(n15241), .ZN(P1_U2829) );
  NOR2_X1 U18643 ( .A1(n14725), .A2(n15242), .ZN(n15243) );
  OR2_X1 U18644 ( .A1(n15165), .A2(n15243), .ZN(n15635) );
  INV_X1 U18645 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15244) );
  NOR2_X1 U18646 ( .A1(n15266), .A2(n15244), .ZN(n15247) );
  INV_X1 U18647 ( .A(n15245), .ZN(n15246) );
  MUX2_X1 U18648 ( .A(n15247), .B(n15246), .S(P1_REIP_REG_10__SCAN_IN), .Z(
        n15248) );
  INV_X1 U18649 ( .A(n15248), .ZN(n15256) );
  INV_X1 U18650 ( .A(n15637), .ZN(n15254) );
  OAI21_X1 U18651 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(n15867) );
  INV_X1 U18652 ( .A(n15867), .ZN(n15320) );
  AOI22_X1 U18653 ( .A1(n15320), .A2(n20627), .B1(n20641), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15252) );
  OAI211_X1 U18654 ( .C1(n20636), .C2(n12959), .A(n15252), .B(n20622), .ZN(
        n15253) );
  AOI21_X1 U18655 ( .B1(n15294), .B2(n15254), .A(n15253), .ZN(n15255) );
  OAI211_X1 U18656 ( .C1(n15635), .C2(n15269), .A(n15256), .B(n15255), .ZN(
        P1_U2830) );
  OAI21_X1 U18657 ( .B1(n20636), .B2(n15257), .A(n20622), .ZN(n15258) );
  AOI21_X1 U18658 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n20641), .A(n15258), .ZN(
        n15259) );
  OAI21_X1 U18659 ( .B1(n20648), .B2(n15877), .A(n15259), .ZN(n15261) );
  NOR2_X1 U18660 ( .A1(n20637), .A2(n15643), .ZN(n15260) );
  AOI211_X1 U18661 ( .C1(n15262), .C2(P1_REIP_REG_9__SCAN_IN), .A(n15261), .B(
        n15260), .ZN(n15265) );
  INV_X1 U18662 ( .A(n15263), .ZN(n15645) );
  NAND2_X1 U18663 ( .A1(n15645), .A2(n20601), .ZN(n15264) );
  OAI211_X1 U18664 ( .C1(n15266), .C2(P1_REIP_REG_9__SCAN_IN), .A(n15265), .B(
        n15264), .ZN(P1_U2831) );
  NAND2_X1 U18665 ( .A1(n9871), .A2(n15267), .ZN(n15268) );
  NAND2_X1 U18666 ( .A1(n15269), .A2(n15268), .ZN(n20635) );
  INV_X1 U18667 ( .A(n20635), .ZN(n15298) );
  OAI211_X1 U18668 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n15281), .B(n15270), .ZN(n15279) );
  NAND2_X1 U18669 ( .A1(n9871), .A2(n15271), .ZN(n20639) );
  INV_X1 U18670 ( .A(n20639), .ZN(n15291) );
  OAI21_X1 U18671 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20645), .A(n20638), .ZN(
        n15283) );
  AOI22_X1 U18672 ( .A1(n20608), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n15283), .ZN(n15273) );
  NAND2_X1 U18673 ( .A1(n20641), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n15272) );
  OAI211_X1 U18674 ( .C1(n20648), .C2(n15274), .A(n15273), .B(n15272), .ZN(
        n15277) );
  NOR2_X1 U18675 ( .A1(n20637), .A2(n15275), .ZN(n15276) );
  AOI211_X1 U18676 ( .C1(n15291), .C2(n21031), .A(n15277), .B(n15276), .ZN(
        n15278) );
  OAI211_X1 U18677 ( .C1(n15298), .C2(n15280), .A(n15279), .B(n15278), .ZN(
        P1_U2837) );
  INV_X1 U18678 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21350) );
  NAND2_X1 U18679 ( .A1(n15281), .A2(n21350), .ZN(n15289) );
  INV_X1 U18680 ( .A(n15282), .ZN(n15287) );
  AOI22_X1 U18681 ( .A1(n20747), .A2(n20627), .B1(n20641), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n15285) );
  AOI22_X1 U18682 ( .A1(n20608), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n15283), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n15284) );
  OAI211_X1 U18683 ( .C1(n21152), .C2(n20639), .A(n15285), .B(n15284), .ZN(
        n15286) );
  AOI21_X1 U18684 ( .B1(n15294), .B2(n15287), .A(n15286), .ZN(n15288) );
  OAI211_X1 U18685 ( .C1(n15298), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        P1_U2838) );
  AOI22_X1 U18686 ( .A1(n20641), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n15291), .B2(
        n20882), .ZN(n15292) );
  OAI21_X1 U18687 ( .B1(n20648), .B2(n20773), .A(n15292), .ZN(n15293) );
  AOI21_X1 U18688 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n20585), .A(n15293), .ZN(
        n15296) );
  OAI21_X1 U18689 ( .B1(n15294), .B2(n20608), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15295) );
  OAI211_X1 U18690 ( .C1(n15298), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        P1_U2840) );
  INV_X1 U18691 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15299) );
  OAI22_X1 U18692 ( .A1(n15300), .A2(n15334), .B1(n20655), .B2(n15299), .ZN(
        P1_U2841) );
  INV_X1 U18693 ( .A(n15435), .ZN(n15343) );
  AOI22_X1 U18694 ( .A1(n15683), .A2(n20650), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15319), .ZN(n15301) );
  OAI21_X1 U18695 ( .B1(n15343), .B2(n15336), .A(n15301), .ZN(P1_U2842) );
  INV_X1 U18696 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21673) );
  OAI222_X1 U18697 ( .A1(n15336), .A2(n15349), .B1(n21673), .B2(n20655), .C1(
        n15700), .C2(n15334), .ZN(P1_U2844) );
  AOI22_X1 U18698 ( .A1(n15705), .A2(n20650), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n15319), .ZN(n15302) );
  OAI21_X1 U18699 ( .B1(n15460), .B2(n15336), .A(n15302), .ZN(P1_U2845) );
  AOI22_X1 U18700 ( .A1(n15719), .A2(n20650), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n15319), .ZN(n15303) );
  OAI21_X1 U18701 ( .B1(n15358), .B2(n15336), .A(n15303), .ZN(P1_U2846) );
  INV_X1 U18702 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15304) );
  OAI222_X1 U18703 ( .A1(n15336), .A2(n15477), .B1(n15304), .B2(n20655), .C1(
        n15732), .C2(n15334), .ZN(P1_U2847) );
  INV_X1 U18704 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15305) );
  OAI222_X1 U18705 ( .A1(n15336), .A2(n15366), .B1(n15305), .B2(n20655), .C1(
        n15733), .C2(n15334), .ZN(P1_U2848) );
  OAI222_X1 U18706 ( .A1(n15336), .A2(n15490), .B1(n21540), .B2(n20655), .C1(
        n15744), .C2(n15334), .ZN(P1_U2849) );
  AOI22_X1 U18707 ( .A1(n15758), .A2(n20650), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15319), .ZN(n15306) );
  OAI21_X1 U18708 ( .B1(n15501), .B2(n15336), .A(n15306), .ZN(P1_U2850) );
  OAI222_X1 U18709 ( .A1(n15336), .A2(n15520), .B1(n15308), .B2(n20655), .C1(
        n15769), .C2(n15334), .ZN(P1_U2851) );
  AOI22_X1 U18710 ( .A1(n15773), .A2(n20650), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n15319), .ZN(n15309) );
  OAI21_X1 U18711 ( .B1(n15525), .B2(n15336), .A(n15309), .ZN(P1_U2852) );
  INV_X1 U18712 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15310) );
  OAI222_X1 U18713 ( .A1(n15536), .A2(n15336), .B1(n15310), .B2(n20655), .C1(
        n15781), .C2(n15334), .ZN(P1_U2853) );
  AOI22_X1 U18714 ( .A1(n15791), .A2(n20650), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n15319), .ZN(n15311) );
  OAI21_X1 U18715 ( .B1(n15545), .B2(n15336), .A(n15311), .ZN(P1_U2854) );
  INV_X1 U18716 ( .A(n15800), .ZN(n15312) );
  OAI222_X1 U18717 ( .A1(n15336), .A2(n15395), .B1(n21516), .B2(n20655), .C1(
        n15312), .C2(n15334), .ZN(P1_U2855) );
  INV_X1 U18718 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15313) );
  OAI222_X1 U18719 ( .A1(n15572), .A2(n15336), .B1(n15313), .B2(n20655), .C1(
        n15334), .C2(n15813), .ZN(P1_U2856) );
  AOI22_X1 U18720 ( .A1(n15819), .A2(n20650), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15319), .ZN(n15314) );
  OAI21_X1 U18721 ( .B1(n15406), .B2(n15336), .A(n15314), .ZN(P1_U2857) );
  AOI22_X1 U18722 ( .A1(n15826), .A2(n20650), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15319), .ZN(n15315) );
  OAI21_X1 U18723 ( .B1(n15591), .B2(n15336), .A(n15315), .ZN(P1_U2858) );
  OAI222_X1 U18724 ( .A1(n15411), .A2(n15336), .B1(n15316), .B2(n20655), .C1(
        n15836), .C2(n15334), .ZN(P1_U2859) );
  AOI22_X1 U18725 ( .A1(n15849), .A2(n20650), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n15319), .ZN(n15317) );
  OAI21_X1 U18726 ( .B1(n15614), .B2(n15336), .A(n15317), .ZN(P1_U2860) );
  INV_X1 U18727 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15318) );
  OAI222_X1 U18728 ( .A1(n15414), .A2(n15336), .B1(n15318), .B2(n20655), .C1(
        n15856), .C2(n15334), .ZN(P1_U2861) );
  AOI22_X1 U18729 ( .A1(n15320), .A2(n20650), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n15319), .ZN(n15321) );
  OAI21_X1 U18730 ( .B1(n15635), .B2(n15336), .A(n15321), .ZN(P1_U2862) );
  AND2_X1 U18731 ( .A1(n15330), .A2(n15322), .ZN(n15324) );
  INV_X1 U18732 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15329) );
  OAI21_X1 U18733 ( .B1(n14617), .B2(n15326), .A(n15325), .ZN(n15328) );
  NAND2_X1 U18734 ( .A1(n15328), .A2(n15327), .ZN(n20589) );
  OAI222_X1 U18735 ( .A1(n15661), .A2(n15336), .B1(n15329), .B2(n20655), .C1(
        n20589), .C2(n15334), .ZN(P1_U2865) );
  INV_X1 U18736 ( .A(n15330), .ZN(n15331) );
  AOI21_X1 U18737 ( .B1(n15333), .B2(n15332), .A(n15331), .ZN(n20602) );
  INV_X1 U18738 ( .A(n20602), .ZN(n15422) );
  INV_X1 U18739 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n15335) );
  OAI222_X1 U18740 ( .A1(n15422), .A2(n15336), .B1(n15335), .B2(n20655), .C1(
        n15334), .C2(n20598), .ZN(P1_U2866) );
  INV_X1 U18741 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n15340) );
  INV_X1 U18742 ( .A(DATAI_14_), .ZN(n15338) );
  NAND2_X1 U18743 ( .A1(n15350), .A2(BUF1_REG_14__SCAN_IN), .ZN(n15337) );
  OAI21_X1 U18744 ( .B1(n15350), .B2(n15338), .A(n15337), .ZN(n20697) );
  AOI22_X1 U18745 ( .A1(n15397), .A2(n20697), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15407), .ZN(n15339) );
  OAI21_X1 U18746 ( .B1(n15340), .B2(n15399), .A(n15339), .ZN(n15341) );
  AOI21_X1 U18747 ( .B1(n15401), .B2(DATAI_30_), .A(n15341), .ZN(n15342) );
  OAI21_X1 U18748 ( .B1(n15343), .B2(n15421), .A(n15342), .ZN(P1_U2874) );
  NAND2_X1 U18749 ( .A1(n15405), .A2(DATAI_12_), .ZN(n15345) );
  NAND2_X1 U18750 ( .A1(n15350), .A2(BUF1_REG_12__SCAN_IN), .ZN(n15344) );
  AND2_X1 U18751 ( .A1(n15345), .A2(n15344), .ZN(n20691) );
  OAI22_X1 U18752 ( .A1(n15390), .A2(n20691), .B1(n15418), .B2(n14326), .ZN(
        n15346) );
  AOI21_X1 U18753 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n15392), .A(n15346), .ZN(
        n15348) );
  NAND2_X1 U18754 ( .A1(n15401), .A2(DATAI_28_), .ZN(n15347) );
  OAI211_X1 U18755 ( .C1(n15349), .C2(n15421), .A(n15348), .B(n15347), .ZN(
        P1_U2876) );
  INV_X1 U18756 ( .A(DATAI_11_), .ZN(n15351) );
  INV_X1 U18757 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n17305) );
  MUX2_X1 U18758 ( .A(n15351), .B(n17305), .S(n15350), .Z(n20688) );
  OAI22_X1 U18759 ( .A1(n15390), .A2(n20688), .B1(n15418), .B2(n14312), .ZN(
        n15352) );
  AOI21_X1 U18760 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n15392), .A(n15352), .ZN(
        n15354) );
  NAND2_X1 U18761 ( .A1(n15401), .A2(DATAI_27_), .ZN(n15353) );
  OAI211_X1 U18762 ( .C1(n15460), .C2(n15421), .A(n15354), .B(n15353), .ZN(
        P1_U2877) );
  OAI22_X1 U18763 ( .A1(n15390), .A2(n15415), .B1(n15418), .B2(n14323), .ZN(
        n15355) );
  AOI21_X1 U18764 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n15392), .A(n15355), .ZN(
        n15357) );
  NAND2_X1 U18765 ( .A1(n15401), .A2(DATAI_26_), .ZN(n15356) );
  OAI211_X1 U18766 ( .C1(n15358), .C2(n15421), .A(n15357), .B(n15356), .ZN(
        P1_U2878) );
  INV_X1 U18767 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n15360) );
  AOI22_X1 U18768 ( .A1(n15397), .A2(n15423), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n15407), .ZN(n15359) );
  OAI21_X1 U18769 ( .B1(n15399), .B2(n15360), .A(n15359), .ZN(n15361) );
  AOI21_X1 U18770 ( .B1(n15401), .B2(DATAI_25_), .A(n15361), .ZN(n15362) );
  OAI21_X1 U18771 ( .B1(n15477), .B2(n15421), .A(n15362), .ZN(P1_U2879) );
  INV_X1 U18772 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U18773 ( .A1(n15397), .A2(n15416), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15407), .ZN(n15363) );
  OAI21_X1 U18774 ( .B1(n15399), .B2(n17284), .A(n15363), .ZN(n15364) );
  AOI21_X1 U18775 ( .B1(n15401), .B2(DATAI_24_), .A(n15364), .ZN(n15365) );
  OAI21_X1 U18776 ( .B1(n15366), .B2(n15421), .A(n15365), .ZN(P1_U2880) );
  OAI22_X1 U18777 ( .A1(n15390), .A2(n20825), .B1(n15418), .B2(n14308), .ZN(
        n15367) );
  AOI21_X1 U18778 ( .B1(n15392), .B2(BUF1_REG_23__SCAN_IN), .A(n15367), .ZN(
        n15369) );
  NAND2_X1 U18779 ( .A1(n15401), .A2(DATAI_23_), .ZN(n15368) );
  OAI211_X1 U18780 ( .C1(n15490), .C2(n15421), .A(n15369), .B(n15368), .ZN(
        P1_U2881) );
  OAI22_X1 U18781 ( .A1(n15390), .A2(n15420), .B1(n15418), .B2(n15370), .ZN(
        n15371) );
  AOI21_X1 U18782 ( .B1(n15392), .B2(BUF1_REG_22__SCAN_IN), .A(n15371), .ZN(
        n15373) );
  NAND2_X1 U18783 ( .A1(n15401), .A2(DATAI_22_), .ZN(n15372) );
  OAI211_X1 U18784 ( .C1(n15501), .C2(n15421), .A(n15373), .B(n15372), .ZN(
        P1_U2882) );
  INV_X1 U18785 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U18786 ( .A1(n15397), .A2(n20816), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15407), .ZN(n15374) );
  OAI21_X1 U18787 ( .B1(n15399), .B2(n17289), .A(n15374), .ZN(n15375) );
  AOI21_X1 U18788 ( .B1(n15401), .B2(DATAI_21_), .A(n15375), .ZN(n15376) );
  OAI21_X1 U18789 ( .B1(n15520), .B2(n15421), .A(n15376), .ZN(P1_U2883) );
  OAI22_X1 U18790 ( .A1(n15390), .A2(n15377), .B1(n15418), .B2(n14314), .ZN(
        n15378) );
  AOI21_X1 U18791 ( .B1(n15392), .B2(BUF1_REG_20__SCAN_IN), .A(n15378), .ZN(
        n15380) );
  NAND2_X1 U18792 ( .A1(n15401), .A2(DATAI_20_), .ZN(n15379) );
  OAI211_X1 U18793 ( .C1(n15525), .C2(n15421), .A(n15380), .B(n15379), .ZN(
        P1_U2884) );
  OAI22_X1 U18794 ( .A1(n15390), .A2(n15382), .B1(n15418), .B2(n15381), .ZN(
        n15383) );
  AOI21_X1 U18795 ( .B1(n15392), .B2(BUF1_REG_19__SCAN_IN), .A(n15383), .ZN(
        n15385) );
  NAND2_X1 U18796 ( .A1(n15401), .A2(DATAI_19_), .ZN(n15384) );
  OAI211_X1 U18797 ( .C1(n15536), .C2(n15421), .A(n15385), .B(n15384), .ZN(
        P1_U2885) );
  INV_X1 U18798 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21578) );
  AOI22_X1 U18799 ( .A1(n15397), .A2(n20803), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15407), .ZN(n15386) );
  OAI21_X1 U18800 ( .B1(n15399), .B2(n21578), .A(n15386), .ZN(n15387) );
  AOI21_X1 U18801 ( .B1(n15401), .B2(DATAI_18_), .A(n15387), .ZN(n15388) );
  OAI21_X1 U18802 ( .B1(n15545), .B2(n15421), .A(n15388), .ZN(P1_U2886) );
  OAI22_X1 U18803 ( .A1(n15390), .A2(n15389), .B1(n15418), .B2(n14320), .ZN(
        n15391) );
  AOI21_X1 U18804 ( .B1(n15392), .B2(BUF1_REG_17__SCAN_IN), .A(n15391), .ZN(
        n15394) );
  NAND2_X1 U18805 ( .A1(n15401), .A2(DATAI_17_), .ZN(n15393) );
  OAI211_X1 U18806 ( .C1(n15395), .C2(n15421), .A(n15394), .B(n15393), .ZN(
        P1_U2887) );
  AOI22_X1 U18807 ( .A1(n15397), .A2(n15396), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15407), .ZN(n15398) );
  OAI21_X1 U18808 ( .B1(n15399), .B2(n19865), .A(n15398), .ZN(n15400) );
  AOI21_X1 U18809 ( .B1(n15401), .B2(DATAI_16_), .A(n15400), .ZN(n15402) );
  OAI21_X1 U18810 ( .B1(n15572), .B2(n15421), .A(n15402), .ZN(P1_U2888) );
  NOR2_X1 U18811 ( .A1(n15405), .A2(n15403), .ZN(n15404) );
  AOI21_X1 U18812 ( .B1(DATAI_15_), .B2(n15405), .A(n15404), .ZN(n15427) );
  INV_X1 U18813 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20656) );
  OAI222_X1 U18814 ( .A1(n15421), .A2(n15406), .B1(n15419), .B2(n15427), .C1(
        n20656), .C2(n15418), .ZN(P1_U2889) );
  AOI22_X1 U18815 ( .A1(n15408), .A2(n20697), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15407), .ZN(n15409) );
  OAI21_X1 U18816 ( .B1(n15591), .B2(n15421), .A(n15409), .ZN(P1_U2890) );
  INV_X1 U18817 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15410) );
  OAI222_X1 U18818 ( .A1(n15421), .A2(n15411), .B1(n20694), .B2(n15419), .C1(
        n15410), .C2(n15418), .ZN(P1_U2891) );
  INV_X1 U18819 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15412) );
  OAI222_X1 U18820 ( .A1(n15614), .A2(n15421), .B1(n20691), .B2(n15419), .C1(
        n15412), .C2(n15418), .ZN(P1_U2892) );
  INV_X1 U18821 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15413) );
  OAI222_X1 U18822 ( .A1(n15421), .A2(n15414), .B1(n20688), .B2(n15419), .C1(
        n15413), .C2(n15418), .ZN(P1_U2893) );
  INV_X1 U18823 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n21726) );
  OAI222_X1 U18824 ( .A1(n15635), .A2(n15421), .B1(n15418), .B2(n21726), .C1(
        n15415), .C2(n15419), .ZN(P1_U2894) );
  INV_X1 U18825 ( .A(n15416), .ZN(n15417) );
  INV_X1 U18826 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21625) );
  OAI222_X1 U18827 ( .A1(n15421), .A2(n15650), .B1(n15417), .B2(n15419), .C1(
        n15418), .C2(n21625), .ZN(P1_U2896) );
  INV_X1 U18828 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20668) );
  OAI222_X1 U18829 ( .A1(n15421), .A2(n15661), .B1(n20825), .B2(n15419), .C1(
        n15418), .C2(n20668), .ZN(P1_U2897) );
  INV_X1 U18830 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20670) );
  OAI222_X1 U18831 ( .A1(n15422), .A2(n15421), .B1(n15420), .B2(n15419), .C1(
        n20670), .C2(n15418), .ZN(P1_U2898) );
  NAND2_X1 U18832 ( .A1(n20698), .A2(n15423), .ZN(n15426) );
  NAND2_X1 U18833 ( .A1(n20706), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n15424) );
  OAI211_X1 U18834 ( .C1(n21622), .C2(n15430), .A(n15426), .B(n15424), .ZN(
        P1_U2946) );
  INV_X1 U18835 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20665) );
  NAND2_X1 U18836 ( .A1(n20706), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n15425) );
  OAI211_X1 U18837 ( .C1(n20665), .C2(n15430), .A(n15426), .B(n15425), .ZN(
        P1_U2961) );
  INV_X1 U18838 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20657) );
  INV_X1 U18839 ( .A(n20698), .ZN(n15428) );
  OAI222_X1 U18840 ( .A1(n15430), .A2(n20656), .B1(n15429), .B2(n20657), .C1(
        n15428), .C2(n15427), .ZN(P1_U2967) );
  NOR2_X1 U18841 ( .A1(n20781), .A2(n15431), .ZN(n15682) );
  AOI21_X1 U18842 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15682), .ZN(n15432) );
  OAI21_X1 U18843 ( .B1(n15433), .B2(n20720), .A(n15432), .ZN(n15434) );
  AOI21_X1 U18844 ( .B1(n15435), .B2(n20715), .A(n15434), .ZN(n15436) );
  OAI21_X1 U18845 ( .B1(n15685), .B2(n15671), .A(n15436), .ZN(P1_U2969) );
  NAND2_X1 U18846 ( .A1(n9689), .A2(n15716), .ZN(n15461) );
  NAND2_X1 U18847 ( .A1(n15438), .A2(n15461), .ZN(n15443) );
  OAI21_X1 U18848 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15439), .A(
        n15443), .ZN(n15442) );
  INV_X1 U18849 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15440) );
  MUX2_X1 U18850 ( .A(n15440), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9689), .Z(n15441) );
  OAI211_X1 U18851 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15443), .A(
        n15442), .B(n15441), .ZN(n15445) );
  XNOR2_X1 U18852 ( .A(n15445), .B(n15444), .ZN(n15704) );
  NOR2_X1 U18853 ( .A1(n20781), .A2(n15446), .ZN(n15699) );
  AOI21_X1 U18854 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15699), .ZN(n15447) );
  OAI21_X1 U18855 ( .B1(n15448), .B2(n20720), .A(n15447), .ZN(n15449) );
  AOI21_X1 U18856 ( .B1(n15450), .B2(n20715), .A(n15449), .ZN(n15451) );
  OAI21_X1 U18857 ( .B1(n15671), .B2(n15704), .A(n15451), .ZN(P1_U2971) );
  NOR2_X1 U18858 ( .A1(n20781), .A2(n15452), .ZN(n15709) );
  NOR2_X1 U18859 ( .A1(n15673), .A2(n21419), .ZN(n15453) );
  AOI211_X1 U18860 ( .C1(n15454), .C2(n15517), .A(n15709), .B(n15453), .ZN(
        n15459) );
  XNOR2_X1 U18861 ( .A(n15457), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15706) );
  NAND2_X1 U18862 ( .A1(n15706), .A2(n20716), .ZN(n15458) );
  OAI211_X1 U18863 ( .C1(n15460), .C2(n15573), .A(n15459), .B(n15458), .ZN(
        P1_U2972) );
  OAI211_X1 U18864 ( .C1(n15621), .C2(n15438), .A(n15462), .B(n15461), .ZN(
        n15463) );
  XOR2_X1 U18865 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15463), .Z(
        n15722) );
  NAND2_X1 U18866 ( .A1(n20727), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15715) );
  NAND2_X1 U18867 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15464) );
  OAI211_X1 U18868 ( .C1(n15465), .C2(n20720), .A(n15715), .B(n15464), .ZN(
        n15466) );
  AOI21_X1 U18869 ( .B1(n15467), .B2(n20715), .A(n15466), .ZN(n15468) );
  OAI21_X1 U18870 ( .B1(n15671), .B2(n15722), .A(n15468), .ZN(P1_U2973) );
  INV_X1 U18871 ( .A(n15438), .ZN(n15469) );
  NAND3_X1 U18872 ( .A1(n15469), .A2(n15748), .A3(n15738), .ZN(n15472) );
  NAND2_X1 U18873 ( .A1(n15481), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15471) );
  MUX2_X1 U18874 ( .A(n15472), .B(n15471), .S(n9689), .Z(n15473) );
  XNOR2_X1 U18875 ( .A(n15473), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15723) );
  NOR2_X1 U18876 ( .A1(n20781), .A2(n21659), .ZN(n15727) );
  AOI21_X1 U18877 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15727), .ZN(n15476) );
  NAND2_X1 U18878 ( .A1(n15517), .A2(n15474), .ZN(n15475) );
  OAI211_X1 U18879 ( .C1(n15477), .C2(n15573), .A(n15476), .B(n15475), .ZN(
        n15478) );
  AOI21_X1 U18880 ( .B1(n20716), .B2(n15723), .A(n15478), .ZN(n15479) );
  INV_X1 U18881 ( .A(n15479), .ZN(P1_U2974) );
  NOR2_X1 U18882 ( .A1(n15481), .A2(n15438), .ZN(n15480) );
  MUX2_X1 U18883 ( .A(n15481), .B(n15480), .S(n15621), .Z(n15482) );
  XNOR2_X1 U18884 ( .A(n15482), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15743) );
  NAND2_X1 U18885 ( .A1(n20727), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15737) );
  INV_X1 U18886 ( .A(n15737), .ZN(n15483) );
  AOI21_X1 U18887 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15483), .ZN(n15484) );
  OAI21_X1 U18888 ( .B1(n20720), .B2(n15485), .A(n15484), .ZN(n15486) );
  AOI21_X1 U18889 ( .B1(n15487), .B2(n20715), .A(n15486), .ZN(n15488) );
  OAI21_X1 U18890 ( .B1(n15671), .B2(n15743), .A(n15488), .ZN(P1_U2975) );
  XNOR2_X1 U18891 ( .A(n9689), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15489) );
  XNOR2_X1 U18892 ( .A(n15438), .B(n15489), .ZN(n15753) );
  INV_X1 U18893 ( .A(n15490), .ZN(n15495) );
  INV_X1 U18894 ( .A(n15491), .ZN(n15493) );
  NOR2_X1 U18895 ( .A1(n20781), .A2(n21373), .ZN(n15745) );
  AOI21_X1 U18896 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15745), .ZN(n15492) );
  OAI21_X1 U18897 ( .B1(n20720), .B2(n15493), .A(n15492), .ZN(n15494) );
  AOI21_X1 U18898 ( .B1(n15495), .B2(n20715), .A(n15494), .ZN(n15496) );
  OAI21_X1 U18899 ( .B1(n15753), .B2(n15671), .A(n15496), .ZN(P1_U2976) );
  NAND2_X1 U18900 ( .A1(n15498), .A2(n15497), .ZN(n15500) );
  XNOR2_X1 U18901 ( .A(n15500), .B(n15499), .ZN(n15761) );
  INV_X1 U18902 ( .A(n15501), .ZN(n15505) );
  NOR2_X1 U18903 ( .A1(n20781), .A2(n21374), .ZN(n15757) );
  AOI21_X1 U18904 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15757), .ZN(n15502) );
  OAI21_X1 U18905 ( .B1(n20720), .B2(n15503), .A(n15502), .ZN(n15504) );
  AOI21_X1 U18906 ( .B1(n15505), .B2(n20715), .A(n15504), .ZN(n15506) );
  OAI21_X1 U18907 ( .B1(n15671), .B2(n15761), .A(n15506), .ZN(P1_U2977) );
  OAI21_X1 U18908 ( .B1(n9689), .B2(n13895), .A(n15507), .ZN(n15535) );
  NAND2_X1 U18909 ( .A1(n15621), .A2(n15508), .ZN(n15533) );
  NAND2_X1 U18910 ( .A1(n9689), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15532) );
  NAND2_X1 U18911 ( .A1(n15521), .A2(n15509), .ZN(n15522) );
  INV_X1 U18912 ( .A(n15532), .ZN(n15510) );
  NAND2_X1 U18913 ( .A1(n15510), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15511) );
  OAI22_X1 U18914 ( .A1(n15522), .A2(n9689), .B1(n15507), .B2(n15511), .ZN(
        n15512) );
  XOR2_X1 U18915 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15512), .Z(
        n15762) );
  NAND2_X1 U18916 ( .A1(n15762), .A2(n20716), .ZN(n15519) );
  NOR2_X1 U18917 ( .A1(n20781), .A2(n15513), .ZN(n15765) );
  NOR2_X1 U18918 ( .A1(n15673), .A2(n15514), .ZN(n15515) );
  AOI211_X1 U18919 ( .C1(n15517), .C2(n15516), .A(n15765), .B(n15515), .ZN(
        n15518) );
  OAI211_X1 U18920 ( .C1(n15573), .C2(n15520), .A(n15519), .B(n15518), .ZN(
        P1_U2978) );
  INV_X1 U18921 ( .A(n15521), .ZN(n15524) );
  INV_X1 U18922 ( .A(n15522), .ZN(n15523) );
  AOI21_X1 U18923 ( .B1(n15524), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15523), .ZN(n15776) );
  INV_X1 U18924 ( .A(n15525), .ZN(n15530) );
  NOR2_X1 U18925 ( .A1(n20781), .A2(n15526), .ZN(n15772) );
  AOI21_X1 U18926 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15772), .ZN(n15527) );
  OAI21_X1 U18927 ( .B1(n20720), .B2(n15528), .A(n15527), .ZN(n15529) );
  AOI21_X1 U18928 ( .B1(n15530), .B2(n20715), .A(n15529), .ZN(n15531) );
  OAI21_X1 U18929 ( .B1(n15776), .B2(n15671), .A(n15531), .ZN(P1_U2979) );
  NAND2_X1 U18930 ( .A1(n15533), .A2(n15532), .ZN(n15534) );
  XNOR2_X1 U18931 ( .A(n15535), .B(n15534), .ZN(n15785) );
  INV_X1 U18932 ( .A(n15536), .ZN(n15541) );
  INV_X1 U18933 ( .A(n15537), .ZN(n15539) );
  NOR2_X1 U18934 ( .A1(n20781), .A2(n21571), .ZN(n15779) );
  AOI21_X1 U18935 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15779), .ZN(n15538) );
  OAI21_X1 U18936 ( .B1(n20720), .B2(n15539), .A(n15538), .ZN(n15540) );
  AOI21_X1 U18937 ( .B1(n15541), .B2(n20715), .A(n15540), .ZN(n15542) );
  OAI21_X1 U18938 ( .B1(n15671), .B2(n15785), .A(n15542), .ZN(P1_U2980) );
  OAI21_X1 U18939 ( .B1(n15544), .B2(n15543), .A(n15507), .ZN(n15794) );
  INV_X1 U18940 ( .A(n15545), .ZN(n15549) );
  INV_X1 U18941 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21369) );
  NOR2_X1 U18942 ( .A1(n20781), .A2(n21369), .ZN(n15789) );
  AOI21_X1 U18943 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15789), .ZN(n15546) );
  OAI21_X1 U18944 ( .B1(n20720), .B2(n15547), .A(n15546), .ZN(n15548) );
  AOI21_X1 U18945 ( .B1(n15549), .B2(n20715), .A(n15548), .ZN(n15550) );
  OAI21_X1 U18946 ( .B1(n15671), .B2(n15794), .A(n15550), .ZN(P1_U2981) );
  INV_X1 U18947 ( .A(n15551), .ZN(n15553) );
  NAND2_X1 U18948 ( .A1(n15553), .A2(n15552), .ZN(n15632) );
  OAI21_X1 U18949 ( .B1(n15621), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15632), .ZN(n15631) );
  NAND2_X1 U18950 ( .A1(n15631), .A2(n15563), .ZN(n15588) );
  OAI21_X1 U18951 ( .B1(n15588), .B2(n15565), .A(n15554), .ZN(n15556) );
  NAND2_X1 U18952 ( .A1(n15556), .A2(n15806), .ZN(n15555) );
  MUX2_X1 U18953 ( .A(n15556), .B(n15555), .S(n15621), .Z(n15557) );
  XOR2_X1 U18954 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15557), .Z(
        n15802) );
  NAND2_X1 U18955 ( .A1(n20727), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15796) );
  NAND2_X1 U18956 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15558) );
  OAI211_X1 U18957 ( .C1(n20720), .C2(n15559), .A(n15796), .B(n15558), .ZN(
        n15560) );
  AOI21_X1 U18958 ( .B1(n15561), .B2(n20715), .A(n15560), .ZN(n15562) );
  OAI21_X1 U18959 ( .B1(n15802), .B2(n15671), .A(n15562), .ZN(P1_U2982) );
  OAI21_X1 U18960 ( .B1(n15631), .B2(n15564), .A(n15563), .ZN(n15575) );
  OAI21_X1 U18961 ( .B1(n15575), .B2(n15565), .A(n15576), .ZN(n15567) );
  XNOR2_X1 U18962 ( .A(n15567), .B(n15566), .ZN(n15803) );
  NAND2_X1 U18963 ( .A1(n15803), .A2(n20716), .ZN(n15571) );
  NOR2_X1 U18964 ( .A1(n20781), .A2(n21367), .ZN(n15808) );
  NOR2_X1 U18965 ( .A1(n20720), .A2(n15568), .ZN(n15569) );
  AOI211_X1 U18966 ( .C1(n20709), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15808), .B(n15569), .ZN(n15570) );
  OAI211_X1 U18967 ( .C1(n15573), .C2(n15572), .A(n15571), .B(n15570), .ZN(
        P1_U2983) );
  NOR2_X1 U18968 ( .A1(n15575), .A2(n10055), .ZN(n15579) );
  NAND2_X1 U18969 ( .A1(n15577), .A2(n15576), .ZN(n15578) );
  XNOR2_X1 U18970 ( .A(n15579), .B(n15578), .ZN(n15821) );
  NAND2_X1 U18971 ( .A1(n20727), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15814) );
  NAND2_X1 U18972 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15580) );
  OAI211_X1 U18973 ( .C1(n20720), .C2(n15581), .A(n15814), .B(n15580), .ZN(
        n15582) );
  AOI21_X1 U18974 ( .B1(n15583), .B2(n20715), .A(n15582), .ZN(n15584) );
  OAI21_X1 U18975 ( .B1(n15821), .B2(n15671), .A(n15584), .ZN(P1_U2984) );
  INV_X1 U18976 ( .A(n15585), .ZN(n15586) );
  AOI21_X1 U18977 ( .B1(n15588), .B2(n15587), .A(n15586), .ZN(n15590) );
  XNOR2_X1 U18978 ( .A(n9689), .B(n21709), .ZN(n15589) );
  XNOR2_X1 U18979 ( .A(n15590), .B(n15589), .ZN(n15831) );
  INV_X1 U18980 ( .A(n15591), .ZN(n15596) );
  INV_X1 U18981 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15592) );
  NOR2_X1 U18982 ( .A1(n20781), .A2(n15592), .ZN(n15825) );
  AOI21_X1 U18983 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15825), .ZN(n15593) );
  OAI21_X1 U18984 ( .B1(n20720), .B2(n15594), .A(n15593), .ZN(n15595) );
  AOI21_X1 U18985 ( .B1(n15596), .B2(n20715), .A(n15595), .ZN(n15597) );
  OAI21_X1 U18986 ( .B1(n15831), .B2(n15671), .A(n15597), .ZN(P1_U2985) );
  INV_X1 U18987 ( .A(n15631), .ZN(n15622) );
  INV_X1 U18988 ( .A(n15598), .ZN(n15599) );
  AOI21_X1 U18989 ( .B1(n15622), .B2(n15600), .A(n15599), .ZN(n15612) );
  AND2_X1 U18990 ( .A1(n15602), .A2(n15601), .ZN(n15611) );
  NAND2_X1 U18991 ( .A1(n15612), .A2(n15611), .ZN(n15610) );
  NAND2_X1 U18992 ( .A1(n15610), .A2(n15601), .ZN(n15603) );
  XNOR2_X1 U18993 ( .A(n15604), .B(n15603), .ZN(n15841) );
  NAND2_X1 U18994 ( .A1(n20727), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15834) );
  NAND2_X1 U18995 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15605) );
  OAI211_X1 U18996 ( .C1(n20720), .C2(n15606), .A(n15834), .B(n15605), .ZN(
        n15607) );
  AOI21_X1 U18997 ( .B1(n15608), .B2(n20715), .A(n15607), .ZN(n15609) );
  OAI21_X1 U18998 ( .B1(n15841), .B2(n15671), .A(n15609), .ZN(P1_U2986) );
  OAI21_X1 U18999 ( .B1(n15612), .B2(n15611), .A(n15610), .ZN(n15613) );
  INV_X1 U19000 ( .A(n15613), .ZN(n15854) );
  INV_X1 U19001 ( .A(n15614), .ZN(n15619) );
  INV_X1 U19002 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15615) );
  NOR2_X1 U19003 ( .A1(n20781), .A2(n15615), .ZN(n15848) );
  AOI21_X1 U19004 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15848), .ZN(n15616) );
  OAI21_X1 U19005 ( .B1(n20720), .B2(n15617), .A(n15616), .ZN(n15618) );
  AOI21_X1 U19006 ( .B1(n15619), .B2(n20715), .A(n15618), .ZN(n15620) );
  OAI21_X1 U19007 ( .B1(n15854), .B2(n15671), .A(n15620), .ZN(P1_U2987) );
  NAND2_X1 U19008 ( .A1(n15621), .A2(n15633), .ZN(n15624) );
  NAND3_X1 U19009 ( .A1(n15622), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9689), .ZN(n15623) );
  OAI21_X1 U19010 ( .B1(n15632), .B2(n15624), .A(n15623), .ZN(n15625) );
  XNOR2_X1 U19011 ( .A(n15625), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15862) );
  NAND2_X1 U19012 ( .A1(n20727), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15855) );
  NAND2_X1 U19013 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15626) );
  OAI211_X1 U19014 ( .C1(n20720), .C2(n15627), .A(n15855), .B(n15626), .ZN(
        n15628) );
  AOI21_X1 U19015 ( .B1(n15629), .B2(n20715), .A(n15628), .ZN(n15630) );
  OAI21_X1 U19016 ( .B1(n15862), .B2(n15671), .A(n15630), .ZN(P1_U2988) );
  MUX2_X1 U19017 ( .A(n15632), .B(n15631), .S(n9689), .Z(n15634) );
  XNOR2_X1 U19018 ( .A(n15634), .B(n15633), .ZN(n15873) );
  INV_X1 U19019 ( .A(n15635), .ZN(n15639) );
  NAND2_X1 U19020 ( .A1(n20727), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15866) );
  NAND2_X1 U19021 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15636) );
  OAI211_X1 U19022 ( .C1(n20720), .C2(n15637), .A(n15866), .B(n15636), .ZN(
        n15638) );
  AOI21_X1 U19023 ( .B1(n15639), .B2(n20715), .A(n15638), .ZN(n15640) );
  OAI21_X1 U19024 ( .B1(n15873), .B2(n15671), .A(n15640), .ZN(P1_U2989) );
  XNOR2_X1 U19025 ( .A(n9689), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15641) );
  XNOR2_X1 U19026 ( .A(n15551), .B(n15641), .ZN(n15882) );
  NAND2_X1 U19027 ( .A1(n20727), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15875) );
  NAND2_X1 U19028 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15642) );
  OAI211_X1 U19029 ( .C1(n20720), .C2(n15643), .A(n15875), .B(n15642), .ZN(
        n15644) );
  AOI21_X1 U19030 ( .B1(n15645), .B2(n20715), .A(n15644), .ZN(n15646) );
  OAI21_X1 U19031 ( .B1(n15882), .B2(n15671), .A(n15646), .ZN(P1_U2990) );
  XNOR2_X1 U19032 ( .A(n15647), .B(n15884), .ZN(n15648) );
  XNOR2_X1 U19033 ( .A(n15649), .B(n15648), .ZN(n15898) );
  INV_X1 U19034 ( .A(n15650), .ZN(n15655) );
  INV_X1 U19035 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15651) );
  NOR2_X1 U19036 ( .A1(n20781), .A2(n15651), .ZN(n15887) );
  AOI21_X1 U19037 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15887), .ZN(n15652) );
  OAI21_X1 U19038 ( .B1(n20720), .B2(n15653), .A(n15652), .ZN(n15654) );
  AOI21_X1 U19039 ( .B1(n15655), .B2(n20715), .A(n15654), .ZN(n15656) );
  OAI21_X1 U19040 ( .B1(n15671), .B2(n15898), .A(n15656), .ZN(P1_U2991) );
  NAND2_X1 U19041 ( .A1(n15658), .A2(n15657), .ZN(n15660) );
  XOR2_X1 U19042 ( .A(n15660), .B(n15659), .Z(n15906) );
  INV_X1 U19043 ( .A(n15661), .ZN(n20592) );
  INV_X1 U19044 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n15662) );
  NOR2_X1 U19045 ( .A1(n20781), .A2(n15662), .ZN(n15899) );
  AOI21_X1 U19046 ( .B1(n20709), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n15899), .ZN(n15663) );
  OAI21_X1 U19047 ( .B1(n20720), .B2(n20586), .A(n15663), .ZN(n15664) );
  AOI21_X1 U19048 ( .B1(n20592), .B2(n20715), .A(n15664), .ZN(n15665) );
  OAI21_X1 U19049 ( .B1(n15906), .B2(n15671), .A(n15665), .ZN(P1_U2992) );
  NAND2_X1 U19050 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15666) );
  OAI211_X1 U19051 ( .C1(n20720), .C2(n20595), .A(n15667), .B(n15666), .ZN(
        n15668) );
  AOI21_X1 U19052 ( .B1(n20602), .B2(n20715), .A(n15668), .ZN(n15669) );
  OAI21_X1 U19053 ( .B1(n15671), .B2(n15670), .A(n15669), .ZN(P1_U2993) );
  NAND2_X1 U19054 ( .A1(n20634), .A2(n20715), .ZN(n15676) );
  OR2_X1 U19055 ( .A1(n15672), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20759) );
  NAND3_X1 U19056 ( .A1(n20759), .A2(n20758), .A3(n20716), .ZN(n15675) );
  NAND2_X1 U19057 ( .A1(n20727), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20762) );
  MUX2_X1 U19058 ( .A(n20720), .B(n15673), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15674) );
  NAND4_X1 U19059 ( .A1(n15676), .A2(n15675), .A3(n20762), .A4(n15674), .ZN(
        P1_U2998) );
  INV_X1 U19060 ( .A(n15677), .ZN(n15678) );
  AOI21_X1 U19061 ( .B1(n15680), .B2(n15679), .A(n15678), .ZN(n15681) );
  AOI211_X1 U19062 ( .C1(n15683), .C2(n20736), .A(n15682), .B(n15681), .ZN(
        n15684) );
  INV_X1 U19063 ( .A(n15686), .ZN(n15693) );
  NAND3_X1 U19064 ( .A1(n15687), .A2(n15696), .A3(n15690), .ZN(n15688) );
  OAI211_X1 U19065 ( .C1(n15691), .C2(n15690), .A(n15689), .B(n15688), .ZN(
        n15692) );
  AOI21_X1 U19066 ( .B1(n15693), .B2(n20736), .A(n15692), .ZN(n15694) );
  OAI21_X1 U19067 ( .B1(n15695), .B2(n20775), .A(n15694), .ZN(P1_U3002) );
  NOR3_X1 U19068 ( .A1(n15707), .A2(n15697), .A3(n15696), .ZN(n15698) );
  AOI211_X1 U19069 ( .C1(n15710), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15699), .B(n15698), .ZN(n15703) );
  INV_X1 U19070 ( .A(n15700), .ZN(n15701) );
  NAND2_X1 U19071 ( .A1(n15701), .A2(n20736), .ZN(n15702) );
  OAI211_X1 U19072 ( .C1(n15704), .C2(n20775), .A(n15703), .B(n15702), .ZN(
        P1_U3003) );
  INV_X1 U19073 ( .A(n15705), .ZN(n15713) );
  NAND2_X1 U19074 ( .A1(n15706), .A2(n20757), .ZN(n15712) );
  NOR2_X1 U19075 ( .A1(n15707), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15708) );
  AOI211_X1 U19076 ( .C1(n15710), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15709), .B(n15708), .ZN(n15711) );
  OAI211_X1 U19077 ( .C1(n20774), .C2(n15713), .A(n15712), .B(n15711), .ZN(
        P1_U3004) );
  INV_X1 U19078 ( .A(n15714), .ZN(n15729) );
  INV_X1 U19079 ( .A(n15715), .ZN(n15718) );
  NOR3_X1 U19080 ( .A1(n15735), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15716), .ZN(n15717) );
  AOI211_X1 U19081 ( .C1(n15729), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15718), .B(n15717), .ZN(n15721) );
  NAND2_X1 U19082 ( .A1(n15719), .A2(n20736), .ZN(n15720) );
  OAI211_X1 U19083 ( .C1(n15722), .C2(n20775), .A(n15721), .B(n15720), .ZN(
        P1_U3005) );
  NAND2_X1 U19084 ( .A1(n15723), .A2(n20757), .ZN(n15731) );
  INV_X1 U19085 ( .A(n15724), .ZN(n15726) );
  OAI21_X1 U19086 ( .B1(n15735), .B2(n15726), .A(n15725), .ZN(n15728) );
  AOI21_X1 U19087 ( .B1(n15729), .B2(n15728), .A(n15727), .ZN(n15730) );
  OAI211_X1 U19088 ( .C1(n20774), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        P1_U3006) );
  INV_X1 U19089 ( .A(n15733), .ZN(n15741) );
  AOI21_X1 U19090 ( .B1(n15845), .B2(n15748), .A(n15734), .ZN(n15739) );
  INV_X1 U19091 ( .A(n15735), .ZN(n15746) );
  NAND3_X1 U19092 ( .A1(n15746), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15738), .ZN(n15736) );
  OAI211_X1 U19093 ( .C1(n15739), .C2(n15738), .A(n15737), .B(n15736), .ZN(
        n15740) );
  AOI21_X1 U19094 ( .B1(n15741), .B2(n20736), .A(n15740), .ZN(n15742) );
  OAI21_X1 U19095 ( .B1(n15743), .B2(n20775), .A(n15742), .ZN(P1_U3007) );
  INV_X1 U19096 ( .A(n15744), .ZN(n15751) );
  AOI21_X1 U19097 ( .B1(n15746), .B2(n15748), .A(n15745), .ZN(n15747) );
  OAI21_X1 U19098 ( .B1(n15749), .B2(n15748), .A(n15747), .ZN(n15750) );
  AOI21_X1 U19099 ( .B1(n15751), .B2(n20736), .A(n15750), .ZN(n15752) );
  OAI21_X1 U19100 ( .B1(n15753), .B2(n20775), .A(n15752), .ZN(P1_U3008) );
  INV_X1 U19101 ( .A(n15754), .ZN(n15763) );
  XNOR2_X1 U19102 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15755) );
  NOR2_X1 U19103 ( .A1(n15763), .A2(n15755), .ZN(n15756) );
  AOI211_X1 U19104 ( .C1(n15766), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15757), .B(n15756), .ZN(n15760) );
  NAND2_X1 U19105 ( .A1(n15758), .A2(n20736), .ZN(n15759) );
  OAI211_X1 U19106 ( .C1(n15761), .C2(n20775), .A(n15760), .B(n15759), .ZN(
        P1_U3009) );
  NAND2_X1 U19107 ( .A1(n15762), .A2(n20757), .ZN(n15768) );
  NOR2_X1 U19108 ( .A1(n15763), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15764) );
  AOI211_X1 U19109 ( .C1(n15766), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15765), .B(n15764), .ZN(n15767) );
  OAI211_X1 U19110 ( .C1(n20774), .C2(n15769), .A(n15768), .B(n15767), .ZN(
        P1_U3010) );
  AOI21_X1 U19111 ( .B1(n15893), .B2(n15786), .A(n15822), .ZN(n15798) );
  OAI21_X1 U19112 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n20761), .A(
        n15798), .ZN(n15780) );
  NOR3_X1 U19113 ( .A1(n15777), .A2(n10939), .A3(n13894), .ZN(n15771) );
  AOI211_X1 U19114 ( .C1(n15780), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15772), .B(n15771), .ZN(n15775) );
  NAND2_X1 U19115 ( .A1(n15773), .A2(n20736), .ZN(n15774) );
  OAI211_X1 U19116 ( .C1(n15776), .C2(n20775), .A(n15775), .B(n15774), .ZN(
        P1_U3011) );
  NOR2_X1 U19117 ( .A1(n15777), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15778) );
  AOI211_X1 U19118 ( .C1(n15780), .C2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15779), .B(n15778), .ZN(n15784) );
  INV_X1 U19119 ( .A(n15781), .ZN(n15782) );
  NAND2_X1 U19120 ( .A1(n15782), .A2(n20736), .ZN(n15783) );
  OAI211_X1 U19121 ( .C1(n15785), .C2(n20775), .A(n15784), .B(n15783), .ZN(
        P1_U3012) );
  INV_X1 U19122 ( .A(n15798), .ZN(n15790) );
  INV_X1 U19123 ( .A(n15810), .ZN(n15787) );
  NOR3_X1 U19124 ( .A1(n15787), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15786), .ZN(n15788) );
  AOI211_X1 U19125 ( .C1(n15790), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15789), .B(n15788), .ZN(n15793) );
  NAND2_X1 U19126 ( .A1(n15791), .A2(n20736), .ZN(n15792) );
  OAI211_X1 U19127 ( .C1(n15794), .C2(n20775), .A(n15793), .B(n15792), .ZN(
        P1_U3013) );
  AOI21_X1 U19128 ( .B1(n15810), .B2(n15795), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15797) );
  OAI21_X1 U19129 ( .B1(n15798), .B2(n15797), .A(n15796), .ZN(n15799) );
  AOI21_X1 U19130 ( .B1(n15800), .B2(n20736), .A(n15799), .ZN(n15801) );
  OAI21_X1 U19131 ( .B1(n15802), .B2(n20775), .A(n15801), .ZN(P1_U3014) );
  NAND2_X1 U19132 ( .A1(n15803), .A2(n20757), .ZN(n15812) );
  NOR2_X1 U19133 ( .A1(n15804), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15809) );
  AOI21_X1 U19134 ( .B1(n21709), .B2(n15893), .A(n15822), .ZN(n15817) );
  AND2_X1 U19135 ( .A1(n15816), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15805) );
  NAND2_X1 U19136 ( .A1(n15810), .A2(n15805), .ZN(n15815) );
  AOI21_X1 U19137 ( .B1(n15817), .B2(n15815), .A(n15806), .ZN(n15807) );
  AOI211_X1 U19138 ( .C1(n15810), .C2(n15809), .A(n15808), .B(n15807), .ZN(
        n15811) );
  OAI211_X1 U19139 ( .C1(n15813), .C2(n20774), .A(n15812), .B(n15811), .ZN(
        P1_U3015) );
  OAI211_X1 U19140 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        n15818) );
  AOI21_X1 U19141 ( .B1(n20736), .B2(n15819), .A(n15818), .ZN(n15820) );
  OAI21_X1 U19142 ( .B1(n15821), .B2(n20775), .A(n15820), .ZN(P1_U3016) );
  INV_X1 U19143 ( .A(n15822), .ZN(n15823) );
  NOR2_X1 U19144 ( .A1(n15823), .A2(n21709), .ZN(n15824) );
  AOI211_X1 U19145 ( .C1(n20736), .C2(n15826), .A(n15825), .B(n15824), .ZN(
        n15830) );
  NOR2_X1 U19146 ( .A1(n15891), .A2(n15827), .ZN(n15880) );
  NAND2_X1 U19147 ( .A1(n15880), .A2(n15869), .ZN(n15857) );
  OR3_X1 U19148 ( .A1(n15857), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15828), .ZN(n15829) );
  OAI211_X1 U19149 ( .C1(n15831), .C2(n20775), .A(n15830), .B(n15829), .ZN(
        P1_U3017) );
  OAI21_X1 U19150 ( .B1(n15832), .B2(n20722), .A(n9889), .ZN(n15839) );
  INV_X1 U19151 ( .A(n15833), .ZN(n15835) );
  OAI21_X1 U19152 ( .B1(n15835), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15834), .ZN(n15838) );
  NOR2_X1 U19153 ( .A1(n15836), .A2(n20774), .ZN(n15837) );
  AOI211_X1 U19154 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15839), .A(
        n15838), .B(n15837), .ZN(n15840) );
  OAI21_X1 U19155 ( .B1(n15841), .B2(n20775), .A(n15840), .ZN(P1_U3018) );
  INV_X1 U19156 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15844) );
  NAND2_X1 U19157 ( .A1(n15893), .A2(n15842), .ZN(n15843) );
  OAI211_X1 U19158 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n20722), .A(
        n15865), .B(n15843), .ZN(n15860) );
  AOI21_X1 U19159 ( .B1(n15845), .B2(n15844), .A(n15860), .ZN(n15846) );
  NOR2_X1 U19160 ( .A1(n15846), .A2(n15850), .ZN(n15847) );
  AOI211_X1 U19161 ( .C1(n20736), .C2(n15849), .A(n15848), .B(n15847), .ZN(
        n15853) );
  NAND4_X1 U19162 ( .A1(n15885), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15851), .A4(n15850), .ZN(n15852) );
  OAI211_X1 U19163 ( .C1(n15854), .C2(n20775), .A(n15853), .B(n15852), .ZN(
        P1_U3019) );
  OAI21_X1 U19164 ( .B1(n15856), .B2(n20774), .A(n15855), .ZN(n15859) );
  NOR2_X1 U19165 ( .A1(n15857), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15858) );
  AOI211_X1 U19166 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15860), .A(
        n15859), .B(n15858), .ZN(n15861) );
  OAI21_X1 U19167 ( .B1(n15862), .B2(n20775), .A(n15861), .ZN(P1_U3020) );
  AOI21_X1 U19168 ( .B1(n15865), .B2(n15864), .A(n15863), .ZN(n15874) );
  OAI21_X1 U19169 ( .B1(n15867), .B2(n20774), .A(n15866), .ZN(n15868) );
  AOI21_X1 U19170 ( .B1(n15874), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15868), .ZN(n15872) );
  INV_X1 U19171 ( .A(n15869), .ZN(n15870) );
  OAI211_X1 U19172 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15880), .B(n15870), .ZN(
        n15871) );
  OAI211_X1 U19173 ( .C1(n15873), .C2(n20775), .A(n15872), .B(n15871), .ZN(
        P1_U3021) );
  NAND2_X1 U19174 ( .A1(n15874), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15876) );
  OAI211_X1 U19175 ( .C1(n20774), .C2(n15877), .A(n15876), .B(n15875), .ZN(
        n15878) );
  AOI21_X1 U19176 ( .B1(n15880), .B2(n15879), .A(n15878), .ZN(n15881) );
  OAI21_X1 U19177 ( .B1(n15882), .B2(n20775), .A(n15881), .ZN(P1_U3022) );
  INV_X1 U19178 ( .A(n15883), .ZN(n15888) );
  AND4_X1 U19179 ( .A1(n15885), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n15884), .ZN(n15886) );
  AOI211_X1 U19180 ( .C1(n20736), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        n15897) );
  NAND2_X1 U19181 ( .A1(n15889), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15890) );
  NOR2_X1 U19182 ( .A1(n15891), .A2(n15890), .ZN(n15903) );
  AND2_X1 U19183 ( .A1(n15893), .A2(n15892), .ZN(n15894) );
  OR2_X1 U19184 ( .A1(n15895), .A2(n15894), .ZN(n15902) );
  OAI21_X1 U19185 ( .B1(n15903), .B2(n15902), .A(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15896) );
  OAI211_X1 U19186 ( .C1(n15898), .C2(n20775), .A(n15897), .B(n15896), .ZN(
        P1_U3023) );
  INV_X1 U19187 ( .A(n15899), .ZN(n15900) );
  OAI21_X1 U19188 ( .B1(n20774), .B2(n20589), .A(n15900), .ZN(n15901) );
  AOI21_X1 U19189 ( .B1(n15902), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15901), .ZN(n15905) );
  INV_X1 U19190 ( .A(n15903), .ZN(n15904) );
  OAI211_X1 U19191 ( .C1(n15906), .C2(n20775), .A(n15905), .B(n15904), .ZN(
        P1_U3024) );
  AND2_X1 U19192 ( .A1(n21008), .A2(n15909), .ZN(n21006) );
  INV_X1 U19193 ( .A(n21006), .ZN(n15913) );
  AOI22_X1 U19194 ( .A1(n15911), .A2(n21270), .B1(n15910), .B2(n21031), .ZN(
        n15912) );
  OAI211_X1 U19195 ( .C1(n21126), .C2(n21266), .A(n15913), .B(n15912), .ZN(
        n15914) );
  MUX2_X1 U19196 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15914), .S(
        n20782), .Z(P1_U3475) );
  INV_X1 U19197 ( .A(n14504), .ZN(n15916) );
  INV_X1 U19198 ( .A(n14178), .ZN(n15915) );
  NAND2_X1 U19199 ( .A1(n15916), .A2(n15915), .ZN(n15921) );
  OAI21_X1 U19200 ( .B1(n15918), .B2(n15921), .A(n15917), .ZN(n15919) );
  AOI21_X1 U19201 ( .B1(n14513), .B2(n15920), .A(n15919), .ZN(n17091) );
  INV_X1 U19202 ( .A(n15921), .ZN(n15924) );
  AOI22_X1 U19203 ( .A1(n17123), .A2(n15924), .B1(n15923), .B2(n15922), .ZN(
        n15925) );
  OAI21_X1 U19204 ( .B1(n17091), .B2(n15931), .A(n15925), .ZN(n15927) );
  INV_X1 U19205 ( .A(n15926), .ZN(n17166) );
  MUX2_X1 U19206 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15927), .S(
        n17166), .Z(P1_U3473) );
  INV_X1 U19207 ( .A(n15928), .ZN(n15930) );
  OAI22_X1 U19208 ( .A1(n15932), .A2(n15931), .B1(n15930), .B2(n15929), .ZN(
        n15933) );
  MUX2_X1 U19209 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15933), .S(
        n17166), .Z(P1_U3469) );
  NAND2_X1 U19210 ( .A1(n15934), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15938) );
  INV_X1 U19211 ( .A(n15935), .ZN(n17199) );
  OAI21_X1 U19212 ( .B1(n20456), .B2(n20393), .A(n17199), .ZN(n15937) );
  NAND3_X1 U19213 ( .A1(n11607), .A2(n11650), .A3(n20198), .ZN(n15936) );
  OAI211_X1 U19214 ( .C1(n15939), .C2(n15938), .A(n15937), .B(n15936), .ZN(
        n15944) );
  OAI22_X1 U19215 ( .A1(n17002), .A2(n10538), .B1(n15940), .B2(n20456), .ZN(
        n15941) );
  NOR2_X1 U19216 ( .A1(n15942), .A2(n15941), .ZN(n15943) );
  MUX2_X1 U19217 ( .A(n15944), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n15943), 
        .Z(P2_U3610) );
  NAND2_X1 U19218 ( .A1(n15948), .A2(n19809), .ZN(n15953) );
  OAI22_X1 U19219 ( .A1(n19774), .A2(n15950), .B1(n15949), .B2(n19812), .ZN(
        n15951) );
  AOI21_X1 U19220 ( .B1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19787), .A(
        n15951), .ZN(n15952) );
  NAND2_X1 U19221 ( .A1(n16481), .A2(n19819), .ZN(n15963) );
  OAI21_X1 U19222 ( .B1(n15954), .B2(n19820), .A(n19826), .ZN(n15960) );
  INV_X1 U19223 ( .A(n15961), .ZN(n16478) );
  NAND3_X1 U19224 ( .A1(n15954), .A2(n9686), .A3(n16478), .ZN(n15956) );
  AOI22_X1 U19225 ( .A1(n19789), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19807), .ZN(n15955) );
  OAI211_X1 U19226 ( .C1(n19815), .C2(n10735), .A(n15956), .B(n15955), .ZN(
        n15959) );
  NOR2_X1 U19227 ( .A1(n15957), .A2(n19791), .ZN(n15958) );
  AOI211_X1 U19228 ( .C1(n15961), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        n15962) );
  OAI211_X1 U19229 ( .C1(n19813), .C2(n16376), .A(n15963), .B(n15962), .ZN(
        P2_U2827) );
  NOR2_X1 U19230 ( .A1(n13788), .A2(n15964), .ZN(n15965) );
  AOI21_X1 U19231 ( .B1(n15967), .B2(n13780), .A(n13622), .ZN(n16724) );
  XOR2_X1 U19232 ( .A(n16490), .B(n15968), .Z(n15972) );
  AOI22_X1 U19233 ( .A1(n19789), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19807), .ZN(n15969) );
  OAI21_X1 U19234 ( .B1(n19815), .B2(n15970), .A(n15969), .ZN(n15971) );
  AOI21_X1 U19235 ( .B1(n15972), .B2(n19782), .A(n15971), .ZN(n15973) );
  OAI21_X1 U19236 ( .B1(n15974), .B2(n19791), .A(n15973), .ZN(n15975) );
  AOI21_X1 U19237 ( .B1(n16724), .B2(n19794), .A(n15975), .ZN(n15976) );
  OAI21_X1 U19238 ( .B1(n16721), .B2(n16238), .A(n15976), .ZN(P2_U2828) );
  OAI21_X1 U19239 ( .B1(n15977), .B2(n19820), .A(n19826), .ZN(n15981) );
  NAND3_X1 U19240 ( .A1(n15977), .A2(n9686), .A3(n13708), .ZN(n15979) );
  AOI22_X1 U19241 ( .A1(n19789), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19807), .ZN(n15978) );
  OAI211_X1 U19242 ( .C1(n19815), .C2(n21655), .A(n15979), .B(n15978), .ZN(
        n15980) );
  AOI21_X1 U19243 ( .B1(n15982), .B2(n15981), .A(n15980), .ZN(n15983) );
  OAI21_X1 U19244 ( .B1(n15984), .B2(n19791), .A(n15983), .ZN(n15985) );
  AOI21_X1 U19245 ( .B1(n16397), .B2(n19794), .A(n15985), .ZN(n15986) );
  OAI21_X1 U19246 ( .B1(n16287), .B2(n16238), .A(n15986), .ZN(P2_U2829) );
  INV_X1 U19247 ( .A(n15987), .ZN(n15988) );
  AND2_X1 U19248 ( .A1(n15988), .A2(n15989), .ZN(n15990) );
  OR2_X1 U19249 ( .A1(n13781), .A2(n15990), .ZN(n16735) );
  AND2_X1 U19250 ( .A1(n15991), .A2(n15992), .ZN(n15993) );
  OR2_X1 U19251 ( .A1(n15993), .A2(n9835), .ZN(n16736) );
  INV_X1 U19252 ( .A(n16736), .ZN(n15994) );
  NAND2_X1 U19253 ( .A1(n15994), .A2(n19819), .ZN(n16003) );
  XOR2_X1 U19254 ( .A(n16502), .B(n15995), .Z(n16001) );
  AOI22_X1 U19255 ( .A1(n19789), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19807), .ZN(n15996) );
  OAI21_X1 U19256 ( .B1(n19815), .B2(n15997), .A(n15996), .ZN(n16000) );
  NOR2_X1 U19257 ( .A1(n15998), .A2(n19791), .ZN(n15999) );
  AOI211_X1 U19258 ( .C1(n19782), .C2(n16001), .A(n16000), .B(n15999), .ZN(
        n16002) );
  OAI211_X1 U19259 ( .C1(n19813), .C2(n16735), .A(n16003), .B(n16002), .ZN(
        P2_U2830) );
  NAND2_X1 U19260 ( .A1(n16022), .A2(n16005), .ZN(n16006) );
  NAND2_X1 U19261 ( .A1(n15991), .A2(n16006), .ZN(n16747) );
  INV_X1 U19262 ( .A(n16010), .ZN(n16007) );
  AOI21_X1 U19263 ( .B1(n16007), .B2(n19782), .A(n16242), .ZN(n16013) );
  INV_X1 U19264 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20501) );
  OAI22_X1 U19265 ( .A1(n19774), .A2(n16008), .B1(n20501), .B2(n19812), .ZN(
        n16009) );
  AOI21_X1 U19266 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19787), .A(
        n16009), .ZN(n16012) );
  NAND3_X1 U19267 ( .A1(n16010), .A2(n19764), .A3(n13704), .ZN(n16011) );
  OAI211_X1 U19268 ( .C1(n16013), .C2(n13704), .A(n16012), .B(n16011), .ZN(
        n16018) );
  NAND2_X1 U19269 ( .A1(n16025), .A2(n16015), .ZN(n16016) );
  NAND2_X1 U19270 ( .A1(n15988), .A2(n16016), .ZN(n16746) );
  NOR2_X1 U19271 ( .A1(n16746), .A2(n19813), .ZN(n16017) );
  AOI211_X1 U19272 ( .C1(n19809), .C2(n16019), .A(n16018), .B(n16017), .ZN(
        n16020) );
  OAI21_X1 U19273 ( .B1(n16747), .B2(n16238), .A(n16020), .ZN(P2_U2831) );
  OAI21_X1 U19274 ( .B1(n16021), .B2(n16023), .A(n16022), .ZN(n16753) );
  OAI21_X1 U19275 ( .B1(n16024), .B2(n16026), .A(n16025), .ZN(n16760) );
  INV_X1 U19276 ( .A(n16760), .ZN(n16419) );
  INV_X1 U19277 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20499) );
  OAI22_X1 U19278 ( .A1(n19774), .A2(n16027), .B1(n20499), .B2(n19812), .ZN(
        n16031) );
  XNOR2_X1 U19279 ( .A(n16028), .B(n16519), .ZN(n16029) );
  NOR2_X1 U19280 ( .A1(n16029), .A2(n19820), .ZN(n16030) );
  AOI211_X1 U19281 ( .C1(n19787), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16031), .B(n16030), .ZN(n16032) );
  OAI21_X1 U19282 ( .B1(n16033), .B2(n19791), .A(n16032), .ZN(n16034) );
  AOI21_X1 U19283 ( .B1(n16419), .B2(n19794), .A(n16034), .ZN(n16035) );
  OAI21_X1 U19284 ( .B1(n16753), .B2(n16238), .A(n16035), .ZN(P2_U2832) );
  AOI21_X1 U19285 ( .B1(n16037), .B2(n16036), .A(n16021), .ZN(n16763) );
  INV_X1 U19286 ( .A(n16763), .ZN(n16309) );
  AOI21_X1 U19287 ( .B1(n9781), .B2(n19782), .A(n16242), .ZN(n16041) );
  INV_X1 U19288 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20497) );
  OAI22_X1 U19289 ( .A1(n19774), .A2(n21506), .B1(n20497), .B2(n19812), .ZN(
        n16039) );
  NOR3_X1 U19290 ( .A1(n9781), .A2(n10519), .A3(n16195), .ZN(n16038) );
  AOI211_X1 U19291 ( .C1(n19787), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16039), .B(n16038), .ZN(n16040) );
  OAI21_X1 U19292 ( .B1(n16041), .B2(n16528), .A(n16040), .ZN(n16046) );
  AND2_X1 U19293 ( .A1(n16043), .A2(n16042), .ZN(n16044) );
  OR2_X1 U19294 ( .A1(n16044), .A2(n16024), .ZN(n16770) );
  NOR2_X1 U19295 ( .A1(n16770), .A2(n19813), .ZN(n16045) );
  AOI211_X1 U19296 ( .C1(n19809), .C2(n16047), .A(n16046), .B(n16045), .ZN(
        n16048) );
  OAI21_X1 U19297 ( .B1(n16309), .B2(n16238), .A(n16048), .ZN(P2_U2833) );
  OAI21_X1 U19298 ( .B1(n16050), .B2(n19820), .A(n19826), .ZN(n16054) );
  OAI22_X1 U19299 ( .A1(n16049), .A2(n19815), .B1(n20495), .B2(n19812), .ZN(
        n16052) );
  NAND2_X1 U19300 ( .A1(n19764), .A2(n16050), .ZN(n16060) );
  OAI22_X1 U19301 ( .A1(n16053), .A2(n16060), .B1(n19774), .B2(n16316), .ZN(
        n16051) );
  AOI211_X1 U19302 ( .C1(n16054), .C2(n16053), .A(n16052), .B(n16051), .ZN(
        n16057) );
  NAND2_X1 U19303 ( .A1(n16055), .A2(n19809), .ZN(n16056) );
  OAI211_X1 U19304 ( .C1(n16429), .C2(n19813), .A(n16057), .B(n16056), .ZN(
        n16058) );
  AOI21_X1 U19305 ( .B1(n16310), .B2(n19819), .A(n16058), .ZN(n16059) );
  INV_X1 U19306 ( .A(n16059), .ZN(P2_U2834) );
  INV_X1 U19307 ( .A(n16060), .ZN(n16061) );
  OAI21_X1 U19308 ( .B1(n16063), .B2(n16062), .A(n16061), .ZN(n16071) );
  NAND2_X1 U19309 ( .A1(n19787), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16066) );
  OAI22_X1 U19310 ( .A1(n19812), .A2(n20493), .B1(n16063), .B2(n19826), .ZN(
        n16064) );
  INV_X1 U19311 ( .A(n16064), .ZN(n16065) );
  OAI211_X1 U19312 ( .C1(n19774), .C2(n16067), .A(n16066), .B(n16065), .ZN(
        n16068) );
  AOI21_X1 U19313 ( .B1(n16069), .B2(n19809), .A(n16068), .ZN(n16070) );
  OAI211_X1 U19314 ( .C1(n16442), .C2(n19813), .A(n16071), .B(n16070), .ZN(
        n16072) );
  AOI21_X1 U19315 ( .B1(n16073), .B2(n19819), .A(n16072), .ZN(n16074) );
  INV_X1 U19316 ( .A(n16074), .ZN(P2_U2835) );
  INV_X1 U19317 ( .A(n16075), .ZN(n16078) );
  INV_X1 U19318 ( .A(n16076), .ZN(n16077) );
  AOI21_X1 U19319 ( .B1(n16078), .B2(n16077), .A(n11818), .ZN(n16782) );
  OAI21_X1 U19320 ( .B1(n16086), .B2(n19820), .A(n19826), .ZN(n16084) );
  OAI21_X1 U19321 ( .B1(n19812), .B2(n16079), .A(n16706), .ZN(n16080) );
  AOI21_X1 U19322 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19807), .A(n16080), .ZN(
        n16081) );
  OAI21_X1 U19323 ( .B1(n16082), .B2(n19815), .A(n16081), .ZN(n16083) );
  AOI21_X1 U19324 ( .B1(n16085), .B2(n16084), .A(n16083), .ZN(n16089) );
  INV_X1 U19325 ( .A(n16085), .ZN(n16087) );
  NAND3_X1 U19326 ( .A1(n16087), .A2(n9686), .A3(n16086), .ZN(n16088) );
  OAI211_X1 U19327 ( .C1(n16090), .C2(n19791), .A(n16089), .B(n16088), .ZN(
        n16091) );
  AOI21_X1 U19328 ( .B1(n16782), .B2(n19794), .A(n16091), .ZN(n16092) );
  OAI21_X1 U19329 ( .B1(n16784), .B2(n16238), .A(n16092), .ZN(P2_U2836) );
  INV_X1 U19330 ( .A(n11901), .ZN(n16093) );
  OAI21_X1 U19331 ( .B1(n16095), .B2(n16094), .A(n16093), .ZN(n16797) );
  AOI21_X1 U19332 ( .B1(n16096), .B2(n19782), .A(n16242), .ZN(n16102) );
  AOI21_X1 U19333 ( .B1(n19789), .B2(P2_REIP_REG_18__SCAN_IN), .A(n19788), 
        .ZN(n16097) );
  OAI21_X1 U19334 ( .B1(n19774), .B2(n16098), .A(n16097), .ZN(n16099) );
  AOI21_X1 U19335 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19787), .A(
        n16099), .ZN(n16101) );
  NAND3_X1 U19336 ( .A1(n16534), .A2(n19764), .A3(n19763), .ZN(n16100) );
  OAI211_X1 U19337 ( .C1(n16102), .C2(n16534), .A(n16101), .B(n16100), .ZN(
        n16103) );
  AOI21_X1 U19338 ( .B1(n16104), .B2(n19809), .A(n16103), .ZN(n16109) );
  AND2_X1 U19339 ( .A1(n16105), .A2(n16106), .ZN(n16107) );
  NOR2_X1 U19340 ( .A1(n16076), .A2(n16107), .ZN(n16794) );
  NAND2_X1 U19341 ( .A1(n16794), .A2(n19794), .ZN(n16108) );
  OAI211_X1 U19342 ( .C1(n16797), .C2(n16238), .A(n16109), .B(n16108), .ZN(
        P2_U2837) );
  NAND2_X1 U19343 ( .A1(n16836), .A2(n19819), .ZN(n16120) );
  INV_X1 U19344 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n21485) );
  INV_X1 U19345 ( .A(n16111), .ZN(n16110) );
  AOI21_X1 U19346 ( .B1(n19782), .B2(n16110), .A(n16242), .ZN(n16113) );
  NAND3_X1 U19347 ( .A1(n9686), .A2(n16111), .A3(n16558), .ZN(n16112) );
  OAI211_X1 U19348 ( .C1(n16113), .C2(n16558), .A(n16706), .B(n16112), .ZN(
        n16114) );
  AOI21_X1 U19349 ( .B1(n19789), .B2(P2_REIP_REG_15__SCAN_IN), .A(n16114), 
        .ZN(n16115) );
  OAI21_X1 U19350 ( .B1(n19774), .B2(n21485), .A(n16115), .ZN(n16118) );
  NOR2_X1 U19351 ( .A1(n16116), .A2(n19791), .ZN(n16117) );
  AOI211_X1 U19352 ( .C1(n19787), .C2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16118), .B(n16117), .ZN(n16119) );
  OAI211_X1 U19353 ( .C1(n19813), .C2(n16833), .A(n16120), .B(n16119), .ZN(
        P2_U2840) );
  NAND2_X1 U19354 ( .A1(n16852), .A2(n19819), .ZN(n16131) );
  AOI21_X1 U19355 ( .B1(n19782), .B2(n16121), .A(n16242), .ZN(n16123) );
  NOR2_X1 U19356 ( .A1(n16195), .A2(n16121), .ZN(n16132) );
  NAND2_X1 U19357 ( .A1(n16132), .A2(n16565), .ZN(n16122) );
  OAI211_X1 U19358 ( .C1(n16565), .C2(n16123), .A(n16122), .B(n16706), .ZN(
        n16124) );
  AOI21_X1 U19359 ( .B1(n19789), .B2(P2_REIP_REG_14__SCAN_IN), .A(n16124), 
        .ZN(n16126) );
  NAND2_X1 U19360 ( .A1(n19787), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16125) );
  OAI211_X1 U19361 ( .C1(n19774), .C2(n16127), .A(n16126), .B(n16125), .ZN(
        n16128) );
  AOI21_X1 U19362 ( .B1(n16129), .B2(n19809), .A(n16128), .ZN(n16130) );
  OAI211_X1 U19363 ( .C1(n19813), .C2(n16850), .A(n16131), .B(n16130), .ZN(
        P2_U2841) );
  INV_X1 U19364 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20483) );
  INV_X1 U19365 ( .A(n16132), .ZN(n16133) );
  AOI21_X1 U19366 ( .B1(n16578), .B2(n16134), .A(n16133), .ZN(n16135) );
  AOI211_X1 U19367 ( .C1(n16578), .C2(n16242), .A(n19788), .B(n16135), .ZN(
        n16136) );
  OAI21_X1 U19368 ( .B1(n19812), .B2(n20483), .A(n16136), .ZN(n16137) );
  AOI21_X1 U19369 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n19807), .A(n16137), .ZN(
        n16138) );
  OAI21_X1 U19370 ( .B1(n21703), .B2(n19815), .A(n16138), .ZN(n16140) );
  NOR2_X1 U19371 ( .A1(n16859), .A2(n19813), .ZN(n16139) );
  OAI21_X1 U19372 ( .B1(n16865), .B2(n16238), .A(n16142), .ZN(P2_U2842) );
  AND2_X1 U19373 ( .A1(n14023), .A2(n16143), .ZN(n16145) );
  OR2_X1 U19374 ( .A1(n16145), .A2(n16144), .ZN(n16348) );
  NAND2_X1 U19375 ( .A1(n16880), .A2(n19819), .ZN(n16158) );
  INV_X1 U19376 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n16153) );
  NAND2_X1 U19377 ( .A1(n16147), .A2(n19782), .ZN(n16146) );
  AOI21_X1 U19378 ( .B1(n19826), .B2(n16146), .A(n16590), .ZN(n16151) );
  INV_X1 U19379 ( .A(n16147), .ZN(n16148) );
  NAND3_X1 U19380 ( .A1(n19764), .A2(n16590), .A3(n16148), .ZN(n16149) );
  NAND2_X1 U19381 ( .A1(n16149), .A2(n16706), .ZN(n16150) );
  AOI211_X1 U19382 ( .C1(n19789), .C2(P2_REIP_REG_12__SCAN_IN), .A(n16151), 
        .B(n16150), .ZN(n16152) );
  OAI21_X1 U19383 ( .B1(n19774), .B2(n16153), .A(n16152), .ZN(n16156) );
  NOR2_X1 U19384 ( .A1(n16154), .A2(n19791), .ZN(n16155) );
  AOI211_X1 U19385 ( .C1(n19787), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16156), .B(n16155), .ZN(n16157) );
  OAI211_X1 U19386 ( .C1(n16878), .C2(n19813), .A(n16158), .B(n16157), .ZN(
        P2_U2843) );
  INV_X1 U19387 ( .A(n16896), .ZN(n16159) );
  NAND2_X1 U19388 ( .A1(n16159), .A2(n19819), .ZN(n16171) );
  AOI21_X1 U19389 ( .B1(n19782), .B2(n16160), .A(n16242), .ZN(n16163) );
  INV_X1 U19390 ( .A(n16160), .ZN(n16161) );
  NAND3_X1 U19391 ( .A1(n16161), .A2(n19764), .A3(n16616), .ZN(n16162) );
  OAI211_X1 U19392 ( .C1(n16163), .C2(n16616), .A(n16706), .B(n16162), .ZN(
        n16164) );
  AOI21_X1 U19393 ( .B1(n19789), .B2(P2_REIP_REG_10__SCAN_IN), .A(n16164), 
        .ZN(n16165) );
  OAI21_X1 U19394 ( .B1(n19774), .B2(n16166), .A(n16165), .ZN(n16169) );
  NOR2_X1 U19395 ( .A1(n16167), .A2(n19791), .ZN(n16168) );
  AOI211_X1 U19396 ( .C1(n19787), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16169), .B(n16168), .ZN(n16170) );
  OAI211_X1 U19397 ( .C1(n19813), .C2(n16903), .A(n16171), .B(n16170), .ZN(
        P2_U2845) );
  INV_X1 U19398 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16630) );
  NAND2_X1 U19399 ( .A1(n16172), .A2(n19809), .ZN(n16178) );
  NAND2_X1 U19400 ( .A1(n9682), .A2(n9795), .ZN(n16173) );
  XOR2_X1 U19401 ( .A(n16633), .B(n16173), .Z(n16175) );
  NAND2_X1 U19402 ( .A1(n19789), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n16174) );
  OAI211_X1 U19403 ( .C1(n19820), .C2(n16175), .A(n16174), .B(n16706), .ZN(
        n16176) );
  AOI21_X1 U19404 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n19807), .A(n16176), .ZN(
        n16177) );
  OAI211_X1 U19405 ( .C1(n19815), .C2(n16630), .A(n16178), .B(n16177), .ZN(
        n16179) );
  AOI21_X1 U19406 ( .B1(n16918), .B2(n19794), .A(n16179), .ZN(n16180) );
  OAI21_X1 U19407 ( .B1(n16915), .B2(n16238), .A(n16180), .ZN(P2_U2846) );
  INV_X1 U19408 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16190) );
  NAND2_X1 U19409 ( .A1(n16181), .A2(n19809), .ZN(n16189) );
  OAI21_X1 U19410 ( .B1(n19820), .B2(n16182), .A(n19826), .ZN(n16185) );
  INV_X1 U19411 ( .A(n16182), .ZN(n16183) );
  NOR3_X1 U19412 ( .A1(n16195), .A2(n16641), .A3(n16183), .ZN(n16184) );
  AOI211_X1 U19413 ( .C1(n16641), .C2(n16185), .A(n19788), .B(n16184), .ZN(
        n16186) );
  OAI21_X1 U19414 ( .B1(n19812), .B2(n20474), .A(n16186), .ZN(n16187) );
  AOI21_X1 U19415 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19807), .A(n16187), .ZN(
        n16188) );
  OAI211_X1 U19416 ( .C1(n19815), .C2(n16190), .A(n16189), .B(n16188), .ZN(
        n16191) );
  AOI21_X1 U19417 ( .B1(n16928), .B2(n19794), .A(n16191), .ZN(n16192) );
  OAI21_X1 U19418 ( .B1(n16930), .B2(n16238), .A(n16192), .ZN(P2_U2847) );
  NAND2_X1 U19419 ( .A1(n19789), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16199) );
  OAI21_X1 U19420 ( .B1(n16193), .B2(n19820), .A(n19826), .ZN(n16197) );
  INV_X1 U19421 ( .A(n16193), .ZN(n16194) );
  NOR3_X1 U19422 ( .A1(n16195), .A2(n16655), .A3(n16194), .ZN(n16196) );
  AOI211_X1 U19423 ( .C1(n16655), .C2(n16197), .A(n19788), .B(n16196), .ZN(
        n16198) );
  OAI211_X1 U19424 ( .C1(n19774), .C2(n11434), .A(n16199), .B(n16198), .ZN(
        n16200) );
  AOI21_X1 U19425 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19787), .A(
        n16200), .ZN(n16201) );
  OAI21_X1 U19426 ( .B1(n16202), .B2(n19791), .A(n16201), .ZN(n16203) );
  AOI21_X1 U19427 ( .B1(n16940), .B2(n19794), .A(n16203), .ZN(n16204) );
  OAI21_X1 U19428 ( .B1(n16942), .B2(n16238), .A(n16204), .ZN(P2_U2848) );
  INV_X1 U19429 ( .A(n16205), .ZN(n16950) );
  AOI21_X1 U19430 ( .B1(n16206), .B2(n19782), .A(n16242), .ZN(n16208) );
  NAND3_X1 U19431 ( .A1(n10525), .A2(n16663), .A3(n9686), .ZN(n16207) );
  OAI211_X1 U19432 ( .C1(n16208), .C2(n16663), .A(n16706), .B(n16207), .ZN(
        n16209) );
  AOI21_X1 U19433 ( .B1(n19789), .B2(P2_REIP_REG_6__SCAN_IN), .A(n16209), .ZN(
        n16210) );
  OAI21_X1 U19434 ( .B1(n19774), .B2(n16211), .A(n16210), .ZN(n16212) );
  AOI21_X1 U19435 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19787), .A(
        n16212), .ZN(n16213) );
  OAI21_X1 U19436 ( .B1(n16214), .B2(n19791), .A(n16213), .ZN(n16215) );
  AOI21_X1 U19437 ( .B1(n16950), .B2(n19794), .A(n16215), .ZN(n16216) );
  OAI21_X1 U19438 ( .B1(n16217), .B2(n16238), .A(n16216), .ZN(P2_U2849) );
  NAND2_X1 U19439 ( .A1(n16971), .A2(n19819), .ZN(n16228) );
  NAND2_X1 U19440 ( .A1(n19807), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n16222) );
  NAND2_X1 U19441 ( .A1(n16218), .A2(n9682), .ZN(n16219) );
  XNOR2_X1 U19442 ( .A(n16219), .B(n16670), .ZN(n16220) );
  AOI21_X1 U19443 ( .B1(n16220), .B2(n19782), .A(n19788), .ZN(n16221) );
  OAI211_X1 U19444 ( .C1(n19812), .C2(n16223), .A(n16222), .B(n16221), .ZN(
        n16226) );
  NOR2_X1 U19445 ( .A1(n16224), .A2(n19791), .ZN(n16225) );
  AOI211_X1 U19446 ( .C1(n19787), .C2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16226), .B(n16225), .ZN(n16227) );
  OAI211_X1 U19447 ( .C1(n16961), .C2(n19813), .A(n16228), .B(n16227), .ZN(
        P2_U2850) );
  AOI21_X1 U19448 ( .B1(n19782), .B2(n16229), .A(n16242), .ZN(n16232) );
  INV_X1 U19449 ( .A(n16229), .ZN(n16230) );
  NAND3_X1 U19450 ( .A1(n19764), .A2(n16709), .A3(n16230), .ZN(n16231) );
  OAI21_X1 U19451 ( .B1(n16232), .B2(n16709), .A(n16231), .ZN(n16234) );
  NOR2_X1 U19452 ( .A1(n19812), .A2(n16705), .ZN(n16233) );
  AOI211_X1 U19453 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19807), .A(n16234), .B(
        n16233), .ZN(n16236) );
  NAND2_X1 U19454 ( .A1(n19787), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16235) );
  OAI211_X1 U19455 ( .C1(n19791), .C2(n16237), .A(n16236), .B(n16235), .ZN(
        n16240) );
  NOR2_X1 U19456 ( .A1(n11180), .A2(n16238), .ZN(n16239) );
  AOI211_X1 U19457 ( .C1(n20529), .C2(n19794), .A(n16240), .B(n16239), .ZN(
        n16241) );
  OAI21_X1 U19458 ( .B1(n20155), .B2(n19796), .A(n16241), .ZN(P2_U2852) );
  NAND2_X1 U19459 ( .A1(n19807), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n16249) );
  AOI21_X1 U19460 ( .B1(n19782), .B2(n17015), .A(n16242), .ZN(n16245) );
  NAND3_X1 U19461 ( .A1(n19764), .A2(n16244), .A3(n10510), .ZN(n16243) );
  OAI21_X1 U19462 ( .B1(n16245), .B2(n16244), .A(n16243), .ZN(n16246) );
  AOI21_X1 U19463 ( .B1(n19809), .B2(n16247), .A(n16246), .ZN(n16248) );
  OAI211_X1 U19464 ( .C1(n19812), .C2(n11130), .A(n16249), .B(n16248), .ZN(
        n16250) );
  AOI21_X1 U19465 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19787), .A(
        n16250), .ZN(n16251) );
  OAI21_X1 U19466 ( .B1(n16252), .B2(n19813), .A(n16251), .ZN(n16253) );
  OAI21_X1 U19467 ( .B1(n16255), .B2(n19796), .A(n16254), .ZN(P2_U2853) );
  AOI22_X1 U19468 ( .A1(n19789), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19794), 
        .B2(n16256), .ZN(n16259) );
  AOI22_X1 U19469 ( .A1(n19809), .A2(n16257), .B1(n19764), .B2(n17012), .ZN(
        n16258) );
  OAI211_X1 U19470 ( .C1(n16260), .C2(n19774), .A(n16259), .B(n16258), .ZN(
        n16263) );
  INV_X1 U19471 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16261) );
  AOI21_X1 U19472 ( .B1(n19815), .B2(n19826), .A(n16261), .ZN(n16262) );
  AOI211_X1 U19473 ( .C1(n19819), .C2(n11168), .A(n16263), .B(n16262), .ZN(
        n16264) );
  OAI21_X1 U19474 ( .B1(n19796), .B2(n17033), .A(n16264), .ZN(P2_U2855) );
  MUX2_X1 U19475 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16265), .S(n19832), .Z(
        P2_U2856) );
  NAND2_X1 U19476 ( .A1(n16267), .A2(n16266), .ZN(n16371) );
  NAND3_X1 U19477 ( .A1(n16373), .A2(n19828), .A3(n16371), .ZN(n16269) );
  NAND2_X1 U19478 ( .A1(n16351), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16268) );
  OAI211_X1 U19479 ( .C1(n15945), .C2(n16351), .A(n16269), .B(n16268), .ZN(
        P2_U2858) );
  NAND2_X1 U19480 ( .A1(n16271), .A2(n16270), .ZN(n16273) );
  XNOR2_X1 U19481 ( .A(n16273), .B(n16272), .ZN(n16384) );
  NOR2_X1 U19482 ( .A1(n16274), .A2(n16351), .ZN(n16275) );
  AOI21_X1 U19483 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16351), .A(n16275), .ZN(
        n16276) );
  OAI21_X1 U19484 ( .B1(n16384), .B2(n16354), .A(n16276), .ZN(P2_U2859) );
  NAND2_X1 U19485 ( .A1(n16385), .A2(n19828), .ZN(n16280) );
  NAND2_X1 U19486 ( .A1(n16351), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16279) );
  OAI211_X1 U19487 ( .C1(n16721), .C2(n16351), .A(n16280), .B(n16279), .ZN(
        P2_U2860) );
  NAND2_X1 U19488 ( .A1(n16281), .A2(n16291), .ZN(n16290) );
  NOR2_X1 U19489 ( .A1(n16282), .A2(n14347), .ZN(n16283) );
  XNOR2_X1 U19490 ( .A(n16284), .B(n16283), .ZN(n16285) );
  XNOR2_X1 U19491 ( .A(n16286), .B(n16285), .ZN(n16399) );
  MUX2_X1 U19492 ( .A(n16288), .B(n16287), .S(n19832), .Z(n16289) );
  OAI21_X1 U19493 ( .B1(n16399), .B2(n16354), .A(n16289), .ZN(P2_U2861) );
  OAI21_X1 U19494 ( .B1(n16281), .B2(n16291), .A(n16290), .ZN(n16406) );
  MUX2_X1 U19495 ( .A(n16736), .B(n16292), .S(n16351), .Z(n16293) );
  OAI21_X1 U19496 ( .B1(n16354), .B2(n16406), .A(n16293), .ZN(P2_U2862) );
  OAI21_X1 U19497 ( .B1(n16296), .B2(n16295), .A(n16294), .ZN(n16413) );
  NOR2_X1 U19498 ( .A1(n16747), .A2(n16351), .ZN(n16297) );
  AOI21_X1 U19499 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16351), .A(n16297), .ZN(
        n16298) );
  OAI21_X1 U19500 ( .B1(n16354), .B2(n16413), .A(n16298), .ZN(P2_U2863) );
  OAI21_X1 U19501 ( .B1(n16299), .B2(n16301), .A(n16300), .ZN(n16421) );
  NOR2_X1 U19502 ( .A1(n16753), .A2(n16351), .ZN(n16303) );
  AOI21_X1 U19503 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16351), .A(n16303), .ZN(
        n16304) );
  OAI21_X1 U19504 ( .B1(n16354), .B2(n16421), .A(n16304), .ZN(P2_U2864) );
  OAI21_X1 U19505 ( .B1(n16313), .B2(n16306), .A(n16305), .ZN(n16427) );
  INV_X1 U19506 ( .A(n16427), .ZN(n16307) );
  AOI22_X1 U19507 ( .A1(n16307), .A2(n19828), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16351), .ZN(n16308) );
  OAI21_X1 U19508 ( .B1(n16309), .B2(n16351), .A(n16308), .ZN(P2_U2865) );
  NAND2_X1 U19509 ( .A1(n16310), .A2(n19832), .ZN(n16315) );
  AND2_X1 U19510 ( .A1(n16318), .A2(n16311), .ZN(n16312) );
  NOR2_X1 U19511 ( .A1(n16313), .A2(n16312), .ZN(n16428) );
  NAND2_X1 U19512 ( .A1(n16428), .A2(n19828), .ZN(n16314) );
  OAI211_X1 U19513 ( .C1(n19832), .C2(n16316), .A(n16315), .B(n16314), .ZN(
        P2_U2866) );
  INV_X1 U19514 ( .A(n16318), .ZN(n16319) );
  AOI21_X1 U19515 ( .B1(n16320), .B2(n16317), .A(n16319), .ZN(n16437) );
  AOI22_X1 U19516 ( .A1(n16437), .A2(n19828), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n16351), .ZN(n16321) );
  OAI21_X1 U19517 ( .B1(n16322), .B2(n16351), .A(n16321), .ZN(P2_U2867) );
  AOI21_X1 U19518 ( .B1(n16324), .B2(n16323), .A(n12293), .ZN(n16447) );
  AOI22_X1 U19519 ( .A1(n16447), .A2(n19828), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16351), .ZN(n16325) );
  OAI21_X1 U19520 ( .B1(n16784), .B2(n16351), .A(n16325), .ZN(P2_U2868) );
  OAI21_X1 U19521 ( .B1(n9850), .B2(n16326), .A(n16323), .ZN(n16460) );
  INV_X1 U19522 ( .A(n16460), .ZN(n16327) );
  AOI22_X1 U19523 ( .A1(n16327), .A2(n19828), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n16351), .ZN(n16328) );
  OAI21_X1 U19524 ( .B1(n16797), .B2(n16351), .A(n16328), .ZN(P2_U2869) );
  XNOR2_X1 U19525 ( .A(n16335), .B(n16330), .ZN(n16815) );
  NAND2_X1 U19526 ( .A1(n16351), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16334) );
  AND2_X1 U19527 ( .A1(n14804), .A2(n16331), .ZN(n16332) );
  NOR2_X1 U19528 ( .A1(n9850), .A2(n16332), .ZN(n16461) );
  NAND2_X1 U19529 ( .A1(n16461), .A2(n19828), .ZN(n16333) );
  OAI211_X1 U19530 ( .C1(n16815), .C2(n16351), .A(n16334), .B(n16333), .ZN(
        P2_U2870) );
  INV_X1 U19531 ( .A(n16335), .ZN(n16336) );
  AOI21_X1 U19532 ( .B1(n16338), .B2(n16337), .A(n16336), .ZN(n19784) );
  NAND2_X1 U19533 ( .A1(n19784), .A2(n19832), .ZN(n16340) );
  NAND2_X1 U19534 ( .A1(n16351), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16339) );
  OAI211_X1 U19535 ( .C1(n16341), .C2(n16354), .A(n16340), .B(n16339), .ZN(
        P2_U2871) );
  INV_X1 U19536 ( .A(n16342), .ZN(n16349) );
  OAI21_X1 U19537 ( .B1(n16350), .B2(n16349), .A(n16343), .ZN(n16345) );
  NAND3_X1 U19538 ( .A1(n16345), .A2(n19828), .A3(n16344), .ZN(n16347) );
  NAND2_X1 U19539 ( .A1(n16351), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n16346) );
  OAI211_X1 U19540 ( .C1(n16348), .C2(n16351), .A(n16347), .B(n16346), .ZN(
        P2_U2875) );
  XNOR2_X1 U19541 ( .A(n16350), .B(n16349), .ZN(n16355) );
  NAND2_X1 U19542 ( .A1(n16351), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n16353) );
  NAND2_X1 U19543 ( .A1(n16892), .A2(n19832), .ZN(n16352) );
  OAI211_X1 U19544 ( .C1(n16355), .C2(n16354), .A(n16353), .B(n16352), .ZN(
        P2_U2876) );
  INV_X1 U19545 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U19546 ( .A1(n16466), .A2(n16356), .B1(n16465), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n16357) );
  OAI21_X1 U19547 ( .B1(n16470), .B2(n16358), .A(n16357), .ZN(n16359) );
  INV_X1 U19548 ( .A(n16359), .ZN(n16361) );
  INV_X1 U19549 ( .A(n16362), .ZN(n16363) );
  OAI21_X1 U19550 ( .B1(n16364), .B2(n16475), .A(n16363), .ZN(P2_U2889) );
  INV_X1 U19551 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16368) );
  NAND2_X1 U19552 ( .A1(n16464), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19553 ( .A1(n16466), .A2(n16365), .B1(n16465), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16366) );
  OAI211_X1 U19554 ( .C1(n16470), .C2(n16368), .A(n16367), .B(n16366), .ZN(
        n16369) );
  AOI21_X1 U19555 ( .B1(n16370), .B2(n16472), .A(n16369), .ZN(n16375) );
  NAND3_X1 U19556 ( .A1(n16373), .A2(n16372), .A3(n16371), .ZN(n16374) );
  NAND2_X1 U19557 ( .A1(n16375), .A2(n16374), .ZN(P2_U2890) );
  INV_X1 U19558 ( .A(n16376), .ZN(n16382) );
  INV_X1 U19559 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U19560 ( .A1(n16464), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16379) );
  AOI22_X1 U19561 ( .A1(n16466), .A2(n16377), .B1(n16465), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16378) );
  OAI211_X1 U19562 ( .C1(n16470), .C2(n16380), .A(n16379), .B(n16378), .ZN(
        n16381) );
  AOI21_X1 U19563 ( .B1(n16382), .B2(n16472), .A(n16381), .ZN(n16383) );
  OAI21_X1 U19564 ( .B1(n16384), .B2(n16475), .A(n16383), .ZN(P2_U2891) );
  INV_X1 U19565 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n16388) );
  NAND2_X1 U19566 ( .A1(n16464), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16387) );
  AOI22_X1 U19567 ( .A1(n16466), .A2(n19833), .B1(n16465), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16386) );
  OAI211_X1 U19568 ( .C1(n16470), .C2(n16388), .A(n16387), .B(n16386), .ZN(
        n16389) );
  AOI21_X1 U19569 ( .B1(n16724), .B2(n16472), .A(n16389), .ZN(n16390) );
  OAI21_X1 U19570 ( .B1(n16475), .B2(n16391), .A(n16390), .ZN(P2_U2892) );
  INV_X1 U19571 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16395) );
  NAND2_X1 U19572 ( .A1(n16464), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16394) );
  AOI22_X1 U19573 ( .A1(n16466), .A2(n16392), .B1(n16465), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16393) );
  OAI211_X1 U19574 ( .C1(n16470), .C2(n16395), .A(n16394), .B(n16393), .ZN(
        n16396) );
  AOI21_X1 U19575 ( .B1(n16397), .B2(n16472), .A(n16396), .ZN(n16398) );
  OAI21_X1 U19576 ( .B1(n16399), .B2(n16475), .A(n16398), .ZN(P2_U2893) );
  INV_X1 U19577 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16402) );
  AOI22_X1 U19578 ( .A1(n16466), .A2(n16400), .B1(n16465), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16401) );
  OAI21_X1 U19579 ( .B1(n16470), .B2(n16402), .A(n16401), .ZN(n16404) );
  NOR2_X1 U19580 ( .A1(n16735), .A2(n16441), .ZN(n16403) );
  AOI211_X1 U19581 ( .C1(n16464), .C2(BUF1_REG_25__SCAN_IN), .A(n16404), .B(
        n16403), .ZN(n16405) );
  OAI21_X1 U19582 ( .B1(n16475), .B2(n16406), .A(n16405), .ZN(P2_U2894) );
  INV_X1 U19583 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16409) );
  AOI22_X1 U19584 ( .A1(n16466), .A2(n16407), .B1(n16465), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16408) );
  OAI21_X1 U19585 ( .B1(n16470), .B2(n16409), .A(n16408), .ZN(n16411) );
  NOR2_X1 U19586 ( .A1(n16746), .A2(n16441), .ZN(n16410) );
  AOI211_X1 U19587 ( .C1(n16464), .C2(BUF1_REG_24__SCAN_IN), .A(n16411), .B(
        n16410), .ZN(n16412) );
  OAI21_X1 U19588 ( .B1(n16475), .B2(n16413), .A(n16412), .ZN(P2_U2895) );
  INV_X1 U19589 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16417) );
  NAND2_X1 U19590 ( .A1(n16464), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16416) );
  AOI22_X1 U19591 ( .A1(n16466), .A2(n16414), .B1(n16465), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16415) );
  OAI211_X1 U19592 ( .C1(n16470), .C2(n16417), .A(n16416), .B(n16415), .ZN(
        n16418) );
  AOI21_X1 U19593 ( .B1(n16419), .B2(n16472), .A(n16418), .ZN(n16420) );
  OAI21_X1 U19594 ( .B1(n16475), .B2(n16421), .A(n16420), .ZN(P2_U2896) );
  AOI22_X1 U19595 ( .A1(n16466), .A2(n16422), .B1(n16465), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16423) );
  OAI21_X1 U19596 ( .B1(n16470), .B2(n21624), .A(n16423), .ZN(n16425) );
  NOR2_X1 U19597 ( .A1(n16770), .A2(n16441), .ZN(n16424) );
  AOI211_X1 U19598 ( .C1(BUF1_REG_22__SCAN_IN), .C2(n16464), .A(n16425), .B(
        n16424), .ZN(n16426) );
  OAI21_X1 U19599 ( .B1(n16475), .B2(n16427), .A(n16426), .ZN(P2_U2897) );
  INV_X1 U19600 ( .A(n16428), .ZN(n16436) );
  INV_X1 U19601 ( .A(n16429), .ZN(n16434) );
  INV_X1 U19602 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16432) );
  NAND2_X1 U19603 ( .A1(n16464), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16431) );
  AOI22_X1 U19604 ( .A1(n16466), .A2(n19880), .B1(n16465), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16430) );
  OAI211_X1 U19605 ( .C1(n16470), .C2(n16432), .A(n16431), .B(n16430), .ZN(
        n16433) );
  AOI21_X1 U19606 ( .B1(n16434), .B2(n16472), .A(n16433), .ZN(n16435) );
  OAI21_X1 U19607 ( .B1(n16475), .B2(n16436), .A(n16435), .ZN(P2_U2898) );
  INV_X1 U19608 ( .A(n16437), .ZN(n16446) );
  INV_X1 U19609 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16440) );
  AOI22_X1 U19610 ( .A1(n16466), .A2(n16438), .B1(n16465), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16439) );
  OAI21_X1 U19611 ( .B1(n16470), .B2(n16440), .A(n16439), .ZN(n16444) );
  NOR2_X1 U19612 ( .A1(n16442), .A2(n16441), .ZN(n16443) );
  AOI211_X1 U19613 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n16464), .A(n16444), .B(
        n16443), .ZN(n16445) );
  OAI21_X1 U19614 ( .B1(n16475), .B2(n16446), .A(n16445), .ZN(P2_U2899) );
  INV_X1 U19615 ( .A(n16447), .ZN(n16454) );
  INV_X1 U19616 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16451) );
  NAND2_X1 U19617 ( .A1(n16464), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16450) );
  AOI22_X1 U19618 ( .A1(n16466), .A2(n16448), .B1(n16465), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16449) );
  OAI211_X1 U19619 ( .C1(n16470), .C2(n16451), .A(n16450), .B(n16449), .ZN(
        n16452) );
  AOI21_X1 U19620 ( .B1(n16782), .B2(n16472), .A(n16452), .ZN(n16453) );
  OAI21_X1 U19621 ( .B1(n16475), .B2(n16454), .A(n16453), .ZN(P2_U2900) );
  INV_X1 U19622 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16457) );
  NAND2_X1 U19623 ( .A1(n16464), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16456) );
  AOI22_X1 U19624 ( .A1(n16466), .A2(n19870), .B1(n16465), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16455) );
  OAI211_X1 U19625 ( .C1(n16470), .C2(n16457), .A(n16456), .B(n16455), .ZN(
        n16458) );
  AOI21_X1 U19626 ( .B1(n16794), .B2(n16472), .A(n16458), .ZN(n16459) );
  OAI21_X1 U19627 ( .B1(n16475), .B2(n16460), .A(n16459), .ZN(P2_U2901) );
  INV_X1 U19628 ( .A(n16461), .ZN(n16474) );
  INV_X1 U19629 ( .A(n16105), .ZN(n16462) );
  AOI21_X1 U19630 ( .B1(n16463), .B2(n14807), .A(n16462), .ZN(n19761) );
  INV_X1 U19631 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16469) );
  NAND2_X1 U19632 ( .A1(n16464), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16468) );
  AOI22_X1 U19633 ( .A1(n16466), .A2(n17046), .B1(n16465), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16467) );
  OAI211_X1 U19634 ( .C1(n16470), .C2(n16469), .A(n16468), .B(n16467), .ZN(
        n16471) );
  AOI21_X1 U19635 ( .B1(n19761), .B2(n16472), .A(n16471), .ZN(n16473) );
  OAI21_X1 U19636 ( .B1(n16475), .B2(n16474), .A(n16473), .ZN(P2_U2902) );
  NAND2_X1 U19637 ( .A1(n16707), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16476) );
  OAI211_X1 U19638 ( .C1(n16710), .C2(n16478), .A(n16477), .B(n16476), .ZN(
        n16480) );
  OAI21_X1 U19639 ( .B1(n16483), .B2(n16680), .A(n16482), .ZN(P2_U2986) );
  XNOR2_X1 U19640 ( .A(n16486), .B(n16719), .ZN(n16487) );
  INV_X1 U19641 ( .A(n16721), .ZN(n16493) );
  INV_X1 U19642 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n16488) );
  OR2_X1 U19643 ( .A1(n16706), .A2(n16488), .ZN(n16717) );
  NAND2_X1 U19644 ( .A1(n16707), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16489) );
  OAI211_X1 U19645 ( .C1(n16710), .C2(n16490), .A(n16717), .B(n16489), .ZN(
        n16492) );
  INV_X1 U19646 ( .A(n16495), .ZN(n16498) );
  NOR2_X1 U19647 ( .A1(n16498), .A2(n16496), .ZN(n16497) );
  INV_X1 U19648 ( .A(n16510), .ZN(n16501) );
  AOI21_X1 U19649 ( .B1(n16732), .B2(n16501), .A(n16500), .ZN(n16739) );
  INV_X1 U19650 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20503) );
  NOR2_X1 U19651 ( .A1(n16706), .A2(n20503), .ZN(n16731) );
  NOR2_X1 U19652 ( .A1(n16710), .A2(n16502), .ZN(n16503) );
  AOI211_X1 U19653 ( .C1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n16707), .A(
        n16731), .B(n16503), .ZN(n16504) );
  OAI21_X1 U19654 ( .B1(n16736), .B2(n16695), .A(n16504), .ZN(n16505) );
  AOI21_X1 U19655 ( .B1(n16697), .B2(n16739), .A(n16505), .ZN(n16506) );
  XNOR2_X1 U19656 ( .A(n16507), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16508) );
  XNOR2_X1 U19657 ( .A(n16509), .B(n16508), .ZN(n16752) );
  AOI21_X1 U19658 ( .B1(n10547), .B2(n16511), .A(n16510), .ZN(n16750) );
  NOR2_X1 U19659 ( .A1(n16706), .A2(n20501), .ZN(n16743) );
  AOI21_X1 U19660 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16743), .ZN(n16514) );
  NAND2_X1 U19661 ( .A1(n16692), .A2(n16512), .ZN(n16513) );
  OAI211_X1 U19662 ( .C1(n16747), .C2(n16695), .A(n16514), .B(n16513), .ZN(
        n16515) );
  AOI21_X1 U19663 ( .B1(n16697), .B2(n16750), .A(n16515), .ZN(n16516) );
  OAI21_X1 U19664 ( .B1(n16752), .B2(n16680), .A(n16516), .ZN(P2_U2990) );
  NOR2_X1 U19665 ( .A1(n16706), .A2(n20499), .ZN(n16758) );
  NOR2_X1 U19666 ( .A1(n16710), .A2(n16519), .ZN(n16520) );
  AOI211_X1 U19667 ( .C1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n16707), .A(
        n16758), .B(n16520), .ZN(n16521) );
  OAI21_X1 U19668 ( .B1(n16753), .B2(n16695), .A(n16521), .ZN(n16522) );
  NOR2_X1 U19669 ( .A1(n16523), .A2(n9876), .ZN(n16524) );
  XNOR2_X1 U19670 ( .A(n16525), .B(n16524), .ZN(n16772) );
  NAND2_X1 U19671 ( .A1(n16763), .A2(n16715), .ZN(n16527) );
  NOR2_X1 U19672 ( .A1(n16706), .A2(n20497), .ZN(n16766) );
  AOI21_X1 U19673 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16766), .ZN(n16526) );
  OAI211_X1 U19674 ( .C1(n16710), .C2(n16528), .A(n16527), .B(n16526), .ZN(
        n16529) );
  AOI21_X1 U19675 ( .B1(n16772), .B2(n11531), .A(n16529), .ZN(n16530) );
  NAND2_X1 U19676 ( .A1(n11525), .A2(n16531), .ZN(n16532) );
  XNOR2_X1 U19677 ( .A(n11909), .B(n16532), .ZN(n16801) );
  INV_X1 U19678 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20490) );
  NOR2_X1 U19679 ( .A1(n16706), .A2(n20490), .ZN(n16792) );
  NOR2_X1 U19680 ( .A1(n16534), .A2(n16710), .ZN(n16535) );
  AOI211_X1 U19681 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n16707), .A(
        n16792), .B(n16535), .ZN(n16536) );
  OAI21_X1 U19682 ( .B1(n16797), .B2(n16695), .A(n16536), .ZN(n16537) );
  AOI21_X1 U19683 ( .B1(n16799), .B2(n16697), .A(n16537), .ZN(n16538) );
  OAI21_X1 U19684 ( .B1(n16680), .B2(n16801), .A(n16538), .ZN(P2_U2996) );
  XOR2_X1 U19685 ( .A(n16540), .B(n16539), .Z(n16817) );
  INV_X1 U19686 ( .A(n16815), .ZN(n19762) );
  NOR2_X1 U19687 ( .A1(n16706), .A2(n20488), .ZN(n16813) );
  AOI21_X1 U19688 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16813), .ZN(n16541) );
  OAI21_X1 U19689 ( .B1(n19765), .B2(n16710), .A(n16541), .ZN(n16542) );
  AOI21_X1 U19690 ( .B1(n19762), .B2(n16715), .A(n16542), .ZN(n16545) );
  OAI211_X1 U19691 ( .C1(n16802), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16543), .B(n16697), .ZN(n16544) );
  OAI211_X1 U19692 ( .C1(n16817), .C2(n16680), .A(n16545), .B(n16544), .ZN(
        P2_U2997) );
  XNOR2_X1 U19693 ( .A(n16559), .B(n16825), .ZN(n16552) );
  XNOR2_X1 U19694 ( .A(n16546), .B(n16547), .ZN(n16822) );
  NAND2_X1 U19695 ( .A1(n16822), .A2(n11531), .ZN(n16551) );
  NAND2_X1 U19696 ( .A1(n19788), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16818) );
  NAND2_X1 U19697 ( .A1(n16707), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16548) );
  OAI211_X1 U19698 ( .C1(n16710), .C2(n19779), .A(n16818), .B(n16548), .ZN(
        n16549) );
  AOI21_X1 U19699 ( .B1(n19784), .B2(n16715), .A(n16549), .ZN(n16550) );
  OAI211_X1 U19700 ( .C1(n16712), .C2(n16552), .A(n16551), .B(n16550), .ZN(
        P2_U2998) );
  NAND2_X1 U19701 ( .A1(n16554), .A2(n16553), .ZN(n16556) );
  XOR2_X1 U19702 ( .A(n16556), .B(n16555), .Z(n16838) );
  NOR2_X1 U19703 ( .A1(n16706), .A2(n20485), .ZN(n16827) );
  AOI21_X1 U19704 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16827), .ZN(n16557) );
  OAI21_X1 U19705 ( .B1(n16710), .B2(n16558), .A(n16557), .ZN(n16560) );
  INV_X1 U19706 ( .A(n16839), .ZN(n16885) );
  INV_X1 U19707 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16888) );
  NAND2_X1 U19708 ( .A1(n16563), .A2(n16562), .ZN(n16856) );
  INV_X1 U19709 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20484) );
  NOR2_X1 U19710 ( .A1(n16706), .A2(n20484), .ZN(n16842) );
  AOI21_X1 U19711 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16842), .ZN(n16564) );
  OAI21_X1 U19712 ( .B1(n16565), .B2(n16710), .A(n16564), .ZN(n16571) );
  OR2_X1 U19713 ( .A1(n16566), .A2(n10584), .ZN(n16570) );
  OAI21_X1 U19714 ( .B1(n16856), .B2(n16712), .A(n16572), .ZN(P2_U3000) );
  XNOR2_X1 U19715 ( .A(n16870), .B(n16857), .ZN(n16869) );
  NOR2_X1 U19716 ( .A1(n16706), .A2(n20483), .ZN(n16861) );
  NOR2_X1 U19717 ( .A1(n16672), .A2(n21703), .ZN(n16577) );
  AOI211_X1 U19718 ( .C1(n16578), .C2(n16692), .A(n16861), .B(n16577), .ZN(
        n16579) );
  OAI21_X1 U19719 ( .B1(n16865), .B2(n16695), .A(n16579), .ZN(n16580) );
  AOI21_X1 U19720 ( .B1(n16867), .B2(n11531), .A(n16580), .ZN(n16581) );
  OAI21_X1 U19721 ( .B1(n16869), .B2(n16712), .A(n16581), .ZN(P2_U3001) );
  INV_X1 U19722 ( .A(n16582), .ZN(n16587) );
  AOI21_X1 U19723 ( .B1(n16586), .B2(n16584), .A(n16583), .ZN(n16585) );
  AOI21_X1 U19724 ( .B1(n16587), .B2(n16586), .A(n16585), .ZN(n16883) );
  NAND2_X1 U19725 ( .A1(n16588), .A2(n16875), .ZN(n16871) );
  NAND3_X1 U19726 ( .A1(n16871), .A2(n16697), .A3(n16870), .ZN(n16593) );
  NOR2_X1 U19727 ( .A1(n16706), .A2(n20481), .ZN(n16874) );
  AOI21_X1 U19728 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16874), .ZN(n16589) );
  OAI21_X1 U19729 ( .B1(n16590), .B2(n16710), .A(n16589), .ZN(n16591) );
  AOI21_X1 U19730 ( .B1(n16880), .B2(n16715), .A(n16591), .ZN(n16592) );
  OAI211_X1 U19731 ( .C1(n16883), .C2(n16680), .A(n16593), .B(n16592), .ZN(
        P2_U3002) );
  XNOR2_X1 U19732 ( .A(n16595), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16596) );
  XNOR2_X1 U19733 ( .A(n16594), .B(n16596), .ZN(n16895) );
  NAND2_X1 U19734 ( .A1(n16692), .A2(n16597), .ZN(n16598) );
  NAND2_X1 U19735 ( .A1(n19788), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16887) );
  OAI211_X1 U19736 ( .C1(n21718), .C2(n16672), .A(n16598), .B(n16887), .ZN(
        n16599) );
  AOI21_X1 U19737 ( .B1(n16892), .B2(n16715), .A(n16599), .ZN(n16600) );
  OAI211_X1 U19738 ( .C1(n16895), .C2(n16680), .A(n16601), .B(n16600), .ZN(
        P2_U3003) );
  INV_X1 U19739 ( .A(n16629), .ZN(n16603) );
  OAI21_X1 U19740 ( .B1(n16603), .B2(n16913), .A(n16602), .ZN(n16605) );
  NAND2_X1 U19741 ( .A1(n16605), .A2(n16604), .ZN(n16908) );
  NAND2_X1 U19742 ( .A1(n16668), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16608) );
  NAND2_X1 U19743 ( .A1(n16608), .A2(n16607), .ZN(n16660) );
  AND2_X1 U19744 ( .A1(n16661), .A2(n16660), .ZN(n16622) );
  OAI21_X1 U19745 ( .B1(n16622), .B2(n16610), .A(n16609), .ZN(n16611) );
  NAND2_X1 U19746 ( .A1(n16611), .A2(n16625), .ZN(n16615) );
  NAND2_X1 U19747 ( .A1(n16613), .A2(n16612), .ZN(n16614) );
  XNOR2_X1 U19748 ( .A(n16615), .B(n16614), .ZN(n16906) );
  INV_X1 U19749 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20478) );
  NOR2_X1 U19750 ( .A1(n16706), .A2(n20478), .ZN(n16897) );
  NOR2_X1 U19751 ( .A1(n16710), .A2(n16616), .ZN(n16617) );
  AOI211_X1 U19752 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n16707), .A(
        n16897), .B(n16617), .ZN(n16618) );
  OAI21_X1 U19753 ( .B1(n16896), .B2(n16695), .A(n16618), .ZN(n16619) );
  AOI21_X1 U19754 ( .B1(n16906), .B2(n11531), .A(n16619), .ZN(n16620) );
  OAI21_X1 U19755 ( .B1(n16908), .B2(n16712), .A(n16620), .ZN(P2_U3004) );
  OAI21_X1 U19756 ( .B1(n16653), .B2(n10302), .A(n16624), .ZN(n16628) );
  NAND2_X1 U19757 ( .A1(n16626), .A2(n16625), .ZN(n16627) );
  XNOR2_X1 U19758 ( .A(n16628), .B(n16627), .ZN(n16921) );
  XNOR2_X1 U19759 ( .A(n16629), .B(n16913), .ZN(n16909) );
  NAND2_X1 U19760 ( .A1(n16909), .A2(n16697), .ZN(n16635) );
  NAND2_X1 U19761 ( .A1(n19788), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n16912) );
  OAI21_X1 U19762 ( .B1(n16672), .B2(n16630), .A(n16912), .ZN(n16632) );
  NOR2_X1 U19763 ( .A1(n16915), .A2(n16695), .ZN(n16631) );
  AOI211_X1 U19764 ( .C1(n16692), .C2(n16633), .A(n16632), .B(n16631), .ZN(
        n16634) );
  OAI211_X1 U19765 ( .C1(n16680), .C2(n16921), .A(n16635), .B(n16634), .ZN(
        P2_U3005) );
  XNOR2_X1 U19766 ( .A(n16636), .B(n16637), .ZN(n16934) );
  NAND2_X1 U19767 ( .A1(n16639), .A2(n16638), .ZN(n16640) );
  NOR2_X1 U19768 ( .A1(n16706), .A2(n20474), .ZN(n16923) );
  AOI21_X1 U19769 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16923), .ZN(n16643) );
  NAND2_X1 U19770 ( .A1(n16692), .A2(n16641), .ZN(n16642) );
  OAI211_X1 U19771 ( .C1(n16930), .C2(n16695), .A(n16643), .B(n16642), .ZN(
        n16644) );
  OAI21_X1 U19772 ( .B1(n16712), .B2(n16934), .A(n16645), .ZN(P2_U3006) );
  NAND2_X1 U19773 ( .A1(n16647), .A2(n16646), .ZN(n16648) );
  XNOR2_X1 U19774 ( .A(n16649), .B(n16648), .ZN(n16947) );
  NAND2_X1 U19775 ( .A1(n16651), .A2(n16650), .ZN(n16652) );
  XNOR2_X1 U19776 ( .A(n16653), .B(n16652), .ZN(n16945) );
  NOR2_X1 U19777 ( .A1(n16706), .A2(n16654), .ZN(n16939) );
  AOI21_X1 U19778 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16939), .ZN(n16657) );
  NAND2_X1 U19779 ( .A1(n16692), .A2(n16655), .ZN(n16656) );
  OAI211_X1 U19780 ( .C1(n16942), .C2(n16695), .A(n16657), .B(n16656), .ZN(
        n16658) );
  AOI21_X1 U19781 ( .B1(n16945), .B2(n11531), .A(n16658), .ZN(n16659) );
  OAI21_X1 U19782 ( .B1(n16947), .B2(n16712), .A(n16659), .ZN(P2_U3007) );
  XNOR2_X1 U19783 ( .A(n16661), .B(n16660), .ZN(n16958) );
  INV_X1 U19784 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20471) );
  NOR2_X1 U19785 ( .A1(n16706), .A2(n20471), .ZN(n16949) );
  AOI21_X1 U19786 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16949), .ZN(n16662) );
  OAI21_X1 U19787 ( .B1(n16663), .B2(n16710), .A(n16662), .ZN(n16666) );
  NOR2_X1 U19788 ( .A1(n16953), .A2(n16712), .ZN(n16665) );
  AOI211_X1 U19789 ( .C1(n16715), .C2(n16956), .A(n16666), .B(n16665), .ZN(
        n16667) );
  OAI21_X1 U19790 ( .B1(n16680), .B2(n16958), .A(n16667), .ZN(P2_U3008) );
  XNOR2_X1 U19791 ( .A(n16668), .B(n16966), .ZN(n16669) );
  INV_X1 U19792 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21589) );
  NAND2_X1 U19793 ( .A1(n16692), .A2(n16670), .ZN(n16671) );
  NAND2_X1 U19794 ( .A1(n19788), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n16960) );
  OAI211_X1 U19795 ( .C1(n21589), .C2(n16672), .A(n16671), .B(n16960), .ZN(
        n16678) );
  NAND2_X1 U19796 ( .A1(n16674), .A2(n16673), .ZN(n16675) );
  XOR2_X1 U19797 ( .A(n16676), .B(n16675), .Z(n16967) );
  NOR2_X1 U19798 ( .A1(n16967), .A2(n16712), .ZN(n16677) );
  AOI211_X1 U19799 ( .C1(n16715), .C2(n16971), .A(n16678), .B(n16677), .ZN(
        n16679) );
  OAI21_X1 U19800 ( .B1(n16680), .B2(n16973), .A(n16679), .ZN(P2_U3009) );
  INV_X1 U19801 ( .A(n16681), .ZN(n16702) );
  NAND2_X1 U19802 ( .A1(n16682), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16700) );
  NOR2_X1 U19803 ( .A1(n16682), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16699) );
  AOI21_X1 U19804 ( .B1(n16702), .B2(n16700), .A(n16699), .ZN(n16684) );
  XNOR2_X1 U19805 ( .A(n19792), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16683) );
  XNOR2_X1 U19806 ( .A(n16684), .B(n16683), .ZN(n16982) );
  XNOR2_X1 U19807 ( .A(n16685), .B(n10042), .ZN(n16686) );
  XNOR2_X1 U19808 ( .A(n16687), .B(n16686), .ZN(n16980) );
  NAND2_X1 U19809 ( .A1(n16689), .A2(n16688), .ZN(n16690) );
  NAND2_X1 U19810 ( .A1(n14655), .A2(n16690), .ZN(n19797) );
  NOR2_X1 U19811 ( .A1(n16706), .A2(n16691), .ZN(n16976) );
  AOI21_X1 U19812 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16976), .ZN(n16694) );
  NAND2_X1 U19813 ( .A1(n16692), .A2(n19802), .ZN(n16693) );
  OAI211_X1 U19814 ( .C1(n19797), .C2(n16695), .A(n16694), .B(n16693), .ZN(
        n16696) );
  AOI21_X1 U19815 ( .B1(n16980), .B2(n16697), .A(n16696), .ZN(n16698) );
  OAI21_X1 U19816 ( .B1(n16982), .B2(n16680), .A(n16698), .ZN(P2_U3010) );
  INV_X1 U19817 ( .A(n16699), .ZN(n16701) );
  NAND2_X1 U19818 ( .A1(n16701), .A2(n16700), .ZN(n16703) );
  XNOR2_X1 U19819 ( .A(n16703), .B(n16702), .ZN(n16996) );
  NOR2_X1 U19820 ( .A1(n16706), .A2(n16705), .ZN(n16988) );
  AOI21_X1 U19821 ( .B1(n16707), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16988), .ZN(n16708) );
  OAI21_X1 U19822 ( .B1(n16710), .B2(n16709), .A(n16708), .ZN(n16714) );
  NOR2_X1 U19823 ( .A1(n16983), .A2(n16712), .ZN(n16713) );
  AOI211_X1 U19824 ( .C1(n16715), .C2(n16704), .A(n16714), .B(n16713), .ZN(
        n16716) );
  OAI21_X1 U19825 ( .B1(n16996), .B2(n16680), .A(n16716), .ZN(P2_U3011) );
  OAI211_X1 U19826 ( .C1(n16720), .C2(n16719), .A(n16718), .B(n16717), .ZN(
        n16723) );
  NOR2_X1 U19827 ( .A1(n16721), .A2(n17185), .ZN(n16722) );
  AOI211_X1 U19828 ( .C1(n16989), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        n16727) );
  OAI211_X1 U19829 ( .C1(n16728), .C2(n17182), .A(n16727), .B(n16726), .ZN(
        P2_U3019) );
  NOR2_X1 U19830 ( .A1(n16729), .A2(n16732), .ZN(n16730) );
  AOI211_X1 U19831 ( .C1(n16733), .C2(n16732), .A(n16731), .B(n16730), .ZN(
        n16734) );
  OAI21_X1 U19832 ( .B1(n16735), .B2(n17180), .A(n16734), .ZN(n16738) );
  NOR2_X1 U19833 ( .A1(n16736), .A2(n17185), .ZN(n16737) );
  AOI211_X1 U19834 ( .C1(n16739), .C2(n16993), .A(n16738), .B(n16737), .ZN(
        n16740) );
  OAI21_X1 U19835 ( .B1(n16741), .B2(n17182), .A(n16740), .ZN(P2_U3021) );
  AOI211_X1 U19836 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16744), .A(
        n16743), .B(n16742), .ZN(n16745) );
  OAI21_X1 U19837 ( .B1(n16746), .B2(n17180), .A(n16745), .ZN(n16749) );
  NOR2_X1 U19838 ( .A1(n16747), .A2(n17185), .ZN(n16748) );
  AOI211_X1 U19839 ( .C1(n16750), .C2(n16993), .A(n16749), .B(n16748), .ZN(
        n16751) );
  OAI21_X1 U19840 ( .B1(n16752), .B2(n17182), .A(n16751), .ZN(P2_U3022) );
  NOR2_X1 U19841 ( .A1(n16753), .A2(n17185), .ZN(n16762) );
  INV_X1 U19842 ( .A(n16754), .ZN(n16767) );
  OAI21_X1 U19843 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16755), .ZN(n16756) );
  NOR2_X1 U19844 ( .A1(n16764), .A2(n16756), .ZN(n16757) );
  AOI211_X1 U19845 ( .C1(n16767), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16758), .B(n16757), .ZN(n16759) );
  OAI21_X1 U19846 ( .B1(n16760), .B2(n17180), .A(n16759), .ZN(n16761) );
  NAND2_X1 U19847 ( .A1(n16763), .A2(n16970), .ZN(n16769) );
  NOR2_X1 U19848 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16765) );
  AOI211_X1 U19849 ( .C1(n16767), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16766), .B(n16765), .ZN(n16768) );
  OAI211_X1 U19850 ( .C1(n17180), .C2(n16770), .A(n16769), .B(n16768), .ZN(
        n16771) );
  AOI21_X1 U19851 ( .B1(n16772), .B2(n16944), .A(n16771), .ZN(n16773) );
  INV_X1 U19852 ( .A(n16776), .ZN(n16778) );
  OAI211_X1 U19853 ( .C1(n16780), .C2(n16779), .A(n16778), .B(n16777), .ZN(
        n16781) );
  AOI21_X1 U19854 ( .B1(n16782), .B2(n16989), .A(n16781), .ZN(n16783) );
  OAI21_X1 U19855 ( .B1(n16784), .B2(n17185), .A(n16783), .ZN(n16785) );
  AOI21_X1 U19856 ( .B1(n16786), .B2(n16993), .A(n16785), .ZN(n16787) );
  OAI21_X1 U19857 ( .B1(n16788), .B2(n17182), .A(n16787), .ZN(P2_U3027) );
  INV_X1 U19858 ( .A(n16790), .ZN(n16789) );
  INV_X1 U19859 ( .A(n16844), .ZN(n16914) );
  OAI21_X1 U19860 ( .B1(n16789), .B2(n16810), .A(n16914), .ZN(n16793) );
  NOR3_X1 U19861 ( .A1(n16884), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16790), .ZN(n16791) );
  AOI211_X1 U19862 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16793), .A(
        n16792), .B(n16791), .ZN(n16796) );
  NAND2_X1 U19863 ( .A1(n16794), .A2(n16989), .ZN(n16795) );
  OAI211_X1 U19864 ( .C1(n16797), .C2(n17185), .A(n16796), .B(n16795), .ZN(
        n16798) );
  AOI21_X1 U19865 ( .B1(n16799), .B2(n16993), .A(n16798), .ZN(n16800) );
  OAI21_X1 U19866 ( .B1(n17182), .B2(n16801), .A(n16800), .ZN(P2_U3028) );
  AOI21_X1 U19867 ( .B1(n17193), .B2(n16803), .A(n16802), .ZN(n16809) );
  INV_X1 U19868 ( .A(n16811), .ZN(n16804) );
  AND2_X1 U19869 ( .A1(n17188), .A2(n16804), .ZN(n16805) );
  OR2_X1 U19870 ( .A1(n16844), .A2(n16805), .ZN(n16830) );
  INV_X1 U19871 ( .A(n16806), .ZN(n16807) );
  AND2_X1 U19872 ( .A1(n16807), .A2(n16828), .ZN(n16808) );
  AND2_X1 U19873 ( .A1(n16910), .A2(n16811), .ZN(n16829) );
  AOI21_X1 U19874 ( .B1(n19761), .B2(n16989), .A(n16813), .ZN(n16814) );
  OAI21_X1 U19875 ( .B1(n16815), .B2(n17185), .A(n16814), .ZN(n16816) );
  OAI21_X1 U19876 ( .B1(n16819), .B2(n17180), .A(n16818), .ZN(n16821) );
  NAND2_X1 U19877 ( .A1(n16822), .A2(n16944), .ZN(n16823) );
  OAI211_X1 U19878 ( .C1(n16826), .C2(n16825), .A(n16824), .B(n16823), .ZN(
        P2_U3030) );
  AOI21_X1 U19879 ( .B1(n16829), .B2(n16828), .A(n16827), .ZN(n16832) );
  NAND2_X1 U19880 ( .A1(n16830), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16831) );
  OAI211_X1 U19881 ( .C1(n16833), .C2(n17180), .A(n16832), .B(n16831), .ZN(
        n16835) );
  OAI21_X1 U19882 ( .B1(n16838), .B2(n17182), .A(n16837), .ZN(P2_U3031) );
  NOR2_X1 U19883 ( .A1(n16839), .A2(n16888), .ZN(n16840) );
  NAND2_X1 U19884 ( .A1(n16910), .A2(n16840), .ZN(n16858) );
  INV_X1 U19885 ( .A(n16858), .ZN(n16876) );
  AND2_X1 U19886 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16846) );
  INV_X1 U19887 ( .A(n16846), .ZN(n16841) );
  NOR2_X1 U19888 ( .A1(n16841), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16843) );
  AOI21_X1 U19889 ( .B1(n16876), .B2(n16843), .A(n16842), .ZN(n16849) );
  OR2_X1 U19890 ( .A1(n16844), .A2(n16913), .ZN(n16900) );
  NAND2_X1 U19891 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16845) );
  OAI22_X1 U19892 ( .A1(n16900), .A2(n16845), .B1(n17188), .B2(n16844), .ZN(
        n16872) );
  OR2_X1 U19893 ( .A1(n16858), .A2(n16846), .ZN(n16847) );
  NAND2_X1 U19894 ( .A1(n16872), .A2(n16847), .ZN(n16863) );
  NAND2_X1 U19895 ( .A1(n16863), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16848) );
  OAI211_X1 U19896 ( .C1(n16850), .C2(n17180), .A(n16849), .B(n16848), .ZN(
        n16851) );
  AOI21_X1 U19897 ( .B1(n16852), .B2(n16970), .A(n16851), .ZN(n16855) );
  OR2_X1 U19898 ( .A1(n16853), .A2(n17182), .ZN(n16854) );
  OAI211_X1 U19899 ( .C1(n16856), .C2(n17193), .A(n16855), .B(n16854), .ZN(
        P2_U3032) );
  OAI21_X1 U19900 ( .B1(n16858), .B2(n16875), .A(n16857), .ZN(n16862) );
  NOR2_X1 U19901 ( .A1(n16859), .A2(n17180), .ZN(n16860) );
  AOI211_X1 U19902 ( .C1(n16863), .C2(n16862), .A(n16861), .B(n16860), .ZN(
        n16864) );
  OAI21_X1 U19903 ( .B1(n17185), .B2(n16865), .A(n16864), .ZN(n16866) );
  AOI21_X1 U19904 ( .B1(n16867), .B2(n16944), .A(n16866), .ZN(n16868) );
  OAI21_X1 U19905 ( .B1(n16869), .B2(n17193), .A(n16868), .ZN(P2_U3033) );
  NAND3_X1 U19906 ( .A1(n16871), .A2(n16993), .A3(n16870), .ZN(n16882) );
  NOR2_X1 U19907 ( .A1(n16872), .A2(n16875), .ZN(n16873) );
  AOI211_X1 U19908 ( .C1(n16876), .C2(n16875), .A(n16874), .B(n16873), .ZN(
        n16877) );
  OAI21_X1 U19909 ( .B1(n16878), .B2(n17180), .A(n16877), .ZN(n16879) );
  AOI21_X1 U19910 ( .B1(n16970), .B2(n16880), .A(n16879), .ZN(n16881) );
  OAI211_X1 U19911 ( .C1(n16883), .C2(n17182), .A(n16882), .B(n16881), .ZN(
        P2_U3034) );
  NOR2_X1 U19912 ( .A1(n19837), .A2(n17180), .ZN(n16891) );
  NOR3_X1 U19913 ( .A1(n16884), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16913), .ZN(n16898) );
  AOI21_X1 U19914 ( .B1(n16899), .B2(n16900), .A(n16898), .ZN(n16889) );
  NAND3_X1 U19915 ( .A1(n16910), .A2(n16885), .A3(n16888), .ZN(n16886) );
  OAI211_X1 U19916 ( .C1(n16889), .C2(n16888), .A(n16887), .B(n16886), .ZN(
        n16890) );
  AOI211_X1 U19917 ( .C1(n16892), .C2(n16970), .A(n16891), .B(n16890), .ZN(
        n16893) );
  OAI211_X1 U19918 ( .C1(n16895), .C2(n17182), .A(n16894), .B(n16893), .ZN(
        P2_U3035) );
  NOR2_X1 U19919 ( .A1(n16896), .A2(n17185), .ZN(n16905) );
  NOR2_X1 U19920 ( .A1(n16898), .A2(n16897), .ZN(n16902) );
  NAND3_X1 U19921 ( .A1(n16900), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16899), .ZN(n16901) );
  OAI211_X1 U19922 ( .C1(n16903), .C2(n17180), .A(n16902), .B(n16901), .ZN(
        n16904) );
  AOI211_X1 U19923 ( .C1(n16906), .C2(n16944), .A(n16905), .B(n16904), .ZN(
        n16907) );
  OAI21_X1 U19924 ( .B1(n16908), .B2(n17193), .A(n16907), .ZN(P2_U3036) );
  NAND2_X1 U19925 ( .A1(n16909), .A2(n16993), .ZN(n16920) );
  NAND2_X1 U19926 ( .A1(n16910), .A2(n16913), .ZN(n16911) );
  OAI211_X1 U19927 ( .C1(n16914), .C2(n16913), .A(n16912), .B(n16911), .ZN(
        n16917) );
  NOR2_X1 U19928 ( .A1(n16915), .A2(n17185), .ZN(n16916) );
  AOI211_X1 U19929 ( .C1(n16989), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        n16919) );
  OAI211_X1 U19930 ( .C1(n16921), .C2(n17182), .A(n16920), .B(n16919), .ZN(
        P2_U3037) );
  OAI211_X1 U19931 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16935), .B(n16922), .ZN(n16925) );
  INV_X1 U19932 ( .A(n16923), .ZN(n16924) );
  OAI211_X1 U19933 ( .C1(n9780), .C2(n16926), .A(n16925), .B(n16924), .ZN(
        n16927) );
  AOI21_X1 U19934 ( .B1(n16928), .B2(n16989), .A(n16927), .ZN(n16929) );
  OAI21_X1 U19935 ( .B1(n16930), .B2(n17185), .A(n16929), .ZN(n16931) );
  AOI21_X1 U19936 ( .B1(n16932), .B2(n16944), .A(n16931), .ZN(n16933) );
  OAI21_X1 U19937 ( .B1(n17193), .B2(n16934), .A(n16933), .ZN(P2_U3038) );
  NAND2_X1 U19938 ( .A1(n16935), .A2(n16937), .ZN(n16936) );
  OAI21_X1 U19939 ( .B1(n9780), .B2(n16937), .A(n16936), .ZN(n16938) );
  AOI211_X1 U19940 ( .C1(n16989), .C2(n16940), .A(n16939), .B(n16938), .ZN(
        n16941) );
  OAI21_X1 U19941 ( .B1(n17185), .B2(n16942), .A(n16941), .ZN(n16943) );
  AOI21_X1 U19942 ( .B1(n16945), .B2(n16944), .A(n16943), .ZN(n16946) );
  OAI21_X1 U19943 ( .B1(n16947), .B2(n17193), .A(n16946), .ZN(P2_U3039) );
  INV_X1 U19944 ( .A(n16974), .ZN(n16964) );
  AOI21_X1 U19945 ( .B1(n16964), .B2(n16948), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16952) );
  AOI21_X1 U19946 ( .B1(n16950), .B2(n16989), .A(n16949), .ZN(n16951) );
  OAI21_X1 U19947 ( .B1(n16952), .B2(n9780), .A(n16951), .ZN(n16955) );
  NOR2_X1 U19948 ( .A1(n16953), .A2(n17193), .ZN(n16954) );
  AOI211_X1 U19949 ( .C1(n16956), .C2(n16970), .A(n16955), .B(n16954), .ZN(
        n16957) );
  OAI21_X1 U19950 ( .B1(n17182), .B2(n16958), .A(n16957), .ZN(P2_U3040) );
  INV_X1 U19951 ( .A(n16959), .ZN(n16975) );
  XNOR2_X1 U19952 ( .A(n10042), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16963) );
  OAI21_X1 U19953 ( .B1(n16961), .B2(n17180), .A(n16960), .ZN(n16962) );
  AOI21_X1 U19954 ( .B1(n16964), .B2(n16963), .A(n16962), .ZN(n16965) );
  OAI21_X1 U19955 ( .B1(n16975), .B2(n16966), .A(n16965), .ZN(n16969) );
  NOR2_X1 U19956 ( .A1(n16967), .A2(n17193), .ZN(n16968) );
  AOI211_X1 U19957 ( .C1(n16971), .C2(n16970), .A(n16969), .B(n16968), .ZN(
        n16972) );
  OAI21_X1 U19958 ( .B1(n17182), .B2(n16973), .A(n16972), .ZN(P2_U3041) );
  MUX2_X1 U19959 ( .A(n16975), .B(n16974), .S(n10042), .Z(n16978) );
  AOI21_X1 U19960 ( .B1(n19795), .B2(n16989), .A(n16976), .ZN(n16977) );
  OAI211_X1 U19961 ( .C1(n19797), .C2(n17185), .A(n16978), .B(n16977), .ZN(
        n16979) );
  AOI21_X1 U19962 ( .B1(n16980), .B2(n16993), .A(n16979), .ZN(n16981) );
  OAI21_X1 U19963 ( .B1(n16982), .B2(n17182), .A(n16981), .ZN(P2_U3042) );
  INV_X1 U19964 ( .A(n16983), .ZN(n16994) );
  INV_X1 U19965 ( .A(n16984), .ZN(n16987) );
  MUX2_X1 U19966 ( .A(n16987), .B(n16986), .S(n16985), .Z(n16991) );
  AOI21_X1 U19967 ( .B1(n16989), .B2(n20529), .A(n16988), .ZN(n16990) );
  OAI211_X1 U19968 ( .C1(n17185), .C2(n11180), .A(n16991), .B(n16990), .ZN(
        n16992) );
  AOI21_X1 U19969 ( .B1(n16994), .B2(n16993), .A(n16992), .ZN(n16995) );
  OAI21_X1 U19970 ( .B1(n16996), .B2(n17182), .A(n16995), .ZN(P2_U3043) );
  INV_X1 U19971 ( .A(n16997), .ZN(n16999) );
  INV_X1 U19972 ( .A(n16998), .ZN(n20303) );
  AOI21_X1 U19973 ( .B1(n17000), .B2(n16999), .A(n20303), .ZN(n17001) );
  OAI21_X1 U19974 ( .B1(n17033), .B2(n17002), .A(n17001), .ZN(n17003) );
  MUX2_X1 U19975 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17003), .S(
        n20540), .Z(P2_U3605) );
  INV_X1 U19976 ( .A(n17004), .ZN(n17005) );
  AOI21_X1 U19977 ( .B1(n17005), .B2(n20300), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n17010) );
  INV_X1 U19978 ( .A(n17012), .ZN(n17006) );
  NAND2_X1 U19979 ( .A1(n9682), .A2(n17006), .ZN(n17008) );
  AOI21_X1 U19980 ( .B1(n19778), .B2(n17189), .A(n11127), .ZN(n17007) );
  OAI22_X1 U19981 ( .A1(n17010), .A2(n17026), .B1(n17009), .B2(n17022), .ZN(
        n17011) );
  MUX2_X1 U19982 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17011), .S(
        n17023), .Z(P2_U3601) );
  AND2_X1 U19983 ( .A1(n17013), .A2(n17012), .ZN(n17014) );
  NOR2_X1 U19984 ( .A1(n17015), .A2(n17014), .ZN(n17016) );
  NAND2_X1 U19985 ( .A1(n9682), .A2(n17016), .ZN(n19821) );
  OAI21_X1 U19986 ( .B1(n9682), .B2(n17017), .A(n19821), .ZN(n17025) );
  INV_X1 U19987 ( .A(n17025), .ZN(n17018) );
  AOI22_X1 U19988 ( .A1(n17020), .A2(n17019), .B1(n17018), .B2(n17026), .ZN(
        n17021) );
  OAI21_X1 U19989 ( .B1(n19998), .B2(n17022), .A(n17021), .ZN(n17024) );
  MUX2_X1 U19990 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17024), .S(
        n17023), .Z(P2_U3600) );
  AOI22_X1 U19991 ( .A1(n20537), .A2(n17200), .B1(n17026), .B2(n17025), .ZN(
        n17031) );
  AOI22_X1 U19992 ( .A1(n17028), .A2(n17027), .B1(n21424), .B2(n17030), .ZN(
        n17029) );
  OAI21_X1 U19993 ( .B1(n17031), .B2(n17030), .A(n17029), .ZN(P2_U3599) );
  INV_X1 U19994 ( .A(n20307), .ZN(n17032) );
  OAI21_X1 U19995 ( .B1(n21746), .B2(n19896), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17034) );
  NAND2_X1 U19996 ( .A1(n17034), .A2(n20528), .ZN(n17045) );
  INV_X1 U19997 ( .A(n17045), .ZN(n17037) );
  OR2_X1 U19998 ( .A1(n19960), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19904) );
  NOR2_X1 U19999 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19904), .ZN(
        n19892) );
  INV_X1 U20000 ( .A(n19892), .ZN(n17051) );
  AND2_X1 U20001 ( .A1(n20400), .A2(n17051), .ZN(n17044) );
  OAI21_X1 U20002 ( .B1(n17035), .B2(n19892), .A(n20403), .ZN(n17036) );
  AOI22_X1 U20003 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19894), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19895), .ZN(n21751) );
  INV_X1 U20004 ( .A(n21751), .ZN(n20310) );
  AOI22_X1 U20005 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19894), .ZN(n20356) );
  OAI22_X1 U20006 ( .A1(n20352), .A2(n17051), .B1(n19929), .B2(n20356), .ZN(
        n17041) );
  AOI21_X1 U20007 ( .B1(n21746), .B2(n20310), .A(n17041), .ZN(n17049) );
  OAI21_X1 U20008 ( .B1(n17042), .B2(n19892), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17043) );
  INV_X1 U20009 ( .A(n17046), .ZN(n17047) );
  NOR2_X2 U20010 ( .A1(n19930), .A2(n17047), .ZN(n21743) );
  NAND2_X1 U20011 ( .A1(n19897), .A2(n21743), .ZN(n17048) );
  OAI211_X1 U20012 ( .C1(n19900), .C2(n17050), .A(n17049), .B(n17048), .ZN(
        P2_U3049) );
  AOI22_X2 U20013 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19894), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19895), .ZN(n20420) );
  INV_X1 U20014 ( .A(n20420), .ZN(n20316) );
  AOI22_X1 U20015 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19894), .ZN(n20363) );
  OAI22_X1 U20016 ( .A1(n20362), .A2(n17051), .B1(n19929), .B2(n20363), .ZN(
        n17052) );
  AOI21_X1 U20017 ( .B1(n21746), .B2(n20316), .A(n17052), .ZN(n17055) );
  NOR2_X2 U20018 ( .A1(n19930), .A2(n17053), .ZN(n20416) );
  NAND2_X1 U20019 ( .A1(n19897), .A2(n20416), .ZN(n17054) );
  OAI211_X1 U20020 ( .C1(n19900), .C2(n17056), .A(n17055), .B(n17054), .ZN(
        P2_U3051) );
  INV_X1 U20021 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17771) );
  INV_X1 U20022 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17474) );
  INV_X1 U20023 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17873) );
  INV_X1 U20024 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17960) );
  INV_X1 U20025 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n18001) );
  INV_X1 U20026 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18122) );
  NAND2_X1 U20027 ( .A1(n19105), .A2(n19091), .ZN(n17058) );
  NAND3_X1 U20028 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18124) );
  INV_X1 U20029 ( .A(n18124), .ZN(n17060) );
  NAND4_X1 U20030 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17061), .ZN(n18126) );
  INV_X1 U20031 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18030) );
  NAND2_X1 U20032 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17985), .ZN(n17984) );
  NOR2_X2 U20033 ( .A1(n17960), .A2(n17984), .ZN(n17973) );
  NAND2_X1 U20034 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17973), .ZN(n17958) );
  INV_X2 U20035 ( .A(n17958), .ZN(n17935) );
  NAND3_X1 U20036 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .ZN(n17878) );
  NOR4_X1 U20037 ( .A1(n17474), .A2(n17873), .A3(n17933), .A4(n17878), .ZN(
        n17062) );
  NAND4_X1 U20038 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(n17062), .ZN(n17770) );
  NOR2_X2 U20039 ( .A1(n17771), .A2(n17770), .ZN(n17872) );
  NAND2_X1 U20040 ( .A1(n18143), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17064) );
  NAND2_X1 U20041 ( .A1(n17872), .A2(n19105), .ZN(n17063) );
  OAI22_X1 U20042 ( .A1(n17872), .A2(n17064), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17063), .ZN(P3_U2672) );
  NAND2_X1 U20043 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19289) );
  AOI221_X1 U20044 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19289), .C1(n17066), 
        .C2(n19289), .A(n17065), .ZN(n19070) );
  NOR2_X1 U20045 ( .A1(n17067), .A2(n19553), .ZN(n17068) );
  OAI21_X1 U20046 ( .B1(n17068), .B2(n19067), .A(n19071), .ZN(n19068) );
  AOI22_X1 U20047 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19070), .B1(
        n19068), .B2(n19557), .ZN(P3_U2865) );
  INV_X1 U20048 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17253) );
  INV_X1 U20049 ( .A(n17070), .ZN(n17071) );
  INV_X1 U20050 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18418) );
  NOR2_X1 U20051 ( .A1(n18573), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17074) );
  INV_X1 U20052 ( .A(n17127), .ZN(n17075) );
  NAND2_X1 U20053 ( .A1(n17128), .A2(n17075), .ZN(n17076) );
  XOR2_X1 U20054 ( .A(n17253), .B(n17076), .Z(n17249) );
  NOR2_X1 U20055 ( .A1(n19049), .A2(n19544), .ZN(n18947) );
  INV_X1 U20056 ( .A(n18947), .ZN(n18954) );
  AND2_X1 U20057 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18877), .ZN(
        n18937) );
  NAND2_X1 U20058 ( .A1(n17077), .A2(n18937), .ZN(n18832) );
  NAND2_X1 U20059 ( .A1(n18780), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17083) );
  AOI221_X1 U20060 ( .B1(n18832), .B2(n19546), .C1(n17083), .C2(n19546), .A(
        n17078), .ZN(n17079) );
  OAI221_X1 U20061 ( .B1(n19548), .B2(n18780), .C1(n19548), .C2(n18857), .A(
        n17079), .ZN(n17132) );
  AOI21_X1 U20062 ( .B1(n10746), .B2(n18954), .A(n17132), .ZN(n17264) );
  INV_X1 U20063 ( .A(n18880), .ZN(n17130) );
  NAND2_X1 U20064 ( .A1(n17130), .A2(n18418), .ZN(n17081) );
  NAND3_X1 U20065 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17131) );
  NOR2_X1 U20066 ( .A1(n17131), .A2(n18415), .ZN(n17237) );
  NAND2_X1 U20067 ( .A1(n17261), .A2(n19039), .ZN(n19060) );
  NOR2_X1 U20068 ( .A1(n17262), .A2(n19060), .ZN(n17257) );
  INV_X1 U20069 ( .A(n17257), .ZN(n18969) );
  OAI22_X1 U20070 ( .A1(n17237), .A2(n18969), .B1(n17236), .B2(n19062), .ZN(
        n17080) );
  OAI221_X1 U20071 ( .B1(n19054), .B2(n17264), .C1(n19054), .C2(n17081), .A(
        n17133), .ZN(n17086) );
  NAND2_X1 U20072 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17082) );
  NOR2_X1 U20073 ( .A1(n18416), .A2(n17082), .ZN(n17265) );
  NOR2_X1 U20074 ( .A1(n17082), .A2(n18415), .ZN(n17263) );
  AOI22_X1 U20075 ( .A1(n19021), .A2(n17265), .B1(n17257), .B2(n17263), .ZN(
        n17085) );
  NOR2_X1 U20076 ( .A1(n19054), .A2(n17083), .ZN(n17268) );
  NAND3_X1 U20077 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17268), .A3(
        n17084), .ZN(n17251) );
  NAND2_X1 U20078 ( .A1(n17085), .A2(n17251), .ZN(n17135) );
  AOI22_X1 U20079 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17086), .B1(
        n17135), .B2(n17253), .ZN(n17087) );
  NAND2_X1 U20080 ( .A1(n18963), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17245) );
  OAI211_X1 U20081 ( .C1(n17249), .C2(n18970), .A(n17087), .B(n17245), .ZN(
        P3_U2833) );
  NOR3_X1 U20082 ( .A1(n17089), .A2(n17088), .A3(n21199), .ZN(n17094) );
  AOI211_X1 U20083 ( .C1(n17094), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17091), .B(n17090), .ZN(n17092) );
  INV_X1 U20084 ( .A(n17092), .ZN(n17093) );
  OAI21_X1 U20085 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17094), .A(
        n17093), .ZN(n17095) );
  AOI222_X1 U20086 ( .A1(n17096), .A2(n17095), .B1(n17096), .B2(n21157), .C1(
        n17095), .C2(n21157), .ZN(n17097) );
  AOI222_X1 U20087 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17098), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17097), .C1(n17098), 
        .C2(n17097), .ZN(n17100) );
  AOI21_X1 U20088 ( .B1(n17100), .B2(n20783), .A(n17099), .ZN(n17109) );
  NOR2_X1 U20089 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n17103) );
  OAI22_X1 U20090 ( .A1(n17104), .A2(n17103), .B1(n17102), .B2(n17101), .ZN(
        n17105) );
  NOR2_X1 U20091 ( .A1(n17106), .A2(n17105), .ZN(n17107) );
  NAND3_X1 U20092 ( .A1(n17109), .A2(n17108), .A3(n17107), .ZN(n17118) );
  NAND4_X1 U20093 ( .A1(n17113), .A2(n17112), .A3(n17111), .A4(n17110), .ZN(
        n17116) );
  OAI21_X1 U20094 ( .B1(n17114), .B2(n21409), .A(n21329), .ZN(n17115) );
  NAND2_X1 U20095 ( .A1(n17116), .A2(n17115), .ZN(n17169) );
  AOI21_X1 U20096 ( .B1(n17119), .B2(n17118), .A(n17117), .ZN(n17121) );
  OAI211_X1 U20097 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21409), .A(n17121), 
        .B(n17120), .ZN(n17122) );
  NOR2_X1 U20098 ( .A1(n17175), .A2(n17122), .ZN(n17126) );
  NAND2_X1 U20099 ( .A1(n21413), .A2(n17123), .ZN(n17124) );
  NAND2_X1 U20100 ( .A1(n17176), .A2(n17124), .ZN(n17125) );
  OAI22_X1 U20101 ( .A1(n17126), .A2(n17176), .B1(n17175), .B2(n17125), .ZN(
        P1_U3161) );
  NAND2_X1 U20102 ( .A1(n17213), .A2(n17216), .ZN(n17129) );
  INV_X1 U20103 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17252) );
  XOR2_X1 U20104 ( .A(n17129), .B(n17252), .Z(n17235) );
  NOR2_X1 U20105 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17131), .ZN(
        n17231) );
  OAI211_X1 U20106 ( .C1(n17132), .C2(n17131), .A(n17130), .B(n19039), .ZN(
        n17250) );
  AOI21_X1 U20107 ( .B1(n17133), .B2(n17250), .A(n17252), .ZN(n17134) );
  AOI21_X1 U20108 ( .B1(n17231), .B2(n17135), .A(n17134), .ZN(n17136) );
  NAND2_X1 U20109 ( .A1(n18963), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17225) );
  OAI211_X1 U20110 ( .C1(n17235), .C2(n18970), .A(n17136), .B(n17225), .ZN(
        P3_U2832) );
  INV_X1 U20111 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17350) );
  NOR2_X1 U20112 ( .A1(n20678), .A2(n17350), .ZN(P1_U2905) );
  NOR2_X1 U20113 ( .A1(n17137), .A2(n20540), .ZN(P2_U3047) );
  NAND3_X1 U20114 ( .A1(n19076), .A2(n19715), .A3(n17138), .ZN(n17139) );
  NAND2_X1 U20115 ( .A1(n19105), .A2(n17142), .ZN(n18281) );
  INV_X1 U20116 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18373) );
  NOR2_X1 U20117 ( .A1(n19547), .A2(n18286), .ZN(n18292) );
  AOI22_X1 U20118 ( .A1(n18292), .A2(BUF2_REG_0__SCAN_IN), .B1(n18255), .B2(
        n18762), .ZN(n17141) );
  OAI221_X1 U20119 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n18281), .C1(n18373), 
        .C2(n17142), .A(n17141), .ZN(P3_U2735) );
  AOI22_X1 U20120 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20727), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17148) );
  OAI21_X1 U20121 ( .B1(n17145), .B2(n17144), .A(n17143), .ZN(n17146) );
  INV_X1 U20122 ( .A(n17146), .ZN(n17158) );
  AOI22_X1 U20123 ( .A1(n20652), .A2(n20715), .B1(n20716), .B2(n17158), .ZN(
        n17147) );
  OAI211_X1 U20124 ( .C1(n20720), .C2(n20611), .A(n17148), .B(n17147), .ZN(
        P1_U2994) );
  NAND2_X1 U20125 ( .A1(n17149), .A2(n20725), .ZN(n17161) );
  INV_X1 U20126 ( .A(n14617), .ZN(n17150) );
  AOI21_X1 U20127 ( .B1(n17152), .B2(n17151), .A(n17150), .ZN(n20649) );
  AOI22_X1 U20128 ( .A1(n20649), .A2(n20736), .B1(n20727), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n17160) );
  NOR2_X1 U20129 ( .A1(n20754), .A2(n20768), .ZN(n17153) );
  AND2_X1 U20130 ( .A1(n20725), .A2(n17153), .ZN(n17154) );
  NOR2_X1 U20131 ( .A1(n20723), .A2(n17154), .ZN(n17155) );
  OR2_X1 U20132 ( .A1(n17156), .A2(n17155), .ZN(n17157) );
  AOI22_X1 U20133 ( .A1(n17158), .A2(n20757), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17157), .ZN(n17159) );
  OAI211_X1 U20134 ( .C1(n17161), .C2(n20737), .A(n17160), .B(n17159), .ZN(
        P1_U3026) );
  NAND3_X1 U20135 ( .A1(n17164), .A2(n17163), .A3(n17162), .ZN(n17165) );
  OAI21_X1 U20136 ( .B1(n17166), .B2(n12920), .A(n17165), .ZN(P1_U3468) );
  NAND4_X1 U20137 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21201), .A4(n21409), .ZN(n17167) );
  NAND2_X1 U20138 ( .A1(n17168), .A2(n17167), .ZN(n21328) );
  OAI21_X1 U20139 ( .B1(n17170), .B2(n21328), .A(n17169), .ZN(n17171) );
  OAI221_X1 U20140 ( .B1(n17172), .B2(n21091), .C1(n17172), .C2(n21409), .A(
        n17171), .ZN(n17173) );
  AOI221_X1 U20141 ( .B1(n17175), .B2(n17174), .C1(n17176), .C2(n17174), .A(
        n17173), .ZN(P1_U3162) );
  NOR2_X1 U20142 ( .A1(n17175), .A2(n17176), .ZN(n17178) );
  OAI22_X1 U20143 ( .A1(n21091), .A2(n17178), .B1(n17177), .B2(n17176), .ZN(
        P1_U3466) );
  OAI22_X1 U20144 ( .A1(n17182), .A2(n17181), .B1(n17180), .B2(n17179), .ZN(
        n17187) );
  OAI22_X1 U20145 ( .A1(n17185), .A2(n17184), .B1(n17183), .B2(n17189), .ZN(
        n17186) );
  AOI211_X1 U20146 ( .C1(n17189), .C2(n17188), .A(n17187), .B(n17186), .ZN(
        n17191) );
  OAI211_X1 U20147 ( .C1(n17193), .C2(n17192), .A(n17191), .B(n17190), .ZN(
        P2_U3046) );
  OAI21_X1 U20148 ( .B1(n17196), .B2(n17195), .A(n17194), .ZN(n17197) );
  NOR2_X1 U20149 ( .A1(n17198), .A2(n17197), .ZN(n17205) );
  OAI21_X1 U20150 ( .B1(n17200), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17199), 
        .ZN(n17202) );
  NAND2_X1 U20151 ( .A1(n19859), .A2(n20456), .ZN(n17201) );
  AOI22_X1 U20152 ( .A1(n17203), .A2(n20547), .B1(n17202), .B2(n17201), .ZN(
        n17204) );
  OAI211_X1 U20153 ( .C1(n17206), .C2(n19736), .A(n17205), .B(n17204), .ZN(
        P2_U3176) );
  NAND2_X2 U20154 ( .A1(n19564), .A2(n19711), .ZN(n17364) );
  NOR2_X4 U20155 ( .A1(n18343), .A2(n17364), .ZN(n18756) );
  INV_X1 U20156 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19675) );
  INV_X1 U20157 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17407) );
  INV_X1 U20158 ( .A(n18639), .ZN(n17633) );
  NAND3_X1 U20159 ( .A1(n17633), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17584) );
  NOR2_X2 U20160 ( .A1(n18740), .A2(n18729), .ZN(n17697) );
  INV_X1 U20161 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18638) );
  NOR2_X1 U20162 ( .A1(n18638), .A2(n18703), .ZN(n17207) );
  INV_X1 U20163 ( .A(n18539), .ZN(n17208) );
  NAND2_X1 U20164 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18460) );
  NOR2_X2 U20165 ( .A1(n18451), .A2(n18460), .ZN(n18440) );
  NAND2_X1 U20166 ( .A1(n18440), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18407) );
  NAND2_X1 U20167 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18410) );
  NOR2_X2 U20168 ( .A1(n18407), .A2(n18410), .ZN(n17241) );
  NOR2_X2 U20169 ( .A1(n17209), .A2(n18768), .ZN(n17224) );
  INV_X1 U20170 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19652) );
  NOR2_X1 U20171 ( .A1(n19652), .A2(n19055), .ZN(n17255) );
  NAND2_X1 U20172 ( .A1(n17380), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18773) );
  OR2_X1 U20173 ( .A1(n17209), .A2(n18588), .ZN(n17227) );
  XNOR2_X1 U20174 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17211) );
  NOR2_X1 U20175 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n9690), .ZN(
        n17239) );
  INV_X1 U20176 ( .A(n18773), .ZN(n18613) );
  NAND2_X1 U20177 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17241), .ZN(
        n17387) );
  AOI22_X1 U20178 ( .A1(n19455), .A2(n17209), .B1(n18613), .B2(n17387), .ZN(
        n17210) );
  NAND2_X1 U20179 ( .A1(n17210), .A2(n18772), .ZN(n17240) );
  NOR2_X1 U20180 ( .A1(n17239), .A2(n17240), .ZN(n17226) );
  OAI22_X1 U20181 ( .A1(n17227), .A2(n17211), .B1(n17226), .B2(n17407), .ZN(
        n17212) );
  AOI211_X1 U20182 ( .C1(n18577), .C2(n17723), .A(n17255), .B(n17212), .ZN(
        n17223) );
  AOI21_X1 U20183 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17214), .A(
        n18573), .ZN(n17215) );
  NAND2_X1 U20184 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18573), .ZN(
        n17219) );
  OAI22_X1 U20185 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18573), .B1(
        n17219), .B2(n17252), .ZN(n17218) );
  NAND2_X1 U20186 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17237), .ZN(
        n17221) );
  XOR2_X1 U20187 ( .A(n19675), .B(n17221), .Z(n17258) );
  INV_X1 U20188 ( .A(n17258), .ZN(n17222) );
  INV_X1 U20189 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17412) );
  XNOR2_X1 U20190 ( .A(n17412), .B(n17224), .ZN(n17410) );
  OAI221_X1 U20191 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17227), .C1(
        n17412), .C2(n17226), .A(n17225), .ZN(n17228) );
  AOI21_X1 U20192 ( .B1(n18577), .B2(n17410), .A(n17228), .ZN(n17234) );
  OAI22_X1 U20193 ( .A1(n17236), .A2(n18777), .B1(n17237), .B2(n18620), .ZN(
        n17232) );
  NOR2_X1 U20194 ( .A1(n18859), .A2(n18474), .ZN(n17229) );
  NAND2_X1 U20195 ( .A1(n9779), .A2(n17229), .ZN(n18487) );
  NAND2_X1 U20196 ( .A1(n18887), .A2(n17229), .ZN(n18486) );
  NOR2_X1 U20197 ( .A1(n18805), .A2(n18486), .ZN(n18800) );
  NOR2_X1 U20198 ( .A1(n18469), .A2(n17230), .ZN(n18436) );
  AOI22_X1 U20199 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17232), .B1(
        n18436), .B2(n17231), .ZN(n17233) );
  OAI211_X1 U20200 ( .C1(n17235), .C2(n18687), .A(n17234), .B(n17233), .ZN(
        P3_U2800) );
  NOR2_X1 U20201 ( .A1(n17236), .A2(n18777), .ZN(n17247) );
  NOR2_X1 U20202 ( .A1(n17237), .A2(n18620), .ZN(n17238) );
  OAI21_X1 U20203 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17263), .A(
        n17238), .ZN(n17244) );
  INV_X1 U20204 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17423) );
  AOI21_X1 U20205 ( .B1(n17423), .B2(n17387), .A(n17224), .ZN(n17422) );
  OAI21_X1 U20206 ( .B1(n17239), .B2(n18577), .A(n17422), .ZN(n17243) );
  OAI221_X1 U20207 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17241), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19455), .A(n17240), .ZN(
        n17242) );
  NAND4_X1 U20208 ( .A1(n17245), .A2(n17244), .A3(n17243), .A4(n17242), .ZN(
        n17246) );
  AOI221_X1 U20209 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17247), 
        .C1(n17265), .C2(n17247), .A(n17246), .ZN(n17248) );
  OAI21_X1 U20210 ( .B1(n17249), .B2(n18687), .A(n17248), .ZN(P3_U2801) );
  NOR2_X1 U20211 ( .A1(n19054), .A2(n18880), .ZN(n19048) );
  INV_X1 U20212 ( .A(n19048), .ZN(n18993) );
  OAI211_X1 U20213 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18993), .A(
        n17250), .B(n19053), .ZN(n17256) );
  NOR4_X1 U20214 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17253), .A3(
        n17252), .A4(n17251), .ZN(n17254) );
  AOI211_X1 U20215 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17256), .A(
        n17255), .B(n17254), .ZN(n17259) );
  NAND2_X1 U20216 ( .A1(n18963), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18411) );
  OAI22_X1 U20217 ( .A1(n18418), .A2(n18673), .B1(n18573), .B2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18421) );
  INV_X1 U20218 ( .A(n17261), .ZN(n19515) );
  OAI211_X1 U20219 ( .C1(n17265), .C2(n18820), .A(n19039), .B(n17264), .ZN(
        n17266) );
  NOR3_X1 U20220 ( .A1(n18419), .A2(n18970), .A3(n17267), .ZN(n17269) );
  OAI211_X1 U20221 ( .C1(n17269), .C2(n18829), .A(n17268), .B(n18418), .ZN(
        n17271) );
  NAND3_X1 U20222 ( .A1(n18962), .A2(n18429), .A3(n18421), .ZN(n17270) );
  NOR3_X1 U20223 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17273) );
  NOR4_X1 U20224 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17272) );
  NAND4_X1 U20225 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17273), .A3(n17272), .A4(
        U215), .ZN(U213) );
  INV_X1 U20226 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19841) );
  NOR2_X2 U20227 ( .A1(n17303), .A2(n17274), .ZN(n17318) );
  OAI222_X1 U20228 ( .A1(U212), .A2(n19841), .B1(n17316), .B2(n19890), .C1(
        U214), .C2(n17350), .ZN(U216) );
  AOI222_X1 U20229 ( .A1(n17313), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17318), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17303), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17275) );
  INV_X1 U20230 ( .A(n17275), .ZN(U217) );
  INV_X1 U20231 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n21537) );
  AOI22_X1 U20232 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17313), .ZN(n17276) );
  OAI21_X1 U20233 ( .B1(n21537), .B2(n17316), .A(n17276), .ZN(U218) );
  INV_X1 U20234 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U20235 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17313), .ZN(n17277) );
  OAI21_X1 U20236 ( .B1(n17278), .B2(n17316), .A(n17277), .ZN(U219) );
  INV_X1 U20237 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20238 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17313), .ZN(n17279) );
  OAI21_X1 U20239 ( .B1(n17280), .B2(n17316), .A(n17279), .ZN(U220) );
  AOI222_X1 U20240 ( .A1(n17303), .A2(P1_DATAO_REG_26__SCAN_IN), .B1(n17318), 
        .B2(BUF1_REG_26__SCAN_IN), .C1(n17313), .C2(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n17281) );
  INV_X1 U20241 ( .A(n17281), .ZN(U221) );
  AOI22_X1 U20242 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17313), .ZN(n17282) );
  OAI21_X1 U20243 ( .B1(n15360), .B2(n17316), .A(n17282), .ZN(U222) );
  AOI22_X1 U20244 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17313), .ZN(n17283) );
  OAI21_X1 U20245 ( .B1(n17284), .B2(n17316), .A(n17283), .ZN(U223) );
  INV_X1 U20246 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20247 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17313), .ZN(n17285) );
  OAI21_X1 U20248 ( .B1(n17286), .B2(n17316), .A(n17285), .ZN(U224) );
  INV_X1 U20249 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U20250 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17313), .ZN(n17287) );
  OAI21_X1 U20251 ( .B1(n19885), .B2(n17316), .A(n17287), .ZN(U225) );
  AOI22_X1 U20252 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17313), .ZN(n17288) );
  OAI21_X1 U20253 ( .B1(n17289), .B2(n17316), .A(n17288), .ZN(U226) );
  AOI222_X1 U20254 ( .A1(n17303), .A2(P1_DATAO_REG_20__SCAN_IN), .B1(n17318), 
        .B2(BUF1_REG_20__SCAN_IN), .C1(n17313), .C2(P2_DATAO_REG_20__SCAN_IN), 
        .ZN(n17290) );
  INV_X1 U20255 ( .A(n17290), .ZN(U227) );
  INV_X1 U20256 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20257 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17313), .ZN(n17291) );
  OAI21_X1 U20258 ( .B1(n17292), .B2(n17316), .A(n17291), .ZN(U228) );
  AOI222_X1 U20259 ( .A1(n17303), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n17318), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n17313), .C2(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n17293) );
  INV_X1 U20260 ( .A(n17293), .ZN(U229) );
  INV_X1 U20261 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20262 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17313), .ZN(n17294) );
  OAI21_X1 U20263 ( .B1(n17295), .B2(n17316), .A(n17294), .ZN(U230) );
  AOI22_X1 U20264 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17313), .ZN(n17296) );
  OAI21_X1 U20265 ( .B1(n19865), .B2(n17316), .A(n17296), .ZN(U231) );
  INV_X1 U20266 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n21633) );
  AOI22_X1 U20267 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17318), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17313), .ZN(n17297) );
  OAI21_X1 U20268 ( .B1(n21633), .B2(U214), .A(n17297), .ZN(U232) );
  INV_X1 U20269 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20270 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17303), .ZN(n17298) );
  OAI21_X1 U20271 ( .B1(n17299), .B2(U212), .A(n17298), .ZN(U233) );
  AOI22_X1 U20272 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17313), .ZN(n17300) );
  OAI21_X1 U20273 ( .B1(n17301), .B2(n17316), .A(n17300), .ZN(U234) );
  INV_X1 U20274 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U20275 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n17303), .ZN(n17302) );
  OAI21_X1 U20276 ( .B1(n17331), .B2(U212), .A(n17302), .ZN(U235) );
  AOI22_X1 U20277 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17303), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17313), .ZN(n17304) );
  OAI21_X1 U20278 ( .B1(n17305), .B2(n17316), .A(n17304), .ZN(U236) );
  INV_X1 U20279 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n21545) );
  AOI22_X1 U20280 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n17318), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17313), .ZN(n17306) );
  OAI21_X1 U20281 ( .B1(n21545), .B2(U214), .A(n17306), .ZN(U237) );
  INV_X1 U20282 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20283 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17303), .ZN(n17307) );
  OAI21_X1 U20284 ( .B1(n17328), .B2(U212), .A(n17307), .ZN(U238) );
  INV_X1 U20285 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20286 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n17303), .ZN(n17308) );
  OAI21_X1 U20287 ( .B1(n17309), .B2(U212), .A(n17308), .ZN(U239) );
  INV_X1 U20288 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20289 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17303), .ZN(n17310) );
  OAI21_X1 U20290 ( .B1(n17326), .B2(U212), .A(n17310), .ZN(U240) );
  INV_X1 U20291 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20292 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17303), .ZN(n17311) );
  OAI21_X1 U20293 ( .B1(n17325), .B2(U212), .A(n17311), .ZN(U241) );
  INV_X1 U20294 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n21649) );
  AOI22_X1 U20295 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17318), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17313), .ZN(n17312) );
  OAI21_X1 U20296 ( .B1(n21649), .B2(U214), .A(n17312), .ZN(U242) );
  INV_X1 U20297 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n20673) );
  AOI22_X1 U20298 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n17318), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17313), .ZN(n17314) );
  OAI21_X1 U20299 ( .B1(n20673), .B2(U214), .A(n17314), .ZN(U243) );
  INV_X1 U20300 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17322) );
  INV_X1 U20301 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17315) );
  INV_X1 U20302 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n20675) );
  OAI222_X1 U20303 ( .A1(U212), .A2(n17322), .B1(n17316), .B2(n17315), .C1(
        U214), .C2(n20675), .ZN(U244) );
  INV_X1 U20304 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17321) );
  INV_X1 U20305 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n21699) );
  INV_X1 U20306 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n20677) );
  OAI222_X1 U20307 ( .A1(U212), .A2(n17321), .B1(n17316), .B2(n21699), .C1(
        U214), .C2(n20677), .ZN(U245) );
  AOI22_X1 U20308 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17303), .ZN(n17317) );
  OAI21_X1 U20309 ( .B1(n14236), .B2(U212), .A(n17317), .ZN(U246) );
  AOI22_X1 U20310 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17318), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17303), .ZN(n17319) );
  OAI21_X1 U20311 ( .B1(n17320), .B2(U212), .A(n17319), .ZN(U247) );
  AOI22_X1 U20312 ( .A1(n17349), .A2(n17320), .B1(n14119), .B2(U215), .ZN(U251) );
  AOI22_X1 U20313 ( .A1(n17349), .A2(n14236), .B1(n14088), .B2(U215), .ZN(U252) );
  AOI22_X1 U20314 ( .A1(n17349), .A2(n17321), .B1(n14082), .B2(U215), .ZN(U253) );
  AOI22_X1 U20315 ( .A1(n17349), .A2(n17322), .B1(n14097), .B2(U215), .ZN(U254) );
  OAI22_X1 U20316 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17349), .ZN(n17323) );
  INV_X1 U20317 ( .A(n17323), .ZN(U255) );
  OAI22_X1 U20318 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17349), .ZN(n17324) );
  INV_X1 U20319 ( .A(n17324), .ZN(U256) );
  AOI22_X1 U20320 ( .A1(n17349), .A2(n17325), .B1(n14069), .B2(U215), .ZN(U257) );
  AOI22_X1 U20321 ( .A1(n17338), .A2(n17326), .B1(n14107), .B2(U215), .ZN(U258) );
  OAI22_X1 U20322 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17349), .ZN(n17327) );
  INV_X1 U20323 ( .A(n17327), .ZN(U259) );
  AOI22_X1 U20324 ( .A1(n17338), .A2(n17328), .B1(n14073), .B2(U215), .ZN(U260) );
  OAI22_X1 U20325 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17338), .ZN(n17329) );
  INV_X1 U20326 ( .A(n17329), .ZN(U261) );
  OAI22_X1 U20327 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17338), .ZN(n17330) );
  INV_X1 U20328 ( .A(n17330), .ZN(U262) );
  AOI22_X1 U20329 ( .A1(n17338), .A2(n17331), .B1(n14092), .B2(U215), .ZN(U263) );
  OAI22_X1 U20330 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17338), .ZN(n17332) );
  INV_X1 U20331 ( .A(n17332), .ZN(U264) );
  OAI22_X1 U20332 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17338), .ZN(n17333) );
  INV_X1 U20333 ( .A(n17333), .ZN(U265) );
  OAI22_X1 U20334 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17338), .ZN(n17334) );
  INV_X1 U20335 ( .A(n17334), .ZN(U266) );
  OAI22_X1 U20336 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17349), .ZN(n17335) );
  INV_X1 U20337 ( .A(n17335), .ZN(U267) );
  OAI22_X1 U20338 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17338), .ZN(n17336) );
  INV_X1 U20339 ( .A(n17336), .ZN(U268) );
  AOI22_X1 U20340 ( .A1(n17349), .A2(n21559), .B1(n16457), .B2(U215), .ZN(U269) );
  OAI22_X1 U20341 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17349), .ZN(n17337) );
  INV_X1 U20342 ( .A(n17337), .ZN(U270) );
  AOI22_X1 U20343 ( .A1(n17338), .A2(n21636), .B1(n16440), .B2(U215), .ZN(U271) );
  OAI22_X1 U20344 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17349), .ZN(n17339) );
  INV_X1 U20345 ( .A(n17339), .ZN(U272) );
  OAI22_X1 U20346 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17349), .ZN(n17340) );
  INV_X1 U20347 ( .A(n17340), .ZN(U273) );
  OAI22_X1 U20348 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17349), .ZN(n17341) );
  INV_X1 U20349 ( .A(n17341), .ZN(U274) );
  OAI22_X1 U20350 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17349), .ZN(n17342) );
  INV_X1 U20351 ( .A(n17342), .ZN(U275) );
  OAI22_X1 U20352 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17349), .ZN(n17343) );
  INV_X1 U20353 ( .A(n17343), .ZN(U276) );
  OAI22_X1 U20354 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17349), .ZN(n17344) );
  INV_X1 U20355 ( .A(n17344), .ZN(U277) );
  OAI22_X1 U20356 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17349), .ZN(n17345) );
  INV_X1 U20357 ( .A(n17345), .ZN(U278) );
  OAI22_X1 U20358 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17349), .ZN(n17346) );
  INV_X1 U20359 ( .A(n17346), .ZN(U279) );
  OAI22_X1 U20360 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17349), .ZN(n17347) );
  INV_X1 U20361 ( .A(n17347), .ZN(U280) );
  AOI22_X1 U20362 ( .A1(n17349), .A2(n17348), .B1(n16358), .B2(U215), .ZN(U281) );
  INV_X1 U20363 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n21561) );
  AOI22_X1 U20364 ( .A1(n17349), .A2(n19841), .B1(n21561), .B2(U215), .ZN(U282) );
  INV_X1 U20365 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18301) );
  AOI222_X1 U20366 ( .A1(n17350), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19841), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n18301), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17351) );
  INV_X2 U20367 ( .A(n17351), .ZN(n17353) );
  INV_X2 U20368 ( .A(n17353), .ZN(n17352) );
  INV_X1 U20369 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19615) );
  INV_X1 U20370 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20479) );
  AOI22_X1 U20371 ( .A1(n17352), .A2(n19615), .B1(n20479), .B2(n17353), .ZN(
        U347) );
  INV_X1 U20372 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19613) );
  INV_X1 U20373 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20477) );
  AOI22_X1 U20374 ( .A1(n17352), .A2(n19613), .B1(n20477), .B2(n17353), .ZN(
        U348) );
  INV_X1 U20375 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19610) );
  INV_X1 U20376 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20475) );
  AOI22_X1 U20377 ( .A1(n17352), .A2(n19610), .B1(n20475), .B2(n17353), .ZN(
        U349) );
  INV_X1 U20378 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n21720) );
  INV_X1 U20379 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20473) );
  AOI22_X1 U20380 ( .A1(n17352), .A2(n21720), .B1(n20473), .B2(n17353), .ZN(
        U350) );
  INV_X1 U20381 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19608) );
  INV_X1 U20382 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20472) );
  AOI22_X1 U20383 ( .A1(n17352), .A2(n19608), .B1(n20472), .B2(n17353), .ZN(
        U351) );
  INV_X1 U20384 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19605) );
  INV_X1 U20385 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20470) );
  AOI22_X1 U20386 ( .A1(n17352), .A2(n19605), .B1(n20470), .B2(n17353), .ZN(
        U352) );
  INV_X1 U20387 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n21501) );
  INV_X1 U20388 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20469) );
  AOI22_X1 U20389 ( .A1(n17352), .A2(n21501), .B1(n20469), .B2(n17353), .ZN(
        U353) );
  INV_X1 U20390 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19604) );
  INV_X1 U20391 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20468) );
  AOI22_X1 U20392 ( .A1(n17352), .A2(n19604), .B1(n20468), .B2(n17353), .ZN(
        U354) );
  INV_X1 U20393 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19653) );
  INV_X1 U20394 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20512) );
  AOI22_X1 U20395 ( .A1(n17352), .A2(n19653), .B1(n20512), .B2(n17353), .ZN(
        U355) );
  INV_X1 U20396 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U20397 ( .A1(n17352), .A2(n19650), .B1(n20510), .B2(n17353), .ZN(
        U356) );
  INV_X1 U20398 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19647) );
  INV_X1 U20399 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20509) );
  AOI22_X1 U20400 ( .A1(n17352), .A2(n19647), .B1(n20509), .B2(n17353), .ZN(
        U357) );
  INV_X1 U20401 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19646) );
  INV_X1 U20402 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20507) );
  AOI22_X1 U20403 ( .A1(n17352), .A2(n19646), .B1(n20507), .B2(n17353), .ZN(
        U358) );
  INV_X1 U20404 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19644) );
  INV_X1 U20405 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20506) );
  AOI22_X1 U20406 ( .A1(n17352), .A2(n19644), .B1(n20506), .B2(n17353), .ZN(
        U359) );
  INV_X1 U20407 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19642) );
  INV_X1 U20408 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20504) );
  AOI22_X1 U20409 ( .A1(n17352), .A2(n19642), .B1(n20504), .B2(n17353), .ZN(
        U360) );
  INV_X1 U20410 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19639) );
  INV_X1 U20411 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20502) );
  AOI22_X1 U20412 ( .A1(n17352), .A2(n19639), .B1(n20502), .B2(n17353), .ZN(
        U361) );
  INV_X1 U20413 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19637) );
  INV_X1 U20414 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20500) );
  AOI22_X1 U20415 ( .A1(n17352), .A2(n19637), .B1(n20500), .B2(n17353), .ZN(
        U362) );
  INV_X1 U20416 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19635) );
  INV_X1 U20417 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20498) );
  AOI22_X1 U20418 ( .A1(n17352), .A2(n19635), .B1(n20498), .B2(n17353), .ZN(
        U363) );
  INV_X1 U20419 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19634) );
  INV_X1 U20420 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20496) );
  AOI22_X1 U20421 ( .A1(n17352), .A2(n19634), .B1(n20496), .B2(n17353), .ZN(
        U364) );
  INV_X1 U20422 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19602) );
  INV_X1 U20423 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20467) );
  AOI22_X1 U20424 ( .A1(n17352), .A2(n19602), .B1(n20467), .B2(n17353), .ZN(
        U365) );
  INV_X1 U20425 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19633) );
  INV_X1 U20426 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20494) );
  AOI22_X1 U20427 ( .A1(n17352), .A2(n19633), .B1(n20494), .B2(n17353), .ZN(
        U366) );
  INV_X1 U20428 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19632) );
  INV_X1 U20429 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20492) );
  AOI22_X1 U20430 ( .A1(n17352), .A2(n19632), .B1(n20492), .B2(n17353), .ZN(
        U367) );
  INV_X1 U20431 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19630) );
  INV_X1 U20432 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20491) );
  AOI22_X1 U20433 ( .A1(n17352), .A2(n19630), .B1(n20491), .B2(n17353), .ZN(
        U368) );
  INV_X1 U20434 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19628) );
  INV_X1 U20435 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20489) );
  AOI22_X1 U20436 ( .A1(n17352), .A2(n19628), .B1(n20489), .B2(n17353), .ZN(
        U369) );
  INV_X1 U20437 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19626) );
  INV_X1 U20438 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n21569) );
  AOI22_X1 U20439 ( .A1(n17352), .A2(n19626), .B1(n21569), .B2(n17353), .ZN(
        U370) );
  INV_X1 U20440 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19624) );
  INV_X1 U20441 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20486) );
  AOI22_X1 U20442 ( .A1(n17352), .A2(n19624), .B1(n20486), .B2(n17353), .ZN(
        U371) );
  INV_X1 U20443 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19622) );
  INV_X1 U20444 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n21680) );
  AOI22_X1 U20445 ( .A1(n17351), .A2(n19622), .B1(n21680), .B2(n17353), .ZN(
        U372) );
  INV_X1 U20446 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19620) );
  INV_X1 U20447 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n21553) );
  AOI22_X1 U20448 ( .A1(n17352), .A2(n19620), .B1(n21553), .B2(n17353), .ZN(
        U373) );
  INV_X1 U20449 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19618) );
  INV_X1 U20450 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20482) );
  AOI22_X1 U20451 ( .A1(n17351), .A2(n19618), .B1(n20482), .B2(n17353), .ZN(
        U374) );
  INV_X1 U20452 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19616) );
  INV_X1 U20453 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20480) );
  AOI22_X1 U20454 ( .A1(n17352), .A2(n19616), .B1(n20480), .B2(n17353), .ZN(
        U375) );
  INV_X1 U20455 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19600) );
  INV_X1 U20456 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20466) );
  AOI22_X1 U20457 ( .A1(n17352), .A2(n19600), .B1(n20466), .B2(n17353), .ZN(
        U376) );
  INV_X1 U20458 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n17354) );
  AND2_X1 U20459 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n17354), .ZN(n17355) );
  MUX2_X1 U20460 ( .A(n19598), .B(n17355), .S(P3_STATE_REG_1__SCAN_IN), .Z(
        n19663) );
  AOI21_X1 U20461 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19663), .ZN(n17356) );
  INV_X1 U20462 ( .A(n17356), .ZN(P3_U2633) );
  INV_X1 U20463 ( .A(n17363), .ZN(n17358) );
  OAI21_X1 U20464 ( .B1(n17358), .B2(n18341), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17359) );
  OAI21_X1 U20465 ( .B1(n17360), .B2(n19578), .A(n17359), .ZN(P3_U2634) );
  AOI21_X1 U20466 ( .B1(n17354), .B2(n19598), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17361) );
  AOI22_X1 U20467 ( .A1(n19723), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17361), 
        .B2(n19724), .ZN(P3_U2635) );
  NOR2_X1 U20468 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21421) );
  OAI21_X1 U20469 ( .B1(n21421), .B2(BS16), .A(n19663), .ZN(n19661) );
  OAI21_X1 U20470 ( .B1(n19663), .B2(n19714), .A(n19661), .ZN(P3_U2636) );
  AND3_X1 U20471 ( .A1(n17363), .A2(n19511), .A3(n17362), .ZN(n19516) );
  NOR2_X1 U20472 ( .A1(n19516), .A2(n19573), .ZN(n19708) );
  OAI21_X1 U20473 ( .B1(n19708), .B2(n19065), .A(n17364), .ZN(P3_U2637) );
  NOR4_X1 U20474 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17368) );
  NOR4_X1 U20475 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n17367) );
  NOR4_X1 U20476 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17366) );
  NOR4_X1 U20477 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17365) );
  NAND4_X1 U20478 ( .A1(n17368), .A2(n17367), .A3(n17366), .A4(n17365), .ZN(
        n17374) );
  NOR4_X1 U20479 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_31__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17372) );
  AOI211_X1 U20480 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_8__SCAN_IN), .B(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17371) );
  NOR4_X1 U20481 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17370) );
  NOR4_X1 U20482 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17369) );
  NAND4_X1 U20483 ( .A1(n17372), .A2(n17371), .A3(n17370), .A4(n17369), .ZN(
        n17373) );
  NOR2_X1 U20484 ( .A1(n17374), .A2(n17373), .ZN(n19702) );
  INV_X1 U20485 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17376) );
  NOR3_X1 U20486 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17377) );
  OAI21_X1 U20487 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17377), .A(n19702), .ZN(
        n17375) );
  OAI21_X1 U20488 ( .B1(n19702), .B2(n17376), .A(n17375), .ZN(P3_U2638) );
  INV_X1 U20489 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19698) );
  INV_X1 U20490 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19662) );
  AOI21_X1 U20491 ( .B1(n19698), .B2(n19662), .A(n17377), .ZN(n17379) );
  INV_X1 U20492 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17378) );
  INV_X1 U20493 ( .A(n19702), .ZN(n19705) );
  AOI22_X1 U20494 ( .A1(n19702), .A2(n17379), .B1(n17378), .B2(n19705), .ZN(
        P3_U2639) );
  NAND3_X1 U20495 ( .A1(n17380), .A2(n19575), .A3(n19714), .ZN(n19583) );
  NOR2_X2 U20496 ( .A1(n19676), .A2(n19583), .ZN(n17745) );
  NOR2_X1 U20497 ( .A1(n19040), .A2(n17745), .ZN(n17655) );
  NAND2_X1 U20498 ( .A1(n19575), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19449) );
  OR2_X1 U20499 ( .A1(n19578), .A2(n19449), .ZN(n19571) );
  AOI211_X1 U20500 ( .C1(n19715), .C2(n19713), .A(n19586), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17382) );
  AOI211_X4 U20501 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18343), .A(n17382), .B(
        n17385), .ZN(n17752) );
  INV_X1 U20502 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19654) );
  INV_X1 U20503 ( .A(n17382), .ZN(n19566) );
  INV_X1 U20504 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19641) );
  INV_X1 U20505 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19636) );
  INV_X1 U20506 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21584) );
  INV_X1 U20507 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19631) );
  INV_X1 U20508 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19629) );
  INV_X1 U20509 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19621) );
  INV_X1 U20510 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19619) );
  INV_X1 U20511 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21642) );
  INV_X1 U20512 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19603) );
  NAND2_X1 U20513 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17721) );
  NOR2_X1 U20514 ( .A1(n19603), .A2(n17721), .ZN(n17714) );
  NAND2_X1 U20515 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17714), .ZN(n17698) );
  NOR2_X1 U20516 ( .A1(n19606), .A2(n17698), .ZN(n17669) );
  NAND4_X1 U20517 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17669), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n17635) );
  NAND2_X1 U20518 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n17623) );
  NOR3_X1 U20519 ( .A1(n21642), .A2(n17635), .A3(n17623), .ZN(n17593) );
  NAND2_X1 U20520 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17593), .ZN(n17598) );
  NOR3_X1 U20521 ( .A1(n19621), .A2(n19619), .A3(n17598), .ZN(n17561) );
  NAND4_X1 U20522 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .A4(n17561), .ZN(n17529) );
  NOR3_X1 U20523 ( .A1(n19631), .A2(n19629), .A3(n17529), .ZN(n17523) );
  NAND2_X1 U20524 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17523), .ZN(n17501) );
  NOR2_X1 U20525 ( .A1(n21584), .A2(n17501), .ZN(n17502) );
  NAND2_X1 U20526 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17502), .ZN(n17488) );
  NOR2_X1 U20527 ( .A1(n19636), .A2(n17488), .ZN(n17476) );
  NAND2_X1 U20528 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17476), .ZN(n17466) );
  NOR2_X1 U20529 ( .A1(n19641), .A2(n17466), .ZN(n17453) );
  NAND2_X1 U20530 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17453), .ZN(n17399) );
  NAND4_X1 U20531 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17438), .ZN(n17401) );
  NOR3_X1 U20532 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19654), .A3(n17401), 
        .ZN(n17383) );
  AOI21_X1 U20533 ( .B1(n17752), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17383), .ZN(
        n17406) );
  NAND2_X1 U20534 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18343), .ZN(n17384) );
  AOI211_X4 U20535 ( .C1(n19714), .C2(n19716), .A(n17385), .B(n17384), .ZN(
        n17731) );
  NAND2_X1 U20536 ( .A1(n17737), .A2(n18125), .ZN(n17730) );
  INV_X1 U20537 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18129) );
  NAND2_X1 U20538 ( .A1(n17710), .A2(n18129), .ZN(n17700) );
  INV_X1 U20539 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17682) );
  NAND2_X1 U20540 ( .A1(n17684), .A2(n17682), .ZN(n17679) );
  NOR2_X2 U20541 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17679), .ZN(n17656) );
  INV_X1 U20542 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17649) );
  NAND2_X1 U20543 ( .A1(n17656), .A2(n17649), .ZN(n17647) );
  NOR2_X2 U20544 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17647), .ZN(n17631) );
  NAND2_X1 U20545 ( .A1(n17631), .A2(n18069), .ZN(n17624) );
  INV_X1 U20546 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17604) );
  NAND2_X1 U20547 ( .A1(n17610), .A2(n17604), .ZN(n17603) );
  INV_X1 U20548 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17581) );
  NAND2_X1 U20549 ( .A1(n17585), .A2(n17581), .ZN(n17580) );
  NOR2_X2 U20550 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17580), .ZN(n17565) );
  INV_X1 U20551 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17552) );
  NAND2_X1 U20552 ( .A1(n17565), .A2(n17552), .ZN(n17555) );
  INV_X1 U20553 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17534) );
  NAND2_X1 U20554 ( .A1(n17541), .A2(n17534), .ZN(n17533) );
  INV_X1 U20555 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17514) );
  NAND2_X1 U20556 ( .A1(n17520), .A2(n17514), .ZN(n17513) );
  INV_X1 U20557 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17492) );
  NAND2_X1 U20558 ( .A1(n17496), .A2(n17492), .ZN(n17491) );
  NAND2_X1 U20559 ( .A1(n17463), .A2(n17474), .ZN(n17457) );
  NOR2_X2 U20560 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17457), .ZN(n17456) );
  INV_X1 U20561 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21705) );
  NAND2_X1 U20562 ( .A1(n17456), .A2(n21705), .ZN(n17448) );
  NOR2_X1 U20563 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17448), .ZN(n17432) );
  INV_X1 U20564 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17881) );
  NAND2_X1 U20565 ( .A1(n17432), .A2(n17881), .ZN(n17408) );
  NOR2_X1 U20566 ( .A1(n17763), .A2(n17408), .ZN(n17417) );
  INV_X1 U20567 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18433) );
  NAND3_X1 U20568 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17386), .A3(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17391) );
  NOR2_X1 U20569 ( .A1(n18460), .A2(n17391), .ZN(n18408) );
  NAND2_X1 U20570 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18408), .ZN(
        n17398) );
  NOR2_X1 U20571 ( .A1(n18433), .A2(n17398), .ZN(n17388) );
  OAI21_X1 U20572 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17388), .A(
        n17387), .ZN(n18413) );
  INV_X1 U20573 ( .A(n18413), .ZN(n17435) );
  AOI21_X1 U20574 ( .B1(n18433), .B2(n17398), .A(n17388), .ZN(n18427) );
  INV_X1 U20575 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17390) );
  INV_X1 U20576 ( .A(n17391), .ZN(n18452) );
  NAND2_X1 U20577 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18452), .ZN(
        n17389) );
  AOI21_X1 U20578 ( .B1(n17390), .B2(n17389), .A(n18408), .ZN(n18453) );
  INV_X1 U20579 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21686) );
  OAI22_X1 U20580 ( .A1(n21686), .A2(n18452), .B1(n17391), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18464) );
  AOI21_X1 U20581 ( .B1(n17386), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18482) );
  NOR2_X1 U20582 ( .A1(n18452), .A2(n18482), .ZN(n18485) );
  INV_X1 U20583 ( .A(n17386), .ZN(n18480) );
  NOR2_X1 U20584 ( .A1(n18768), .A2(n9782), .ZN(n17393) );
  OAI22_X1 U20585 ( .A1(n18768), .A2(n18480), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17393), .ZN(n17392) );
  INV_X1 U20586 ( .A(n17392), .ZN(n18500) );
  NAND2_X1 U20587 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18496), .ZN(
        n17394) );
  AOI21_X1 U20588 ( .B1(n10690), .B2(n17394), .A(n17393), .ZN(n18512) );
  NOR3_X1 U20589 ( .A1(n18768), .A2(n18564), .A3(n18565), .ZN(n18537) );
  NAND3_X1 U20590 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n18537), .ZN(n18494) );
  AOI22_X1 U20591 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18496), .B1(
        n21610), .B2(n18494), .ZN(n18522) );
  INV_X1 U20592 ( .A(n18494), .ZN(n17397) );
  INV_X1 U20593 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18592) );
  NOR2_X1 U20594 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18768), .ZN(
        n17746) );
  NAND2_X1 U20595 ( .A1(n17395), .A2(n17746), .ZN(n17574) );
  NOR2_X1 U20596 ( .A1(n18592), .A2(n17574), .ZN(n17562) );
  NOR2_X1 U20597 ( .A1(n18522), .A2(n17519), .ZN(n17518) );
  NOR2_X1 U20598 ( .A1(n17518), .A2(n17696), .ZN(n17508) );
  NOR2_X1 U20599 ( .A1(n18512), .A2(n17508), .ZN(n17507) );
  NOR2_X1 U20600 ( .A1(n17507), .A2(n17696), .ZN(n17498) );
  NOR2_X1 U20601 ( .A1(n18500), .A2(n17498), .ZN(n17497) );
  NOR2_X1 U20602 ( .A1(n17497), .A2(n17696), .ZN(n17486) );
  NOR2_X1 U20603 ( .A1(n18485), .A2(n17486), .ZN(n17485) );
  NOR2_X1 U20604 ( .A1(n17485), .A2(n17696), .ZN(n17479) );
  NOR2_X1 U20605 ( .A1(n18464), .A2(n17479), .ZN(n17478) );
  NOR2_X1 U20606 ( .A1(n17478), .A2(n17696), .ZN(n17465) );
  NOR2_X1 U20607 ( .A1(n18453), .A2(n17465), .ZN(n17464) );
  OAI21_X1 U20608 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18408), .A(
        n17398), .ZN(n18443) );
  AOI21_X1 U20609 ( .B1(n17464), .B2(n18443), .A(n17696), .ZN(n17444) );
  NOR2_X1 U20610 ( .A1(n18427), .A2(n17444), .ZN(n17443) );
  NOR2_X1 U20611 ( .A1(n17443), .A2(n17696), .ZN(n17434) );
  NOR2_X1 U20612 ( .A1(n17435), .A2(n17434), .ZN(n17433) );
  NOR2_X1 U20613 ( .A1(n17433), .A2(n17696), .ZN(n17421) );
  NOR2_X1 U20614 ( .A1(n17422), .A2(n17421), .ZN(n17420) );
  NOR2_X1 U20615 ( .A1(n17420), .A2(n17696), .ZN(n17409) );
  NAND2_X1 U20616 ( .A1(n17723), .A2(n17745), .ZN(n17754) );
  NOR3_X1 U20617 ( .A1(n17410), .A2(n17409), .A3(n17754), .ZN(n17404) );
  NAND3_X1 U20618 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n17400) );
  AND2_X1 U20619 ( .A1(n17736), .A2(n17399), .ZN(n17452) );
  NOR2_X1 U20620 ( .A1(n17751), .A2(n17452), .ZN(n17451) );
  INV_X1 U20621 ( .A(n17451), .ZN(n17460) );
  AOI21_X1 U20622 ( .B1(n17736), .B2(n17400), .A(n17460), .ZN(n17431) );
  NOR2_X1 U20623 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17401), .ZN(n17413) );
  INV_X1 U20624 ( .A(n17413), .ZN(n17402) );
  AOI21_X1 U20625 ( .B1(n17431), .B2(n17402), .A(n19652), .ZN(n17403) );
  OAI211_X1 U20626 ( .C1(n17407), .C2(n17753), .A(n17406), .B(n17405), .ZN(
        P3_U2640) );
  NAND2_X1 U20627 ( .A1(n17731), .A2(n17408), .ZN(n17427) );
  INV_X1 U20628 ( .A(n17409), .ZN(n17411) );
  OAI22_X1 U20629 ( .A1(n17431), .A2(n19654), .B1(n17412), .B2(n17753), .ZN(
        n17414) );
  OAI21_X1 U20630 ( .B1(n17752), .B2(n17417), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17418) );
  OAI211_X1 U20631 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17427), .A(n17419), .B(
        n17418), .ZN(P3_U2641) );
  INV_X1 U20632 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19649) );
  AOI211_X1 U20633 ( .C1(n17422), .C2(n17421), .A(n17420), .B(n19581), .ZN(
        n17426) );
  NAND3_X1 U20634 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17438), .ZN(n17424) );
  OAI22_X1 U20635 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17424), .B1(n17423), 
        .B2(n17753), .ZN(n17425) );
  AOI211_X1 U20636 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17752), .A(n17426), .B(
        n17425), .ZN(n17430) );
  INV_X1 U20637 ( .A(n17427), .ZN(n17428) );
  OAI21_X1 U20638 ( .B1(n17432), .B2(n17881), .A(n17428), .ZN(n17429) );
  OAI211_X1 U20639 ( .C1(n17431), .C2(n19649), .A(n17430), .B(n17429), .ZN(
        P3_U2642) );
  AOI22_X1 U20640 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17715), .B1(
        n17752), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17442) );
  AOI211_X1 U20641 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17448), .A(n17432), .B(
        n17763), .ZN(n17437) );
  AOI211_X1 U20642 ( .C1(n17435), .C2(n17434), .A(n17433), .B(n19581), .ZN(
        n17436) );
  NOR2_X1 U20643 ( .A1(n17437), .A2(n17436), .ZN(n17441) );
  INV_X1 U20644 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19645) );
  AND2_X1 U20645 ( .A1(n19645), .A2(n17438), .ZN(n17447) );
  OAI21_X1 U20646 ( .B1(n17447), .B2(n17460), .A(P3_REIP_REG_28__SCAN_IN), 
        .ZN(n17440) );
  INV_X1 U20647 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21470) );
  NAND3_X1 U20648 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17438), .A3(n21470), 
        .ZN(n17439) );
  NAND4_X1 U20649 ( .A1(n17442), .A2(n17441), .A3(n17440), .A4(n17439), .ZN(
        P3_U2643) );
  AOI211_X1 U20650 ( .C1(n18427), .C2(n17444), .A(n17443), .B(n19581), .ZN(
        n17446) );
  OAI22_X1 U20651 ( .A1(n18433), .A2(n17753), .B1(n17764), .B2(n21705), .ZN(
        n17445) );
  NOR3_X1 U20652 ( .A1(n17447), .A2(n17446), .A3(n17445), .ZN(n17450) );
  OAI211_X1 U20653 ( .C1(n17456), .C2(n21705), .A(n17731), .B(n17448), .ZN(
        n17449) );
  OAI211_X1 U20654 ( .C1(n17451), .C2(n19645), .A(n17450), .B(n17449), .ZN(
        P3_U2644) );
  INV_X1 U20655 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21556) );
  AOI22_X1 U20656 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17715), .B1(
        n17453), .B2(n17452), .ZN(n17462) );
  OR2_X1 U20657 ( .A1(n17696), .A2(n17464), .ZN(n17455) );
  OAI21_X1 U20658 ( .B1(n18443), .B2(n17455), .A(n17745), .ZN(n17454) );
  AOI21_X1 U20659 ( .B1(n18443), .B2(n17455), .A(n17454), .ZN(n17459) );
  AOI211_X1 U20660 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17457), .A(n17456), .B(
        n17763), .ZN(n17458) );
  AOI211_X1 U20661 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17460), .A(n17459), 
        .B(n17458), .ZN(n17461) );
  OAI211_X1 U20662 ( .C1(n17764), .C2(n21556), .A(n17462), .B(n17461), .ZN(
        P3_U2645) );
  OR2_X1 U20663 ( .A1(n17763), .A2(n17463), .ZN(n17477) );
  AOI21_X1 U20664 ( .B1(n17731), .B2(n17463), .A(n17752), .ZN(n17473) );
  AOI211_X1 U20665 ( .C1(n18453), .C2(n17465), .A(n17464), .B(n19581), .ZN(
        n17471) );
  NOR2_X1 U20666 ( .A1(n17757), .A2(n17466), .ZN(n17469) );
  INV_X1 U20667 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19640) );
  OAI21_X1 U20668 ( .B1(n17476), .B2(n17757), .A(n17767), .ZN(n17484) );
  AOI21_X1 U20669 ( .B1(n17736), .B2(n19640), .A(n17484), .ZN(n17467) );
  INV_X1 U20670 ( .A(n17467), .ZN(n17468) );
  MUX2_X1 U20671 ( .A(n17469), .B(n17468), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n17470) );
  AOI211_X1 U20672 ( .C1(n17715), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17471), .B(n17470), .ZN(n17472) );
  OAI221_X1 U20673 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17477), .C1(n17474), 
        .C2(n17473), .A(n17472), .ZN(P3_U2646) );
  NOR2_X1 U20674 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17757), .ZN(n17475) );
  AOI22_X1 U20675 ( .A1(n17752), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17476), 
        .B2(n17475), .ZN(n17483) );
  AOI21_X1 U20676 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17491), .A(n17477), .ZN(
        n17481) );
  AOI211_X1 U20677 ( .C1(n18464), .C2(n17479), .A(n17478), .B(n19581), .ZN(
        n17480) );
  AOI211_X1 U20678 ( .C1(n17484), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17481), 
        .B(n17480), .ZN(n17482) );
  OAI211_X1 U20679 ( .C1(n21686), .C2(n17753), .A(n17483), .B(n17482), .ZN(
        P3_U2647) );
  INV_X1 U20680 ( .A(n17484), .ZN(n17495) );
  AOI211_X1 U20681 ( .C1(n18485), .C2(n17486), .A(n17485), .B(n19581), .ZN(
        n17490) );
  NAND2_X1 U20682 ( .A1(n17736), .A2(n19636), .ZN(n17487) );
  OAI22_X1 U20683 ( .A1(n17764), .A2(n17492), .B1(n17488), .B2(n17487), .ZN(
        n17489) );
  AOI211_X1 U20684 ( .C1(n17715), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17490), .B(n17489), .ZN(n17494) );
  OAI211_X1 U20685 ( .C1(n17496), .C2(n17492), .A(n17731), .B(n17491), .ZN(
        n17493) );
  OAI211_X1 U20686 ( .C1(n17495), .C2(n19636), .A(n17494), .B(n17493), .ZN(
        P3_U2648) );
  AOI22_X1 U20687 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17715), .B1(
        n17752), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n17506) );
  AOI211_X1 U20688 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17513), .A(n17496), .B(
        n17763), .ZN(n17500) );
  AOI211_X1 U20689 ( .C1(n18500), .C2(n17498), .A(n17497), .B(n19581), .ZN(
        n17499) );
  NOR2_X1 U20690 ( .A1(n17500), .A2(n17499), .ZN(n17505) );
  NOR3_X1 U20691 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17757), .A3(n17501), 
        .ZN(n17512) );
  AND2_X1 U20692 ( .A1(n17736), .A2(n17501), .ZN(n17524) );
  NOR2_X1 U20693 ( .A1(n17751), .A2(n17524), .ZN(n17527) );
  INV_X1 U20694 ( .A(n17527), .ZN(n17511) );
  OAI21_X1 U20695 ( .B1(n17512), .B2(n17511), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n17504) );
  INV_X1 U20696 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21609) );
  NAND3_X1 U20697 ( .A1(n17736), .A2(n17502), .A3(n21609), .ZN(n17503) );
  NAND4_X1 U20698 ( .A1(n17506), .A2(n17505), .A3(n17504), .A4(n17503), .ZN(
        P3_U2649) );
  AOI211_X1 U20699 ( .C1(n18512), .C2(n17508), .A(n17507), .B(n19581), .ZN(
        n17510) );
  OAI22_X1 U20700 ( .A1(n10690), .A2(n17753), .B1(n17764), .B2(n17514), .ZN(
        n17509) );
  AOI211_X1 U20701 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n17511), .A(n17510), 
        .B(n17509), .ZN(n17517) );
  INV_X1 U20702 ( .A(n17512), .ZN(n17516) );
  OAI211_X1 U20703 ( .C1(n17520), .C2(n17514), .A(n17731), .B(n17513), .ZN(
        n17515) );
  NAND3_X1 U20704 ( .A1(n17517), .A2(n17516), .A3(n17515), .ZN(P3_U2650) );
  INV_X1 U20705 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21658) );
  AOI22_X1 U20706 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17715), .B1(
        n17752), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n17526) );
  AOI211_X1 U20707 ( .C1(n18522), .C2(n17519), .A(n17518), .B(n19581), .ZN(
        n17522) );
  AOI211_X1 U20708 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17533), .A(n17520), .B(
        n17763), .ZN(n17521) );
  AOI211_X1 U20709 ( .C1(n17524), .C2(n17523), .A(n17522), .B(n17521), .ZN(
        n17525) );
  OAI211_X1 U20710 ( .C1(n17527), .C2(n21658), .A(n17526), .B(n17525), .ZN(
        P3_U2651) );
  AOI22_X1 U20711 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17715), .B1(
        n17752), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17537) );
  INV_X1 U20712 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18553) );
  INV_X1 U20713 ( .A(n18537), .ZN(n17549) );
  NOR2_X1 U20714 ( .A1(n18553), .A2(n17549), .ZN(n17528) );
  OAI21_X1 U20715 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17528), .A(
        n18494), .ZN(n18541) );
  INV_X1 U20716 ( .A(n17562), .ZN(n17548) );
  INV_X1 U20717 ( .A(n17528), .ZN(n17538) );
  OAI21_X1 U20718 ( .B1(n17548), .B2(n17538), .A(n17723), .ZN(n17540) );
  XOR2_X1 U20719 ( .A(n18541), .B(n17540), .Z(n17532) );
  INV_X1 U20720 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19625) );
  NOR4_X1 U20721 ( .A1(n17757), .A2(n19621), .A3(n19619), .A4(n17598), .ZN(
        n17572) );
  NAND2_X1 U20722 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17572), .ZN(n17571) );
  NOR2_X1 U20723 ( .A1(n19625), .A2(n17571), .ZN(n17547) );
  NAND2_X1 U20724 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17547), .ZN(n17546) );
  XOR2_X1 U20725 ( .A(P3_REIP_REG_19__SCAN_IN), .B(n19629), .Z(n17530) );
  AOI21_X1 U20726 ( .B1(n17736), .B2(n17529), .A(n17751), .ZN(n17559) );
  OAI22_X1 U20727 ( .A1(n17546), .A2(n17530), .B1(n19631), .B2(n17559), .ZN(
        n17531) );
  AOI21_X1 U20728 ( .B1(n17532), .B2(n17745), .A(n17531), .ZN(n17536) );
  OAI211_X1 U20729 ( .C1(n17541), .C2(n17534), .A(n17731), .B(n17533), .ZN(
        n17535) );
  NAND4_X1 U20730 ( .A1(n17537), .A2(n17536), .A3(n19055), .A4(n17535), .ZN(
        P3_U2652) );
  OAI21_X1 U20731 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18537), .A(
        n17538), .ZN(n18550) );
  NAND2_X1 U20732 ( .A1(n17745), .A2(n17696), .ZN(n17741) );
  OAI221_X1 U20733 ( .B1(n18550), .B2(n17562), .C1(n18550), .C2(n18553), .A(
        n17745), .ZN(n17539) );
  AOI22_X1 U20734 ( .A1(n17540), .A2(n18550), .B1(n17741), .B2(n17539), .ZN(
        n17544) );
  AOI211_X1 U20735 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17555), .A(n17541), .B(
        n17763), .ZN(n17543) );
  OAI22_X1 U20736 ( .A1(n18553), .A2(n17753), .B1(n17764), .B2(n17960), .ZN(
        n17542) );
  NOR4_X1 U20737 ( .A1(n19040), .A2(n17544), .A3(n17543), .A4(n17542), .ZN(
        n17545) );
  OAI221_X1 U20738 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17546), .C1(n19629), 
        .C2(n17559), .A(n17545), .ZN(P3_U2653) );
  NOR2_X1 U20739 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17547), .ZN(n17560) );
  AOI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17715), .A(
        n19040), .ZN(n17558) );
  INV_X1 U20741 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17566) );
  INV_X1 U20742 ( .A(n17395), .ZN(n18587) );
  NOR2_X1 U20743 ( .A1(n18768), .A2(n18587), .ZN(n18575) );
  NAND2_X1 U20744 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18575), .ZN(
        n17573) );
  NOR2_X1 U20745 ( .A1(n18768), .A2(n18564), .ZN(n17550) );
  AOI21_X1 U20746 ( .B1(n17566), .B2(n17573), .A(n17550), .ZN(n18576) );
  OAI21_X1 U20747 ( .B1(n17548), .B2(n18576), .A(n17723), .ZN(n17551) );
  OAI21_X1 U20748 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17550), .A(
        n17549), .ZN(n18568) );
  XOR2_X1 U20749 ( .A(n17551), .B(n18568), .Z(n17556) );
  NOR2_X1 U20750 ( .A1(n17565), .A2(n17552), .ZN(n17553) );
  OAI22_X1 U20751 ( .A1(n17763), .A2(n17553), .B1(n17764), .B2(n17552), .ZN(
        n17554) );
  AOI22_X1 U20752 ( .A1(n17556), .A2(n17745), .B1(n17555), .B2(n17554), .ZN(
        n17557) );
  OAI211_X1 U20753 ( .C1(n17560), .C2(n17559), .A(n17558), .B(n17557), .ZN(
        P3_U2654) );
  INV_X1 U20754 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19623) );
  NAND2_X1 U20755 ( .A1(n17561), .A2(n17767), .ZN(n17586) );
  NAND2_X1 U20756 ( .A1(n17757), .A2(n17767), .ZN(n17765) );
  OAI21_X1 U20757 ( .B1(n19623), .B2(n17586), .A(n17765), .ZN(n17577) );
  NOR2_X1 U20758 ( .A1(n17562), .A2(n17696), .ZN(n17564) );
  NOR2_X1 U20759 ( .A1(n18576), .A2(n17564), .ZN(n17563) );
  AOI211_X1 U20760 ( .C1(n18576), .C2(n17564), .A(n17563), .B(n19581), .ZN(
        n17569) );
  AOI211_X1 U20761 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17580), .A(n17565), .B(
        n17763), .ZN(n17568) );
  OAI22_X1 U20762 ( .A1(n17566), .A2(n17753), .B1(n17764), .B2(n18001), .ZN(
        n17567) );
  NOR4_X1 U20763 ( .A1(n19040), .A2(n17569), .A3(n17568), .A4(n17567), .ZN(
        n17570) );
  OAI221_X1 U20764 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n17571), .C1(n19625), 
        .C2(n17577), .A(n17570), .ZN(P3_U2655) );
  NOR2_X1 U20765 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17572), .ZN(n17578) );
  OAI21_X1 U20766 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18575), .A(
        n17573), .ZN(n18589) );
  NAND2_X1 U20767 ( .A1(n17723), .A2(n17574), .ZN(n17575) );
  XNOR2_X1 U20768 ( .A(n18589), .B(n17575), .ZN(n17576) );
  OAI22_X1 U20769 ( .A1(n17578), .A2(n17577), .B1(n19581), .B2(n17576), .ZN(
        n17579) );
  AOI211_X1 U20770 ( .C1(n17752), .C2(P3_EBX_REG_15__SCAN_IN), .A(n19040), .B(
        n17579), .ZN(n17583) );
  OAI211_X1 U20771 ( .C1(n17585), .C2(n17581), .A(n17731), .B(n17580), .ZN(
        n17582) );
  OAI211_X1 U20772 ( .C1(n17753), .C2(n18592), .A(n17583), .B(n17582), .ZN(
        P3_U2656) );
  INV_X1 U20773 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17607) );
  INV_X1 U20774 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17755) );
  INV_X1 U20775 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n21679) );
  INV_X1 U20776 ( .A(n17659), .ZN(n18675) );
  NAND2_X1 U20777 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18675), .ZN(
        n17685) );
  NOR2_X1 U20778 ( .A1(n17584), .A2(n17685), .ZN(n17620) );
  INV_X1 U20779 ( .A(n17620), .ZN(n18612) );
  NOR2_X1 U20780 ( .A1(n21679), .A2(n18612), .ZN(n17608) );
  NAND2_X1 U20781 ( .A1(n17755), .A2(n17608), .ZN(n17595) );
  OAI21_X1 U20782 ( .B1(n17607), .B2(n17595), .A(n17723), .ZN(n17597) );
  NAND3_X1 U20783 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(n17620), .ZN(n17594) );
  AOI21_X1 U20784 ( .B1(n18602), .B2(n17594), .A(n18575), .ZN(n18604) );
  XOR2_X1 U20785 ( .A(n17597), .B(n18604), .Z(n17592) );
  AOI211_X1 U20786 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17603), .A(n17585), .B(
        n17763), .ZN(n17590) );
  NOR3_X1 U20787 ( .A1(n17757), .A2(n19619), .A3(n17598), .ZN(n17587) );
  OAI211_X1 U20788 ( .C1(n17587), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17765), 
        .B(n17586), .ZN(n17588) );
  OAI211_X1 U20789 ( .C1(n17764), .C2(n18030), .A(n19055), .B(n17588), .ZN(
        n17589) );
  AOI211_X1 U20790 ( .C1(n17715), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17590), .B(n17589), .ZN(n17591) );
  OAI21_X1 U20791 ( .B1(n19581), .B2(n17592), .A(n17591), .ZN(P3_U2657) );
  INV_X1 U20792 ( .A(n17593), .ZN(n17615) );
  AOI21_X1 U20793 ( .B1(n17736), .B2(n17615), .A(n17751), .ZN(n17622) );
  INV_X1 U20794 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19617) );
  NAND2_X1 U20795 ( .A1(n17736), .A2(n19617), .ZN(n17614) );
  AOI21_X1 U20796 ( .B1(n17622), .B2(n17614), .A(n19619), .ZN(n17602) );
  OAI21_X1 U20797 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17608), .A(
        n17594), .ZN(n18615) );
  INV_X1 U20798 ( .A(n17595), .ZN(n17609) );
  OAI21_X1 U20799 ( .B1(n17609), .B2(n18615), .A(n17745), .ZN(n17596) );
  AOI22_X1 U20800 ( .A1(n18615), .A2(n17597), .B1(n17741), .B2(n17596), .ZN(
        n17601) );
  OR2_X1 U20801 ( .A1(n17757), .A2(n17598), .ZN(n17599) );
  OAI22_X1 U20802 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17599), .B1(n17764), 
        .B2(n17604), .ZN(n17600) );
  NOR4_X1 U20803 ( .A1(n19040), .A2(n17602), .A3(n17601), .A4(n17600), .ZN(
        n17606) );
  OAI211_X1 U20804 ( .C1(n17610), .C2(n17604), .A(n17731), .B(n17603), .ZN(
        n17605) );
  OAI211_X1 U20805 ( .C1(n17753), .C2(n17607), .A(n17606), .B(n17605), .ZN(
        P3_U2658) );
  AOI21_X1 U20806 ( .B1(n21679), .B2(n18612), .A(n17608), .ZN(n17613) );
  NOR3_X1 U20807 ( .A1(n17613), .A2(n17609), .A3(n17754), .ZN(n17612) );
  AOI211_X1 U20808 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17624), .A(n17610), .B(
        n17763), .ZN(n17611) );
  AOI211_X1 U20809 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17752), .A(n17612), .B(
        n17611), .ZN(n17619) );
  AOI21_X1 U20810 ( .B1(n17723), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19581), .ZN(n17760) );
  INV_X1 U20811 ( .A(n17613), .ZN(n18625) );
  AOI21_X1 U20812 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17723), .A(
        n18625), .ZN(n17617) );
  OAI22_X1 U20813 ( .A1(n21679), .A2(n17753), .B1(n17615), .B2(n17614), .ZN(
        n17616) );
  AOI211_X1 U20814 ( .C1(n17760), .C2(n17617), .A(n18963), .B(n17616), .ZN(
        n17618) );
  OAI211_X1 U20815 ( .C1(n19617), .C2(n17622), .A(n17619), .B(n17618), .ZN(
        P3_U2659) );
  INV_X1 U20816 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17626) );
  NOR2_X1 U20817 ( .A1(n18639), .A2(n17685), .ZN(n17642) );
  NAND2_X1 U20818 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17642), .ZN(
        n17634) );
  AOI21_X1 U20819 ( .B1(n17626), .B2(n17634), .A(n17620), .ZN(n18644) );
  OAI21_X1 U20820 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17634), .A(
        n17723), .ZN(n17621) );
  XNOR2_X1 U20821 ( .A(n18644), .B(n17621), .ZN(n17629) );
  NAND2_X1 U20822 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17675) );
  NAND2_X1 U20823 ( .A1(n17736), .A2(n17669), .ZN(n17674) );
  NOR2_X1 U20824 ( .A1(n17675), .A2(n17674), .ZN(n17665) );
  NAND2_X1 U20825 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17665), .ZN(n17636) );
  AOI221_X1 U20826 ( .B1(n17623), .B2(n21642), .C1(n17636), .C2(n21642), .A(
        n17622), .ZN(n17628) );
  OAI211_X1 U20827 ( .C1(n17631), .C2(n18069), .A(n17731), .B(n17624), .ZN(
        n17625) );
  OAI21_X1 U20828 ( .B1(n17753), .B2(n17626), .A(n17625), .ZN(n17627) );
  AOI211_X1 U20829 ( .C1(n17745), .C2(n17629), .A(n17628), .B(n17627), .ZN(
        n17630) );
  OAI211_X1 U20830 ( .C1(n17764), .C2(n18069), .A(n17630), .B(n19055), .ZN(
        P3_U2660) );
  AOI211_X1 U20831 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17647), .A(n17631), .B(
        n17763), .ZN(n17632) );
  AOI211_X1 U20832 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n17715), .A(
        n18963), .B(n17632), .ZN(n17641) );
  NOR2_X1 U20833 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17685), .ZN(
        n17670) );
  AOI21_X1 U20834 ( .B1(n17633), .B2(n17670), .A(n17696), .ZN(n17646) );
  OAI21_X1 U20835 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17642), .A(
        n17634), .ZN(n18652) );
  XNOR2_X1 U20836 ( .A(n17646), .B(n18652), .ZN(n17639) );
  INV_X1 U20837 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19612) );
  NOR3_X1 U20838 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n19612), .A3(n17636), 
        .ZN(n17638) );
  AOI21_X1 U20839 ( .B1(n17736), .B2(n17635), .A(n17751), .ZN(n17658) );
  OR2_X1 U20840 ( .A1(n17636), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17652) );
  INV_X1 U20841 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19614) );
  AOI21_X1 U20842 ( .B1(n17658), .B2(n17652), .A(n19614), .ZN(n17637) );
  AOI211_X1 U20843 ( .C1(n17745), .C2(n17639), .A(n17638), .B(n17637), .ZN(
        n17640) );
  OAI211_X1 U20844 ( .C1(n17764), .C2(n18072), .A(n17641), .B(n17640), .ZN(
        P3_U2661) );
  NOR2_X1 U20845 ( .A1(n18676), .A2(n17685), .ZN(n17660) );
  INV_X1 U20846 ( .A(n17642), .ZN(n17643) );
  OAI21_X1 U20847 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17660), .A(
        n17643), .ZN(n18664) );
  INV_X1 U20848 ( .A(n17670), .ZN(n17644) );
  NOR3_X1 U20849 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18676), .A3(
        n17644), .ZN(n17645) );
  AOI211_X1 U20850 ( .C1(n17646), .C2(n18664), .A(n19040), .B(n17645), .ZN(
        n17654) );
  OAI22_X1 U20851 ( .A1(n19612), .A2(n17658), .B1(n18664), .B2(n17741), .ZN(
        n17651) );
  OAI211_X1 U20852 ( .C1(n17656), .C2(n17649), .A(n17731), .B(n17647), .ZN(
        n17648) );
  OAI21_X1 U20853 ( .B1(n17649), .B2(n17764), .A(n17648), .ZN(n17650) );
  AOI211_X1 U20854 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17715), .A(
        n17651), .B(n17650), .ZN(n17653) );
  OAI211_X1 U20855 ( .C1(n17655), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        P3_U2662) );
  AOI211_X1 U20856 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17679), .A(n17656), .B(
        n17763), .ZN(n17657) );
  AOI211_X1 U20857 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17715), .A(
        n19040), .B(n17657), .ZN(n17668) );
  INV_X1 U20858 ( .A(n17658), .ZN(n17666) );
  INV_X1 U20859 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19611) );
  INV_X1 U20860 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18690) );
  NOR2_X1 U20861 ( .A1(n17659), .A2(n18690), .ZN(n18677) );
  AND2_X1 U20862 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18677), .ZN(
        n17671) );
  INV_X1 U20863 ( .A(n17660), .ZN(n17661) );
  OAI21_X1 U20864 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17671), .A(
        n17661), .ZN(n18679) );
  AOI21_X1 U20865 ( .B1(n17746), .B2(n18677), .A(n17696), .ZN(n17662) );
  INV_X1 U20866 ( .A(n17662), .ZN(n17673) );
  OAI21_X1 U20867 ( .B1(n18679), .B2(n17673), .A(n17745), .ZN(n17663) );
  AOI21_X1 U20868 ( .B1(n18679), .B2(n17673), .A(n17663), .ZN(n17664) );
  AOI221_X1 U20869 ( .B1(n17666), .B2(P3_REIP_REG_8__SCAN_IN), .C1(n17665), 
        .C2(n19611), .A(n17664), .ZN(n17667) );
  OAI211_X1 U20870 ( .C1(n17764), .C2(n18122), .A(n17668), .B(n17667), .ZN(
        P3_U2663) );
  OAI21_X1 U20871 ( .B1(n17669), .B2(n17757), .A(n17767), .ZN(n17704) );
  NOR2_X1 U20872 ( .A1(n17670), .A2(n17696), .ZN(n17687) );
  AOI21_X1 U20873 ( .B1(n18690), .B2(n17685), .A(n17671), .ZN(n18696) );
  INV_X1 U20874 ( .A(n18696), .ZN(n17672) );
  AOI221_X1 U20875 ( .B1(n17687), .B2(n18696), .C1(n17673), .C2(n17672), .A(
        n19581), .ZN(n17678) );
  INV_X1 U20876 ( .A(n17674), .ZN(n17683) );
  OAI211_X1 U20877 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n17683), .B(n17675), .ZN(n17676) );
  OAI211_X1 U20878 ( .C1(n18690), .C2(n17753), .A(n19055), .B(n17676), .ZN(
        n17677) );
  AOI211_X1 U20879 ( .C1(n17704), .C2(P3_REIP_REG_7__SCAN_IN), .A(n17678), .B(
        n17677), .ZN(n17681) );
  OAI211_X1 U20880 ( .C1(n17684), .C2(n17682), .A(n17731), .B(n17679), .ZN(
        n17680) );
  OAI211_X1 U20881 ( .C1(n17682), .C2(n17764), .A(n17681), .B(n17680), .ZN(
        P3_U2664) );
  INV_X1 U20882 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19607) );
  AOI22_X1 U20883 ( .A1(n17752), .A2(P3_EBX_REG_6__SCAN_IN), .B1(n17683), .B2(
        n19607), .ZN(n17694) );
  AOI211_X1 U20884 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17700), .A(n17684), .B(
        n17763), .ZN(n17690) );
  INV_X1 U20885 ( .A(n17697), .ZN(n18716) );
  NOR2_X1 U20886 ( .A1(n18768), .A2(n18716), .ZN(n17695) );
  INV_X1 U20887 ( .A(n17695), .ZN(n17707) );
  NOR2_X1 U20888 ( .A1(n18638), .A2(n17707), .ZN(n17686) );
  OAI21_X1 U20889 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17686), .A(
        n17685), .ZN(n18709) );
  NAND3_X1 U20890 ( .A1(n17745), .A2(n17687), .A3(n18709), .ZN(n17688) );
  OAI21_X1 U20891 ( .B1(n17753), .B2(n18703), .A(n17688), .ZN(n17689) );
  AOI211_X1 U20892 ( .C1(n17704), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17690), .B(
        n17689), .ZN(n17693) );
  INV_X1 U20893 ( .A(n18709), .ZN(n17691) );
  OAI211_X1 U20894 ( .C1(n18703), .C2(n17696), .A(n17691), .B(n17760), .ZN(
        n17692) );
  NAND4_X1 U20895 ( .A1(n17694), .A2(n17693), .A3(n19055), .A4(n17692), .ZN(
        P3_U2665) );
  AOI22_X1 U20896 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17707), .B1(
        n17695), .B2(n18638), .ZN(n18720) );
  AOI21_X1 U20897 ( .B1(n17697), .B2(n17746), .A(n17696), .ZN(n17708) );
  XOR2_X1 U20898 ( .A(n18720), .B(n17708), .Z(n17706) );
  NOR3_X1 U20899 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17757), .A3(n17698), .ZN(
        n17699) );
  AOI211_X1 U20900 ( .C1(n17752), .C2(P3_EBX_REG_5__SCAN_IN), .A(n19040), .B(
        n17699), .ZN(n17702) );
  OAI211_X1 U20901 ( .C1(n17710), .C2(n18129), .A(n17731), .B(n17700), .ZN(
        n17701) );
  OAI211_X1 U20902 ( .C1(n17753), .C2(n18638), .A(n17702), .B(n17701), .ZN(
        n17703) );
  AOI21_X1 U20903 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17704), .A(n17703), .ZN(
        n17705) );
  OAI21_X1 U20904 ( .B1(n19581), .B2(n17706), .A(n17705), .ZN(P3_U2666) );
  NOR2_X1 U20905 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18740), .ZN(
        n18724) );
  NOR2_X1 U20906 ( .A1(n18768), .A2(n18740), .ZN(n17722) );
  OAI21_X1 U20907 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17722), .A(
        n17707), .ZN(n18730) );
  AOI22_X1 U20908 ( .A1(n17746), .A2(n18724), .B1(n17708), .B2(n18730), .ZN(
        n17720) );
  OAI21_X1 U20909 ( .B1(n17714), .B2(n17757), .A(n17767), .ZN(n17729) );
  NAND2_X1 U20910 ( .A1(n19076), .A2(n17709), .ZN(n19730) );
  AOI21_X1 U20911 ( .B1(n9778), .B2(n19519), .A(n19730), .ZN(n17712) );
  AOI211_X1 U20912 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17730), .A(n17710), .B(
        n17763), .ZN(n17711) );
  AOI211_X1 U20913 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17752), .A(n17712), .B(
        n17711), .ZN(n17717) );
  NOR2_X1 U20914 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17757), .ZN(n17713) );
  AOI22_X1 U20915 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17715), .B1(
        n17714), .B2(n17713), .ZN(n17716) );
  OAI211_X1 U20916 ( .C1(n18730), .C2(n17741), .A(n17717), .B(n17716), .ZN(
        n17718) );
  AOI21_X1 U20917 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17729), .A(n17718), .ZN(
        n17719) );
  OAI211_X1 U20918 ( .C1(n17720), .C2(n19581), .A(n17719), .B(n19055), .ZN(
        P3_U2667) );
  INV_X1 U20919 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18743) );
  OAI21_X1 U20920 ( .B1(n17757), .B2(n17721), .A(n19603), .ZN(n17728) );
  NAND2_X1 U20921 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17735) );
  AOI21_X1 U20922 ( .B1(n18743), .B2(n17735), .A(n17722), .ZN(n18746) );
  OAI21_X1 U20923 ( .B1(n17735), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17723), .ZN(n17724) );
  INV_X1 U20924 ( .A(n17724), .ZN(n17744) );
  OAI21_X1 U20925 ( .B1(n18746), .B2(n17744), .A(n17745), .ZN(n17725) );
  AOI21_X1 U20926 ( .B1(n18746), .B2(n17744), .A(n17725), .ZN(n17727) );
  AOI21_X1 U20927 ( .B1(n19530), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n9692), .ZN(n19667) );
  OAI22_X1 U20928 ( .A1(n19667), .A2(n19730), .B1(n17764), .B2(n18125), .ZN(
        n17726) );
  AOI211_X1 U20929 ( .C1(n17729), .C2(n17728), .A(n17727), .B(n17726), .ZN(
        n17733) );
  OAI211_X1 U20930 ( .C1(n17737), .C2(n18125), .A(n17731), .B(n17730), .ZN(
        n17732) );
  OAI211_X1 U20931 ( .C1(n17753), .C2(n18743), .A(n17733), .B(n17732), .ZN(
        P3_U2668) );
  AOI21_X1 U20932 ( .B1(n17736), .B2(n19698), .A(n17751), .ZN(n17749) );
  INV_X1 U20933 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19601) );
  INV_X1 U20934 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17734) );
  NAND2_X1 U20935 ( .A1(n12161), .A2(n19536), .ZN(n19527) );
  OAI21_X1 U20936 ( .B1(n19533), .B2(n19696), .A(n19527), .ZN(n19677) );
  OAI22_X1 U20937 ( .A1(n17734), .A2(n17753), .B1(n19677), .B2(n19730), .ZN(
        n17743) );
  OAI21_X1 U20938 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17735), .ZN(n18760) );
  NAND3_X1 U20939 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17736), .A3(n19601), 
        .ZN(n17740) );
  OR2_X1 U20940 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n17756) );
  AOI211_X1 U20941 ( .C1(n17756), .C2(P3_EBX_REG_2__SCAN_IN), .A(n17763), .B(
        n17737), .ZN(n17738) );
  INV_X1 U20942 ( .A(n17738), .ZN(n17739) );
  OAI211_X1 U20943 ( .C1(n17741), .C2(n18760), .A(n17740), .B(n17739), .ZN(
        n17742) );
  AOI211_X1 U20944 ( .C1(n17752), .C2(P3_EBX_REG_2__SCAN_IN), .A(n17743), .B(
        n17742), .ZN(n17748) );
  OAI211_X1 U20945 ( .C1(n17746), .C2(n18760), .A(n17745), .B(n17744), .ZN(
        n17747) );
  OAI211_X1 U20946 ( .C1(n17749), .C2(n19601), .A(n17748), .B(n17747), .ZN(
        P3_U2669) );
  NAND2_X1 U20947 ( .A1(n17750), .A2(n19536), .ZN(n19682) );
  AOI22_X1 U20948 ( .A1(n17752), .A2(P3_EBX_REG_1__SCAN_IN), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n17751), .ZN(n17762) );
  OAI21_X1 U20949 ( .B1(n17755), .B2(n17754), .A(n17753), .ZN(n17759) );
  NAND2_X1 U20950 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18140) );
  NAND2_X1 U20951 ( .A1(n17756), .A2(n18140), .ZN(n18146) );
  OAI22_X1 U20952 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17757), .B1(n17763), 
        .B2(n18146), .ZN(n17758) );
  AOI221_X1 U20953 ( .B1(n17760), .B2(n18768), .C1(n17759), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17758), .ZN(n17761) );
  OAI211_X1 U20954 ( .C1(n19682), .C2(n19730), .A(n17762), .B(n17761), .ZN(
        P3_U2670) );
  NAND2_X1 U20955 ( .A1(n17764), .A2(n17763), .ZN(n17766) );
  AOI22_X1 U20956 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17766), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17765), .ZN(n17769) );
  NAND3_X1 U20957 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19726), .A3(
        n17767), .ZN(n17768) );
  NAND2_X1 U20958 ( .A1(n17771), .A2(n17770), .ZN(n17772) );
  NAND2_X1 U20959 ( .A1(n17772), .A2(n18143), .ZN(n17871) );
  AOI22_X1 U20960 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U20961 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17776) );
  AOI22_X1 U20962 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U20963 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17774) );
  NAND4_X1 U20964 ( .A1(n17777), .A2(n17776), .A3(n17775), .A4(n17774), .ZN(
        n17783) );
  AOI22_X1 U20965 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U20966 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U20967 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U20968 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17778) );
  NAND4_X1 U20969 ( .A1(n17781), .A2(n17780), .A3(n17779), .A4(n17778), .ZN(
        n17782) );
  NOR2_X1 U20970 ( .A1(n17783), .A2(n17782), .ZN(n17883) );
  AOI22_X1 U20971 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U20972 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17786) );
  AOI22_X1 U20973 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17785) );
  AOI22_X1 U20974 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17784) );
  NAND4_X1 U20975 ( .A1(n17787), .A2(n17786), .A3(n17785), .A4(n17784), .ZN(
        n17794) );
  AOI22_X1 U20976 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17792) );
  AOI22_X1 U20977 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17791) );
  AOI22_X1 U20978 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17790) );
  AOI22_X1 U20979 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9692), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17789) );
  NAND4_X1 U20980 ( .A1(n17792), .A2(n17791), .A3(n17790), .A4(n17789), .ZN(
        n17793) );
  NOR2_X1 U20981 ( .A1(n17794), .A2(n17793), .ZN(n17893) );
  AOI22_X1 U20982 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12075), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17798) );
  AOI22_X1 U20983 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18075), .B1(
        n9692), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17797) );
  AOI22_X1 U20984 ( .A1(n18104), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17796) );
  AOI22_X1 U20985 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17795) );
  NAND4_X1 U20986 ( .A1(n17798), .A2(n17797), .A3(n17796), .A4(n17795), .ZN(
        n17804) );
  AOI22_X1 U20987 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17802) );
  AOI22_X1 U20988 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18095), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17801) );
  AOI22_X1 U20989 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9688), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17800) );
  AOI22_X1 U20990 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18106), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17799) );
  NAND4_X1 U20991 ( .A1(n17802), .A2(n17801), .A3(n17800), .A4(n17799), .ZN(
        n17803) );
  NOR2_X1 U20992 ( .A1(n17804), .A2(n17803), .ZN(n17902) );
  AOI22_X1 U20993 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17816) );
  AOI22_X1 U20994 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U20995 ( .A1(n18104), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17805) );
  OAI21_X1 U20996 ( .B1(n11976), .B2(n21634), .A(n17805), .ZN(n17813) );
  AOI22_X1 U20997 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U20998 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17810) );
  AOI22_X1 U20999 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U21000 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17808) );
  NAND4_X1 U21001 ( .A1(n17811), .A2(n17810), .A3(n17809), .A4(n17808), .ZN(
        n17812) );
  AOI211_X1 U21002 ( .C1(n18105), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17813), .B(n17812), .ZN(n17814) );
  NAND3_X1 U21003 ( .A1(n17816), .A2(n17815), .A3(n17814), .ZN(n17906) );
  AOI22_X1 U21004 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U21005 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17826) );
  AOI22_X1 U21006 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17818) );
  OAI21_X1 U21007 ( .B1(n11976), .B2(n21618), .A(n17818), .ZN(n17824) );
  AOI22_X1 U21008 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U21009 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U21010 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U21011 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17819) );
  NAND4_X1 U21012 ( .A1(n17822), .A2(n17821), .A3(n17820), .A4(n17819), .ZN(
        n17823) );
  AOI211_X1 U21013 ( .C1(n18105), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17824), .B(n17823), .ZN(n17825) );
  NAND3_X1 U21014 ( .A1(n17827), .A2(n17826), .A3(n17825), .ZN(n17907) );
  NAND2_X1 U21015 ( .A1(n17906), .A2(n17907), .ZN(n17905) );
  NOR2_X1 U21016 ( .A1(n17902), .A2(n17905), .ZN(n17898) );
  AOI22_X1 U21017 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U21018 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U21019 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17828) );
  OAI21_X1 U21020 ( .B1(n17817), .B2(n21639), .A(n17828), .ZN(n17834) );
  AOI22_X1 U21021 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U21022 ( .A1(n18104), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U21023 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17830) );
  AOI22_X1 U21024 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17829) );
  NAND4_X1 U21025 ( .A1(n17832), .A2(n17831), .A3(n17830), .A4(n17829), .ZN(
        n17833) );
  AOI211_X1 U21026 ( .C1(n18043), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n17834), .B(n17833), .ZN(n17835) );
  NAND3_X1 U21027 ( .A1(n17837), .A2(n17836), .A3(n17835), .ZN(n17897) );
  NAND2_X1 U21028 ( .A1(n17898), .A2(n17897), .ZN(n17896) );
  NOR2_X1 U21029 ( .A1(n17893), .A2(n17896), .ZN(n17890) );
  AOI22_X1 U21030 ( .A1(n18104), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17847) );
  AOI22_X1 U21031 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17846) );
  AOI22_X1 U21032 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17838) );
  OAI21_X1 U21033 ( .B1(n11969), .B2(n21691), .A(n17838), .ZN(n17844) );
  AOI22_X1 U21034 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17842) );
  AOI22_X1 U21035 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U21036 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17840) );
  AOI22_X1 U21037 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17839) );
  NAND4_X1 U21038 ( .A1(n17842), .A2(n17841), .A3(n17840), .A4(n17839), .ZN(
        n17843) );
  AOI211_X1 U21039 ( .C1(n12071), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17844), .B(n17843), .ZN(n17845) );
  NAND3_X1 U21040 ( .A1(n17847), .A2(n17846), .A3(n17845), .ZN(n17889) );
  NAND2_X1 U21041 ( .A1(n17890), .A2(n17889), .ZN(n17888) );
  NOR2_X1 U21042 ( .A1(n17883), .A2(n17888), .ZN(n17882) );
  INV_X1 U21043 ( .A(n17882), .ZN(n17876) );
  AOI22_X1 U21044 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17851) );
  AOI22_X1 U21045 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17850) );
  AOI22_X1 U21046 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17849) );
  AOI22_X1 U21047 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17848) );
  NAND4_X1 U21048 ( .A1(n17851), .A2(n17850), .A3(n17849), .A4(n17848), .ZN(
        n17858) );
  AOI22_X1 U21049 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17856) );
  AOI22_X1 U21050 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17855) );
  AOI22_X1 U21051 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U21052 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17853) );
  NAND4_X1 U21053 ( .A1(n17856), .A2(n17855), .A3(n17854), .A4(n17853), .ZN(
        n17857) );
  NOR2_X1 U21054 ( .A1(n17858), .A2(n17857), .ZN(n17875) );
  NOR2_X1 U21055 ( .A1(n17876), .A2(n17875), .ZN(n17870) );
  AOI22_X1 U21056 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17862) );
  AOI22_X1 U21057 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17861) );
  AOI22_X1 U21058 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17860) );
  AOI22_X1 U21059 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17859) );
  NAND4_X1 U21060 ( .A1(n17862), .A2(n17861), .A3(n17860), .A4(n17859), .ZN(
        n17868) );
  AOI22_X1 U21061 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17866) );
  AOI22_X1 U21062 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17865) );
  AOI22_X1 U21063 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17864) );
  AOI22_X1 U21064 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17863) );
  NAND4_X1 U21065 ( .A1(n17866), .A2(n17865), .A3(n17864), .A4(n17863), .ZN(
        n17867) );
  NOR2_X1 U21066 ( .A1(n17868), .A2(n17867), .ZN(n17869) );
  XOR2_X1 U21067 ( .A(n17870), .B(n17869), .Z(n18163) );
  OAI22_X1 U21068 ( .A1(n17872), .A2(n17871), .B1(n18163), .B2(n18143), .ZN(
        P3_U2673) );
  NOR2_X1 U21069 ( .A1(n18197), .A2(n18147), .ZN(n18123) );
  NAND2_X1 U21070 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17874) );
  XOR2_X1 U21071 ( .A(n17876), .B(n17875), .Z(n18164) );
  INV_X1 U21072 ( .A(n17877), .ZN(n17900) );
  NOR2_X1 U21073 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17878), .ZN(n17879) );
  AOI22_X1 U21074 ( .A1(n18148), .A2(n18164), .B1(n17900), .B2(n17879), .ZN(
        n17880) );
  OAI21_X1 U21075 ( .B1(n17887), .B2(n17881), .A(n17880), .ZN(P3_U2674) );
  INV_X1 U21076 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17886) );
  AOI21_X1 U21077 ( .B1(n17883), .B2(n17888), .A(n17882), .ZN(n18168) );
  NOR2_X1 U21078 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21705), .ZN(n17884) );
  AOI22_X1 U21079 ( .A1(n18148), .A2(n18168), .B1(n17891), .B2(n17884), .ZN(
        n17885) );
  OAI21_X1 U21080 ( .B1(n17890), .B2(n17889), .A(n17888), .ZN(n18176) );
  AOI22_X1 U21081 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17894), .B1(n17891), 
        .B2(n21705), .ZN(n17892) );
  OAI21_X1 U21082 ( .B1(n18143), .B2(n18176), .A(n17892), .ZN(P3_U2676) );
  XNOR2_X1 U21083 ( .A(n17893), .B(n17896), .ZN(n18180) );
  OAI21_X1 U21084 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17900), .A(n17894), .ZN(
        n17895) );
  OAI21_X1 U21085 ( .B1(n18180), .B2(n18143), .A(n17895), .ZN(P3_U2677) );
  AOI21_X1 U21086 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18143), .A(n17904), .ZN(
        n17899) );
  OAI21_X1 U21087 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n18185) );
  OAI22_X1 U21088 ( .A1(n17900), .A2(n17899), .B1(n18143), .B2(n18185), .ZN(
        P3_U2678) );
  INV_X1 U21089 ( .A(n17901), .ZN(n17909) );
  AOI21_X1 U21090 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18143), .A(n17909), .ZN(
        n17903) );
  XNOR2_X1 U21091 ( .A(n17902), .B(n17905), .ZN(n18190) );
  OAI22_X1 U21092 ( .A1(n17904), .A2(n17903), .B1(n18143), .B2(n18190), .ZN(
        P3_U2679) );
  AOI22_X1 U21093 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18143), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n17910), .ZN(n17908) );
  OAI21_X1 U21094 ( .B1(n17907), .B2(n17906), .A(n17905), .ZN(n18195) );
  OAI22_X1 U21095 ( .A1(n17909), .A2(n17908), .B1(n18143), .B2(n18195), .ZN(
        P3_U2680) );
  AOI22_X1 U21096 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17915) );
  AOI22_X1 U21097 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17914) );
  AOI22_X1 U21098 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17911), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U21099 ( .A1(n12071), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17912) );
  NAND4_X1 U21100 ( .A1(n17915), .A2(n17914), .A3(n17913), .A4(n17912), .ZN(
        n17921) );
  AOI22_X1 U21101 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17919) );
  AOI22_X1 U21102 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U21103 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U21104 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17916) );
  NAND4_X1 U21105 ( .A1(n17919), .A2(n17918), .A3(n17917), .A4(n17916), .ZN(
        n17920) );
  NOR2_X1 U21106 ( .A1(n17921), .A2(n17920), .ZN(n18198) );
  NAND3_X1 U21107 ( .A1(n10704), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18143), 
        .ZN(n17922) );
  OAI221_X1 U21108 ( .B1(n10704), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18143), 
        .C2(n18198), .A(n17922), .ZN(P3_U2681) );
  AOI22_X1 U21109 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17926) );
  AOI22_X1 U21110 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U21111 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U21112 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17923) );
  NAND4_X1 U21113 ( .A1(n17926), .A2(n17925), .A3(n17924), .A4(n17923), .ZN(
        n17932) );
  AOI22_X1 U21114 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17930) );
  AOI22_X1 U21115 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U21116 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U21117 ( .A1(n9702), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17927) );
  NAND4_X1 U21118 ( .A1(n17930), .A2(n17929), .A3(n17928), .A4(n17927), .ZN(
        n17931) );
  NOR2_X1 U21119 ( .A1(n17932), .A2(n17931), .ZN(n18203) );
  OAI21_X1 U21120 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17947), .A(n17933), .ZN(
        n17934) );
  AOI22_X1 U21121 ( .A1(n18148), .A2(n18203), .B1(n17934), .B2(n18143), .ZN(
        P3_U2682) );
  OAI21_X1 U21122 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17935), .A(n18143), .ZN(
        n17946) );
  AOI22_X1 U21123 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17939) );
  AOI22_X1 U21124 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17938) );
  AOI22_X1 U21125 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U21126 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17936) );
  NAND4_X1 U21127 ( .A1(n17939), .A2(n17938), .A3(n17937), .A4(n17936), .ZN(
        n17945) );
  AOI22_X1 U21128 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9695), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17943) );
  AOI22_X1 U21129 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17942) );
  AOI22_X1 U21130 ( .A1(n9702), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17941) );
  AOI22_X1 U21131 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17940) );
  NAND4_X1 U21132 ( .A1(n17943), .A2(n17942), .A3(n17941), .A4(n17940), .ZN(
        n17944) );
  NOR2_X1 U21133 ( .A1(n17945), .A2(n17944), .ZN(n18209) );
  OAI22_X1 U21134 ( .A1(n17947), .A2(n17946), .B1(n18209), .B2(n18143), .ZN(
        P3_U2683) );
  AOI22_X1 U21135 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U21136 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U21137 ( .A1(n18104), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17949) );
  AOI22_X1 U21138 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17948) );
  NAND4_X1 U21139 ( .A1(n17951), .A2(n17950), .A3(n17949), .A4(n17948), .ZN(
        n17957) );
  AOI22_X1 U21140 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17955) );
  AOI22_X1 U21141 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U21142 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17953) );
  AOI22_X1 U21143 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17952) );
  NAND4_X1 U21144 ( .A1(n17955), .A2(n17954), .A3(n17953), .A4(n17952), .ZN(
        n17956) );
  NOR2_X1 U21145 ( .A1(n17957), .A2(n17956), .ZN(n18216) );
  OAI21_X1 U21146 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17973), .A(n17958), .ZN(
        n17959) );
  AOI22_X1 U21147 ( .A1(n18148), .A2(n18216), .B1(n17959), .B2(n18143), .ZN(
        P3_U2684) );
  AOI21_X1 U21148 ( .B1(n17960), .B2(n17984), .A(n18148), .ZN(n17961) );
  INV_X1 U21149 ( .A(n17961), .ZN(n17972) );
  AOI22_X1 U21150 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17807), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17965) );
  AOI22_X1 U21151 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17964) );
  AOI22_X1 U21152 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17963) );
  AOI22_X1 U21153 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17962) );
  NAND4_X1 U21154 ( .A1(n17965), .A2(n17964), .A3(n17963), .A4(n17962), .ZN(
        n17971) );
  AOI22_X1 U21155 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U21156 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17968) );
  AOI22_X1 U21157 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17967) );
  AOI22_X1 U21158 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17966) );
  NAND4_X1 U21159 ( .A1(n17969), .A2(n17968), .A3(n17967), .A4(n17966), .ZN(
        n17970) );
  NOR2_X1 U21160 ( .A1(n17971), .A2(n17970), .ZN(n18221) );
  OAI22_X1 U21161 ( .A1(n17973), .A2(n17972), .B1(n18221), .B2(n18143), .ZN(
        P3_U2685) );
  AOI22_X1 U21162 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18106), .ZN(n17977) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18104), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12075), .ZN(n17976) );
  AOI22_X1 U21164 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18095), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18073), .ZN(n17975) );
  AOI22_X1 U21165 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9701), .ZN(n17974) );
  NAND4_X1 U21166 ( .A1(n17977), .A2(n17976), .A3(n17975), .A4(n17974), .ZN(
        n17983) );
  AOI22_X1 U21167 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18043), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n9688), .ZN(n17981) );
  AOI22_X1 U21168 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n18075), .ZN(n17980) );
  AOI22_X1 U21169 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17979) );
  AOI22_X1 U21170 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18107), .ZN(n17978) );
  NAND4_X1 U21171 ( .A1(n17981), .A2(n17980), .A3(n17979), .A4(n17978), .ZN(
        n17982) );
  NOR2_X1 U21172 ( .A1(n17983), .A2(n17982), .ZN(n18227) );
  OAI21_X1 U21173 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17985), .A(n17984), .ZN(
        n17986) );
  AOI22_X1 U21174 ( .A1(n18148), .A2(n18227), .B1(n17986), .B2(n18143), .ZN(
        P3_U2686) );
  NAND2_X1 U21175 ( .A1(n18143), .A2(n17998), .ZN(n18013) );
  AOI22_X1 U21176 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17997) );
  AOI22_X1 U21177 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U21178 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17987) );
  OAI21_X1 U21179 ( .B1(n17988), .B2(n21634), .A(n17987), .ZN(n17994) );
  AOI22_X1 U21180 ( .A1(n9702), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U21181 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U21182 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17990) );
  AOI22_X1 U21183 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17989) );
  NAND4_X1 U21184 ( .A1(n17992), .A2(n17991), .A3(n17990), .A4(n17989), .ZN(
        n17993) );
  AOI211_X1 U21185 ( .C1(n9692), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17994), .B(n17993), .ZN(n17995) );
  NAND3_X1 U21186 ( .A1(n17997), .A2(n17996), .A3(n17995), .ZN(n18228) );
  NOR3_X1 U21187 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18197), .A3(n17998), .ZN(
        n17999) );
  AOI21_X1 U21188 ( .B1(n18148), .B2(n18228), .A(n17999), .ZN(n18000) );
  OAI21_X1 U21189 ( .B1(n18001), .B2(n18013), .A(n18000), .ZN(P3_U2687) );
  AOI22_X1 U21190 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U21191 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18004) );
  AOI22_X1 U21192 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18003) );
  AOI22_X1 U21193 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18002) );
  NAND4_X1 U21194 ( .A1(n18005), .A2(n18004), .A3(n18003), .A4(n18002), .ZN(
        n18012) );
  AOI22_X1 U21195 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18010) );
  AOI22_X1 U21196 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U21197 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18008) );
  AOI22_X1 U21198 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9693), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18007) );
  NAND4_X1 U21199 ( .A1(n18010), .A2(n18009), .A3(n18008), .A4(n18007), .ZN(
        n18011) );
  NOR2_X1 U21200 ( .A1(n18012), .A2(n18011), .ZN(n18237) );
  NOR2_X1 U21201 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n9881), .ZN(n18014) );
  OAI22_X1 U21202 ( .A1(n18237), .A2(n18143), .B1(n18014), .B2(n18013), .ZN(
        P3_U2688) );
  NAND2_X1 U21203 ( .A1(n18143), .A2(n18027), .ZN(n18041) );
  AOI22_X1 U21204 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18026) );
  AOI22_X1 U21205 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18025) );
  INV_X1 U21206 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21523) );
  AOI22_X1 U21207 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18015) );
  OAI21_X1 U21208 ( .B1(n18016), .B2(n21523), .A(n18015), .ZN(n18023) );
  AOI22_X1 U21209 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U21210 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18020) );
  AOI22_X1 U21211 ( .A1(n17852), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U21212 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18018) );
  NAND4_X1 U21213 ( .A1(n18021), .A2(n18020), .A3(n18019), .A4(n18018), .ZN(
        n18022) );
  AOI211_X1 U21214 ( .C1(n9695), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n18023), .B(n18022), .ZN(n18024) );
  NAND3_X1 U21215 ( .A1(n18026), .A2(n18025), .A3(n18024), .ZN(n18240) );
  NOR3_X1 U21216 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18197), .A3(n18027), .ZN(
        n18028) );
  AOI21_X1 U21217 ( .B1(n18148), .B2(n18240), .A(n18028), .ZN(n18029) );
  OAI21_X1 U21218 ( .B1(n18030), .B2(n18041), .A(n18029), .ZN(P3_U2689) );
  AOI22_X1 U21219 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U21220 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18033) );
  AOI22_X1 U21221 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9696), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18032) );
  AOI22_X1 U21222 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9701), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18031) );
  NAND4_X1 U21223 ( .A1(n18034), .A2(n18033), .A3(n18032), .A4(n18031), .ZN(
        n18040) );
  AOI22_X1 U21224 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18038) );
  AOI22_X1 U21225 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18037) );
  AOI22_X1 U21226 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U21227 ( .A1(n9693), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18035) );
  NAND4_X1 U21228 ( .A1(n18038), .A2(n18037), .A3(n18036), .A4(n18035), .ZN(
        n18039) );
  NOR2_X1 U21229 ( .A1(n18040), .A2(n18039), .ZN(n18244) );
  NOR2_X1 U21230 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18055), .ZN(n18042) );
  OAI22_X1 U21231 ( .A1(n18244), .A2(n18143), .B1(n18042), .B2(n18041), .ZN(
        P3_U2690) );
  OAI21_X1 U21232 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18068), .A(n18143), .ZN(
        n18054) );
  AOI22_X1 U21233 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18047) );
  AOI22_X1 U21234 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18046) );
  AOI22_X1 U21235 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18045) );
  AOI22_X1 U21236 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18044) );
  NAND4_X1 U21237 ( .A1(n18047), .A2(n18046), .A3(n18045), .A4(n18044), .ZN(
        n18053) );
  AOI22_X1 U21238 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9693), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18051) );
  AOI22_X1 U21239 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U21240 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U21241 ( .A1(n18094), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18048) );
  NAND4_X1 U21242 ( .A1(n18051), .A2(n18050), .A3(n18049), .A4(n18048), .ZN(
        n18052) );
  NOR2_X1 U21243 ( .A1(n18053), .A2(n18052), .ZN(n18248) );
  OAI22_X1 U21244 ( .A1(n18055), .A2(n18054), .B1(n18248), .B2(n18143), .ZN(
        P3_U2691) );
  AOI22_X1 U21245 ( .A1(n9713), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18113), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18067) );
  AOI22_X1 U21246 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U21247 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18057) );
  OAI21_X1 U21248 ( .B1(n18058), .B2(n21702), .A(n18057), .ZN(n18064) );
  AOI22_X1 U21249 ( .A1(n18006), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18062) );
  AOI22_X1 U21250 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18061) );
  AOI22_X1 U21251 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12075), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U21252 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18059) );
  NAND4_X1 U21253 ( .A1(n18062), .A2(n18061), .A3(n18060), .A4(n18059), .ZN(
        n18063) );
  AOI211_X1 U21254 ( .C1(n9688), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n18064), .B(n18063), .ZN(n18065) );
  NAND3_X1 U21255 ( .A1(n18067), .A2(n18066), .A3(n18065), .ZN(n18251) );
  AOI21_X1 U21256 ( .B1(n18069), .B2(n18087), .A(n18068), .ZN(n18070) );
  OAI22_X1 U21257 ( .A1(n18143), .A2(n18251), .B1(n18070), .B2(n18148), .ZN(
        n18071) );
  INV_X1 U21258 ( .A(n18071), .ZN(P3_U2692) );
  AOI21_X1 U21259 ( .B1(n18072), .B2(n18102), .A(n18148), .ZN(n18086) );
  AOI22_X1 U21260 ( .A1(n18073), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18085) );
  AOI22_X1 U21261 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U21262 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18074) );
  OAI21_X1 U21263 ( .B1(n9778), .B2(n21639), .A(n18074), .ZN(n18082) );
  AOI22_X1 U21264 ( .A1(n18075), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U21265 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U21266 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U21267 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18077) );
  NAND4_X1 U21268 ( .A1(n18080), .A2(n18079), .A3(n18078), .A4(n18077), .ZN(
        n18081) );
  AOI211_X1 U21269 ( .C1(n18104), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n18082), .B(n18081), .ZN(n18083) );
  NAND3_X1 U21270 ( .A1(n18085), .A2(n18084), .A3(n18083), .ZN(n18254) );
  AOI22_X1 U21271 ( .A1(n18087), .A2(n18086), .B1(n18254), .B2(n18148), .ZN(
        n18088) );
  INV_X1 U21272 ( .A(n18088), .ZN(P3_U2693) );
  AOI22_X1 U21273 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18093) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12075), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n18104), .ZN(n18092) );
  AOI22_X1 U21275 ( .A1(n9695), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18006), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18091) );
  AOI22_X1 U21276 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12071), .ZN(n18090) );
  NAND4_X1 U21277 ( .A1(n18093), .A2(n18092), .A3(n18091), .A4(n18090), .ZN(
        n18101) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17852), .B1(
        n9696), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18099) );
  AOI22_X1 U21279 ( .A1(n18113), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18075), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U21280 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n18095), .ZN(n18097) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18106), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9693), .ZN(n18096) );
  NAND4_X1 U21282 ( .A1(n18099), .A2(n18098), .A3(n18097), .A4(n18096), .ZN(
        n18100) );
  NOR2_X1 U21283 ( .A1(n18101), .A2(n18100), .ZN(n18259) );
  OAI21_X1 U21284 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18120), .A(n18102), .ZN(
        n18103) );
  AOI22_X1 U21285 ( .A1(n18148), .A2(n18259), .B1(n18103), .B2(n18143), .ZN(
        P3_U2694) );
  AND2_X1 U21286 ( .A1(n18143), .A2(n18126), .ZN(n18121) );
  AOI22_X1 U21287 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18104), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18111) );
  AOI22_X1 U21288 ( .A1(n9692), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U21289 ( .A1(n9696), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9693), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18109) );
  AOI22_X1 U21290 ( .A1(n12075), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12071), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18108) );
  NAND4_X1 U21291 ( .A1(n18111), .A2(n18110), .A3(n18109), .A4(n18108), .ZN(
        n18119) );
  AOI22_X1 U21292 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9702), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18117) );
  AOI22_X1 U21293 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18116) );
  AOI22_X1 U21294 ( .A1(n18017), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18073), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U21295 ( .A1(n18076), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18094), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18114) );
  NAND4_X1 U21296 ( .A1(n18117), .A2(n18116), .A3(n18115), .A4(n18114), .ZN(
        n18118) );
  NOR2_X1 U21297 ( .A1(n18119), .A2(n18118), .ZN(n18266) );
  AOI222_X1 U21298 ( .A1(n18122), .A2(n18121), .B1(n18148), .B2(n18266), .C1(
        n19105), .C2(n18120), .ZN(P3_U2695) );
  INV_X1 U21299 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19109) );
  INV_X1 U21300 ( .A(n18123), .ZN(n18150) );
  NOR2_X1 U21301 ( .A1(n18124), .A2(n18150), .ZN(n18136) );
  INV_X1 U21302 ( .A(n18136), .ZN(n18141) );
  NOR2_X1 U21303 ( .A1(n18125), .A2(n18141), .ZN(n18138) );
  NAND2_X1 U21304 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18138), .ZN(n18128) );
  INV_X1 U21305 ( .A(n18128), .ZN(n18135) );
  AND3_X1 U21306 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n18135), .ZN(n18131) );
  OAI211_X1 U21307 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n18131), .A(n18126), .B(
        n18143), .ZN(n18127) );
  OAI21_X1 U21308 ( .B1(n18143), .B2(n19109), .A(n18127), .ZN(P3_U2696) );
  NOR2_X1 U21309 ( .A1(n18129), .A2(n18128), .ZN(n18133) );
  AOI21_X1 U21310 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18143), .A(n18133), .ZN(
        n18130) );
  INV_X1 U21311 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19102) );
  OAI22_X1 U21312 ( .A1(n18131), .A2(n18130), .B1(n19102), .B2(n18143), .ZN(
        P3_U2697) );
  AOI21_X1 U21313 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18143), .A(n18135), .ZN(
        n18132) );
  INV_X1 U21314 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19098) );
  OAI22_X1 U21315 ( .A1(n18133), .A2(n18132), .B1(n19098), .B2(n18143), .ZN(
        P3_U2698) );
  AOI21_X1 U21316 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18143), .A(n18138), .ZN(
        n18134) );
  INV_X1 U21317 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19094) );
  OAI22_X1 U21318 ( .A1(n18135), .A2(n18134), .B1(n19094), .B2(n18143), .ZN(
        P3_U2699) );
  AOI21_X1 U21319 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18143), .A(n18136), .ZN(
        n18137) );
  INV_X1 U21320 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19090) );
  OAI22_X1 U21321 ( .A1(n18138), .A2(n18137), .B1(n19090), .B2(n18143), .ZN(
        P3_U2700) );
  INV_X1 U21322 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19086) );
  INV_X1 U21323 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18139) );
  OAI21_X1 U21324 ( .B1(n18147), .B2(n18140), .A(n18139), .ZN(n18142) );
  NAND3_X1 U21325 ( .A1(n18143), .A2(n18142), .A3(n18141), .ZN(n18144) );
  OAI21_X1 U21326 ( .B1(n18143), .B2(n19086), .A(n18144), .ZN(P3_U2701) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18148), .B1(
        P3_EBX_REG_1__SCAN_IN), .B2(n18147), .ZN(n18145) );
  OAI21_X1 U21328 ( .B1(n18150), .B2(n18146), .A(n18145), .ZN(P3_U2702) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18148), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18147), .ZN(n18149) );
  OAI21_X1 U21330 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18150), .A(n18149), .ZN(
        P3_U2703) );
  INV_X1 U21331 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18363) );
  INV_X1 U21332 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18380) );
  NAND4_X1 U21333 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n18277) );
  NOR2_X1 U21334 ( .A1(n18380), .A2(n18277), .ZN(n18151) );
  NAND4_X1 U21335 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n18151), .ZN(n18238) );
  NAND2_X1 U21336 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n18152) );
  INV_X1 U21337 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18394) );
  INV_X1 U21338 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18392) );
  INV_X1 U21339 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18390) );
  NOR4_X1 U21340 ( .A1(n18152), .A2(n18394), .A3(n18392), .A4(n18390), .ZN(
        n18153) );
  INV_X1 U21341 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18406) );
  INV_X1 U21342 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18354) );
  INV_X1 U21343 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18352) );
  NAND4_X1 U21344 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(n18155), .ZN(n18196) );
  INV_X1 U21345 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18356) );
  NAND2_X1 U21346 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18192), .ZN(n18191) );
  NAND2_X1 U21347 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18186), .ZN(n18187) );
  INV_X1 U21348 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18367) );
  NAND2_X1 U21349 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18169), .ZN(n18165) );
  INV_X1 U21350 ( .A(n18165), .ZN(n18160) );
  NAND2_X1 U21351 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18160), .ZN(n18159) );
  NAND3_X1 U21352 ( .A1(n18286), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n18159), 
        .ZN(n18158) );
  NAND2_X1 U21353 ( .A1(n18156), .A2(n18263), .ZN(n18233) );
  NAND2_X1 U21354 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18222), .ZN(n18157) );
  OAI211_X1 U21355 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n18159), .A(n18158), .B(
        n18157), .ZN(P3_U2704) );
  NAND2_X1 U21356 ( .A1(n19095), .A2(n18263), .ZN(n18207) );
  AOI22_X1 U21357 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18222), .ZN(n18162) );
  OAI211_X1 U21358 ( .C1(n18160), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18286), .B(
        n18159), .ZN(n18161) );
  OAI211_X1 U21359 ( .C1(n18163), .C2(n18297), .A(n18162), .B(n18161), .ZN(
        P3_U2705) );
  AOI22_X1 U21360 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18222), .B1(n18164), .B2(
        n18255), .ZN(n18167) );
  OAI211_X1 U21361 ( .C1(n18169), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18286), .B(
        n18165), .ZN(n18166) );
  OAI211_X1 U21362 ( .C1(n18207), .C2(n18400), .A(n18167), .B(n18166), .ZN(
        P3_U2706) );
  AOI22_X1 U21363 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18222), .B1(n18168), .B2(
        n18255), .ZN(n18172) );
  AOI211_X1 U21364 ( .C1(n18367), .C2(n18173), .A(n18169), .B(n18263), .ZN(
        n18170) );
  INV_X1 U21365 ( .A(n18170), .ZN(n18171) );
  OAI211_X1 U21366 ( .C1(n18207), .C2(n14092), .A(n18172), .B(n18171), .ZN(
        P3_U2707) );
  AOI22_X1 U21367 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18222), .ZN(n18175) );
  OAI211_X1 U21368 ( .C1(n9785), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18286), .B(
        n18173), .ZN(n18174) );
  OAI211_X1 U21369 ( .C1(n18297), .C2(n18176), .A(n18175), .B(n18174), .ZN(
        P3_U2708) );
  AOI22_X1 U21370 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18222), .ZN(n18179) );
  AOI211_X1 U21371 ( .C1(n18363), .C2(n18181), .A(n9785), .B(n18263), .ZN(
        n18177) );
  INV_X1 U21372 ( .A(n18177), .ZN(n18178) );
  OAI211_X1 U21373 ( .C1(n18297), .C2(n18180), .A(n18179), .B(n18178), .ZN(
        P3_U2709) );
  AOI22_X1 U21374 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18222), .ZN(n18184) );
  OAI211_X1 U21375 ( .C1(n18182), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18286), .B(
        n18181), .ZN(n18183) );
  OAI211_X1 U21376 ( .C1(n18185), .C2(n18297), .A(n18184), .B(n18183), .ZN(
        P3_U2710) );
  AOI22_X1 U21377 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18222), .ZN(n18189) );
  OAI211_X1 U21378 ( .C1(n18186), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18286), .B(
        n18187), .ZN(n18188) );
  OAI211_X1 U21379 ( .C1(n18190), .C2(n18297), .A(n18189), .B(n18188), .ZN(
        P3_U2711) );
  AOI22_X1 U21380 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18222), .ZN(n18194) );
  OAI211_X1 U21381 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18192), .A(n18286), .B(
        n18191), .ZN(n18193) );
  OAI211_X1 U21382 ( .C1(n18195), .C2(n18297), .A(n18194), .B(n18193), .ZN(
        P3_U2712) );
  INV_X1 U21383 ( .A(n18281), .ZN(n18294) );
  INV_X1 U21384 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18348) );
  NOR2_X1 U21385 ( .A1(n18197), .A2(n18230), .ZN(n18224) );
  NAND2_X1 U21386 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18224), .ZN(n18223) );
  NAND2_X1 U21387 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18217), .ZN(n18213) );
  NOR2_X1 U21388 ( .A1(n18352), .A2(n18213), .ZN(n18205) );
  NOR2_X1 U21389 ( .A1(n18263), .A2(n18205), .ZN(n18208) );
  AOI21_X1 U21390 ( .B1(n18294), .B2(n18354), .A(n18208), .ZN(n18202) );
  NOR3_X1 U21391 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18197), .A3(n18196), .ZN(
        n18200) );
  OAI22_X1 U21392 ( .A1(n18198), .A2(n18297), .B1(n21624), .B2(n18233), .ZN(
        n18199) );
  AOI211_X1 U21393 ( .C1(n18229), .C2(BUF2_REG_6__SCAN_IN), .A(n18200), .B(
        n18199), .ZN(n18201) );
  OAI21_X1 U21394 ( .B1(n18202), .B2(n18356), .A(n18201), .ZN(P3_U2713) );
  OAI22_X1 U21395 ( .A1(n18203), .A2(n18297), .B1(n16432), .B2(n18233), .ZN(
        n18204) );
  AOI221_X1 U21396 ( .B1(n18208), .B2(P3_EAX_REG_21__SCAN_IN), .C1(n18205), 
        .C2(n18354), .A(n18204), .ZN(n18206) );
  OAI21_X1 U21397 ( .B1(n14101), .B2(n18207), .A(n18206), .ZN(P3_U2714) );
  INV_X1 U21398 ( .A(n18208), .ZN(n18212) );
  OAI22_X1 U21399 ( .A1(n18209), .A2(n18297), .B1(n16440), .B2(n18233), .ZN(
        n18210) );
  AOI21_X1 U21400 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n18229), .A(n18210), .ZN(
        n18211) );
  OAI221_X1 U21401 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n18213), .C1(n18352), 
        .C2(n18212), .A(n18211), .ZN(P3_U2715) );
  AOI22_X1 U21402 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18222), .ZN(n18215) );
  OAI211_X1 U21403 ( .C1(n18217), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18286), .B(
        n18213), .ZN(n18214) );
  OAI211_X1 U21404 ( .C1(n18216), .C2(n18297), .A(n18215), .B(n18214), .ZN(
        P3_U2716) );
  AOI22_X1 U21405 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18222), .ZN(n18220) );
  AOI211_X1 U21406 ( .C1(n18348), .C2(n18223), .A(n18217), .B(n18263), .ZN(
        n18218) );
  INV_X1 U21407 ( .A(n18218), .ZN(n18219) );
  OAI211_X1 U21408 ( .C1(n18221), .C2(n18297), .A(n18220), .B(n18219), .ZN(
        P3_U2717) );
  AOI22_X1 U21409 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18229), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18222), .ZN(n18226) );
  OAI211_X1 U21410 ( .C1(n18224), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18286), .B(
        n18223), .ZN(n18225) );
  OAI211_X1 U21411 ( .C1(n18227), .C2(n18297), .A(n18226), .B(n18225), .ZN(
        P3_U2718) );
  INV_X1 U21412 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U21413 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18229), .B1(n18255), .B2(
        n18228), .ZN(n18232) );
  OAI211_X1 U21414 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18234), .A(n18230), .B(
        n18286), .ZN(n18231) );
  OAI211_X1 U21415 ( .C1(n18233), .C2(n19864), .A(n18232), .B(n18231), .ZN(
        P3_U2719) );
  AOI211_X1 U21416 ( .C1(n18406), .C2(n18239), .A(n18263), .B(n18234), .ZN(
        n18235) );
  AOI21_X1 U21417 ( .B1(n18292), .B2(BUF2_REG_15__SCAN_IN), .A(n18235), .ZN(
        n18236) );
  OAI21_X1 U21418 ( .B1(n18237), .B2(n18297), .A(n18236), .ZN(P3_U2720) );
  NAND3_X1 U21419 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n18269), .ZN(n18257) );
  INV_X1 U21420 ( .A(n18257), .ZN(n18261) );
  NAND2_X1 U21421 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18261), .ZN(n18253) );
  NOR2_X1 U21422 ( .A1(n18394), .A2(n18253), .ZN(n18247) );
  NAND2_X1 U21423 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18250), .ZN(n18243) );
  INV_X1 U21424 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21486) );
  NAND2_X1 U21425 ( .A1(n18286), .A2(n18239), .ZN(n18242) );
  AOI22_X1 U21426 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18292), .B1(n18255), .B2(
        n18240), .ZN(n18241) );
  OAI221_X1 U21427 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18243), .C1(n21486), 
        .C2(n18242), .A(n18241), .ZN(P3_U2721) );
  INV_X1 U21428 ( .A(n18243), .ZN(n18246) );
  AOI21_X1 U21429 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18286), .A(n18250), .ZN(
        n18245) );
  OAI222_X1 U21430 ( .A1(n18290), .A2(n18400), .B1(n18246), .B2(n18245), .C1(
        n18297), .C2(n18244), .ZN(P3_U2722) );
  AOI21_X1 U21431 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18286), .A(n18247), .ZN(
        n18249) );
  OAI222_X1 U21432 ( .A1(n18290), .A2(n14092), .B1(n18250), .B2(n18249), .C1(
        n18297), .C2(n18248), .ZN(P3_U2723) );
  NAND2_X1 U21433 ( .A1(n18286), .A2(n18253), .ZN(n18258) );
  AOI22_X1 U21434 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18292), .B1(n18255), .B2(
        n18251), .ZN(n18252) );
  OAI221_X1 U21435 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18253), .C1(n18394), 
        .C2(n18258), .A(n18252), .ZN(P3_U2724) );
  AOI22_X1 U21436 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18292), .B1(n18255), .B2(
        n18254), .ZN(n18256) );
  OAI221_X1 U21437 ( .B1(n18258), .B2(n18392), .C1(n18258), .C2(n18257), .A(
        n18256), .ZN(P3_U2725) );
  AOI22_X1 U21438 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18269), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n18286), .ZN(n18260) );
  OAI222_X1 U21439 ( .A1(n18290), .A2(n14073), .B1(n18261), .B2(n18260), .C1(
        n18297), .C2(n18259), .ZN(P3_U2726) );
  INV_X1 U21440 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21518) );
  AOI22_X1 U21441 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18292), .B1(n18269), .B2(
        n21518), .ZN(n18265) );
  OR3_X1 U21442 ( .A1(n18263), .A2(n18262), .A3(n21518), .ZN(n18264) );
  OAI211_X1 U21443 ( .C1(n18266), .C2(n18297), .A(n18265), .B(n18264), .ZN(
        P3_U2727) );
  INV_X1 U21444 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18384) );
  NOR3_X1 U21445 ( .A1(n18380), .A2(n18277), .A3(n18281), .ZN(n18279) );
  NAND2_X1 U21446 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18279), .ZN(n18270) );
  NOR2_X1 U21447 ( .A1(n18384), .A2(n18270), .ZN(n18272) );
  AOI21_X1 U21448 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18286), .A(n18272), .ZN(
        n18268) );
  OAI222_X1 U21449 ( .A1(n18290), .A2(n14107), .B1(n18269), .B2(n18268), .C1(
        n18297), .C2(n18267), .ZN(P3_U2728) );
  INV_X1 U21450 ( .A(n18270), .ZN(n18275) );
  AOI21_X1 U21451 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18286), .A(n18275), .ZN(
        n18273) );
  OAI222_X1 U21452 ( .A1(n18290), .A2(n14069), .B1(n18273), .B2(n18272), .C1(
        n18297), .C2(n18271), .ZN(P3_U2729) );
  AOI21_X1 U21453 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18286), .A(n18279), .ZN(
        n18276) );
  OAI222_X1 U21454 ( .A1(n18290), .A2(n14101), .B1(n18276), .B2(n18275), .C1(
        n18297), .C2(n18274), .ZN(P3_U2730) );
  NOR2_X1 U21455 ( .A1(n18277), .A2(n18281), .ZN(n18283) );
  AOI21_X1 U21456 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18286), .A(n18283), .ZN(
        n18280) );
  OAI222_X1 U21457 ( .A1(n18290), .A2(n14104), .B1(n18280), .B2(n18279), .C1(
        n18297), .C2(n18278), .ZN(P3_U2731) );
  INV_X1 U21458 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18375) );
  NOR3_X1 U21459 ( .A1(n18375), .A2(n18373), .A3(n18281), .ZN(n18285) );
  AND2_X1 U21460 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18285), .ZN(n18289) );
  AOI21_X1 U21461 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18286), .A(n18289), .ZN(
        n18284) );
  OAI222_X1 U21462 ( .A1(n18290), .A2(n14097), .B1(n18284), .B2(n18283), .C1(
        n18297), .C2(n12124), .ZN(P3_U2732) );
  AOI21_X1 U21463 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18286), .A(n18285), .ZN(
        n18288) );
  OAI222_X1 U21464 ( .A1(n14082), .A2(n18290), .B1(n18289), .B2(n18288), .C1(
        n18297), .C2(n18287), .ZN(P3_U2733) );
  AOI22_X1 U21465 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18292), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n18291), .ZN(n18296) );
  NAND2_X1 U21466 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n18293) );
  OAI211_X1 U21467 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n18294), .B(n18293), .ZN(n18295) );
  OAI211_X1 U21468 ( .C1(n18298), .C2(n18297), .A(n18296), .B(n18295), .ZN(
        P3_U2734) );
  NAND2_X1 U21469 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18613), .ZN(n18335) );
  NOR2_X1 U21470 ( .A1(n18322), .A2(n18301), .ZN(P3_U2736) );
  INV_X1 U21471 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18371) );
  INV_X1 U21472 ( .A(n18340), .ZN(n18333) );
  INV_X2 U21473 ( .A(n18335), .ZN(n18338) );
  AOI22_X1 U21474 ( .A1(n18338), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18303) );
  OAI21_X1 U21475 ( .B1(n18371), .B2(n18318), .A(n18303), .ZN(P3_U2737) );
  INV_X1 U21476 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U21477 ( .A1(n18338), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18304) );
  OAI21_X1 U21478 ( .B1(n18369), .B2(n18318), .A(n18304), .ZN(P3_U2738) );
  AOI22_X1 U21479 ( .A1(n18338), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18305) );
  OAI21_X1 U21480 ( .B1(n18367), .B2(n18318), .A(n18305), .ZN(P3_U2739) );
  INV_X1 U21481 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18365) );
  AOI22_X1 U21482 ( .A1(n18338), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18306) );
  OAI21_X1 U21483 ( .B1(n18365), .B2(n18318), .A(n18306), .ZN(P3_U2740) );
  AOI22_X1 U21484 ( .A1(n18338), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18307) );
  OAI21_X1 U21485 ( .B1(n18363), .B2(n18318), .A(n18307), .ZN(P3_U2741) );
  AOI22_X1 U21486 ( .A1(n18338), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18308) );
  OAI21_X1 U21487 ( .B1(n10411), .B2(n18318), .A(n18308), .ZN(P3_U2742) );
  INV_X1 U21488 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18360) );
  AOI22_X1 U21489 ( .A1(n18338), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18309) );
  OAI21_X1 U21490 ( .B1(n18360), .B2(n18318), .A(n18309), .ZN(P3_U2743) );
  INV_X1 U21491 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18358) );
  AOI22_X1 U21492 ( .A1(n18338), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18310) );
  OAI21_X1 U21493 ( .B1(n18358), .B2(n18318), .A(n18310), .ZN(P3_U2744) );
  AOI22_X1 U21494 ( .A1(n18338), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18311) );
  OAI21_X1 U21495 ( .B1(n18356), .B2(n18318), .A(n18311), .ZN(P3_U2745) );
  AOI22_X1 U21496 ( .A1(n18338), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18312) );
  OAI21_X1 U21497 ( .B1(n18354), .B2(n18318), .A(n18312), .ZN(P3_U2746) );
  AOI22_X1 U21498 ( .A1(n18338), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18313) );
  OAI21_X1 U21499 ( .B1(n18352), .B2(n18318), .A(n18313), .ZN(P3_U2747) );
  INV_X1 U21500 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U21501 ( .A1(n18338), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18314) );
  OAI21_X1 U21502 ( .B1(n18350), .B2(n18318), .A(n18314), .ZN(P3_U2748) );
  AOI22_X1 U21503 ( .A1(n18338), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18315) );
  OAI21_X1 U21504 ( .B1(n18348), .B2(n18318), .A(n18315), .ZN(P3_U2749) );
  INV_X1 U21505 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U21506 ( .A1(n18338), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18316) );
  OAI21_X1 U21507 ( .B1(n18346), .B2(n18318), .A(n18316), .ZN(P3_U2750) );
  INV_X1 U21508 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n21640) );
  AOI22_X1 U21509 ( .A1(n18338), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18317) );
  OAI21_X1 U21510 ( .B1(n21640), .B2(n18318), .A(n18317), .ZN(P3_U2751) );
  AOI22_X1 U21511 ( .A1(n18338), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18319) );
  OAI21_X1 U21512 ( .B1(n18406), .B2(n18340), .A(n18319), .ZN(P3_U2752) );
  AOI22_X1 U21513 ( .A1(n18338), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18320) );
  OAI21_X1 U21514 ( .B1(n21486), .B2(n18340), .A(n18320), .ZN(P3_U2753) );
  INV_X1 U21515 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n21555) );
  AOI22_X1 U21516 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18333), .B1(n18338), 
        .B2(P3_LWORD_REG_13__SCAN_IN), .ZN(n18321) );
  OAI21_X1 U21517 ( .B1(n21555), .B2(n18322), .A(n18321), .ZN(P3_U2754) );
  INV_X1 U21518 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18396) );
  AOI22_X1 U21519 ( .A1(P3_LWORD_REG_12__SCAN_IN), .A2(n18338), .B1(n18329), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18323) );
  OAI21_X1 U21520 ( .B1(n18396), .B2(n18340), .A(n18323), .ZN(P3_U2755) );
  AOI22_X1 U21521 ( .A1(n18338), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18324) );
  OAI21_X1 U21522 ( .B1(n18394), .B2(n18340), .A(n18324), .ZN(P3_U2756) );
  AOI22_X1 U21523 ( .A1(n18338), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18325) );
  OAI21_X1 U21524 ( .B1(n18392), .B2(n18340), .A(n18325), .ZN(P3_U2757) );
  AOI22_X1 U21525 ( .A1(n18338), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18326) );
  OAI21_X1 U21526 ( .B1(n18390), .B2(n18340), .A(n18326), .ZN(P3_U2758) );
  AOI22_X1 U21527 ( .A1(P3_LWORD_REG_8__SCAN_IN), .A2(n18338), .B1(n18329), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18327) );
  OAI21_X1 U21528 ( .B1(n21518), .B2(n18340), .A(n18327), .ZN(P3_U2759) );
  INV_X1 U21529 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18386) );
  AOI22_X1 U21530 ( .A1(n18338), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18328) );
  OAI21_X1 U21531 ( .B1(n18386), .B2(n18340), .A(n18328), .ZN(P3_U2760) );
  AOI22_X1 U21532 ( .A1(n18338), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18330) );
  OAI21_X1 U21533 ( .B1(n18384), .B2(n18340), .A(n18330), .ZN(P3_U2761) );
  INV_X1 U21534 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18382) );
  AOI22_X1 U21535 ( .A1(n18338), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18331) );
  OAI21_X1 U21536 ( .B1(n18382), .B2(n18340), .A(n18331), .ZN(P3_U2762) );
  AOI22_X1 U21537 ( .A1(n18338), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18332) );
  OAI21_X1 U21538 ( .B1(n18380), .B2(n18340), .A(n18332), .ZN(P3_U2763) );
  INV_X1 U21539 ( .A(P3_LWORD_REG_3__SCAN_IN), .ZN(n21536) );
  AOI22_X1 U21540 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18333), .B1(n18329), .B2(
        P3_DATAO_REG_3__SCAN_IN), .ZN(n18334) );
  OAI21_X1 U21541 ( .B1(n21536), .B2(n18335), .A(n18334), .ZN(P3_U2764) );
  INV_X1 U21542 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18377) );
  AOI22_X1 U21543 ( .A1(n18338), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18336) );
  OAI21_X1 U21544 ( .B1(n18377), .B2(n18340), .A(n18336), .ZN(P3_U2765) );
  AOI22_X1 U21545 ( .A1(n18338), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18337) );
  OAI21_X1 U21546 ( .B1(n18375), .B2(n18340), .A(n18337), .ZN(P3_U2766) );
  AOI22_X1 U21547 ( .A1(n18338), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18329), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18339) );
  OAI21_X1 U21548 ( .B1(n18373), .B2(n18340), .A(n18339), .ZN(P3_U2767) );
  NAND2_X1 U21549 ( .A1(n18343), .A2(n18388), .ZN(n18399) );
  INV_X2 U21550 ( .A(n18388), .ZN(n18402) );
  AOI22_X1 U21551 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18402), .ZN(n18344) );
  OAI21_X1 U21552 ( .B1(n21640), .B2(n18405), .A(n18344), .ZN(P3_U2768) );
  AOI22_X1 U21553 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18402), .ZN(n18345) );
  OAI21_X1 U21554 ( .B1(n18346), .B2(n18405), .A(n18345), .ZN(P3_U2769) );
  AOI22_X1 U21555 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18402), .ZN(n18347) );
  OAI21_X1 U21556 ( .B1(n18348), .B2(n18405), .A(n18347), .ZN(P3_U2770) );
  AOI22_X1 U21557 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18402), .ZN(n18349) );
  OAI21_X1 U21558 ( .B1(n18350), .B2(n18405), .A(n18349), .ZN(P3_U2771) );
  AOI22_X1 U21559 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18402), .ZN(n18351) );
  OAI21_X1 U21560 ( .B1(n18352), .B2(n18405), .A(n18351), .ZN(P3_U2772) );
  AOI22_X1 U21561 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18402), .ZN(n18353) );
  OAI21_X1 U21562 ( .B1(n18354), .B2(n18405), .A(n18353), .ZN(P3_U2773) );
  AOI22_X1 U21563 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18402), .ZN(n18355) );
  OAI21_X1 U21564 ( .B1(n18356), .B2(n18405), .A(n18355), .ZN(P3_U2774) );
  AOI22_X1 U21565 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18402), .ZN(n18357) );
  OAI21_X1 U21566 ( .B1(n18358), .B2(n18405), .A(n18357), .ZN(P3_U2775) );
  AOI22_X1 U21567 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18402), .ZN(n18359) );
  OAI21_X1 U21568 ( .B1(n18360), .B2(n18405), .A(n18359), .ZN(P3_U2776) );
  AOI22_X1 U21569 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18402), .ZN(n18361) );
  OAI21_X1 U21570 ( .B1(n10411), .B2(n18405), .A(n18361), .ZN(P3_U2777) );
  AOI22_X1 U21571 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18402), .ZN(n18362) );
  OAI21_X1 U21572 ( .B1(n18363), .B2(n18405), .A(n18362), .ZN(P3_U2778) );
  AOI22_X1 U21573 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18402), .ZN(n18364) );
  OAI21_X1 U21574 ( .B1(n18365), .B2(n18405), .A(n18364), .ZN(P3_U2779) );
  AOI22_X1 U21575 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18402), .ZN(n18366) );
  OAI21_X1 U21576 ( .B1(n18367), .B2(n18405), .A(n18366), .ZN(P3_U2780) );
  AOI22_X1 U21577 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18402), .ZN(n18368) );
  OAI21_X1 U21578 ( .B1(n18369), .B2(n18405), .A(n18368), .ZN(P3_U2781) );
  AOI22_X1 U21579 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18403), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18402), .ZN(n18370) );
  OAI21_X1 U21580 ( .B1(n18371), .B2(n18405), .A(n18370), .ZN(P3_U2782) );
  AOI22_X1 U21581 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18402), .ZN(n18372) );
  OAI21_X1 U21582 ( .B1(n18373), .B2(n18405), .A(n18372), .ZN(P3_U2783) );
  AOI22_X1 U21583 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18402), .ZN(n18374) );
  OAI21_X1 U21584 ( .B1(n18375), .B2(n18405), .A(n18374), .ZN(P3_U2784) );
  AOI22_X1 U21585 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18402), .ZN(n18376) );
  OAI21_X1 U21586 ( .B1(n18377), .B2(n18405), .A(n18376), .ZN(P3_U2785) );
  AOI22_X1 U21587 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18403), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n18397), .ZN(n18378) );
  OAI21_X1 U21588 ( .B1(n18388), .B2(n21536), .A(n18378), .ZN(P3_U2786) );
  AOI22_X1 U21589 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18402), .ZN(n18379) );
  OAI21_X1 U21590 ( .B1(n18380), .B2(n18405), .A(n18379), .ZN(P3_U2787) );
  AOI22_X1 U21591 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18402), .ZN(n18381) );
  OAI21_X1 U21592 ( .B1(n18382), .B2(n18405), .A(n18381), .ZN(P3_U2788) );
  AOI22_X1 U21593 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18402), .ZN(n18383) );
  OAI21_X1 U21594 ( .B1(n18384), .B2(n18405), .A(n18383), .ZN(P3_U2789) );
  AOI22_X1 U21595 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18402), .ZN(n18385) );
  OAI21_X1 U21596 ( .B1(n18386), .B2(n18405), .A(n18385), .ZN(P3_U2790) );
  INV_X1 U21597 ( .A(P3_LWORD_REG_8__SCAN_IN), .ZN(n21527) );
  AOI22_X1 U21598 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18403), .B1(
        P3_EAX_REG_8__SCAN_IN), .B2(n18397), .ZN(n18387) );
  OAI21_X1 U21599 ( .B1(n18388), .B2(n21527), .A(n18387), .ZN(P3_U2791) );
  AOI22_X1 U21600 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18402), .ZN(n18389) );
  OAI21_X1 U21601 ( .B1(n18390), .B2(n18405), .A(n18389), .ZN(P3_U2792) );
  AOI22_X1 U21602 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18402), .ZN(n18391) );
  OAI21_X1 U21603 ( .B1(n18392), .B2(n18405), .A(n18391), .ZN(P3_U2793) );
  AOI22_X1 U21604 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18402), .ZN(n18393) );
  OAI21_X1 U21605 ( .B1(n18394), .B2(n18405), .A(n18393), .ZN(P3_U2794) );
  AOI22_X1 U21606 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18402), .ZN(n18395) );
  OAI21_X1 U21607 ( .B1(n18396), .B2(n18405), .A(n18395), .ZN(P3_U2795) );
  AOI22_X1 U21608 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18397), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18402), .ZN(n18398) );
  OAI21_X1 U21609 ( .B1(n18400), .B2(n18399), .A(n18398), .ZN(P3_U2796) );
  AOI22_X1 U21610 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18402), .ZN(n18401) );
  OAI21_X1 U21611 ( .B1(n21486), .B2(n18405), .A(n18401), .ZN(P3_U2797) );
  AOI22_X1 U21612 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18403), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18402), .ZN(n18404) );
  OAI21_X1 U21613 ( .B1(n18406), .B2(n18405), .A(n18404), .ZN(P3_U2798) );
  OAI21_X1 U21614 ( .B1(n18408), .B2(n18773), .A(n18772), .ZN(n18409) );
  AOI21_X1 U21615 ( .B1(n18741), .B2(n18407), .A(n18409), .ZN(n18442) );
  OAI21_X1 U21616 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n9690), .A(
        n18442), .ZN(n18428) );
  NOR2_X1 U21617 ( .A1(n18588), .A2(n18407), .ZN(n18434) );
  OAI211_X1 U21618 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18434), .B(n18410), .ZN(n18412) );
  OAI211_X1 U21619 ( .C1(n18626), .C2(n18413), .A(n18412), .B(n18411), .ZN(
        n18414) );
  AOI21_X1 U21620 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18428), .A(
        n18414), .ZN(n18426) );
  NOR2_X1 U21621 ( .A1(n18756), .A2(n18684), .ZN(n18529) );
  INV_X1 U21622 ( .A(n18529), .ZN(n18417) );
  AOI22_X1 U21623 ( .A1(n18756), .A2(n18416), .B1(n18684), .B2(n18415), .ZN(
        n18446) );
  NAND2_X1 U21624 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18446), .ZN(
        n18435) );
  NAND3_X1 U21625 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18417), .A3(
        n18435), .ZN(n18425) );
  NAND3_X1 U21626 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18436), .A3(
        n18418), .ZN(n18424) );
  AOI211_X1 U21627 ( .C1(n18421), .C2(n18420), .A(n18687), .B(n18419), .ZN(
        n18422) );
  INV_X1 U21628 ( .A(n18422), .ZN(n18423) );
  NAND4_X1 U21629 ( .A1(n18426), .A2(n18425), .A3(n18424), .A4(n18423), .ZN(
        P3_U2802) );
  AOI22_X1 U21630 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18428), .B1(
        n18577), .B2(n18427), .ZN(n18439) );
  INV_X1 U21631 ( .A(n18429), .ZN(n18431) );
  NAND2_X1 U21632 ( .A1(n18431), .A2(n18430), .ZN(n18432) );
  XOR2_X1 U21633 ( .A(n18573), .B(n18432), .Z(n18781) );
  AOI22_X1 U21634 ( .A1(n18669), .A2(n18781), .B1(n18434), .B2(n18433), .ZN(
        n18438) );
  OAI21_X1 U21635 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18436), .A(
        n18435), .ZN(n18437) );
  NAND2_X1 U21636 ( .A1(n18963), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18782) );
  NAND4_X1 U21637 ( .A1(n18439), .A2(n18438), .A3(n18437), .A4(n18782), .ZN(
        P3_U2803) );
  AOI21_X1 U21638 ( .B1(n19455), .B2(n18440), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18441) );
  OAI22_X1 U21639 ( .A1(n18761), .A2(n18443), .B1(n18442), .B2(n18441), .ZN(
        n18448) );
  OAI22_X1 U21640 ( .A1(n18446), .A2(n18445), .B1(n18444), .B2(n18687), .ZN(
        n18447) );
  AOI211_X1 U21641 ( .C1(n18963), .C2(P3_REIP_REG_26__SCAN_IN), .A(n18448), 
        .B(n18447), .ZN(n18449) );
  OAI21_X1 U21642 ( .B1(n18469), .B2(n18450), .A(n18449), .ZN(P3_U2804) );
  NAND2_X1 U21643 ( .A1(n19455), .A2(n18451), .ZN(n18479) );
  OAI211_X1 U21644 ( .C1(n18452), .C2(n18773), .A(n18772), .B(n18479), .ZN(
        n18478) );
  AOI22_X1 U21645 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18478), .B1(
        n18577), .B2(n18453), .ZN(n18463) );
  AOI21_X1 U21646 ( .B1(n18455), .B2(n18673), .A(n18454), .ZN(n18456) );
  XOR2_X1 U21647 ( .A(n18456), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18798) );
  NAND3_X1 U21648 ( .A1(n18806), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n9779), .ZN(n18457) );
  XOR2_X1 U21649 ( .A(n18457), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18795) );
  NAND3_X1 U21650 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18887), .A3(
        n18806), .ZN(n18458) );
  XOR2_X1 U21651 ( .A(n18458), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18794) );
  OAI22_X1 U21652 ( .A1(n18777), .A2(n18795), .B1(n18620), .B2(n18794), .ZN(
        n18459) );
  AOI21_X1 U21653 ( .B1(n18669), .B2(n18798), .A(n18459), .ZN(n18462) );
  NAND2_X1 U21654 ( .A1(n18963), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18792) );
  NOR2_X1 U21655 ( .A1(n18588), .A2(n18451), .ZN(n18466) );
  OAI211_X1 U21656 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18466), .B(n18460), .ZN(n18461) );
  NAND4_X1 U21657 ( .A1(n18463), .A2(n18462), .A3(n18792), .A4(n18461), .ZN(
        P3_U2805) );
  INV_X1 U21658 ( .A(n18464), .ZN(n18473) );
  NOR2_X1 U21659 ( .A1(n19055), .A2(n19640), .ZN(n18465) );
  AOI221_X1 U21660 ( .B1(n18466), .B2(n21686), .C1(n18478), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18465), .ZN(n18472) );
  NOR2_X1 U21661 ( .A1(n18800), .A2(n18620), .ZN(n18491) );
  NOR2_X1 U21662 ( .A1(n18802), .A2(n18777), .ZN(n18489) );
  AOI21_X1 U21663 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18468), .A(
        n18467), .ZN(n18808) );
  OAI22_X1 U21664 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18469), .B1(
        n18808), .B2(n18687), .ZN(n18470) );
  AOI221_X1 U21665 ( .B1(n18491), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), 
        .C1(n18489), .C2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n18470), .ZN(
        n18471) );
  OAI211_X1 U21666 ( .C1(n18626), .C2(n18473), .A(n18472), .B(n18471), .ZN(
        P3_U2806) );
  INV_X1 U21667 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18828) );
  OAI21_X1 U21668 ( .B1(n18557), .B2(n18474), .A(n18501), .ZN(n18475) );
  OAI211_X1 U21669 ( .C1(n18573), .C2(n18828), .A(n18476), .B(n18475), .ZN(
        n18477) );
  XOR2_X1 U21670 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18477), .Z(
        n18815) );
  NOR2_X1 U21671 ( .A1(n19055), .A2(n19636), .ZN(n18484) );
  OAI21_X1 U21672 ( .B1(n18521), .B2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n18478), .ZN(n18481) );
  OAI22_X1 U21673 ( .A1(n18482), .A2(n18481), .B1(n18480), .B2(n18479), .ZN(
        n18483) );
  AOI211_X1 U21674 ( .C1(n18577), .C2(n18485), .A(n18484), .B(n18483), .ZN(
        n18493) );
  NAND2_X1 U21675 ( .A1(n18805), .A2(n18486), .ZN(n18490) );
  NAND2_X1 U21676 ( .A1(n18805), .A2(n18487), .ZN(n18488) );
  AOI22_X1 U21677 ( .A1(n18491), .A2(n18490), .B1(n18489), .B2(n18488), .ZN(
        n18492) );
  OAI211_X1 U21678 ( .C1(n18687), .C2(n18815), .A(n18493), .B(n18492), .ZN(
        P3_U2807) );
  INV_X1 U21679 ( .A(n18741), .ZN(n18674) );
  NAND2_X1 U21680 ( .A1(n18613), .A2(n18494), .ZN(n18495) );
  OAI211_X1 U21681 ( .C1(n18496), .C2(n18674), .A(n18772), .B(n18495), .ZN(
        n18527) );
  AOI21_X1 U21682 ( .B1(n18521), .B2(n21610), .A(n18527), .ZN(n18510) );
  INV_X1 U21683 ( .A(n18588), .ZN(n18624) );
  NAND3_X1 U21684 ( .A1(n18496), .A2(n18624), .A3(n10690), .ZN(n18509) );
  AOI21_X1 U21685 ( .B1(n18510), .B2(n18509), .A(n18497), .ZN(n18499) );
  NOR3_X1 U21686 ( .A1(n18588), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(
        n9782), .ZN(n18498) );
  AOI211_X1 U21687 ( .C1(n18500), .C2(n18577), .A(n18499), .B(n18498), .ZN(
        n18506) );
  OAI22_X1 U21688 ( .A1(n18777), .A2(n9779), .B1(n18620), .B2(n18887), .ZN(
        n18581) );
  INV_X1 U21689 ( .A(n18581), .ZN(n18528) );
  OAI21_X1 U21690 ( .B1(n18529), .B2(n18821), .A(n18528), .ZN(n18517) );
  AOI221_X1 U21691 ( .B1(n18502), .B2(n18501), .C1(n18823), .C2(n18501), .A(
        n18530), .ZN(n18503) );
  XOR2_X1 U21692 ( .A(n18503), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n18826) );
  AOI22_X1 U21693 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18517), .B1(
        n18669), .B2(n18826), .ZN(n18505) );
  NAND2_X1 U21694 ( .A1(n19040), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18827) );
  NAND3_X1 U21695 ( .A1(n18821), .A2(n9722), .A3(n18828), .ZN(n18504) );
  NAND4_X1 U21696 ( .A1(n18506), .A2(n18505), .A3(n18827), .A4(n18504), .ZN(
        P3_U2808) );
  NAND2_X1 U21697 ( .A1(n18838), .A2(n18516), .ZN(n18843) );
  NAND2_X1 U21698 ( .A1(n18507), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18817) );
  INV_X1 U21699 ( .A(n18817), .ZN(n18833) );
  NAND2_X1 U21700 ( .A1(n18833), .A2(n9722), .ZN(n18549) );
  NAND2_X1 U21701 ( .A1(n19040), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18508) );
  OAI211_X1 U21702 ( .C1(n18510), .C2(n10690), .A(n18509), .B(n18508), .ZN(
        n18511) );
  AOI21_X1 U21703 ( .B1(n18577), .B2(n18512), .A(n18511), .ZN(n18519) );
  NAND3_X1 U21704 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18573), .A3(
        n18513), .ZN(n18531) );
  INV_X1 U21705 ( .A(n18531), .ZN(n18543) );
  AOI22_X1 U21706 ( .A1(n18838), .A2(n18543), .B1(n18557), .B2(n18514), .ZN(
        n18515) );
  XOR2_X1 U21707 ( .A(n18516), .B(n18515), .Z(n18830) );
  AOI22_X1 U21708 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18517), .B1(
        n18669), .B2(n18830), .ZN(n18518) );
  OAI211_X1 U21709 ( .C1(n18843), .C2(n18549), .A(n18519), .B(n18518), .ZN(
        P3_U2809) );
  NAND2_X1 U21710 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21613), .ZN(
        n18850) );
  OAI21_X1 U21711 ( .B1(n19221), .B2(n18520), .A(n21610), .ZN(n18526) );
  NOR2_X1 U21712 ( .A1(n19055), .A2(n21658), .ZN(n18525) );
  INV_X1 U21713 ( .A(n18522), .ZN(n18523) );
  AOI21_X1 U21714 ( .B1(n18626), .B2(n9690), .A(n18523), .ZN(n18524) );
  AOI211_X1 U21715 ( .C1(n18527), .C2(n18526), .A(n18525), .B(n18524), .ZN(
        n18535) );
  NOR2_X1 U21716 ( .A1(n18545), .A2(n18817), .ZN(n18845) );
  OAI21_X1 U21717 ( .B1(n18529), .B2(n18845), .A(n18528), .ZN(n18546) );
  AOI221_X1 U21718 ( .B1(n18545), .B2(n18532), .C1(n18531), .C2(n18532), .A(
        n18530), .ZN(n18533) );
  XNOR2_X1 U21719 ( .A(n21613), .B(n18533), .ZN(n18844) );
  AOI22_X1 U21720 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18546), .B1(
        n18669), .B2(n18844), .ZN(n18534) );
  OAI211_X1 U21721 ( .C1(n18850), .C2(n18549), .A(n18535), .B(n18534), .ZN(
        P3_U2810) );
  INV_X1 U21722 ( .A(n18536), .ZN(n18538) );
  AOI21_X1 U21723 ( .B1(n18741), .B2(n18538), .A(n18728), .ZN(n18563) );
  OAI21_X1 U21724 ( .B1(n18537), .B2(n18773), .A(n18563), .ZN(n18552) );
  NAND2_X1 U21725 ( .A1(n19040), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18853) );
  NOR2_X1 U21726 ( .A1(n18588), .A2(n18538), .ZN(n18554) );
  OAI211_X1 U21727 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18554), .B(n18539), .ZN(n18540) );
  OAI211_X1 U21728 ( .C1(n18626), .C2(n18541), .A(n18853), .B(n18540), .ZN(
        n18542) );
  AOI21_X1 U21729 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18552), .A(
        n18542), .ZN(n18548) );
  AOI21_X1 U21730 ( .B1(n18555), .B2(n18557), .A(n18543), .ZN(n18544) );
  XOR2_X1 U21731 ( .A(n18545), .B(n18544), .Z(n18851) );
  AOI22_X1 U21732 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18546), .B1(
        n18669), .B2(n18851), .ZN(n18547) );
  OAI211_X1 U21733 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18549), .A(
        n18548), .B(n18547), .ZN(P3_U2811) );
  AOI21_X1 U21734 ( .B1(n9722), .B2(n18859), .A(n18581), .ZN(n18567) );
  INV_X1 U21735 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18560) );
  OAI22_X1 U21736 ( .A1(n19055), .A2(n19629), .B1(n18626), .B2(n18550), .ZN(
        n18551) );
  AOI221_X1 U21737 ( .B1(n18554), .B2(n18553), .C1(n18552), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18551), .ZN(n18559) );
  AOI21_X1 U21738 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18573), .A(
        n18555), .ZN(n18556) );
  XOR2_X1 U21739 ( .A(n18557), .B(n18556), .Z(n18867) );
  NOR2_X1 U21740 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18859), .ZN(
        n18866) );
  AOI22_X1 U21741 ( .A1(n18669), .A2(n18867), .B1(n18866), .B2(n9722), .ZN(
        n18558) );
  OAI211_X1 U21742 ( .C1(n18567), .C2(n18560), .A(n18559), .B(n18558), .ZN(
        P3_U2812) );
  AOI21_X1 U21743 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18562), .A(
        n18561), .ZN(n18874) );
  AOI221_X1 U21744 ( .B1(n19221), .B2(n18565), .C1(n18564), .C2(n18565), .A(
        n18563), .ZN(n18570) );
  AOI21_X1 U21745 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n9722), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18566) );
  OAI22_X1 U21746 ( .A1(n18761), .A2(n18568), .B1(n18567), .B2(n18566), .ZN(
        n18569) );
  AOI211_X1 U21747 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n19040), .A(n18570), 
        .B(n18569), .ZN(n18571) );
  OAI21_X1 U21748 ( .B1(n18874), .B2(n18687), .A(n18571), .ZN(P3_U2813) );
  NAND2_X1 U21749 ( .A1(n18573), .A2(n18943), .ZN(n18659) );
  OAI22_X1 U21750 ( .A1(n18573), .A2(n18572), .B1(n18659), .B2(n18865), .ZN(
        n18574) );
  XOR2_X1 U21751 ( .A(n18881), .B(n18574), .Z(n18886) );
  OAI211_X1 U21752 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17395), .B(n18624), .ZN(n18579) );
  AOI21_X1 U21753 ( .B1(n18741), .B2(n18587), .A(n18728), .ZN(n18600) );
  OAI21_X1 U21754 ( .B1(n18575), .B2(n18773), .A(n18600), .ZN(n18591) );
  AOI22_X1 U21755 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18591), .B1(
        n18577), .B2(n18576), .ZN(n18578) );
  NAND2_X1 U21756 ( .A1(n18963), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18884) );
  OAI211_X1 U21757 ( .C1(n10937), .C2(n18579), .A(n18578), .B(n18884), .ZN(
        n18580) );
  AOI221_X1 U21758 ( .B1(n9722), .B2(n18881), .C1(n18581), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18580), .ZN(n18582) );
  OAI21_X1 U21759 ( .B1(n18886), .B2(n18687), .A(n18582), .ZN(P3_U2814) );
  INV_X1 U21760 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18929) );
  NOR3_X1 U21761 ( .A1(n18910), .A2(n18920), .A3(n18645), .ZN(n18584) );
  NAND2_X1 U21762 ( .A1(n9746), .A2(n18673), .ZN(n18660) );
  NOR2_X1 U21763 ( .A1(n18583), .A2(n18660), .ZN(n18631) );
  AOI22_X1 U21764 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18584), .B1(
        n18631), .B2(n18905), .ZN(n18585) );
  AOI221_X1 U21765 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18929), 
        .C1(n18673), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18585), .ZN(
        n18586) );
  XOR2_X1 U21766 ( .A(n18900), .B(n18586), .Z(n18893) );
  NOR2_X1 U21767 ( .A1(n18588), .A2(n18587), .ZN(n18593) );
  OAI22_X1 U21768 ( .A1(n19055), .A2(n19623), .B1(n18626), .B2(n18589), .ZN(
        n18590) );
  AOI221_X1 U21769 ( .B1(n18593), .B2(n18592), .C1(n18591), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18590), .ZN(n18597) );
  NOR2_X1 U21770 ( .A1(n18887), .A2(n18620), .ZN(n18595) );
  NOR2_X1 U21771 ( .A1(n10766), .A2(n18645), .ZN(n18599) );
  NAND2_X1 U21772 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18599), .ZN(
        n18598) );
  NAND2_X1 U21773 ( .A1(n18900), .A2(n18598), .ZN(n18891) );
  NOR2_X1 U21774 ( .A1(n9779), .A2(n18777), .ZN(n18594) );
  OR2_X1 U21775 ( .A1(n18605), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18896) );
  AOI22_X1 U21776 ( .A1(n18595), .A2(n18891), .B1(n18594), .B2(n18896), .ZN(
        n18596) );
  OAI211_X1 U21777 ( .C1(n18687), .C2(n18893), .A(n18597), .B(n18596), .ZN(
        P3_U2815) );
  OAI21_X1 U21778 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18599), .A(
        n18598), .ZN(n18917) );
  AOI221_X1 U21779 ( .B1(n19221), .B2(n18602), .C1(n18601), .C2(n18602), .A(
        n18600), .ZN(n18603) );
  NOR2_X1 U21780 ( .A1(n19055), .A2(n19621), .ZN(n18912) );
  AOI211_X1 U21781 ( .C1(n18604), .C2(n18767), .A(n18603), .B(n18912), .ZN(
        n18611) );
  AOI21_X1 U21782 ( .B1(n18910), .B2(n18606), .A(n18605), .ZN(n18913) );
  INV_X1 U21783 ( .A(n18607), .ZN(n18608) );
  OAI22_X1 U21784 ( .A1(n10766), .A2(n18659), .B1(n18608), .B2(n18660), .ZN(
        n18609) );
  XOR2_X1 U21785 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18609), .Z(
        n18914) );
  AOI22_X1 U21786 ( .A1(n18756), .A2(n18913), .B1(n18669), .B2(n18914), .ZN(
        n18610) );
  OAI211_X1 U21787 ( .C1(n18620), .C2(n18917), .A(n18611), .B(n18610), .ZN(
        P3_U2816) );
  INV_X1 U21788 ( .A(n18619), .ZN(n18901) );
  NAND2_X1 U21789 ( .A1(n18901), .A2(n18905), .ZN(n18928) );
  AOI21_X1 U21790 ( .B1(n18613), .B2(n18612), .A(n18728), .ZN(n18614) );
  OAI21_X1 U21791 ( .B1(n18641), .B2(n18674), .A(n18614), .ZN(n18628) );
  NOR2_X1 U21792 ( .A1(n19055), .A2(n19619), .ZN(n18618) );
  OAI211_X1 U21793 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18641), .B(n18624), .ZN(n18616) );
  OAI22_X1 U21794 ( .A1(n9721), .A2(n18616), .B1(n18615), .B2(n18626), .ZN(
        n18617) );
  AOI211_X1 U21795 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18628), .A(
        n18618), .B(n18617), .ZN(n18623) );
  NOR2_X1 U21796 ( .A1(n18619), .A2(n18645), .ZN(n18924) );
  NOR2_X1 U21797 ( .A1(n18619), .A2(n18940), .ZN(n18919) );
  OAI22_X1 U21798 ( .A1(n18924), .A2(n18620), .B1(n18919), .B2(n18777), .ZN(
        n18633) );
  NOR2_X1 U21799 ( .A1(n18920), .A2(n18659), .ZN(n18630) );
  AOI22_X1 U21800 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18630), .B1(
        n18631), .B2(n18929), .ZN(n18621) );
  XOR2_X1 U21801 ( .A(n18905), .B(n18621), .Z(n18918) );
  AOI22_X1 U21802 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18633), .B1(
        n18669), .B2(n18918), .ZN(n18622) );
  OAI211_X1 U21803 ( .C1(n18672), .C2(n18928), .A(n18623), .B(n18622), .ZN(
        P3_U2817) );
  NAND2_X1 U21804 ( .A1(n18948), .A2(n18929), .ZN(n18636) );
  AND2_X1 U21805 ( .A1(n18624), .A2(n18641), .ZN(n18629) );
  NAND2_X1 U21806 ( .A1(n18963), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18933) );
  OAI21_X1 U21807 ( .B1(n18626), .B2(n18625), .A(n18933), .ZN(n18627) );
  AOI221_X1 U21808 ( .B1(n18629), .B2(n21679), .C1(n18628), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18627), .ZN(n18635) );
  NOR2_X1 U21809 ( .A1(n18631), .A2(n18630), .ZN(n18632) );
  XOR2_X1 U21810 ( .A(n18632), .B(n18929), .Z(n18932) );
  AOI22_X1 U21811 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18633), .B1(
        n18669), .B2(n18932), .ZN(n18634) );
  OAI211_X1 U21812 ( .C1(n18672), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2818) );
  NAND2_X1 U21813 ( .A1(n18946), .A2(n18637), .ZN(n18953) );
  NOR3_X1 U21814 ( .A1(n19221), .A2(n18716), .A3(n18638), .ZN(n18704) );
  NAND2_X1 U21815 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18704), .ZN(
        n18662) );
  NOR2_X1 U21816 ( .A1(n18639), .A2(n18662), .ZN(n18666) );
  NAND2_X1 U21817 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18666), .ZN(
        n18650) );
  INV_X1 U21818 ( .A(n18699), .ZN(n18769) );
  NAND2_X1 U21819 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18769), .ZN(
        n18640) );
  AOI22_X1 U21820 ( .A1(n19455), .A2(n18641), .B1(n18650), .B2(n18640), .ZN(
        n18643) );
  NOR2_X1 U21821 ( .A1(n19055), .A2(n21642), .ZN(n18642) );
  AOI211_X1 U21822 ( .C1(n18644), .C2(n18767), .A(n18643), .B(n18642), .ZN(
        n18649) );
  AOI22_X1 U21823 ( .A1(n18756), .A2(n18940), .B1(n18684), .B2(n18645), .ZN(
        n18671) );
  OAI21_X1 U21824 ( .B1(n18946), .B2(n18672), .A(n18671), .ZN(n18647) );
  OAI33_X1 U21825 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n18660), .B1(n21474), .B2(
        n18659), .B3(n18966), .ZN(n18646) );
  XOR2_X1 U21826 ( .A(n18646), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18936) );
  AOI22_X1 U21827 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18647), .B1(
        n18669), .B2(n18936), .ZN(n18648) );
  OAI211_X1 U21828 ( .C1(n18672), .C2(n18953), .A(n18649), .B(n18648), .ZN(
        P3_U2819) );
  OAI211_X1 U21829 ( .C1(n18666), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18769), .B(n18650), .ZN(n18651) );
  OAI21_X1 U21830 ( .B1(n18761), .B2(n18652), .A(n18651), .ZN(n18653) );
  AOI21_X1 U21831 ( .B1(n18963), .B2(P3_REIP_REG_10__SCAN_IN), .A(n18653), 
        .ZN(n18658) );
  AOI22_X1 U21832 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18659), .B1(
        n18660), .B2(n18966), .ZN(n18654) );
  XOR2_X1 U21833 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18654), .Z(
        n18957) );
  AOI21_X1 U21834 ( .B1(n21474), .B2(n18966), .A(n18946), .ZN(n18656) );
  AOI22_X1 U21835 ( .A1(n18669), .A2(n18957), .B1(n18656), .B2(n18655), .ZN(
        n18657) );
  OAI211_X1 U21836 ( .C1(n18671), .C2(n21474), .A(n18658), .B(n18657), .ZN(
        P3_U2820) );
  NAND2_X1 U21837 ( .A1(n18660), .A2(n18659), .ZN(n18661) );
  XOR2_X1 U21838 ( .A(n18661), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18961) );
  NOR2_X1 U21839 ( .A1(n19055), .A2(n19612), .ZN(n18668) );
  INV_X1 U21840 ( .A(n18662), .ZN(n18691) );
  AOI22_X1 U21841 ( .A1(n18663), .A2(n18691), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18769), .ZN(n18665) );
  OAI22_X1 U21842 ( .A1(n18666), .A2(n18665), .B1(n18761), .B2(n18664), .ZN(
        n18667) );
  AOI211_X1 U21843 ( .C1(n18669), .C2(n18961), .A(n18668), .B(n18667), .ZN(
        n18670) );
  OAI221_X1 U21844 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18672), .C1(
        n18966), .C2(n18671), .A(n18670), .ZN(P3_U2821) );
  NOR2_X1 U21845 ( .A1(n18943), .A2(n9746), .ZN(n18683) );
  INV_X1 U21846 ( .A(n18683), .ZN(n18968) );
  XOR2_X1 U21847 ( .A(n18968), .B(n18673), .Z(n18971) );
  OAI21_X1 U21848 ( .B1(n18675), .B2(n18674), .A(n18772), .ZN(n18692) );
  OAI211_X1 U21849 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18677), .A(
        n19455), .B(n18676), .ZN(n18678) );
  NAND2_X1 U21850 ( .A1(n18963), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18981) );
  OAI211_X1 U21851 ( .C1(n18761), .C2(n18679), .A(n18678), .B(n18981), .ZN(
        n18680) );
  AOI21_X1 U21852 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18692), .A(
        n18680), .ZN(n18686) );
  AOI21_X1 U21853 ( .B1(n18682), .B2(n10759), .A(n18681), .ZN(n18973) );
  AOI22_X1 U21854 ( .A1(n18756), .A2(n18973), .B1(n18684), .B2(n18683), .ZN(
        n18685) );
  OAI211_X1 U21855 ( .C1(n18971), .C2(n18687), .A(n18686), .B(n18685), .ZN(
        P3_U2822) );
  OAI21_X1 U21856 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18689), .A(
        n18688), .ZN(n18992) );
  INV_X1 U21857 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19609) );
  NOR2_X1 U21858 ( .A1(n19055), .A2(n19609), .ZN(n18983) );
  AOI221_X1 U21859 ( .B1(n18692), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18691), .C2(n18690), .A(n18983), .ZN(n18698) );
  NAND2_X1 U21860 ( .A1(n18694), .A2(n18693), .ZN(n18695) );
  XOR2_X1 U21861 ( .A(n18695), .B(n18984), .Z(n18989) );
  AOI22_X1 U21862 ( .A1(n18756), .A2(n18989), .B1(n18696), .B2(n18767), .ZN(
        n18697) );
  OAI211_X1 U21863 ( .C1(n18776), .C2(n18992), .A(n18698), .B(n18697), .ZN(
        P3_U2823) );
  NOR2_X1 U21864 ( .A1(n18699), .A2(n18704), .ZN(n18717) );
  OAI22_X1 U21865 ( .A1(n18776), .A2(n19001), .B1(n19055), .B2(n19607), .ZN(
        n18702) );
  AOI221_X1 U21866 ( .B1(n18717), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C1(
        n18704), .C2(n18703), .A(n18702), .ZN(n18708) );
  AOI21_X1 U21867 ( .B1(n18997), .B2(n18706), .A(n18705), .ZN(n18996) );
  NAND2_X1 U21868 ( .A1(n18756), .A2(n18996), .ZN(n18707) );
  OAI211_X1 U21869 ( .C1(n18761), .C2(n18709), .A(n18708), .B(n18707), .ZN(
        P3_U2824) );
  AOI21_X1 U21870 ( .B1(n18712), .B2(n18711), .A(n18710), .ZN(n19007) );
  OAI21_X1 U21871 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18714), .A(
        n18713), .ZN(n19010) );
  OAI22_X1 U21872 ( .A1(n18776), .A2(n19010), .B1(n19055), .B2(n19606), .ZN(
        n18715) );
  AOI21_X1 U21873 ( .B1(n18756), .B2(n19007), .A(n18715), .ZN(n18719) );
  OAI221_X1 U21874 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17697), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18772), .A(n18717), .ZN(n18718) );
  OAI211_X1 U21875 ( .C1(n18761), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2825) );
  OAI21_X1 U21876 ( .B1(n18723), .B2(n18722), .A(n18721), .ZN(n19012) );
  AOI22_X1 U21877 ( .A1(n18963), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n19455), 
        .B2(n18724), .ZN(n18733) );
  AOI21_X1 U21878 ( .B1(n18727), .B2(n18726), .A(n18725), .ZN(n19014) );
  AOI21_X1 U21879 ( .B1(n18741), .B2(n18740), .A(n18728), .ZN(n18744) );
  OAI22_X1 U21880 ( .A1(n18761), .A2(n18730), .B1(n18744), .B2(n18729), .ZN(
        n18731) );
  AOI21_X1 U21881 ( .B1(n18756), .B2(n19014), .A(n18731), .ZN(n18732) );
  OAI211_X1 U21882 ( .C1(n18776), .C2(n19012), .A(n18733), .B(n18732), .ZN(
        P3_U2826) );
  XOR2_X1 U21883 ( .A(n18736), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n19018) );
  AOI21_X1 U21884 ( .B1(n18739), .B2(n18738), .A(n18737), .ZN(n19020) );
  AOI22_X1 U21885 ( .A1(n18756), .A2(n19020), .B1(n19040), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18748) );
  NAND2_X1 U21886 ( .A1(n18741), .A2(n18740), .ZN(n18742) );
  NAND2_X1 U21887 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18772), .ZN(
        n18757) );
  OAI22_X1 U21888 ( .A1(n18744), .A2(n18743), .B1(n18742), .B2(n18757), .ZN(
        n18745) );
  AOI21_X1 U21889 ( .B1(n18746), .B2(n18767), .A(n18745), .ZN(n18747) );
  OAI211_X1 U21890 ( .C1(n18776), .C2(n19018), .A(n18748), .B(n18747), .ZN(
        P3_U2827) );
  AOI21_X1 U21891 ( .B1(n18751), .B2(n18750), .A(n18749), .ZN(n19033) );
  OAI21_X1 U21892 ( .B1(n18754), .B2(n18753), .A(n18752), .ZN(n19043) );
  OAI22_X1 U21893 ( .A1(n18776), .A2(n19043), .B1(n19055), .B2(n19601), .ZN(
        n18755) );
  AOI21_X1 U21894 ( .B1(n18756), .B2(n19033), .A(n18755), .ZN(n18759) );
  OAI21_X1 U21895 ( .B1(n19455), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n18757), .ZN(n18758) );
  OAI211_X1 U21896 ( .C1(n18761), .C2(n18760), .A(n18759), .B(n18758), .ZN(
        P3_U2828) );
  NOR2_X1 U21897 ( .A1(n18762), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18763) );
  XNOR2_X1 U21898 ( .A(n18763), .B(n18765), .ZN(n19052) );
  OAI21_X1 U21899 ( .B1(n18765), .B2(n18771), .A(n18764), .ZN(n19045) );
  OAI22_X1 U21900 ( .A1(n18776), .A2(n19045), .B1(n19055), .B2(n19698), .ZN(
        n18766) );
  AOI221_X1 U21901 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18769), .C1(
        n18768), .C2(n18767), .A(n18766), .ZN(n18770) );
  OAI21_X1 U21902 ( .B1(n19052), .B2(n18777), .A(n18770), .ZN(P3_U2829) );
  AOI21_X1 U21903 ( .B1(n9952), .B2(n19693), .A(n18771), .ZN(n19063) );
  INV_X1 U21904 ( .A(n19063), .ZN(n19061) );
  NAND3_X1 U21905 ( .A1(n19676), .A2(n18773), .A3(n18772), .ZN(n18774) );
  AOI22_X1 U21906 ( .A1(n18963), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18774), .ZN(n18775) );
  OAI221_X1 U21907 ( .B1(n19063), .B2(n18777), .C1(n19061), .C2(n18776), .A(
        n18775), .ZN(P3_U2830) );
  OAI211_X1 U21908 ( .C1(n19548), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18778), .ZN(n18779) );
  OAI221_X1 U21909 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18780), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18829), .A(n18779), .ZN(
        n18784) );
  AOI22_X1 U21910 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n19047), .B1(
        n18962), .B2(n18781), .ZN(n18783) );
  OAI211_X1 U21911 ( .C1(n19054), .C2(n18784), .A(n18783), .B(n18782), .ZN(
        P3_U2835) );
  AOI21_X1 U21912 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n19027), .A(
        n18785), .ZN(n18790) );
  NAND2_X1 U21913 ( .A1(n18806), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18786) );
  OAI21_X1 U21914 ( .B1(n18787), .B2(n18786), .A(n18793), .ZN(n18788) );
  OAI211_X1 U21915 ( .C1(n18790), .C2(n18789), .A(n19039), .B(n18788), .ZN(
        n18791) );
  OAI211_X1 U21916 ( .C1(n19053), .C2(n18793), .A(n18792), .B(n18791), .ZN(
        n18797) );
  OAI22_X1 U21917 ( .A1(n19062), .A2(n18795), .B1(n18969), .B2(n18794), .ZN(
        n18796) );
  AOI211_X1 U21918 ( .C1(n18962), .C2(n18798), .A(n18797), .B(n18796), .ZN(
        n18799) );
  INV_X1 U21919 ( .A(n18799), .ZN(P3_U2837) );
  OAI21_X1 U21920 ( .B1(n19544), .B2(n18805), .A(n18804), .ZN(n18811) );
  NAND4_X1 U21921 ( .A1(n18806), .A2(n19039), .A3(n10592), .A4(n18829), .ZN(
        n18807) );
  NAND2_X1 U21922 ( .A1(n18821), .A2(n18829), .ZN(n18824) );
  NOR2_X1 U21923 ( .A1(n18824), .A2(n19047), .ZN(n18809) );
  AOI21_X1 U21924 ( .B1(n18809), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18810) );
  AOI211_X1 U21925 ( .C1(n18812), .C2(n18811), .A(n19040), .B(n18810), .ZN(
        n18813) );
  AOI21_X1 U21926 ( .B1(n19040), .B2(P3_REIP_REG_23__SCAN_IN), .A(n18813), 
        .ZN(n18814) );
  OAI21_X1 U21927 ( .B1(n18970), .B2(n18815), .A(n18814), .ZN(P3_U2839) );
  OAI221_X1 U21928 ( .B1(n19548), .B2(n18857), .C1(n19548), .C2(n18845), .A(
        n18819), .ZN(n18831) );
  NAND2_X1 U21929 ( .A1(n18820), .A2(n18942), .ZN(n18858) );
  OAI22_X1 U21930 ( .A1(n19548), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18821), .B2(n18945), .ZN(n18840) );
  OAI22_X1 U21931 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18947), .B1(
        n18838), .B2(n19027), .ZN(n18822) );
  OAI21_X1 U21932 ( .B1(n18832), .B2(n18823), .A(n19546), .ZN(n18825) );
  NAND3_X1 U21933 ( .A1(n19039), .A2(n18833), .A3(n18829), .ZN(n18855) );
  AOI22_X1 U21934 ( .A1(n18963), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18962), 
        .B2(n18830), .ZN(n18842) );
  NAND2_X1 U21935 ( .A1(n19027), .A2(n18949), .ZN(n18904) );
  INV_X1 U21936 ( .A(n18904), .ZN(n19044) );
  INV_X1 U21937 ( .A(n18831), .ZN(n18837) );
  INV_X1 U21938 ( .A(n18832), .ZN(n18875) );
  AOI21_X1 U21939 ( .B1(n18875), .B2(n18833), .A(n18949), .ZN(n18834) );
  INV_X1 U21940 ( .A(n18834), .ZN(n18835) );
  AND2_X1 U21941 ( .A1(n18835), .A2(n19039), .ZN(n18836) );
  OAI21_X1 U21942 ( .B1(n18838), .B2(n19044), .A(n18846), .ZN(n18839) );
  OAI211_X1 U21943 ( .C1(n18840), .C2(n18839), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n19055), .ZN(n18841) );
  OAI211_X1 U21944 ( .C1(n18843), .C2(n18855), .A(n18842), .B(n18841), .ZN(
        P3_U2841) );
  AOI22_X1 U21945 ( .A1(n18963), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18962), 
        .B2(n18844), .ZN(n18849) );
  NOR3_X1 U21946 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19044), .A3(
        n19575), .ZN(n18847) );
  OAI21_X1 U21947 ( .B1(n18852), .B2(n18847), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18848) );
  OAI211_X1 U21948 ( .C1(n18850), .C2(n18855), .A(n18849), .B(n18848), .ZN(
        P3_U2842) );
  AOI22_X1 U21949 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18852), .B1(
        n18962), .B2(n18851), .ZN(n18854) );
  OAI211_X1 U21950 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18855), .A(
        n18854), .B(n18853), .ZN(P3_U2843) );
  NOR2_X1 U21951 ( .A1(n19054), .A2(n18856), .ZN(n18879) );
  NAND3_X1 U21952 ( .A1(n18857), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18975), .ZN(n18860) );
  AOI22_X1 U21953 ( .A1(n19030), .A2(n18860), .B1(n18859), .B2(n18858), .ZN(
        n18861) );
  OAI211_X1 U21954 ( .C1(n18862), .C2(n19027), .A(n18879), .B(n18861), .ZN(
        n18870) );
  INV_X1 U21955 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18871) );
  OAI221_X1 U21956 ( .B1(n18870), .B2(n19030), .C1(n18870), .C2(n18871), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18869) );
  NAND2_X1 U21957 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18977) );
  OAI22_X1 U21958 ( .A1(n18974), .A2(n19027), .B1(n18977), .B2(n19031), .ZN(
        n19023) );
  NAND2_X1 U21959 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19023), .ZN(
        n18985) );
  NAND2_X1 U21960 ( .A1(n18864), .A2(n18907), .ZN(n18931) );
  NAND2_X1 U21961 ( .A1(n19039), .A2(n18931), .ZN(n18967) );
  NOR2_X1 U21962 ( .A1(n18865), .A2(n18967), .ZN(n18882) );
  AOI22_X1 U21963 ( .A1(n18962), .A2(n18867), .B1(n18882), .B2(n18866), .ZN(
        n18868) );
  OAI221_X1 U21964 ( .B1(n18963), .B2(n18869), .C1(n19055), .C2(n19629), .A(
        n18868), .ZN(P3_U2844) );
  OAI221_X1 U21965 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n19055), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n19040), .A(n18870), .ZN(
        n18873) );
  NAND3_X1 U21966 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18882), .A3(
        n18871), .ZN(n18872) );
  OAI211_X1 U21967 ( .C1(n18874), .C2(n18970), .A(n18873), .B(n18872), .ZN(
        P3_U2845) );
  AOI21_X1 U21968 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18949), .A(
        n18875), .ZN(n18878) );
  OAI22_X1 U21969 ( .A1(n19548), .A2(n18877), .B1(n18876), .B2(n19027), .ZN(
        n18939) );
  AOI211_X1 U21970 ( .C1(n18889), .C2(n18954), .A(n18878), .B(n18939), .ZN(
        n18888) );
  AOI221_X1 U21971 ( .B1(n18880), .B2(n18879), .C1(n18888), .C2(n18879), .A(
        n18963), .ZN(n18883) );
  AOI22_X1 U21972 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18883), .B1(
        n18882), .B2(n18881), .ZN(n18885) );
  OAI211_X1 U21973 ( .C1(n18886), .C2(n18970), .A(n18885), .B(n18884), .ZN(
        P3_U2846) );
  NOR2_X1 U21974 ( .A1(n9779), .A2(n19062), .ZN(n18897) );
  NOR2_X1 U21975 ( .A1(n18887), .A2(n18942), .ZN(n18892) );
  AOI221_X1 U21976 ( .B1(n18889), .B2(n18900), .C1(n18907), .C2(n18900), .A(
        n18888), .ZN(n18890) );
  AOI21_X1 U21977 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(n18894) );
  OAI22_X1 U21978 ( .A1(n18894), .A2(n19054), .B1(n18970), .B2(n18893), .ZN(
        n18895) );
  AOI21_X1 U21979 ( .B1(n18897), .B2(n18896), .A(n18895), .ZN(n18899) );
  NAND2_X1 U21980 ( .A1(n19040), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18898) );
  OAI211_X1 U21981 ( .C1(n19053), .C2(n18900), .A(n18899), .B(n18898), .ZN(
        P3_U2847) );
  AOI21_X1 U21982 ( .B1(n18937), .B2(n18901), .A(n18949), .ZN(n18902) );
  NOR2_X1 U21983 ( .A1(n18902), .A2(n18939), .ZN(n18923) );
  OAI211_X1 U21984 ( .C1(n18903), .C2(n18947), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18923), .ZN(n18906) );
  OAI221_X1 U21985 ( .B1(n18906), .B2(n18905), .C1(n18906), .C2(n18904), .A(
        n19039), .ZN(n18909) );
  OR2_X1 U21986 ( .A1(n10766), .A2(n18907), .ZN(n18908) );
  AOI222_X1 U21987 ( .A1(n18910), .A2(n18909), .B1(n18910), .B2(n18908), .C1(
        n18909), .C2(n19053), .ZN(n18911) );
  AOI211_X1 U21988 ( .C1(n18913), .C2(n19021), .A(n18912), .B(n18911), .ZN(
        n18916) );
  NAND2_X1 U21989 ( .A1(n18962), .A2(n18914), .ZN(n18915) );
  OAI211_X1 U21990 ( .C1(n18917), .C2(n18969), .A(n18916), .B(n18915), .ZN(
        P3_U2848) );
  AOI22_X1 U21991 ( .A1(n18963), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18962), 
        .B2(n18918), .ZN(n18927) );
  INV_X1 U21992 ( .A(n18919), .ZN(n18921) );
  AOI22_X1 U21993 ( .A1(n19509), .A2(n18921), .B1(n18920), .B2(n18954), .ZN(
        n18922) );
  OAI211_X1 U21994 ( .C1(n18924), .C2(n18942), .A(n18923), .B(n18922), .ZN(
        n18930) );
  OAI21_X1 U21995 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18947), .A(
        n19039), .ZN(n18925) );
  OAI211_X1 U21996 ( .C1(n18930), .C2(n18925), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19055), .ZN(n18926) );
  OAI211_X1 U21997 ( .C1(n18967), .C2(n18928), .A(n18927), .B(n18926), .ZN(
        P3_U2849) );
  OAI222_X1 U21998 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18948), 
        .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18931), .C1(n18930), 
        .C2(n18929), .ZN(n18935) );
  AOI22_X1 U21999 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19047), .B1(
        n18962), .B2(n18932), .ZN(n18934) );
  OAI211_X1 U22000 ( .C1(n19054), .C2(n18935), .A(n18934), .B(n18933), .ZN(
        P3_U2850) );
  AOI22_X1 U22001 ( .A1(n18963), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18962), 
        .B2(n18936), .ZN(n18952) );
  OAI21_X1 U22002 ( .B1(n18949), .B2(n18937), .A(n19039), .ZN(n18938) );
  AOI211_X1 U22003 ( .C1(n19509), .C2(n18940), .A(n18939), .B(n18938), .ZN(
        n18941) );
  OAI21_X1 U22004 ( .B1(n18943), .B2(n18942), .A(n18941), .ZN(n18960) );
  AOI21_X1 U22005 ( .B1(n19546), .B2(n18966), .A(n18960), .ZN(n18944) );
  OAI21_X1 U22006 ( .B1(n18946), .B2(n18945), .A(n18944), .ZN(n18955) );
  OAI22_X1 U22007 ( .A1(n18949), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18948), .B2(n18947), .ZN(n18950) );
  OAI211_X1 U22008 ( .C1(n18955), .C2(n18950), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19055), .ZN(n18951) );
  OAI211_X1 U22009 ( .C1(n18953), .C2(n18967), .A(n18952), .B(n18951), .ZN(
        P3_U2851) );
  OAI221_X1 U22010 ( .B1(n18955), .B2(n18966), .C1(n18955), .C2(n18954), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18959) );
  NOR3_X1 U22011 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18966), .A3(
        n18967), .ZN(n18956) );
  AOI21_X1 U22012 ( .B1(n18962), .B2(n18957), .A(n18956), .ZN(n18958) );
  OAI221_X1 U22013 ( .B1(n19040), .B2(n18959), .C1(n19055), .C2(n19614), .A(
        n18958), .ZN(P3_U2852) );
  NAND2_X1 U22014 ( .A1(n19055), .A2(n18960), .ZN(n18965) );
  AOI22_X1 U22015 ( .A1(n18963), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18962), 
        .B2(n18961), .ZN(n18964) );
  OAI221_X1 U22016 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18967), .C1(
        n18966), .C2(n18965), .A(n18964), .ZN(P3_U2853) );
  OAI22_X1 U22017 ( .A1(n18971), .A2(n18970), .B1(n18969), .B2(n18968), .ZN(
        n18972) );
  AOI21_X1 U22018 ( .B1(n19021), .B2(n18973), .A(n18972), .ZN(n18982) );
  NAND2_X1 U22019 ( .A1(n19544), .A2(n18974), .ZN(n19034) );
  NAND3_X1 U22020 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18975), .A3(
        n19034), .ZN(n18976) );
  AOI21_X1 U22021 ( .B1(n19030), .B2(n18977), .A(n18976), .ZN(n19011) );
  AOI21_X1 U22022 ( .B1(n18978), .B2(n19011), .A(n18993), .ZN(n18988) );
  OAI21_X1 U22023 ( .B1(n19047), .B2(n18988), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18980) );
  NOR2_X1 U22024 ( .A1(n19054), .A2(n18985), .ZN(n19002) );
  NAND3_X1 U22025 ( .A1(n18978), .A2(n19002), .A3(n10759), .ZN(n18979) );
  NAND4_X1 U22026 ( .A1(n18982), .A2(n18981), .A3(n18980), .A4(n18979), .ZN(
        P3_U2854) );
  AOI21_X1 U22027 ( .B1(n19047), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18983), .ZN(n18991) );
  OAI21_X1 U22028 ( .B1(n18986), .B2(n18985), .A(n18984), .ZN(n18987) );
  AOI22_X1 U22029 ( .A1(n19021), .A2(n18989), .B1(n18988), .B2(n18987), .ZN(
        n18990) );
  OAI211_X1 U22030 ( .C1(n19060), .C2(n18992), .A(n18991), .B(n18990), .ZN(
        P3_U2855) );
  AOI21_X1 U22031 ( .B1(n19011), .B2(n18998), .A(n18993), .ZN(n18994) );
  NOR2_X1 U22032 ( .A1(n19047), .A2(n18994), .ZN(n19003) );
  OAI22_X1 U22033 ( .A1(n19003), .A2(n18997), .B1(n19055), .B2(n19607), .ZN(
        n18995) );
  AOI21_X1 U22034 ( .B1(n19021), .B2(n18996), .A(n18995), .ZN(n19000) );
  NAND3_X1 U22035 ( .A1(n18998), .A2(n19002), .A3(n18997), .ZN(n18999) );
  OAI211_X1 U22036 ( .C1(n19001), .C2(n19060), .A(n19000), .B(n18999), .ZN(
        P3_U2856) );
  INV_X1 U22037 ( .A(n19002), .ZN(n19017) );
  NOR2_X1 U22038 ( .A1(n12128), .A2(n19017), .ZN(n19005) );
  INV_X1 U22039 ( .A(n19003), .ZN(n19004) );
  MUX2_X1 U22040 ( .A(n19005), .B(n19004), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n19006) );
  AOI21_X1 U22041 ( .B1(n19021), .B2(n19007), .A(n19006), .ZN(n19009) );
  NAND2_X1 U22042 ( .A1(n19040), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n19008) );
  OAI211_X1 U22043 ( .C1(n19060), .C2(n19010), .A(n19009), .B(n19008), .ZN(
        P3_U2857) );
  INV_X1 U22044 ( .A(n19011), .ZN(n19022) );
  AOI21_X1 U22045 ( .B1(n19048), .B2(n19022), .A(n19047), .ZN(n19016) );
  INV_X1 U22046 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n21656) );
  OAI22_X1 U22047 ( .A1(n19055), .A2(n21656), .B1(n19060), .B2(n19012), .ZN(
        n19013) );
  AOI21_X1 U22048 ( .B1(n19021), .B2(n19014), .A(n19013), .ZN(n19015) );
  OAI221_X1 U22049 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19017), .C1(
        n12128), .C2(n19016), .A(n19015), .ZN(P3_U2858) );
  OAI22_X1 U22050 ( .A1(n19055), .A2(n19603), .B1(n19060), .B2(n19018), .ZN(
        n19019) );
  AOI21_X1 U22051 ( .B1(n19021), .B2(n19020), .A(n19019), .ZN(n19025) );
  OAI211_X1 U22052 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19023), .A(
        n19039), .B(n19022), .ZN(n19024) );
  OAI211_X1 U22053 ( .C1(n19053), .C2(n19026), .A(n19025), .B(n19024), .ZN(
        P3_U2859) );
  NOR3_X1 U22054 ( .A1(n19027), .A2(n19693), .A3(n19674), .ZN(n19029) );
  AOI211_X1 U22055 ( .C1(n19030), .C2(n19674), .A(n19029), .B(n19028), .ZN(
        n19037) );
  NOR3_X1 U22056 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19674), .A3(
        n19031), .ZN(n19032) );
  AOI21_X1 U22057 ( .B1(n19033), .B2(n19509), .A(n19032), .ZN(n19035) );
  OAI211_X1 U22058 ( .C1(n19037), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        n19038) );
  AOI22_X1 U22059 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19047), .B1(
        n19039), .B2(n19038), .ZN(n19042) );
  NAND2_X1 U22060 ( .A1(n19040), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19041) );
  OAI211_X1 U22061 ( .C1(n19060), .C2(n19043), .A(n19042), .B(n19041), .ZN(
        P3_U2860) );
  NOR3_X1 U22062 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19044), .A3(
        n19054), .ZN(n19057) );
  OAI22_X1 U22063 ( .A1(n19055), .A2(n19698), .B1(n19060), .B2(n19045), .ZN(
        n19046) );
  AOI221_X1 U22064 ( .B1(n19047), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n19057), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19046), .ZN(
        n19051) );
  OAI211_X1 U22065 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19049), .A(
        n19048), .B(n19674), .ZN(n19050) );
  OAI211_X1 U22066 ( .C1(n19052), .C2(n19062), .A(n19051), .B(n19050), .ZN(
        P3_U2861) );
  OAI21_X1 U22067 ( .B1(n19548), .B2(n19054), .A(n19053), .ZN(n19058) );
  INV_X1 U22068 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19704) );
  NOR2_X1 U22069 ( .A1(n19055), .A2(n19704), .ZN(n19056) );
  AOI211_X1 U22070 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19058), .A(
        n19057), .B(n19056), .ZN(n19059) );
  OAI221_X1 U22071 ( .B1(n19063), .B2(n19062), .C1(n19061), .C2(n19060), .A(
        n19059), .ZN(P3_U2862) );
  AOI211_X1 U22072 ( .C1(n19065), .C2(n19064), .A(n19575), .B(n19676), .ZN(
        n19568) );
  OAI21_X1 U22073 ( .B1(n19568), .B2(n19110), .A(n19071), .ZN(n19066) );
  OAI221_X1 U22074 ( .B1(n19072), .B2(n19710), .C1(n19072), .C2(n19071), .A(
        n19066), .ZN(P3_U2863) );
  INV_X1 U22075 ( .A(n19340), .ZN(n19339) );
  NAND2_X1 U22076 ( .A1(n19067), .A2(n19339), .ZN(n19363) );
  AND2_X1 U22077 ( .A1(n19219), .A2(n19363), .ZN(n19069) );
  OAI22_X1 U22078 ( .A1(n19070), .A2(n19560), .B1(n19069), .B2(n19068), .ZN(
        P3_U2866) );
  INV_X1 U22079 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21539) );
  NOR2_X1 U22080 ( .A1(n21539), .A2(n19071), .ZN(P3_U2867) );
  INV_X1 U22081 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19079) );
  NAND2_X1 U22082 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19418) );
  NAND2_X1 U22083 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19553), .ZN(
        n19292) );
  NAND2_X1 U22084 ( .A1(n19316), .A2(n19292), .ZN(n19315) );
  INV_X1 U22085 ( .A(n19315), .ZN(n19364) );
  INV_X1 U22086 ( .A(n19246), .ZN(n19552) );
  NOR2_X2 U22087 ( .A1(n19552), .A2(n19418), .ZN(n19502) );
  NOR2_X1 U22088 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19173) );
  NAND2_X1 U22089 ( .A1(n19173), .A2(n19152), .ZN(n19167) );
  NOR2_X1 U22090 ( .A1(n19502), .A2(n19169), .ZN(n19130) );
  OAI33_X1 U22091 ( .A1(n19418), .A2(n19364), .A3(n19221), .B1(n19220), .B2(
        n19130), .B3(n19073), .ZN(n19108) );
  NOR2_X1 U22092 ( .A1(n19418), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19454) );
  NAND2_X1 U22093 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19454), .ZN(
        n19497) );
  INV_X1 U22094 ( .A(n19497), .ZN(n19501) );
  NAND2_X1 U22095 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19455), .ZN(n19459) );
  INV_X1 U22096 ( .A(n19459), .ZN(n19419) );
  NOR2_X2 U22097 ( .A1(n19220), .A2(n14119), .ZN(n19450) );
  INV_X1 U22098 ( .A(n19449), .ZN(n19576) );
  NOR2_X1 U22099 ( .A1(n19576), .A2(n19130), .ZN(n19103) );
  AOI22_X1 U22100 ( .A1(n19501), .A2(n19419), .B1(n19450), .B2(n19103), .ZN(
        n19078) );
  NOR2_X2 U22101 ( .A1(n19418), .A2(n19316), .ZN(n19444) );
  NAND2_X1 U22102 ( .A1(n19455), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19392) );
  INV_X1 U22103 ( .A(n19392), .ZN(n19451) );
  NAND2_X1 U22104 ( .A1(n19075), .A2(n19074), .ZN(n19104) );
  NOR2_X2 U22105 ( .A1(n19076), .A2(n19104), .ZN(n19456) );
  AOI22_X1 U22106 ( .A1(n19444), .A2(n19451), .B1(n19456), .B2(n19169), .ZN(
        n19077) );
  OAI211_X1 U22107 ( .C1(n19079), .C2(n19108), .A(n19078), .B(n19077), .ZN(
        P3_U2868) );
  INV_X1 U22108 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19082) );
  NAND2_X1 U22109 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19455), .ZN(n19465) );
  INV_X1 U22110 ( .A(n19465), .ZN(n19422) );
  NOR2_X2 U22111 ( .A1(n19220), .A2(n14088), .ZN(n19460) );
  AOI22_X1 U22112 ( .A1(n19501), .A2(n19422), .B1(n19460), .B2(n19103), .ZN(
        n19081) );
  AND2_X1 U22113 ( .A1(n19455), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19461) );
  NOR2_X1 U22114 ( .A1(n19715), .A2(n19104), .ZN(n19462) );
  AOI22_X1 U22115 ( .A1(n19444), .A2(n19461), .B1(n19462), .B2(n19169), .ZN(
        n19080) );
  OAI211_X1 U22116 ( .C1(n19082), .C2(n19108), .A(n19081), .B(n19080), .ZN(
        P3_U2869) );
  NAND2_X1 U22117 ( .A1(n19455), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19471) );
  INV_X1 U22118 ( .A(n19471), .ZN(n19426) );
  NOR2_X2 U22119 ( .A1(n19220), .A2(n14082), .ZN(n19466) );
  AOI22_X1 U22120 ( .A1(n19444), .A2(n19426), .B1(n19466), .B2(n19103), .ZN(
        n19085) );
  NAND2_X1 U22121 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19455), .ZN(n19429) );
  INV_X1 U22122 ( .A(n19429), .ZN(n19467) );
  NOR2_X2 U22123 ( .A1(n19083), .A2(n19104), .ZN(n19468) );
  AOI22_X1 U22124 ( .A1(n19501), .A2(n19467), .B1(n19468), .B2(n19169), .ZN(
        n19084) );
  OAI211_X1 U22125 ( .C1(n19086), .C2(n19108), .A(n19085), .B(n19084), .ZN(
        P3_U2870) );
  NAND2_X1 U22126 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19455), .ZN(n19477) );
  NOR2_X2 U22127 ( .A1(n14097), .A2(n19220), .ZN(n19472) );
  AOI22_X1 U22128 ( .A1(n19501), .A2(n19430), .B1(n19472), .B2(n19103), .ZN(
        n19089) );
  NOR2_X1 U22129 ( .A1(n16451), .A2(n19221), .ZN(n19473) );
  NOR2_X2 U22130 ( .A1(n19087), .A2(n19104), .ZN(n19474) );
  AOI22_X1 U22131 ( .A1(n19444), .A2(n19473), .B1(n19474), .B2(n19169), .ZN(
        n19088) );
  OAI211_X1 U22132 ( .C1(n19090), .C2(n19108), .A(n19089), .B(n19088), .ZN(
        P3_U2871) );
  NOR2_X2 U22133 ( .A1(n16440), .A2(n19221), .ZN(n19479) );
  NOR2_X2 U22134 ( .A1(n14104), .A2(n19220), .ZN(n19478) );
  AOI22_X1 U22135 ( .A1(n19444), .A2(n19479), .B1(n19478), .B2(n19103), .ZN(
        n19093) );
  NAND2_X1 U22136 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19455), .ZN(n19483) );
  INV_X1 U22137 ( .A(n19483), .ZN(n19434) );
  NOR2_X2 U22138 ( .A1(n19091), .A2(n19104), .ZN(n19480) );
  AOI22_X1 U22139 ( .A1(n19501), .A2(n19434), .B1(n19480), .B2(n19169), .ZN(
        n19092) );
  OAI211_X1 U22140 ( .C1(n19094), .C2(n9915), .A(n19093), .B(n19092), .ZN(
        P3_U2872) );
  NAND2_X1 U22141 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19455), .ZN(n19306) );
  INV_X1 U22142 ( .A(n19306), .ZN(n19485) );
  NOR2_X2 U22143 ( .A1(n14101), .A2(n19220), .ZN(n19484) );
  AOI22_X1 U22144 ( .A1(n19501), .A2(n19485), .B1(n19484), .B2(n19103), .ZN(
        n19097) );
  NOR2_X1 U22145 ( .A1(n16432), .A2(n19221), .ZN(n19303) );
  NOR2_X2 U22146 ( .A1(n19095), .A2(n19104), .ZN(n19486) );
  AOI22_X1 U22147 ( .A1(n19444), .A2(n19303), .B1(n19486), .B2(n19169), .ZN(
        n19096) );
  OAI211_X1 U22148 ( .C1(n19098), .C2(n9915), .A(n19097), .B(n19096), .ZN(
        P3_U2873) );
  NOR2_X1 U22149 ( .A1(n21624), .A2(n19221), .ZN(n19404) );
  NOR2_X2 U22150 ( .A1(n14069), .A2(n19220), .ZN(n19490) );
  AOI22_X1 U22151 ( .A1(n19444), .A2(n19404), .B1(n19490), .B2(n19103), .ZN(
        n19101) );
  NAND2_X1 U22152 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19455), .ZN(n19407) );
  INV_X1 U22153 ( .A(n19407), .ZN(n19491) );
  NOR2_X2 U22154 ( .A1(n19099), .A2(n19104), .ZN(n19493) );
  AOI22_X1 U22155 ( .A1(n19501), .A2(n19491), .B1(n19493), .B2(n19169), .ZN(
        n19100) );
  OAI211_X1 U22156 ( .C1(n19102), .C2(n9915), .A(n19101), .B(n19100), .ZN(
        P3_U2874) );
  NOR2_X1 U22157 ( .A1(n21561), .A2(n19221), .ZN(n19384) );
  NOR2_X2 U22158 ( .A1(n14107), .A2(n19220), .ZN(n19499) );
  AOI22_X1 U22159 ( .A1(n19501), .A2(n19384), .B1(n19499), .B2(n19103), .ZN(
        n19107) );
  NAND2_X1 U22160 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19455), .ZN(n19387) );
  INV_X1 U22161 ( .A(n19387), .ZN(n19500) );
  NOR2_X2 U22162 ( .A1(n19105), .A2(n19104), .ZN(n19503) );
  AOI22_X1 U22163 ( .A1(n19444), .A2(n19500), .B1(n19503), .B2(n19169), .ZN(
        n19106) );
  OAI211_X1 U22164 ( .C1(n19109), .C2(n9915), .A(n19107), .B(n19106), .ZN(
        P3_U2875) );
  INV_X1 U22165 ( .A(n19444), .ZN(n19129) );
  INV_X1 U22166 ( .A(n19152), .ZN(n19196) );
  AOI22_X1 U22167 ( .A1(n19451), .A2(n19502), .B1(n19450), .B2(n19125), .ZN(
        n19112) );
  NOR2_X1 U22168 ( .A1(n19560), .A2(n19289), .ZN(n19452) );
  NOR2_X1 U22169 ( .A1(n19220), .A2(n19110), .ZN(n19453) );
  INV_X1 U22170 ( .A(n19453), .ZN(n19151) );
  NOR2_X1 U22171 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19151), .ZN(
        n19197) );
  AOI22_X1 U22172 ( .A1(n19455), .A2(n19452), .B1(n19152), .B2(n19197), .ZN(
        n19126) );
  NOR2_X2 U22173 ( .A1(n19292), .A2(n19196), .ZN(n19192) );
  AOI22_X1 U22174 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19126), .B1(
        n19456), .B2(n19192), .ZN(n19111) );
  OAI211_X1 U22175 ( .C1(n19129), .C2(n19459), .A(n19112), .B(n19111), .ZN(
        P3_U2876) );
  AOI22_X1 U22176 ( .A1(n19461), .A2(n19502), .B1(n19460), .B2(n19125), .ZN(
        n19114) );
  AOI22_X1 U22177 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19126), .B1(
        n19462), .B2(n19192), .ZN(n19113) );
  OAI211_X1 U22178 ( .C1(n19129), .C2(n19465), .A(n19114), .B(n19113), .ZN(
        P3_U2877) );
  INV_X1 U22179 ( .A(n19502), .ZN(n19146) );
  AOI22_X1 U22180 ( .A1(n19444), .A2(n19467), .B1(n19466), .B2(n19125), .ZN(
        n19116) );
  AOI22_X1 U22181 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19126), .B1(
        n19468), .B2(n19192), .ZN(n19115) );
  OAI211_X1 U22182 ( .C1(n19471), .C2(n19146), .A(n19116), .B(n19115), .ZN(
        P3_U2878) );
  AOI22_X1 U22183 ( .A1(n19473), .A2(n19502), .B1(n19472), .B2(n19125), .ZN(
        n19118) );
  AOI22_X1 U22184 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19126), .B1(
        n19474), .B2(n19192), .ZN(n19117) );
  OAI211_X1 U22185 ( .C1(n19129), .C2(n19477), .A(n19118), .B(n19117), .ZN(
        P3_U2879) );
  AOI22_X1 U22186 ( .A1(n19479), .A2(n19502), .B1(n19478), .B2(n19125), .ZN(
        n19120) );
  AOI22_X1 U22187 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19126), .B1(
        n19480), .B2(n19192), .ZN(n19119) );
  OAI211_X1 U22188 ( .C1(n19129), .C2(n19483), .A(n19120), .B(n19119), .ZN(
        P3_U2880) );
  AOI22_X1 U22189 ( .A1(n19444), .A2(n19485), .B1(n19484), .B2(n19125), .ZN(
        n19122) );
  AOI22_X1 U22190 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19126), .B1(
        n19486), .B2(n19192), .ZN(n19121) );
  OAI211_X1 U22191 ( .C1(n19489), .C2(n19146), .A(n19122), .B(n19121), .ZN(
        P3_U2881) );
  AOI22_X1 U22192 ( .A1(n19404), .A2(n19502), .B1(n19490), .B2(n19125), .ZN(
        n19124) );
  AOI22_X1 U22193 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19126), .B1(
        n19493), .B2(n19192), .ZN(n19123) );
  OAI211_X1 U22194 ( .C1(n19129), .C2(n19407), .A(n19124), .B(n19123), .ZN(
        P3_U2882) );
  INV_X1 U22195 ( .A(n19384), .ZN(n19507) );
  AOI22_X1 U22196 ( .A1(n19499), .A2(n19125), .B1(n19500), .B2(n19502), .ZN(
        n19128) );
  AOI22_X1 U22197 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19126), .B1(
        n19503), .B2(n19192), .ZN(n19127) );
  OAI211_X1 U22198 ( .C1(n19129), .C2(n19507), .A(n19128), .B(n19127), .ZN(
        P3_U2883) );
  NOR2_X2 U22199 ( .A1(n19316), .A2(n19196), .ZN(n19215) );
  INV_X1 U22200 ( .A(n19220), .ZN(n19415) );
  NOR2_X1 U22201 ( .A1(n19192), .A2(n19215), .ZN(n19174) );
  OAI21_X1 U22202 ( .B1(n19130), .B2(n19414), .A(n19174), .ZN(n19131) );
  OAI211_X1 U22203 ( .C1(n19215), .C2(n19666), .A(n19415), .B(n19131), .ZN(
        n19148) );
  NOR2_X1 U22204 ( .A1(n19576), .A2(n19174), .ZN(n19147) );
  AOI22_X1 U22205 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19148), .B1(
        n19450), .B2(n19147), .ZN(n19133) );
  AOI22_X1 U22206 ( .A1(n19451), .A2(n19169), .B1(n19456), .B2(n19215), .ZN(
        n19132) );
  OAI211_X1 U22207 ( .C1(n19459), .C2(n19146), .A(n19133), .B(n19132), .ZN(
        P3_U2884) );
  INV_X1 U22208 ( .A(n19462), .ZN(n19345) );
  AOI22_X1 U22209 ( .A1(n19460), .A2(n19147), .B1(n19422), .B2(n19502), .ZN(
        n19135) );
  AOI22_X1 U22210 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19148), .B1(
        n19461), .B2(n19169), .ZN(n19134) );
  OAI211_X1 U22211 ( .C1(n19345), .C2(n19211), .A(n19135), .B(n19134), .ZN(
        P3_U2885) );
  AOI22_X1 U22212 ( .A1(n19467), .A2(n19502), .B1(n19466), .B2(n19147), .ZN(
        n19137) );
  AOI22_X1 U22213 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19148), .B1(
        n19468), .B2(n19215), .ZN(n19136) );
  OAI211_X1 U22214 ( .C1(n19471), .C2(n19167), .A(n19137), .B(n19136), .ZN(
        P3_U2886) );
  AOI22_X1 U22215 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19148), .B1(
        n19472), .B2(n19147), .ZN(n19139) );
  AOI22_X1 U22216 ( .A1(n19474), .A2(n19215), .B1(n19430), .B2(n19502), .ZN(
        n19138) );
  OAI211_X1 U22217 ( .C1(n19433), .C2(n19167), .A(n19139), .B(n19138), .ZN(
        P3_U2887) );
  AOI22_X1 U22218 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19148), .B1(
        n19478), .B2(n19147), .ZN(n19141) );
  AOI22_X1 U22219 ( .A1(n19479), .A2(n19169), .B1(n19480), .B2(n19215), .ZN(
        n19140) );
  OAI211_X1 U22220 ( .C1(n19483), .C2(n19146), .A(n19141), .B(n19140), .ZN(
        P3_U2888) );
  AOI22_X1 U22221 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19148), .B1(
        n19484), .B2(n19147), .ZN(n19143) );
  AOI22_X1 U22222 ( .A1(n19486), .A2(n19215), .B1(n19485), .B2(n19502), .ZN(
        n19142) );
  OAI211_X1 U22223 ( .C1(n19489), .C2(n19167), .A(n19143), .B(n19142), .ZN(
        P3_U2889) );
  AOI22_X1 U22224 ( .A1(n19404), .A2(n19169), .B1(n19490), .B2(n19147), .ZN(
        n19145) );
  AOI22_X1 U22225 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19148), .B1(
        n19493), .B2(n19215), .ZN(n19144) );
  OAI211_X1 U22226 ( .C1(n19407), .C2(n19146), .A(n19145), .B(n19144), .ZN(
        P3_U2890) );
  AOI22_X1 U22227 ( .A1(n19384), .A2(n19502), .B1(n19499), .B2(n19147), .ZN(
        n19150) );
  AOI22_X1 U22228 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19148), .B1(
        n19503), .B2(n19215), .ZN(n19149) );
  OAI211_X1 U22229 ( .C1(n19387), .C2(n19167), .A(n19150), .B(n19149), .ZN(
        P3_U2891) );
  AOI22_X1 U22230 ( .A1(n19451), .A2(n19192), .B1(n19450), .B2(n19168), .ZN(
        n19154) );
  AOI21_X1 U22231 ( .B1(n19553), .B2(n19414), .A(n19151), .ZN(n19244) );
  NAND2_X1 U22232 ( .A1(n19152), .A2(n19244), .ZN(n19170) );
  NAND2_X1 U22233 ( .A1(n19246), .A2(n19152), .ZN(n19243) );
  INV_X1 U22234 ( .A(n19243), .ZN(n19228) );
  AOI22_X1 U22235 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19170), .B1(
        n19456), .B2(n19228), .ZN(n19153) );
  OAI211_X1 U22236 ( .C1(n19459), .C2(n19167), .A(n19154), .B(n19153), .ZN(
        P3_U2892) );
  AOI22_X1 U22237 ( .A1(n19460), .A2(n19168), .B1(n19422), .B2(n19169), .ZN(
        n19156) );
  AOI22_X1 U22238 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19170), .B1(
        n19461), .B2(n19192), .ZN(n19155) );
  OAI211_X1 U22239 ( .C1(n19345), .C2(n19243), .A(n19156), .B(n19155), .ZN(
        P3_U2893) );
  AOI22_X1 U22240 ( .A1(n19466), .A2(n19168), .B1(n19426), .B2(n19192), .ZN(
        n19158) );
  AOI22_X1 U22241 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19170), .B1(
        n19468), .B2(n19228), .ZN(n19157) );
  OAI211_X1 U22242 ( .C1(n19429), .C2(n19167), .A(n19158), .B(n19157), .ZN(
        P3_U2894) );
  INV_X1 U22243 ( .A(n19192), .ZN(n19190) );
  AOI22_X1 U22244 ( .A1(n19472), .A2(n19168), .B1(n19430), .B2(n19169), .ZN(
        n19160) );
  AOI22_X1 U22245 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19170), .B1(
        n19474), .B2(n19228), .ZN(n19159) );
  OAI211_X1 U22246 ( .C1(n19433), .C2(n19190), .A(n19160), .B(n19159), .ZN(
        P3_U2895) );
  INV_X1 U22247 ( .A(n19479), .ZN(n19437) );
  AOI22_X1 U22248 ( .A1(n19434), .A2(n19169), .B1(n19478), .B2(n19168), .ZN(
        n19162) );
  AOI22_X1 U22249 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19170), .B1(
        n19480), .B2(n19228), .ZN(n19161) );
  OAI211_X1 U22250 ( .C1(n19437), .C2(n19190), .A(n19162), .B(n19161), .ZN(
        P3_U2896) );
  AOI22_X1 U22251 ( .A1(n19484), .A2(n19168), .B1(n19485), .B2(n19169), .ZN(
        n19164) );
  AOI22_X1 U22252 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19170), .B1(
        n19486), .B2(n19228), .ZN(n19163) );
  OAI211_X1 U22253 ( .C1(n19489), .C2(n19190), .A(n19164), .B(n19163), .ZN(
        P3_U2897) );
  AOI22_X1 U22254 ( .A1(n19404), .A2(n19192), .B1(n19490), .B2(n19168), .ZN(
        n19166) );
  AOI22_X1 U22255 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19170), .B1(
        n19493), .B2(n19228), .ZN(n19165) );
  OAI211_X1 U22256 ( .C1(n19407), .C2(n19167), .A(n19166), .B(n19165), .ZN(
        P3_U2898) );
  AOI22_X1 U22257 ( .A1(n19384), .A2(n19169), .B1(n19499), .B2(n19168), .ZN(
        n19172) );
  AOI22_X1 U22258 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19170), .B1(
        n19503), .B2(n19228), .ZN(n19171) );
  OAI211_X1 U22259 ( .C1(n19387), .C2(n19190), .A(n19172), .B(n19171), .ZN(
        P3_U2899) );
  INV_X1 U22260 ( .A(n19173), .ZN(n19554) );
  NOR2_X2 U22261 ( .A1(n19554), .A2(n19219), .ZN(n19263) );
  AOI21_X1 U22262 ( .B1(n19243), .B2(n19261), .A(n19576), .ZN(n19191) );
  AOI22_X1 U22263 ( .A1(n19419), .A2(n19192), .B1(n19450), .B2(n19191), .ZN(
        n19177) );
  AOI221_X1 U22264 ( .B1(n19174), .B2(n19243), .C1(n19414), .C2(n19243), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19175) );
  OAI21_X1 U22265 ( .B1(n19263), .B2(n19175), .A(n19415), .ZN(n19193) );
  AOI22_X1 U22266 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19193), .B1(
        n19456), .B2(n19263), .ZN(n19176) );
  OAI211_X1 U22267 ( .C1(n19392), .C2(n19211), .A(n19177), .B(n19176), .ZN(
        P3_U2900) );
  AOI22_X1 U22268 ( .A1(n19460), .A2(n19191), .B1(n19422), .B2(n19192), .ZN(
        n19179) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19193), .B1(
        n19461), .B2(n19215), .ZN(n19178) );
  OAI211_X1 U22270 ( .C1(n19345), .C2(n19261), .A(n19179), .B(n19178), .ZN(
        P3_U2901) );
  AOI22_X1 U22271 ( .A1(n19467), .A2(n19192), .B1(n19466), .B2(n19191), .ZN(
        n19181) );
  AOI22_X1 U22272 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19193), .B1(
        n19468), .B2(n19263), .ZN(n19180) );
  OAI211_X1 U22273 ( .C1(n19471), .C2(n19211), .A(n19181), .B(n19180), .ZN(
        P3_U2902) );
  AOI22_X1 U22274 ( .A1(n19472), .A2(n19191), .B1(n19430), .B2(n19192), .ZN(
        n19183) );
  AOI22_X1 U22275 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19193), .B1(
        n19474), .B2(n19263), .ZN(n19182) );
  OAI211_X1 U22276 ( .C1(n19433), .C2(n19211), .A(n19183), .B(n19182), .ZN(
        P3_U2903) );
  AOI22_X1 U22277 ( .A1(n19479), .A2(n19215), .B1(n19478), .B2(n19191), .ZN(
        n19185) );
  AOI22_X1 U22278 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19193), .B1(
        n19480), .B2(n19263), .ZN(n19184) );
  OAI211_X1 U22279 ( .C1(n19483), .C2(n19190), .A(n19185), .B(n19184), .ZN(
        P3_U2904) );
  AOI22_X1 U22280 ( .A1(n19303), .A2(n19215), .B1(n19484), .B2(n19191), .ZN(
        n19187) );
  AOI22_X1 U22281 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19193), .B1(
        n19486), .B2(n19263), .ZN(n19186) );
  OAI211_X1 U22282 ( .C1(n19306), .C2(n19190), .A(n19187), .B(n19186), .ZN(
        P3_U2905) );
  AOI22_X1 U22283 ( .A1(n19404), .A2(n19215), .B1(n19490), .B2(n19191), .ZN(
        n19189) );
  AOI22_X1 U22284 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19193), .B1(
        n19493), .B2(n19263), .ZN(n19188) );
  OAI211_X1 U22285 ( .C1(n19407), .C2(n19190), .A(n19189), .B(n19188), .ZN(
        P3_U2906) );
  AOI22_X1 U22286 ( .A1(n19384), .A2(n19192), .B1(n19499), .B2(n19191), .ZN(
        n19195) );
  AOI22_X1 U22287 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19193), .B1(
        n19503), .B2(n19263), .ZN(n19194) );
  OAI211_X1 U22288 ( .C1(n19387), .C2(n19211), .A(n19195), .B(n19194), .ZN(
        P3_U2907) );
  AOI22_X1 U22289 ( .A1(n19419), .A2(n19215), .B1(n19450), .B2(n19214), .ZN(
        n19200) );
  NOR2_X1 U22290 ( .A1(n19553), .A2(n19196), .ZN(n19198) );
  INV_X1 U22291 ( .A(n19219), .ZN(n19245) );
  AOI22_X1 U22292 ( .A1(n19455), .A2(n19198), .B1(n19197), .B2(n19245), .ZN(
        n19216) );
  NOR2_X2 U22293 ( .A1(n19292), .A2(n19219), .ZN(n19281) );
  AOI22_X1 U22294 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19216), .B1(
        n19456), .B2(n19281), .ZN(n19199) );
  OAI211_X1 U22295 ( .C1(n19392), .C2(n19243), .A(n19200), .B(n19199), .ZN(
        P3_U2908) );
  AOI22_X1 U22296 ( .A1(n19461), .A2(n19228), .B1(n19460), .B2(n19214), .ZN(
        n19202) );
  AOI22_X1 U22297 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19216), .B1(
        n19462), .B2(n19281), .ZN(n19201) );
  OAI211_X1 U22298 ( .C1(n19465), .C2(n19211), .A(n19202), .B(n19201), .ZN(
        P3_U2909) );
  AOI22_X1 U22299 ( .A1(n19467), .A2(n19215), .B1(n19466), .B2(n19214), .ZN(
        n19204) );
  AOI22_X1 U22300 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19216), .B1(
        n19468), .B2(n19281), .ZN(n19203) );
  OAI211_X1 U22301 ( .C1(n19471), .C2(n19243), .A(n19204), .B(n19203), .ZN(
        P3_U2910) );
  AOI22_X1 U22302 ( .A1(n19473), .A2(n19228), .B1(n19472), .B2(n19214), .ZN(
        n19206) );
  AOI22_X1 U22303 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19216), .B1(
        n19474), .B2(n19281), .ZN(n19205) );
  OAI211_X1 U22304 ( .C1(n19477), .C2(n19211), .A(n19206), .B(n19205), .ZN(
        P3_U2911) );
  AOI22_X1 U22305 ( .A1(n19479), .A2(n19228), .B1(n19478), .B2(n19214), .ZN(
        n19208) );
  AOI22_X1 U22306 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19216), .B1(
        n19480), .B2(n19281), .ZN(n19207) );
  OAI211_X1 U22307 ( .C1(n19483), .C2(n19211), .A(n19208), .B(n19207), .ZN(
        P3_U2912) );
  AOI22_X1 U22308 ( .A1(n19303), .A2(n19228), .B1(n19484), .B2(n19214), .ZN(
        n19210) );
  AOI22_X1 U22309 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19216), .B1(
        n19486), .B2(n19281), .ZN(n19209) );
  OAI211_X1 U22310 ( .C1(n19306), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P3_U2913) );
  INV_X1 U22311 ( .A(n19404), .ZN(n19496) );
  AOI22_X1 U22312 ( .A1(n19491), .A2(n19215), .B1(n19490), .B2(n19214), .ZN(
        n19213) );
  AOI22_X1 U22313 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19216), .B1(
        n19493), .B2(n19281), .ZN(n19212) );
  OAI211_X1 U22314 ( .C1(n19496), .C2(n19243), .A(n19213), .B(n19212), .ZN(
        P3_U2914) );
  AOI22_X1 U22315 ( .A1(n19384), .A2(n19215), .B1(n19499), .B2(n19214), .ZN(
        n19218) );
  AOI22_X1 U22316 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19216), .B1(
        n19503), .B2(n19281), .ZN(n19217) );
  OAI211_X1 U22317 ( .C1(n19387), .C2(n19243), .A(n19218), .B(n19217), .ZN(
        P3_U2915) );
  NOR2_X2 U22318 ( .A1(n19316), .A2(n19219), .ZN(n19311) );
  NOR2_X1 U22319 ( .A1(n19281), .A2(n19311), .ZN(n19267) );
  NOR2_X1 U22320 ( .A1(n19576), .A2(n19267), .ZN(n19239) );
  AOI22_X1 U22321 ( .A1(n19419), .A2(n19228), .B1(n19450), .B2(n19239), .ZN(
        n19225) );
  NOR2_X1 U22322 ( .A1(n19228), .A2(n19263), .ZN(n19222) );
  OAI22_X1 U22323 ( .A1(n19222), .A2(n19221), .B1(n19267), .B2(n19220), .ZN(
        n19223) );
  OAI21_X1 U22324 ( .B1(n19311), .B2(n19666), .A(n19223), .ZN(n19240) );
  AOI22_X1 U22325 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19240), .B1(
        n19456), .B2(n19311), .ZN(n19224) );
  OAI211_X1 U22326 ( .C1(n19392), .C2(n19261), .A(n19225), .B(n19224), .ZN(
        P3_U2916) );
  AOI22_X1 U22327 ( .A1(n19461), .A2(n19263), .B1(n19460), .B2(n19239), .ZN(
        n19227) );
  AOI22_X1 U22328 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19240), .B1(
        n19462), .B2(n19311), .ZN(n19226) );
  OAI211_X1 U22329 ( .C1(n19465), .C2(n19243), .A(n19227), .B(n19226), .ZN(
        P3_U2917) );
  AOI22_X1 U22330 ( .A1(n19467), .A2(n19228), .B1(n19466), .B2(n19239), .ZN(
        n19230) );
  AOI22_X1 U22331 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19240), .B1(
        n19468), .B2(n19311), .ZN(n19229) );
  OAI211_X1 U22332 ( .C1(n19471), .C2(n19261), .A(n19230), .B(n19229), .ZN(
        P3_U2918) );
  AOI22_X1 U22333 ( .A1(n19473), .A2(n19263), .B1(n19472), .B2(n19239), .ZN(
        n19232) );
  AOI22_X1 U22334 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19240), .B1(
        n19474), .B2(n19311), .ZN(n19231) );
  OAI211_X1 U22335 ( .C1(n19477), .C2(n19243), .A(n19232), .B(n19231), .ZN(
        P3_U2919) );
  AOI22_X1 U22336 ( .A1(n19479), .A2(n19263), .B1(n19478), .B2(n19239), .ZN(
        n19234) );
  AOI22_X1 U22337 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19240), .B1(
        n19480), .B2(n19311), .ZN(n19233) );
  OAI211_X1 U22338 ( .C1(n19483), .C2(n19243), .A(n19234), .B(n19233), .ZN(
        P3_U2920) );
  AOI22_X1 U22339 ( .A1(n19303), .A2(n19263), .B1(n19484), .B2(n19239), .ZN(
        n19236) );
  AOI22_X1 U22340 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19240), .B1(
        n19486), .B2(n19311), .ZN(n19235) );
  OAI211_X1 U22341 ( .C1(n19306), .C2(n19243), .A(n19236), .B(n19235), .ZN(
        P3_U2921) );
  AOI22_X1 U22342 ( .A1(n19404), .A2(n19263), .B1(n19490), .B2(n19239), .ZN(
        n19238) );
  AOI22_X1 U22343 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19240), .B1(
        n19493), .B2(n19311), .ZN(n19237) );
  OAI211_X1 U22344 ( .C1(n19407), .C2(n19243), .A(n19238), .B(n19237), .ZN(
        P3_U2922) );
  AOI22_X1 U22345 ( .A1(n19499), .A2(n19239), .B1(n19500), .B2(n19263), .ZN(
        n19242) );
  AOI22_X1 U22346 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19240), .B1(
        n19503), .B2(n19311), .ZN(n19241) );
  OAI211_X1 U22347 ( .C1(n19507), .C2(n19243), .A(n19242), .B(n19241), .ZN(
        P3_U2923) );
  INV_X1 U22348 ( .A(n19281), .ZN(n19288) );
  AOI22_X1 U22349 ( .A1(n19419), .A2(n19263), .B1(n19450), .B2(n19262), .ZN(
        n19248) );
  NAND2_X1 U22350 ( .A1(n19244), .A2(n19245), .ZN(n19264) );
  NAND2_X1 U22351 ( .A1(n19246), .A2(n19245), .ZN(n19329) );
  INV_X1 U22352 ( .A(n19329), .ZN(n19335) );
  AOI22_X1 U22353 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19264), .B1(
        n19456), .B2(n19335), .ZN(n19247) );
  OAI211_X1 U22354 ( .C1(n19392), .C2(n19288), .A(n19248), .B(n19247), .ZN(
        P3_U2924) );
  AOI22_X1 U22355 ( .A1(n19461), .A2(n19281), .B1(n19460), .B2(n19262), .ZN(
        n19250) );
  AOI22_X1 U22356 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19264), .B1(
        n19462), .B2(n19335), .ZN(n19249) );
  OAI211_X1 U22357 ( .C1(n19465), .C2(n19261), .A(n19250), .B(n19249), .ZN(
        P3_U2925) );
  AOI22_X1 U22358 ( .A1(n19466), .A2(n19262), .B1(n19426), .B2(n19281), .ZN(
        n19252) );
  AOI22_X1 U22359 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19264), .B1(
        n19468), .B2(n19335), .ZN(n19251) );
  OAI211_X1 U22360 ( .C1(n19429), .C2(n19261), .A(n19252), .B(n19251), .ZN(
        P3_U2926) );
  AOI22_X1 U22361 ( .A1(n19473), .A2(n19281), .B1(n19472), .B2(n19262), .ZN(
        n19254) );
  AOI22_X1 U22362 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19264), .B1(
        n19474), .B2(n19335), .ZN(n19253) );
  OAI211_X1 U22363 ( .C1(n19477), .C2(n19261), .A(n19254), .B(n19253), .ZN(
        P3_U2927) );
  AOI22_X1 U22364 ( .A1(n19479), .A2(n19281), .B1(n19478), .B2(n19262), .ZN(
        n19256) );
  AOI22_X1 U22365 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19264), .B1(
        n19480), .B2(n19335), .ZN(n19255) );
  OAI211_X1 U22366 ( .C1(n19483), .C2(n19261), .A(n19256), .B(n19255), .ZN(
        P3_U2928) );
  AOI22_X1 U22367 ( .A1(n19484), .A2(n19262), .B1(n19485), .B2(n19263), .ZN(
        n19258) );
  AOI22_X1 U22368 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19264), .B1(
        n19486), .B2(n19335), .ZN(n19257) );
  OAI211_X1 U22369 ( .C1(n19489), .C2(n19288), .A(n19258), .B(n19257), .ZN(
        P3_U2929) );
  AOI22_X1 U22370 ( .A1(n19404), .A2(n19281), .B1(n19490), .B2(n19262), .ZN(
        n19260) );
  AOI22_X1 U22371 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19264), .B1(
        n19493), .B2(n19335), .ZN(n19259) );
  OAI211_X1 U22372 ( .C1(n19407), .C2(n19261), .A(n19260), .B(n19259), .ZN(
        P3_U2930) );
  AOI22_X1 U22373 ( .A1(n19384), .A2(n19263), .B1(n19499), .B2(n19262), .ZN(
        n19266) );
  AOI22_X1 U22374 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19264), .B1(
        n19503), .B2(n19335), .ZN(n19265) );
  OAI211_X1 U22375 ( .C1(n19387), .C2(n19288), .A(n19266), .B(n19265), .ZN(
        P3_U2931) );
  NOR2_X1 U22376 ( .A1(n19554), .A2(n19340), .ZN(n19350) );
  INV_X1 U22377 ( .A(n19350), .ZN(n19362) );
  AOI21_X1 U22378 ( .B1(n19329), .B2(n19362), .A(n19576), .ZN(n19284) );
  AOI22_X1 U22379 ( .A1(n19419), .A2(n19281), .B1(n19450), .B2(n19284), .ZN(
        n19270) );
  AOI221_X1 U22380 ( .B1(n19267), .B2(n19329), .C1(n19414), .C2(n19329), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19268) );
  OAI21_X1 U22381 ( .B1(n19355), .B2(n19268), .A(n19415), .ZN(n19285) );
  AOI22_X1 U22382 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19285), .B1(
        n19456), .B2(n19350), .ZN(n19269) );
  OAI211_X1 U22383 ( .C1(n19392), .C2(n19309), .A(n19270), .B(n19269), .ZN(
        P3_U2932) );
  AOI22_X1 U22384 ( .A1(n19461), .A2(n19311), .B1(n19460), .B2(n19284), .ZN(
        n19272) );
  AOI22_X1 U22385 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19285), .B1(
        n19462), .B2(n19355), .ZN(n19271) );
  OAI211_X1 U22386 ( .C1(n19465), .C2(n19288), .A(n19272), .B(n19271), .ZN(
        P3_U2933) );
  AOI22_X1 U22387 ( .A1(n19466), .A2(n19284), .B1(n19426), .B2(n19311), .ZN(
        n19274) );
  AOI22_X1 U22388 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19285), .B1(
        n19468), .B2(n19355), .ZN(n19273) );
  OAI211_X1 U22389 ( .C1(n19429), .C2(n19288), .A(n19274), .B(n19273), .ZN(
        P3_U2934) );
  AOI22_X1 U22390 ( .A1(n19472), .A2(n19284), .B1(n19430), .B2(n19281), .ZN(
        n19276) );
  AOI22_X1 U22391 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19285), .B1(
        n19474), .B2(n19350), .ZN(n19275) );
  OAI211_X1 U22392 ( .C1(n19433), .C2(n19309), .A(n19276), .B(n19275), .ZN(
        P3_U2935) );
  AOI22_X1 U22393 ( .A1(n19434), .A2(n19281), .B1(n19478), .B2(n19284), .ZN(
        n19278) );
  AOI22_X1 U22394 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19285), .B1(
        n19480), .B2(n19350), .ZN(n19277) );
  OAI211_X1 U22395 ( .C1(n19437), .C2(n19309), .A(n19278), .B(n19277), .ZN(
        P3_U2936) );
  AOI22_X1 U22396 ( .A1(n19303), .A2(n19311), .B1(n19484), .B2(n19284), .ZN(
        n19280) );
  AOI22_X1 U22397 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19285), .B1(
        n19486), .B2(n19355), .ZN(n19279) );
  OAI211_X1 U22398 ( .C1(n19306), .C2(n19288), .A(n19280), .B(n19279), .ZN(
        P3_U2937) );
  AOI22_X1 U22399 ( .A1(n19491), .A2(n19281), .B1(n19490), .B2(n19284), .ZN(
        n19283) );
  AOI22_X1 U22400 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19285), .B1(
        n19493), .B2(n19355), .ZN(n19282) );
  OAI211_X1 U22401 ( .C1(n19496), .C2(n19309), .A(n19283), .B(n19282), .ZN(
        P3_U2938) );
  AOI22_X1 U22402 ( .A1(n19499), .A2(n19284), .B1(n19500), .B2(n19311), .ZN(
        n19287) );
  AOI22_X1 U22403 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19285), .B1(
        n19503), .B2(n19350), .ZN(n19286) );
  OAI211_X1 U22404 ( .C1(n19507), .C2(n19288), .A(n19287), .B(n19286), .ZN(
        P3_U2939) );
  NOR2_X1 U22405 ( .A1(n19340), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19290) );
  AND2_X1 U22406 ( .A1(n19449), .A2(n19290), .ZN(n19310) );
  AOI22_X1 U22407 ( .A1(n19419), .A2(n19311), .B1(n19450), .B2(n19310), .ZN(
        n19294) );
  NOR2_X1 U22408 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19289), .ZN(
        n19291) );
  AOI22_X1 U22409 ( .A1(n19455), .A2(n19291), .B1(n19453), .B2(n19290), .ZN(
        n19312) );
  NOR2_X2 U22410 ( .A1(n19340), .A2(n19292), .ZN(n19383) );
  AOI22_X1 U22411 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19312), .B1(
        n19456), .B2(n19383), .ZN(n19293) );
  OAI211_X1 U22412 ( .C1(n19392), .C2(n19329), .A(n19294), .B(n19293), .ZN(
        P3_U2940) );
  AOI22_X1 U22413 ( .A1(n19460), .A2(n19310), .B1(n19422), .B2(n19311), .ZN(
        n19296) );
  AOI22_X1 U22414 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19312), .B1(
        n19461), .B2(n19335), .ZN(n19295) );
  OAI211_X1 U22415 ( .C1(n19345), .C2(n19376), .A(n19296), .B(n19295), .ZN(
        P3_U2941) );
  AOI22_X1 U22416 ( .A1(n19466), .A2(n19310), .B1(n19426), .B2(n19335), .ZN(
        n19298) );
  AOI22_X1 U22417 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19312), .B1(
        n19468), .B2(n19383), .ZN(n19297) );
  OAI211_X1 U22418 ( .C1(n19429), .C2(n19309), .A(n19298), .B(n19297), .ZN(
        P3_U2942) );
  AOI22_X1 U22419 ( .A1(n19473), .A2(n19335), .B1(n19472), .B2(n19310), .ZN(
        n19300) );
  AOI22_X1 U22420 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19312), .B1(
        n19474), .B2(n19383), .ZN(n19299) );
  OAI211_X1 U22421 ( .C1(n19477), .C2(n19309), .A(n19300), .B(n19299), .ZN(
        P3_U2943) );
  AOI22_X1 U22422 ( .A1(n19479), .A2(n19335), .B1(n19478), .B2(n19310), .ZN(
        n19302) );
  AOI22_X1 U22423 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19312), .B1(
        n19480), .B2(n19383), .ZN(n19301) );
  OAI211_X1 U22424 ( .C1(n19483), .C2(n19309), .A(n19302), .B(n19301), .ZN(
        P3_U2944) );
  AOI22_X1 U22425 ( .A1(n19303), .A2(n19335), .B1(n19484), .B2(n19310), .ZN(
        n19305) );
  AOI22_X1 U22426 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19312), .B1(
        n19486), .B2(n19383), .ZN(n19304) );
  OAI211_X1 U22427 ( .C1(n19306), .C2(n19309), .A(n19305), .B(n19304), .ZN(
        P3_U2945) );
  AOI22_X1 U22428 ( .A1(n19404), .A2(n19335), .B1(n19490), .B2(n19310), .ZN(
        n19308) );
  AOI22_X1 U22429 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19312), .B1(
        n19493), .B2(n19383), .ZN(n19307) );
  OAI211_X1 U22430 ( .C1(n19407), .C2(n19309), .A(n19308), .B(n19307), .ZN(
        P3_U2946) );
  AOI22_X1 U22431 ( .A1(n19384), .A2(n19311), .B1(n19499), .B2(n19310), .ZN(
        n19314) );
  AOI22_X1 U22432 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19312), .B1(
        n19503), .B2(n19383), .ZN(n19313) );
  OAI211_X1 U22433 ( .C1(n19387), .C2(n19329), .A(n19314), .B(n19313), .ZN(
        P3_U2947) );
  NAND2_X1 U22434 ( .A1(n19449), .A2(n19315), .ZN(n19417) );
  NOR2_X1 U22435 ( .A1(n19340), .A2(n19417), .ZN(n19334) );
  AOI22_X1 U22436 ( .A1(n19451), .A2(n19350), .B1(n19450), .B2(n19334), .ZN(
        n19320) );
  NOR2_X2 U22437 ( .A1(n19316), .A2(n19340), .ZN(n19401) );
  NOR2_X1 U22438 ( .A1(n19335), .A2(n19355), .ZN(n19317) );
  AOI221_X1 U22439 ( .B1(n19317), .B2(n19376), .C1(n19414), .C2(n19376), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19318) );
  OAI21_X1 U22440 ( .B1(n19401), .B2(n19318), .A(n19415), .ZN(n19336) );
  AOI22_X1 U22441 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19336), .B1(
        n19456), .B2(n19401), .ZN(n19319) );
  OAI211_X1 U22442 ( .C1(n19459), .C2(n19329), .A(n19320), .B(n19319), .ZN(
        P3_U2948) );
  AOI22_X1 U22443 ( .A1(n19460), .A2(n19334), .B1(n19422), .B2(n19335), .ZN(
        n19322) );
  AOI22_X1 U22444 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19336), .B1(
        n19461), .B2(n19350), .ZN(n19321) );
  OAI211_X1 U22445 ( .C1(n19345), .C2(n19412), .A(n19322), .B(n19321), .ZN(
        P3_U2949) );
  AOI22_X1 U22446 ( .A1(n19466), .A2(n19334), .B1(n19426), .B2(n19355), .ZN(
        n19324) );
  AOI22_X1 U22447 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19336), .B1(
        n19468), .B2(n19401), .ZN(n19323) );
  OAI211_X1 U22448 ( .C1(n19429), .C2(n19329), .A(n19324), .B(n19323), .ZN(
        P3_U2950) );
  AOI22_X1 U22449 ( .A1(n19473), .A2(n19355), .B1(n19472), .B2(n19334), .ZN(
        n19326) );
  AOI22_X1 U22450 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19336), .B1(
        n19474), .B2(n19401), .ZN(n19325) );
  OAI211_X1 U22451 ( .C1(n19477), .C2(n19329), .A(n19326), .B(n19325), .ZN(
        P3_U2951) );
  AOI22_X1 U22452 ( .A1(n19479), .A2(n19355), .B1(n19478), .B2(n19334), .ZN(
        n19328) );
  AOI22_X1 U22453 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19336), .B1(
        n19480), .B2(n19401), .ZN(n19327) );
  OAI211_X1 U22454 ( .C1(n19483), .C2(n19329), .A(n19328), .B(n19327), .ZN(
        P3_U2952) );
  AOI22_X1 U22455 ( .A1(n19484), .A2(n19334), .B1(n19485), .B2(n19335), .ZN(
        n19331) );
  AOI22_X1 U22456 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19336), .B1(
        n19486), .B2(n19401), .ZN(n19330) );
  OAI211_X1 U22457 ( .C1(n19489), .C2(n19362), .A(n19331), .B(n19330), .ZN(
        P3_U2953) );
  AOI22_X1 U22458 ( .A1(n19491), .A2(n19335), .B1(n19490), .B2(n19334), .ZN(
        n19333) );
  AOI22_X1 U22459 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19336), .B1(
        n19493), .B2(n19401), .ZN(n19332) );
  OAI211_X1 U22460 ( .C1(n19496), .C2(n19362), .A(n19333), .B(n19332), .ZN(
        P3_U2954) );
  AOI22_X1 U22461 ( .A1(n19384), .A2(n19335), .B1(n19499), .B2(n19334), .ZN(
        n19338) );
  AOI22_X1 U22462 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19336), .B1(
        n19503), .B2(n19401), .ZN(n19337) );
  OAI211_X1 U22463 ( .C1(n19387), .C2(n19362), .A(n19338), .B(n19337), .ZN(
        P3_U2955) );
  NOR2_X1 U22464 ( .A1(n19553), .A2(n19340), .ZN(n19389) );
  AND2_X1 U22465 ( .A1(n19449), .A2(n19389), .ZN(n19358) );
  AOI22_X1 U22466 ( .A1(n19451), .A2(n19383), .B1(n19450), .B2(n19358), .ZN(
        n19342) );
  OAI211_X1 U22467 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19455), .A(
        n19453), .B(n19339), .ZN(n19359) );
  NOR2_X2 U22468 ( .A1(n19552), .A2(n19340), .ZN(n19440) );
  AOI22_X1 U22469 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19456), .ZN(n19341) );
  OAI211_X1 U22470 ( .C1(n19459), .C2(n19362), .A(n19342), .B(n19341), .ZN(
        P3_U2956) );
  INV_X1 U22471 ( .A(n19440), .ZN(n19448) );
  AOI22_X1 U22472 ( .A1(n19460), .A2(n19358), .B1(n19422), .B2(n19355), .ZN(
        n19344) );
  AOI22_X1 U22473 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19359), .B1(
        n19461), .B2(n19383), .ZN(n19343) );
  OAI211_X1 U22474 ( .C1(n19448), .C2(n19345), .A(n19344), .B(n19343), .ZN(
        P3_U2957) );
  AOI22_X1 U22475 ( .A1(n19467), .A2(n19350), .B1(n19466), .B2(n19358), .ZN(
        n19347) );
  AOI22_X1 U22476 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19468), .ZN(n19346) );
  OAI211_X1 U22477 ( .C1(n19471), .C2(n19376), .A(n19347), .B(n19346), .ZN(
        P3_U2958) );
  AOI22_X1 U22478 ( .A1(n19472), .A2(n19358), .B1(n19430), .B2(n19350), .ZN(
        n19349) );
  AOI22_X1 U22479 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19474), .ZN(n19348) );
  OAI211_X1 U22480 ( .C1(n19433), .C2(n19376), .A(n19349), .B(n19348), .ZN(
        P3_U2959) );
  AOI22_X1 U22481 ( .A1(n19434), .A2(n19350), .B1(n19478), .B2(n19358), .ZN(
        n19352) );
  AOI22_X1 U22482 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19480), .ZN(n19351) );
  OAI211_X1 U22483 ( .C1(n19437), .C2(n19376), .A(n19352), .B(n19351), .ZN(
        P3_U2960) );
  AOI22_X1 U22484 ( .A1(n19484), .A2(n19358), .B1(n19485), .B2(n19355), .ZN(
        n19354) );
  AOI22_X1 U22485 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19486), .ZN(n19353) );
  OAI211_X1 U22486 ( .C1(n19489), .C2(n19376), .A(n19354), .B(n19353), .ZN(
        P3_U2961) );
  AOI22_X1 U22487 ( .A1(n19491), .A2(n19355), .B1(n19490), .B2(n19358), .ZN(
        n19357) );
  AOI22_X1 U22488 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19493), .ZN(n19356) );
  OAI211_X1 U22489 ( .C1(n19496), .C2(n19376), .A(n19357), .B(n19356), .ZN(
        P3_U2962) );
  AOI22_X1 U22490 ( .A1(n19499), .A2(n19358), .B1(n19500), .B2(n19383), .ZN(
        n19361) );
  AOI22_X1 U22491 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19359), .B1(
        n19440), .B2(n19503), .ZN(n19360) );
  OAI211_X1 U22492 ( .C1(n19507), .C2(n19362), .A(n19361), .B(n19360), .ZN(
        P3_U2963) );
  INV_X1 U22493 ( .A(n19454), .ZN(n19388) );
  NOR2_X2 U22494 ( .A1(n19388), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19492) );
  NOR2_X1 U22495 ( .A1(n19492), .A2(n19440), .ZN(n19413) );
  NOR2_X1 U22496 ( .A1(n19576), .A2(n19413), .ZN(n19381) );
  AOI22_X1 U22497 ( .A1(n19419), .A2(n19383), .B1(n19450), .B2(n19381), .ZN(
        n19367) );
  OAI21_X1 U22498 ( .B1(n19364), .B2(n19363), .A(n19413), .ZN(n19365) );
  OAI211_X1 U22499 ( .C1(n19492), .C2(n19666), .A(n19415), .B(n19365), .ZN(
        n19382) );
  AOI22_X1 U22500 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19382), .B1(
        n19492), .B2(n19456), .ZN(n19366) );
  OAI211_X1 U22501 ( .C1(n19392), .C2(n19412), .A(n19367), .B(n19366), .ZN(
        P3_U2964) );
  AOI22_X1 U22502 ( .A1(n19461), .A2(n19401), .B1(n19460), .B2(n19381), .ZN(
        n19369) );
  AOI22_X1 U22503 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19382), .B1(
        n19492), .B2(n19462), .ZN(n19368) );
  OAI211_X1 U22504 ( .C1(n19465), .C2(n19376), .A(n19369), .B(n19368), .ZN(
        P3_U2965) );
  AOI22_X1 U22505 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19382), .B1(
        n19466), .B2(n19381), .ZN(n19371) );
  AOI22_X1 U22506 ( .A1(n19492), .A2(n19468), .B1(n19467), .B2(n19383), .ZN(
        n19370) );
  OAI211_X1 U22507 ( .C1(n19471), .C2(n19412), .A(n19371), .B(n19370), .ZN(
        P3_U2966) );
  AOI22_X1 U22508 ( .A1(n19472), .A2(n19381), .B1(n19430), .B2(n19383), .ZN(
        n19373) );
  AOI22_X1 U22509 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19382), .B1(
        n19492), .B2(n19474), .ZN(n19372) );
  OAI211_X1 U22510 ( .C1(n19433), .C2(n19412), .A(n19373), .B(n19372), .ZN(
        P3_U2967) );
  AOI22_X1 U22511 ( .A1(n19479), .A2(n19401), .B1(n19478), .B2(n19381), .ZN(
        n19375) );
  AOI22_X1 U22512 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19382), .B1(
        n19492), .B2(n19480), .ZN(n19374) );
  OAI211_X1 U22513 ( .C1(n19483), .C2(n19376), .A(n19375), .B(n19374), .ZN(
        P3_U2968) );
  AOI22_X1 U22514 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19382), .B1(
        n19484), .B2(n19381), .ZN(n19378) );
  AOI22_X1 U22515 ( .A1(n19492), .A2(n19486), .B1(n19485), .B2(n19383), .ZN(
        n19377) );
  OAI211_X1 U22516 ( .C1(n19489), .C2(n19412), .A(n19378), .B(n19377), .ZN(
        P3_U2969) );
  AOI22_X1 U22517 ( .A1(n19491), .A2(n19383), .B1(n19490), .B2(n19381), .ZN(
        n19380) );
  AOI22_X1 U22518 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19382), .B1(
        n19492), .B2(n19493), .ZN(n19379) );
  OAI211_X1 U22519 ( .C1(n19496), .C2(n19412), .A(n19380), .B(n19379), .ZN(
        P3_U2970) );
  AOI22_X1 U22520 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19382), .B1(
        n19499), .B2(n19381), .ZN(n19386) );
  AOI22_X1 U22521 ( .A1(n19492), .A2(n19503), .B1(n19384), .B2(n19383), .ZN(
        n19385) );
  OAI211_X1 U22522 ( .C1(n19387), .C2(n19412), .A(n19386), .B(n19385), .ZN(
        P3_U2971) );
  NOR2_X1 U22523 ( .A1(n19576), .A2(n19388), .ZN(n19408) );
  AOI22_X1 U22524 ( .A1(n19419), .A2(n19401), .B1(n19450), .B2(n19408), .ZN(
        n19391) );
  AOI22_X1 U22525 ( .A1(n19455), .A2(n19389), .B1(n19454), .B2(n19453), .ZN(
        n19409) );
  AOI22_X1 U22526 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19456), .ZN(n19390) );
  OAI211_X1 U22527 ( .C1(n19448), .C2(n19392), .A(n19391), .B(n19390), .ZN(
        P3_U2972) );
  AOI22_X1 U22528 ( .A1(n19440), .A2(n19461), .B1(n19460), .B2(n19408), .ZN(
        n19394) );
  AOI22_X1 U22529 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19462), .ZN(n19393) );
  OAI211_X1 U22530 ( .C1(n19465), .C2(n19412), .A(n19394), .B(n19393), .ZN(
        P3_U2973) );
  AOI22_X1 U22531 ( .A1(n19467), .A2(n19401), .B1(n19466), .B2(n19408), .ZN(
        n19396) );
  AOI22_X1 U22532 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19468), .ZN(n19395) );
  OAI211_X1 U22533 ( .C1(n19448), .C2(n19471), .A(n19396), .B(n19395), .ZN(
        P3_U2974) );
  AOI22_X1 U22534 ( .A1(n19440), .A2(n19473), .B1(n19472), .B2(n19408), .ZN(
        n19398) );
  AOI22_X1 U22535 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19474), .ZN(n19397) );
  OAI211_X1 U22536 ( .C1(n19477), .C2(n19412), .A(n19398), .B(n19397), .ZN(
        P3_U2975) );
  AOI22_X1 U22537 ( .A1(n19440), .A2(n19479), .B1(n19478), .B2(n19408), .ZN(
        n19400) );
  AOI22_X1 U22538 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19480), .ZN(n19399) );
  OAI211_X1 U22539 ( .C1(n19483), .C2(n19412), .A(n19400), .B(n19399), .ZN(
        P3_U2976) );
  AOI22_X1 U22540 ( .A1(n19484), .A2(n19408), .B1(n19485), .B2(n19401), .ZN(
        n19403) );
  AOI22_X1 U22541 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19486), .ZN(n19402) );
  OAI211_X1 U22542 ( .C1(n19448), .C2(n19489), .A(n19403), .B(n19402), .ZN(
        P3_U2977) );
  AOI22_X1 U22543 ( .A1(n19440), .A2(n19404), .B1(n19490), .B2(n19408), .ZN(
        n19406) );
  AOI22_X1 U22544 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19493), .ZN(n19405) );
  OAI211_X1 U22545 ( .C1(n19407), .C2(n19412), .A(n19406), .B(n19405), .ZN(
        P3_U2978) );
  AOI22_X1 U22546 ( .A1(n19440), .A2(n19500), .B1(n19499), .B2(n19408), .ZN(
        n19411) );
  AOI22_X1 U22547 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19409), .B1(
        n19501), .B2(n19503), .ZN(n19410) );
  OAI211_X1 U22548 ( .C1(n19507), .C2(n19412), .A(n19411), .B(n19410), .ZN(
        P3_U2979) );
  AOI221_X1 U22549 ( .B1(n19497), .B2(n19414), .C1(n19497), .C2(n19413), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19416) );
  OAI21_X1 U22550 ( .B1(n19444), .B2(n19416), .A(n19415), .ZN(n19445) );
  INV_X1 U22551 ( .A(n19445), .ZN(n19425) );
  NOR2_X1 U22552 ( .A1(n19418), .A2(n19417), .ZN(n19443) );
  AOI22_X1 U22553 ( .A1(n19440), .A2(n19419), .B1(n19450), .B2(n19443), .ZN(
        n19421) );
  AOI22_X1 U22554 ( .A1(n19444), .A2(n19456), .B1(n19492), .B2(n19451), .ZN(
        n19420) );
  OAI211_X1 U22555 ( .C1(n19425), .C2(n21634), .A(n19421), .B(n19420), .ZN(
        P3_U2980) );
  AOI22_X1 U22556 ( .A1(n19440), .A2(n19422), .B1(n19443), .B2(n19460), .ZN(
        n19424) );
  AOI22_X1 U22557 ( .A1(n19444), .A2(n19462), .B1(n19492), .B2(n19461), .ZN(
        n19423) );
  OAI211_X1 U22558 ( .C1(n19425), .C2(n21495), .A(n19424), .B(n19423), .ZN(
        P3_U2981) );
  AOI22_X1 U22559 ( .A1(n19492), .A2(n19426), .B1(n19443), .B2(n19466), .ZN(
        n19428) );
  AOI22_X1 U22560 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19445), .B1(
        n19444), .B2(n19468), .ZN(n19427) );
  OAI211_X1 U22561 ( .C1(n19448), .C2(n19429), .A(n19428), .B(n19427), .ZN(
        P3_U2982) );
  INV_X1 U22562 ( .A(n19492), .ZN(n19508) );
  AOI22_X1 U22563 ( .A1(n19440), .A2(n19430), .B1(n19443), .B2(n19472), .ZN(
        n19432) );
  AOI22_X1 U22564 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19445), .B1(
        n19444), .B2(n19474), .ZN(n19431) );
  OAI211_X1 U22565 ( .C1(n19508), .C2(n19433), .A(n19432), .B(n19431), .ZN(
        P3_U2983) );
  AOI22_X1 U22566 ( .A1(n19440), .A2(n19434), .B1(n19443), .B2(n19478), .ZN(
        n19436) );
  AOI22_X1 U22567 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19445), .B1(
        n19444), .B2(n19480), .ZN(n19435) );
  OAI211_X1 U22568 ( .C1(n19508), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P3_U2984) );
  AOI22_X1 U22569 ( .A1(n19440), .A2(n19485), .B1(n19443), .B2(n19484), .ZN(
        n19439) );
  AOI22_X1 U22570 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19445), .B1(
        n19444), .B2(n19486), .ZN(n19438) );
  OAI211_X1 U22571 ( .C1(n19508), .C2(n19489), .A(n19439), .B(n19438), .ZN(
        P3_U2985) );
  AOI22_X1 U22572 ( .A1(n19440), .A2(n19491), .B1(n19443), .B2(n19490), .ZN(
        n19442) );
  AOI22_X1 U22573 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19445), .B1(
        n19444), .B2(n19493), .ZN(n19441) );
  OAI211_X1 U22574 ( .C1(n19508), .C2(n19496), .A(n19442), .B(n19441), .ZN(
        P3_U2986) );
  AOI22_X1 U22575 ( .A1(n19492), .A2(n19500), .B1(n19443), .B2(n19499), .ZN(
        n19447) );
  AOI22_X1 U22576 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19445), .B1(
        n19444), .B2(n19503), .ZN(n19446) );
  OAI211_X1 U22577 ( .C1(n19448), .C2(n19507), .A(n19447), .B(n19446), .ZN(
        P3_U2987) );
  AND2_X1 U22578 ( .A1(n19449), .A2(n19452), .ZN(n19498) );
  AOI22_X1 U22579 ( .A1(n19501), .A2(n19451), .B1(n19450), .B2(n19498), .ZN(
        n19458) );
  AOI22_X1 U22580 ( .A1(n19455), .A2(n19454), .B1(n19453), .B2(n19452), .ZN(
        n19504) );
  AOI22_X1 U22581 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19504), .B1(
        n19456), .B2(n19502), .ZN(n19457) );
  OAI211_X1 U22582 ( .C1(n19508), .C2(n19459), .A(n19458), .B(n19457), .ZN(
        P3_U2988) );
  AOI22_X1 U22583 ( .A1(n19501), .A2(n19461), .B1(n19460), .B2(n19498), .ZN(
        n19464) );
  AOI22_X1 U22584 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19504), .B1(
        n19462), .B2(n19502), .ZN(n19463) );
  OAI211_X1 U22585 ( .C1(n19508), .C2(n19465), .A(n19464), .B(n19463), .ZN(
        P3_U2989) );
  AOI22_X1 U22586 ( .A1(n19492), .A2(n19467), .B1(n19466), .B2(n19498), .ZN(
        n19470) );
  AOI22_X1 U22587 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19504), .B1(
        n19468), .B2(n19502), .ZN(n19469) );
  OAI211_X1 U22588 ( .C1(n19497), .C2(n19471), .A(n19470), .B(n19469), .ZN(
        P3_U2990) );
  AOI22_X1 U22589 ( .A1(n19501), .A2(n19473), .B1(n19472), .B2(n19498), .ZN(
        n19476) );
  AOI22_X1 U22590 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19504), .B1(
        n19474), .B2(n19502), .ZN(n19475) );
  OAI211_X1 U22591 ( .C1(n19508), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P3_U2991) );
  AOI22_X1 U22592 ( .A1(n19501), .A2(n19479), .B1(n19478), .B2(n19498), .ZN(
        n19482) );
  AOI22_X1 U22593 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19504), .B1(
        n19480), .B2(n19502), .ZN(n19481) );
  OAI211_X1 U22594 ( .C1(n19508), .C2(n19483), .A(n19482), .B(n19481), .ZN(
        P3_U2992) );
  AOI22_X1 U22595 ( .A1(n19492), .A2(n19485), .B1(n19484), .B2(n19498), .ZN(
        n19488) );
  AOI22_X1 U22596 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19504), .B1(
        n19486), .B2(n19502), .ZN(n19487) );
  OAI211_X1 U22597 ( .C1(n19497), .C2(n19489), .A(n19488), .B(n19487), .ZN(
        P3_U2993) );
  AOI22_X1 U22598 ( .A1(n19492), .A2(n19491), .B1(n19490), .B2(n19498), .ZN(
        n19495) );
  AOI22_X1 U22599 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19504), .B1(
        n19493), .B2(n19502), .ZN(n19494) );
  OAI211_X1 U22600 ( .C1(n19497), .C2(n19496), .A(n19495), .B(n19494), .ZN(
        P3_U2994) );
  AOI22_X1 U22601 ( .A1(n19501), .A2(n19500), .B1(n19499), .B2(n19498), .ZN(
        n19506) );
  AOI22_X1 U22602 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19502), .ZN(n19505) );
  OAI211_X1 U22603 ( .C1(n19508), .C2(n19507), .A(n19506), .B(n19505), .ZN(
        P3_U2995) );
  NOR2_X1 U22604 ( .A1(n19544), .A2(n19509), .ZN(n19512) );
  OAI222_X1 U22605 ( .A1(n19515), .A2(n19514), .B1(n19513), .B2(n19512), .C1(
        n19511), .C2(n19510), .ZN(n19709) );
  OAI21_X1 U22606 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19516), .ZN(n19517) );
  OAI211_X1 U22607 ( .C1(n19545), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        n19563) );
  NAND2_X1 U22608 ( .A1(n19535), .A2(n19521), .ZN(n19549) );
  AOI22_X1 U22609 ( .A1(n19528), .A2(n19549), .B1(n19544), .B2(n19527), .ZN(
        n19522) );
  NOR2_X1 U22610 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19522), .ZN(
        n19669) );
  AOI21_X1 U22611 ( .B1(n19525), .B2(n19524), .A(n19523), .ZN(n19526) );
  INV_X1 U22612 ( .A(n19526), .ZN(n19538) );
  OAI21_X1 U22613 ( .B1(n19528), .B2(n19548), .A(n19527), .ZN(n19529) );
  AOI21_X1 U22614 ( .B1(n19538), .B2(n19530), .A(n19529), .ZN(n19670) );
  NAND2_X1 U22615 ( .A1(n19545), .A2(n19670), .ZN(n19531) );
  AOI22_X1 U22616 ( .A1(n19545), .A2(n19669), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19531), .ZN(n19562) );
  INV_X1 U22617 ( .A(n19545), .ZN(n19556) );
  OAI211_X1 U22618 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n19533), .B(n19532), .ZN(
        n19534) );
  INV_X1 U22619 ( .A(n19534), .ZN(n19543) );
  NOR2_X1 U22620 ( .A1(n19535), .A2(n19689), .ZN(n19541) );
  OAI221_X1 U22621 ( .B1(n19538), .B2(n19689), .C1(n19538), .C2(n19537), .A(
        n19536), .ZN(n19539) );
  INV_X1 U22622 ( .A(n19539), .ZN(n19540) );
  MUX2_X1 U22623 ( .A(n19541), .B(n19540), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n19542) );
  AOI211_X1 U22624 ( .C1(n19544), .C2(n19677), .A(n19543), .B(n19542), .ZN(
        n19679) );
  AOI22_X1 U22625 ( .A1(n19556), .A2(n12161), .B1(n19679), .B2(n19545), .ZN(
        n19559) );
  NOR2_X1 U22626 ( .A1(n19547), .A2(n19546), .ZN(n19551) );
  INV_X1 U22627 ( .A(n19549), .ZN(n19550) );
  OAI22_X1 U22628 ( .A1(n19551), .A2(n19682), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19550), .ZN(n19687) );
  AOI222_X1 U22629 ( .A1(n19691), .A2(n19687), .B1(n19691), .B2(n19553), .C1(
        n19687), .C2(n19552), .ZN(n19555) );
  OAI21_X1 U22630 ( .B1(n19556), .B2(n19555), .A(n19554), .ZN(n19558) );
  AOI21_X1 U22631 ( .B1(n21539), .B2(n19560), .A(n19559), .ZN(n19561) );
  INV_X1 U22632 ( .A(n19678), .ZN(n19690) );
  NAND2_X1 U22633 ( .A1(n19676), .A2(n19575), .ZN(n19584) );
  INV_X1 U22634 ( .A(n19584), .ZN(n19718) );
  AOI22_X1 U22635 ( .A1(n19690), .A2(n19718), .B1(n19586), .B2(n18338), .ZN(
        n19565) );
  INV_X1 U22636 ( .A(n19565), .ZN(n19570) );
  OAI211_X1 U22637 ( .C1(n19567), .C2(n19566), .A(n19711), .B(n19574), .ZN(
        n19665) );
  OAI21_X1 U22638 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19716), .A(n19665), 
        .ZN(n19577) );
  NOR2_X1 U22639 ( .A1(n19568), .A2(n19577), .ZN(n19569) );
  MUX2_X1 U22640 ( .A(n19570), .B(n19569), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19572) );
  OAI211_X1 U22641 ( .C1(n19574), .C2(n19573), .A(n19572), .B(n19571), .ZN(
        P3_U2996) );
  NAND2_X1 U22642 ( .A1(n19586), .A2(n18338), .ZN(n19580) );
  NAND4_X1 U22643 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19586), .A4(n19575), .ZN(n19582) );
  OR3_X1 U22644 ( .A1(n19578), .A2(n19577), .A3(n19576), .ZN(n19579) );
  NAND4_X1 U22645 ( .A1(n19581), .A2(n19580), .A3(n19582), .A4(n19579), .ZN(
        P3_U2997) );
  AND4_X1 U22646 ( .A1(n19584), .A2(n19583), .A3(n19582), .A4(n19664), .ZN(
        P3_U2998) );
  INV_X1 U22647 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21590) );
  NOR2_X1 U22648 ( .A1(n21590), .A2(n19663), .ZN(P3_U2999) );
  AND2_X1 U22649 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19585), .ZN(
        P3_U3000) );
  AND2_X1 U22650 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19585), .ZN(
        P3_U3001) );
  AND2_X1 U22651 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19585), .ZN(
        P3_U3002) );
  AND2_X1 U22652 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19585), .ZN(
        P3_U3003) );
  AND2_X1 U22653 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19585), .ZN(
        P3_U3004) );
  AND2_X1 U22654 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19585), .ZN(
        P3_U3005) );
  AND2_X1 U22655 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19585), .ZN(
        P3_U3006) );
  AND2_X1 U22656 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19585), .ZN(
        P3_U3007) );
  AND2_X1 U22657 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19585), .ZN(
        P3_U3008) );
  AND2_X1 U22658 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19585), .ZN(
        P3_U3009) );
  AND2_X1 U22659 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19585), .ZN(
        P3_U3010) );
  INV_X1 U22660 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21652) );
  NOR2_X1 U22661 ( .A1(n21652), .A2(n19663), .ZN(P3_U3011) );
  AND2_X1 U22662 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19585), .ZN(
        P3_U3012) );
  AND2_X1 U22663 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19585), .ZN(
        P3_U3013) );
  AND2_X1 U22664 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19585), .ZN(
        P3_U3014) );
  AND2_X1 U22665 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19585), .ZN(
        P3_U3015) );
  AND2_X1 U22666 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19585), .ZN(
        P3_U3016) );
  AND2_X1 U22667 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19585), .ZN(
        P3_U3017) );
  AND2_X1 U22668 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19585), .ZN(
        P3_U3018) );
  AND2_X1 U22669 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19585), .ZN(
        P3_U3019) );
  AND2_X1 U22670 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19585), .ZN(
        P3_U3020) );
  AND2_X1 U22671 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19585), .ZN(P3_U3021) );
  INV_X1 U22672 ( .A(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21700) );
  NOR2_X1 U22673 ( .A1(n21700), .A2(n19663), .ZN(P3_U3022) );
  AND2_X1 U22674 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19585), .ZN(P3_U3023) );
  INV_X1 U22675 ( .A(P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n21650) );
  NOR2_X1 U22676 ( .A1(n21650), .A2(n19663), .ZN(P3_U3024) );
  AND2_X1 U22677 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19585), .ZN(P3_U3025) );
  INV_X1 U22678 ( .A(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21577) );
  NOR2_X1 U22679 ( .A1(n21577), .A2(n19663), .ZN(P3_U3026) );
  AND2_X1 U22680 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19585), .ZN(P3_U3027) );
  AND2_X1 U22681 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19585), .ZN(P3_U3028) );
  NOR2_X1 U22682 ( .A1(n17354), .A2(n21335), .ZN(n19596) );
  INV_X1 U22683 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21492) );
  AOI211_X1 U22684 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n19596), .B(
        n21492), .ZN(n19588) );
  NAND2_X1 U22685 ( .A1(n19586), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19594) );
  INV_X1 U22686 ( .A(n19594), .ZN(n19592) );
  OAI21_X1 U22687 ( .B1(n19592), .B2(n19598), .A(n17354), .ZN(n19587) );
  INV_X1 U22688 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21574) );
  NAND3_X1 U22689 ( .A1(NA), .A2(n21574), .A3(n19598), .ZN(n19593) );
  OAI211_X1 U22690 ( .C1(n19723), .C2(n19588), .A(n19587), .B(n19593), .ZN(
        P3_U3029) );
  NOR2_X1 U22691 ( .A1(n19596), .A2(n21492), .ZN(n19590) );
  NOR2_X1 U22692 ( .A1(n21574), .A2(n21335), .ZN(n19589) );
  AOI22_X1 U22693 ( .A1(n19590), .A2(P3_STATE_REG_0__SCAN_IN), .B1(n19589), 
        .B2(n17354), .ZN(n19591) );
  NAND3_X1 U22694 ( .A1(n19591), .A2(n19713), .A3(n19594), .ZN(P3_U3030) );
  AOI21_X1 U22695 ( .B1(n19598), .B2(n19593), .A(n19592), .ZN(n19599) );
  OAI22_X1 U22696 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19594), .ZN(n19595) );
  OAI22_X1 U22697 ( .A1(n19596), .A2(n19595), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19597) );
  OAI22_X1 U22698 ( .A1(n19599), .A2(n17354), .B1(n19598), .B2(n19597), .ZN(
        P3_U3031) );
  NAND2_X1 U22699 ( .A1(n19723), .A2(n17354), .ZN(n19638) );
  CLKBUF_X1 U22700 ( .A(n19638), .Z(n19651) );
  OAI222_X1 U22701 ( .A1(n19698), .A2(n19648), .B1(n19600), .B2(n19723), .C1(
        n19601), .C2(n19651), .ZN(P3_U3032) );
  OAI222_X1 U22702 ( .A1(n19638), .A2(n19603), .B1(n19602), .B2(n19723), .C1(
        n19601), .C2(n19648), .ZN(P3_U3033) );
  OAI222_X1 U22703 ( .A1(n19638), .A2(n21656), .B1(n19604), .B2(n19723), .C1(
        n19603), .C2(n19648), .ZN(P3_U3034) );
  OAI222_X1 U22704 ( .A1(n19638), .A2(n19606), .B1(n21501), .B2(n19723), .C1(
        n21656), .C2(n19648), .ZN(P3_U3035) );
  OAI222_X1 U22705 ( .A1(n19606), .A2(n19648), .B1(n19605), .B2(n19723), .C1(
        n19607), .C2(n19651), .ZN(P3_U3036) );
  OAI222_X1 U22706 ( .A1(n19638), .A2(n19609), .B1(n19608), .B2(n19723), .C1(
        n19607), .C2(n19648), .ZN(P3_U3037) );
  OAI222_X1 U22707 ( .A1(n19638), .A2(n19611), .B1(n21720), .B2(n19723), .C1(
        n19609), .C2(n19648), .ZN(P3_U3038) );
  OAI222_X1 U22708 ( .A1(n19611), .A2(n19648), .B1(n19610), .B2(n19723), .C1(
        n19612), .C2(n19651), .ZN(P3_U3039) );
  OAI222_X1 U22709 ( .A1(n19638), .A2(n19614), .B1(n19613), .B2(n19723), .C1(
        n19612), .C2(n19648), .ZN(P3_U3040) );
  OAI222_X1 U22710 ( .A1(n19638), .A2(n21642), .B1(n19615), .B2(n19723), .C1(
        n19614), .C2(n19648), .ZN(P3_U3041) );
  OAI222_X1 U22711 ( .A1(n19651), .A2(n19617), .B1(n19616), .B2(n19723), .C1(
        n21642), .C2(n19648), .ZN(P3_U3042) );
  OAI222_X1 U22712 ( .A1(n19651), .A2(n19619), .B1(n19618), .B2(n19723), .C1(
        n19617), .C2(n19648), .ZN(P3_U3043) );
  OAI222_X1 U22713 ( .A1(n19651), .A2(n19621), .B1(n19620), .B2(n19723), .C1(
        n19619), .C2(n19648), .ZN(P3_U3044) );
  OAI222_X1 U22714 ( .A1(n19651), .A2(n19623), .B1(n19622), .B2(n19723), .C1(
        n19621), .C2(n19655), .ZN(P3_U3045) );
  OAI222_X1 U22715 ( .A1(n19651), .A2(n19625), .B1(n19624), .B2(n19723), .C1(
        n19623), .C2(n19655), .ZN(P3_U3046) );
  INV_X1 U22716 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19627) );
  OAI222_X1 U22717 ( .A1(n19651), .A2(n19627), .B1(n19626), .B2(n19723), .C1(
        n19625), .C2(n19655), .ZN(P3_U3047) );
  OAI222_X1 U22718 ( .A1(n19638), .A2(n19629), .B1(n19628), .B2(n19723), .C1(
        n19627), .C2(n19655), .ZN(P3_U3048) );
  OAI222_X1 U22719 ( .A1(n19638), .A2(n19631), .B1(n19630), .B2(n19723), .C1(
        n19629), .C2(n19655), .ZN(P3_U3049) );
  OAI222_X1 U22720 ( .A1(n19638), .A2(n21658), .B1(n19632), .B2(n19723), .C1(
        n19631), .C2(n19655), .ZN(P3_U3050) );
  OAI222_X1 U22721 ( .A1(n21658), .A2(n19648), .B1(n19633), .B2(n19723), .C1(
        n21584), .C2(n19651), .ZN(P3_U3051) );
  OAI222_X1 U22722 ( .A1(n21584), .A2(n19648), .B1(n19634), .B2(n19723), .C1(
        n21609), .C2(n19651), .ZN(P3_U3052) );
  OAI222_X1 U22723 ( .A1(n19638), .A2(n19636), .B1(n19635), .B2(n19723), .C1(
        n21609), .C2(n19655), .ZN(P3_U3053) );
  OAI222_X1 U22724 ( .A1(n19638), .A2(n19640), .B1(n19637), .B2(n19723), .C1(
        n19636), .C2(n19655), .ZN(P3_U3054) );
  OAI222_X1 U22725 ( .A1(n19640), .A2(n19648), .B1(n19639), .B2(n19723), .C1(
        n19641), .C2(n19651), .ZN(P3_U3055) );
  INV_X1 U22726 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19643) );
  OAI222_X1 U22727 ( .A1(n19651), .A2(n19643), .B1(n19642), .B2(n19723), .C1(
        n19641), .C2(n19648), .ZN(P3_U3056) );
  OAI222_X1 U22728 ( .A1(n19651), .A2(n19645), .B1(n19644), .B2(n19723), .C1(
        n19643), .C2(n19648), .ZN(P3_U3057) );
  OAI222_X1 U22729 ( .A1(n19651), .A2(n21470), .B1(n19646), .B2(n19723), .C1(
        n19645), .C2(n19655), .ZN(P3_U3058) );
  OAI222_X1 U22730 ( .A1(n21470), .A2(n19648), .B1(n19647), .B2(n19723), .C1(
        n19649), .C2(n19651), .ZN(P3_U3059) );
  OAI222_X1 U22731 ( .A1(n19651), .A2(n19654), .B1(n19650), .B2(n19723), .C1(
        n19649), .C2(n19648), .ZN(P3_U3060) );
  OAI222_X1 U22732 ( .A1(n19655), .A2(n19654), .B1(n19653), .B2(n19723), .C1(
        n19652), .C2(n19651), .ZN(P3_U3061) );
  OAI22_X1 U22733 ( .A1(n19724), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19723), .ZN(n19656) );
  INV_X1 U22734 ( .A(n19656), .ZN(P3_U3274) );
  OAI22_X1 U22735 ( .A1(n19724), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19723), .ZN(n19657) );
  INV_X1 U22736 ( .A(n19657), .ZN(P3_U3275) );
  OAI22_X1 U22737 ( .A1(n19724), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19723), .ZN(n19658) );
  INV_X1 U22738 ( .A(n19658), .ZN(P3_U3276) );
  OAI22_X1 U22739 ( .A1(n19724), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19723), .ZN(n19659) );
  INV_X1 U22740 ( .A(n19659), .ZN(P3_U3277) );
  OAI21_X1 U22741 ( .B1(n19663), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19661), 
        .ZN(n19660) );
  INV_X1 U22742 ( .A(n19660), .ZN(P3_U3280) );
  OAI21_X1 U22743 ( .B1(n19663), .B2(n19662), .A(n19661), .ZN(P3_U3281) );
  OAI221_X1 U22744 ( .B1(n19666), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19666), 
        .C2(n19665), .A(n19664), .ZN(P3_U3282) );
  INV_X1 U22745 ( .A(n19726), .ZN(n19692) );
  INV_X1 U22746 ( .A(n19667), .ZN(n19668) );
  AOI22_X1 U22747 ( .A1(n19692), .A2(n19669), .B1(n19690), .B2(n19668), .ZN(
        n19673) );
  INV_X1 U22748 ( .A(n19697), .ZN(n19694) );
  OAI21_X1 U22749 ( .B1(n19726), .B2(n19670), .A(n19694), .ZN(n19671) );
  INV_X1 U22750 ( .A(n19671), .ZN(n19672) );
  OAI22_X1 U22751 ( .A1(n19697), .A2(n19673), .B1(n19672), .B2(n12163), .ZN(
        P3_U3285) );
  OAI22_X1 U22752 ( .A1(n19675), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19674), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19683) );
  NOR2_X1 U22753 ( .A1(n19676), .A2(n19693), .ZN(n19684) );
  OAI22_X1 U22754 ( .A1(n19679), .A2(n19726), .B1(n19678), .B2(n19677), .ZN(
        n19680) );
  AOI21_X1 U22755 ( .B1(n19683), .B2(n19684), .A(n19680), .ZN(n19681) );
  AOI22_X1 U22756 ( .A1(n19697), .A2(n12161), .B1(n19681), .B2(n19694), .ZN(
        P3_U3288) );
  INV_X1 U22757 ( .A(n19682), .ZN(n19686) );
  INV_X1 U22758 ( .A(n19683), .ZN(n19685) );
  AOI222_X1 U22759 ( .A1(n19687), .A2(n19692), .B1(n19690), .B2(n19686), .C1(
        n19685), .C2(n19684), .ZN(n19688) );
  AOI22_X1 U22760 ( .A1(n19697), .A2(n19689), .B1(n19688), .B2(n19694), .ZN(
        P3_U3289) );
  AOI222_X1 U22761 ( .A1(n19693), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19692), 
        .B2(n19691), .C1(n19696), .C2(n19690), .ZN(n19695) );
  AOI22_X1 U22762 ( .A1(n19697), .A2(n19696), .B1(n19695), .B2(n19694), .ZN(
        P3_U3290) );
  AOI21_X1 U22763 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19699) );
  AOI22_X1 U22764 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19699), .B2(n19698), .ZN(n19701) );
  INV_X1 U22765 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19700) );
  AOI22_X1 U22766 ( .A1(n19702), .A2(n19701), .B1(n19700), .B2(n19705), .ZN(
        P3_U3292) );
  INV_X1 U22767 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19706) );
  NOR2_X1 U22768 ( .A1(n19705), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U22769 ( .A1(n19706), .A2(n19705), .B1(n19704), .B2(n19703), .ZN(
        P3_U3293) );
  INV_X1 U22770 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19707) );
  AOI22_X1 U22771 ( .A1(n19723), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19707), 
        .B2(n19724), .ZN(P3_U3294) );
  MUX2_X1 U22772 ( .A(P3_MORE_REG_SCAN_IN), .B(n19709), .S(n19708), .Z(
        P3_U3295) );
  OAI21_X1 U22773 ( .B1(n19711), .B2(n19710), .A(n19728), .ZN(n19712) );
  AOI21_X1 U22774 ( .B1(n18338), .B2(n19716), .A(n19712), .ZN(n19722) );
  AOI21_X1 U22775 ( .B1(n19715), .B2(n19714), .A(n19713), .ZN(n19717) );
  OAI211_X1 U22776 ( .C1(n19727), .C2(n19717), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19716), .ZN(n19719) );
  AOI21_X1 U22777 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19719), .A(n19718), 
        .ZN(n19721) );
  NAND2_X1 U22778 ( .A1(n19722), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19720) );
  OAI21_X1 U22779 ( .B1(n19722), .B2(n19721), .A(n19720), .ZN(P3_U3296) );
  OAI22_X1 U22780 ( .A1(n19724), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19723), .ZN(n19725) );
  INV_X1 U22781 ( .A(n19725), .ZN(P3_U3297) );
  OAI21_X1 U22782 ( .B1(n19726), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19728), 
        .ZN(n19731) );
  OAI22_X1 U22783 ( .A1(n19731), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19728), 
        .B2(n19727), .ZN(n19729) );
  INV_X1 U22784 ( .A(n19729), .ZN(P3_U3298) );
  OAI21_X1 U22785 ( .B1(n19731), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19730), 
        .ZN(n19732) );
  INV_X1 U22786 ( .A(n19732), .ZN(P3_U3299) );
  NAND2_X1 U22787 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20464), .ZN(n20453) );
  AOI22_X1 U22788 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20453), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19734), .ZN(n20520) );
  AOI21_X1 U22789 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20520), .ZN(n19733) );
  INV_X1 U22790 ( .A(n19733), .ZN(P2_U2815) );
  INV_X2 U22791 ( .A(n20557), .ZN(n20556) );
  AOI21_X1 U22792 ( .B1(n19734), .B2(n20464), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19735) );
  AOI22_X1 U22793 ( .A1(n20556), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19735), 
        .B2(n20557), .ZN(P2_U2817) );
  INV_X1 U22794 ( .A(n20459), .ZN(n20446) );
  OAI21_X1 U22795 ( .B1(n20446), .B2(BS16), .A(n20520), .ZN(n20518) );
  OAI21_X1 U22796 ( .B1(n20520), .B2(n20198), .A(n20518), .ZN(P2_U2818) );
  NOR2_X1 U22797 ( .A1(n19737), .A2(n19736), .ZN(n20554) );
  OAI21_X1 U22798 ( .B1(n20554), .B2(n14459), .A(n19738), .ZN(P2_U2819) );
  NOR4_X1 U22799 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19742) );
  NOR4_X1 U22800 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19741) );
  NOR4_X1 U22801 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19740) );
  NOR4_X1 U22802 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19739) );
  NAND4_X1 U22803 ( .A1(n19742), .A2(n19741), .A3(n19740), .A4(n19739), .ZN(
        n19748) );
  NOR4_X1 U22804 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19746) );
  AOI211_X1 U22805 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19745) );
  NOR4_X1 U22806 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19744) );
  NOR4_X1 U22807 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19743) );
  NAND4_X1 U22808 ( .A1(n19746), .A2(n19745), .A3(n19744), .A4(n19743), .ZN(
        n19747) );
  NOR2_X1 U22809 ( .A1(n19748), .A2(n19747), .ZN(n19757) );
  INV_X1 U22810 ( .A(n19757), .ZN(n19756) );
  NOR2_X1 U22811 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19756), .ZN(n19751) );
  INV_X1 U22812 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U22813 ( .A1(n19751), .A2(n14353), .B1(n19756), .B2(n19749), .ZN(
        P2_U2820) );
  OR3_X1 U22814 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19755) );
  INV_X1 U22815 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U22816 ( .A1(n19751), .A2(n19755), .B1(n19756), .B2(n19750), .ZN(
        P2_U2821) );
  INV_X1 U22817 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20519) );
  NAND2_X1 U22818 ( .A1(n19751), .A2(n20519), .ZN(n19754) );
  OAI21_X1 U22819 ( .B1(n14353), .B2(n20465), .A(n19757), .ZN(n19752) );
  OAI21_X1 U22820 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19757), .A(n19752), 
        .ZN(n19753) );
  OAI221_X1 U22821 ( .B1(n19754), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19754), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19753), .ZN(P2_U2822) );
  INV_X1 U22822 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21471) );
  OAI221_X1 U22823 ( .B1(n19757), .B2(n21471), .C1(n19756), .C2(n19755), .A(
        n19754), .ZN(P2_U2823) );
  AOI22_X1 U22824 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19787), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19807), .ZN(n19770) );
  AOI21_X1 U22825 ( .B1(n19789), .B2(P2_REIP_REG_17__SCAN_IN), .A(n19788), 
        .ZN(n19758) );
  OAI21_X1 U22826 ( .B1(n19765), .B2(n19826), .A(n19758), .ZN(n19759) );
  AOI21_X1 U22827 ( .B1(n19760), .B2(n19809), .A(n19759), .ZN(n19769) );
  AOI22_X1 U22828 ( .A1(n19819), .A2(n19762), .B1(n19761), .B2(n19794), .ZN(
        n19768) );
  OAI211_X1 U22829 ( .C1(n19766), .C2(n19765), .A(n19764), .B(n19763), .ZN(
        n19767) );
  NAND4_X1 U22830 ( .A1(n19770), .A2(n19769), .A3(n19768), .A4(n19767), .ZN(
        P2_U2838) );
  INV_X1 U22831 ( .A(n19771), .ZN(n19776) );
  INV_X1 U22832 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19773) );
  AOI21_X1 U22833 ( .B1(n19789), .B2(P2_REIP_REG_16__SCAN_IN), .A(n19788), 
        .ZN(n19772) );
  OAI21_X1 U22834 ( .B1(n19774), .B2(n19773), .A(n19772), .ZN(n19775) );
  AOI21_X1 U22835 ( .B1(n19776), .B2(n19809), .A(n19775), .ZN(n19786) );
  NOR2_X1 U22836 ( .A1(n19778), .A2(n19777), .ZN(n19780) );
  XNOR2_X1 U22837 ( .A(n19780), .B(n19779), .ZN(n19781) );
  AOI222_X1 U22838 ( .A1(n19784), .A2(n19819), .B1(n19783), .B2(n19794), .C1(
        n19782), .C2(n19781), .ZN(n19785) );
  OAI211_X1 U22839 ( .C1(n10723), .C2(n19815), .A(n19786), .B(n19785), .ZN(
        P2_U2839) );
  AOI22_X1 U22840 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19787), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19807), .ZN(n19806) );
  AOI21_X1 U22841 ( .B1(n19789), .B2(P2_REIP_REG_4__SCAN_IN), .A(n19788), .ZN(
        n19790) );
  OAI21_X1 U22842 ( .B1(n19792), .B2(n19791), .A(n19790), .ZN(n19793) );
  AOI21_X1 U22843 ( .B1(n19795), .B2(n19794), .A(n19793), .ZN(n19805) );
  INV_X1 U22844 ( .A(n19796), .ZN(n19823) );
  INV_X1 U22845 ( .A(n19797), .ZN(n19827) );
  AOI22_X1 U22846 ( .A1(n19829), .A2(n19823), .B1(n19819), .B2(n19827), .ZN(
        n19804) );
  AND2_X1 U22847 ( .A1(n19799), .A2(n9682), .ZN(n19801) );
  AOI21_X1 U22848 ( .B1(n19801), .B2(n19802), .A(n19820), .ZN(n19800) );
  OAI21_X1 U22849 ( .B1(n19802), .B2(n19801), .A(n19800), .ZN(n19803) );
  NAND4_X1 U22850 ( .A1(n19806), .A2(n19805), .A3(n19804), .A4(n19803), .ZN(
        P2_U2851) );
  NAND2_X1 U22851 ( .A1(n19807), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19811) );
  NAND2_X1 U22852 ( .A1(n19809), .A2(n19808), .ZN(n19810) );
  OAI211_X1 U22853 ( .C1(n19812), .C2(n20465), .A(n19811), .B(n19810), .ZN(
        n19817) );
  OAI22_X1 U22854 ( .A1(n19815), .A2(n21708), .B1(n19814), .B2(n19813), .ZN(
        n19816) );
  AOI211_X1 U22855 ( .C1(n19819), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        n19825) );
  NOR2_X1 U22856 ( .A1(n19821), .A2(n19820), .ZN(n19822) );
  AOI21_X1 U22857 ( .B1(n20524), .B2(n19823), .A(n19822), .ZN(n19824) );
  OAI211_X1 U22858 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19826), .A(
        n19825), .B(n19824), .ZN(P2_U2854) );
  INV_X1 U22859 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U22860 ( .A1(n19829), .A2(n19828), .B1(n19832), .B2(n19827), .ZN(
        n19830) );
  OAI21_X1 U22861 ( .B1(n19832), .B2(n19831), .A(n19830), .ZN(P2_U2883) );
  INV_X1 U22862 ( .A(n19833), .ZN(n19835) );
  OAI22_X1 U22863 ( .A1(n19837), .A2(n19836), .B1(n19835), .B2(n19834), .ZN(
        n19838) );
  INV_X1 U22864 ( .A(n19838), .ZN(n19839) );
  OAI21_X1 U22865 ( .B1(n19840), .B2(n19850), .A(n19839), .ZN(P2_U2908) );
  NOR2_X1 U22866 ( .A1(n19842), .A2(n19841), .ZN(P2_U2920) );
  AOI22_X1 U22867 ( .A1(n19860), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19843) );
  OAI21_X1 U22868 ( .B1(n14048), .B2(n19862), .A(n19843), .ZN(P2_U2936) );
  AOI22_X1 U22869 ( .A1(n19860), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19844) );
  OAI21_X1 U22870 ( .B1(n19845), .B2(n19862), .A(n19844), .ZN(P2_U2937) );
  AOI22_X1 U22871 ( .A1(n19860), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19846) );
  OAI21_X1 U22872 ( .B1(n19847), .B2(n19862), .A(n19846), .ZN(P2_U2938) );
  AOI22_X1 U22873 ( .A1(n19860), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19848) );
  OAI21_X1 U22874 ( .B1(n14141), .B2(n19862), .A(n19848), .ZN(P2_U2939) );
  AOI22_X1 U22875 ( .A1(n19860), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19849) );
  OAI21_X1 U22876 ( .B1(n19850), .B2(n19862), .A(n19849), .ZN(P2_U2940) );
  AOI22_X1 U22877 ( .A1(n19860), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19851) );
  OAI21_X1 U22878 ( .B1(n14136), .B2(n19862), .A(n19851), .ZN(P2_U2941) );
  AOI22_X1 U22879 ( .A1(n19860), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19852) );
  OAI21_X1 U22880 ( .B1(n14131), .B2(n19862), .A(n19852), .ZN(P2_U2942) );
  AOI22_X1 U22881 ( .A1(n19860), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n19853) );
  OAI21_X1 U22882 ( .B1(n14128), .B2(n19862), .A(n19853), .ZN(P2_U2943) );
  AOI22_X1 U22883 ( .A1(n19860), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19854) );
  OAI21_X1 U22884 ( .B1(n14276), .B2(n19862), .A(n19854), .ZN(P2_U2944) );
  AOI22_X1 U22885 ( .A1(n19860), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19855) );
  OAI21_X1 U22886 ( .B1(n14290), .B2(n19862), .A(n19855), .ZN(P2_U2945) );
  AOI22_X1 U22887 ( .A1(n19860), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19856) );
  OAI21_X1 U22888 ( .B1(n14117), .B2(n19862), .A(n19856), .ZN(P2_U2947) );
  AOI22_X1 U22889 ( .A1(n19860), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n19857) );
  OAI21_X1 U22890 ( .B1(n19858), .B2(n19862), .A(n19857), .ZN(P2_U2948) );
  AOI22_X1 U22891 ( .A1(n19860), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n19859), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n19861) );
  OAI21_X1 U22892 ( .B1(n14112), .B2(n19862), .A(n19861), .ZN(P2_U2949) );
  AOI22_X2 U22893 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19894), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19895), .ZN(n20408) );
  INV_X1 U22894 ( .A(n20408), .ZN(n20238) );
  AOI22_X1 U22895 ( .A1(n21746), .A2(n20238), .B1(n19892), .B2(n9869), .ZN(
        n19867) );
  NOR2_X2 U22896 ( .A1(n19930), .A2(n19863), .ZN(n20395) );
  OAI22_X2 U22897 ( .A1(n19865), .A2(n19889), .B1(n19864), .B2(n19888), .ZN(
        n20405) );
  AOI22_X1 U22898 ( .A1(n20395), .A2(n19897), .B1(n19896), .B2(n20405), .ZN(
        n19866) );
  OAI211_X1 U22899 ( .C1(n19900), .C2(n19868), .A(n19867), .B(n19866), .ZN(
        P2_U3048) );
  AOI22_X1 U22900 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19894), .ZN(n20414) );
  INV_X1 U22901 ( .A(n20414), .ZN(n20313) );
  OR2_X1 U22902 ( .A1(n19891), .A2(n19869), .ZN(n20357) );
  AOI22_X1 U22903 ( .A1(n21746), .A2(n20313), .B1(n19892), .B2(n20409), .ZN(
        n19873) );
  INV_X1 U22904 ( .A(n19870), .ZN(n19871) );
  NOR2_X2 U22905 ( .A1(n19930), .A2(n19871), .ZN(n20410) );
  AOI22_X1 U22906 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19894), .ZN(n20361) );
  INV_X1 U22907 ( .A(n20361), .ZN(n20411) );
  AOI22_X1 U22908 ( .A1(n20410), .A2(n19897), .B1(n19896), .B2(n20411), .ZN(
        n19872) );
  OAI211_X1 U22909 ( .C1(n19900), .C2(n19874), .A(n19873), .B(n19872), .ZN(
        P2_U3050) );
  AOI22_X2 U22910 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19894), .ZN(n20426) );
  INV_X1 U22911 ( .A(n20426), .ZN(n20248) );
  OR2_X1 U22912 ( .A1(n19891), .A2(n19875), .ZN(n20367) );
  AOI22_X1 U22913 ( .A1(n21746), .A2(n20248), .B1(n19892), .B2(n20421), .ZN(
        n19878) );
  NOR2_X2 U22914 ( .A1(n19930), .A2(n19876), .ZN(n20422) );
  AOI22_X1 U22915 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19894), .ZN(n20371) );
  AOI22_X1 U22916 ( .A1(n20422), .A2(n19897), .B1(n19896), .B2(n20423), .ZN(
        n19877) );
  OAI211_X1 U22917 ( .C1(n19900), .C2(n14651), .A(n19878), .B(n19877), .ZN(
        P2_U3052) );
  AOI22_X1 U22918 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19894), .ZN(n20432) );
  INV_X1 U22919 ( .A(n20432), .ZN(n20322) );
  AOI22_X1 U22920 ( .A1(n21746), .A2(n20322), .B1(n19892), .B2(n20427), .ZN(
        n19883) );
  INV_X1 U22921 ( .A(n19880), .ZN(n19881) );
  NOR2_X2 U22922 ( .A1(n19930), .A2(n19881), .ZN(n20428) );
  AOI22_X1 U22923 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19894), .ZN(n20376) );
  INV_X1 U22924 ( .A(n20376), .ZN(n20429) );
  AOI22_X1 U22925 ( .A1(n20428), .A2(n19897), .B1(n19896), .B2(n20429), .ZN(
        n19882) );
  OAI211_X1 U22926 ( .C1(n19900), .C2(n14732), .A(n19883), .B(n19882), .ZN(
        P2_U3053) );
  AOI22_X1 U22927 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19894), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19895), .ZN(n20438) );
  INV_X1 U22928 ( .A(n20438), .ZN(n20325) );
  OR2_X1 U22929 ( .A1(n19891), .A2(n12213), .ZN(n20144) );
  AOI22_X1 U22930 ( .A1(n21746), .A2(n20325), .B1(n19892), .B2(n20433), .ZN(
        n19887) );
  NOR2_X2 U22931 ( .A1(n19930), .A2(n19884), .ZN(n20434) );
  OAI22_X2 U22932 ( .A1(n19885), .A2(n19889), .B1(n21624), .B2(n19888), .ZN(
        n20435) );
  AOI22_X1 U22933 ( .A1(n20434), .A2(n19897), .B1(n19896), .B2(n20435), .ZN(
        n19886) );
  OAI211_X1 U22934 ( .C1(n19900), .C2(n21603), .A(n19887), .B(n19886), .ZN(
        P2_U3054) );
  OR2_X1 U22935 ( .A1(n19891), .A2(n9691), .ZN(n20381) );
  AOI22_X1 U22936 ( .A1(n21746), .A2(n20331), .B1(n19892), .B2(n20439), .ZN(
        n19899) );
  NOR2_X2 U22937 ( .A1(n19930), .A2(n19893), .ZN(n20440) );
  AOI22_X1 U22938 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19895), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19894), .ZN(n20383) );
  INV_X1 U22939 ( .A(n20383), .ZN(n20441) );
  AOI22_X1 U22940 ( .A1(n20440), .A2(n19897), .B1(n19896), .B2(n20441), .ZN(
        n19898) );
  OAI211_X1 U22941 ( .C1(n19900), .C2(n21653), .A(n19899), .B(n19898), .ZN(
        P2_U3055) );
  OR2_X1 U22942 ( .A1(n20297), .A2(n19960), .ZN(n19905) );
  AND2_X1 U22943 ( .A1(n19905), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19901) );
  NAND2_X1 U22944 ( .A1(n19902), .A2(n19901), .ZN(n19907) );
  INV_X1 U22945 ( .A(n19907), .ZN(n19903) );
  AOI211_X2 U22946 ( .C1(n19904), .C2(n20393), .A(n20298), .B(n19903), .ZN(
        n19925) );
  INV_X1 U22947 ( .A(n19905), .ZN(n19924) );
  AOI22_X1 U22948 ( .A1(n19925), .A2(n20395), .B1(n9869), .B2(n19924), .ZN(
        n19911) );
  NAND2_X1 U22949 ( .A1(n20155), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20090) );
  OAI21_X1 U22950 ( .B1(n20090), .B2(n19909), .A(n19904), .ZN(n19908) );
  NAND2_X1 U22951 ( .A1(n19905), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19906) );
  NAND4_X1 U22952 ( .A1(n19908), .A2(n20403), .A3(n19907), .A4(n19906), .ZN(
        n19926) );
  AOI22_X1 U22953 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20405), .ZN(n19910) );
  OAI211_X1 U22954 ( .C1(n20408), .C2(n19929), .A(n19911), .B(n19910), .ZN(
        P2_U3056) );
  AOI22_X1 U22955 ( .A1(n19925), .A2(n21743), .B1(n21741), .B2(n19924), .ZN(
        n19913) );
  INV_X1 U22956 ( .A(n20356), .ZN(n21745) );
  AOI22_X1 U22957 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n21745), .ZN(n19912) );
  OAI211_X1 U22958 ( .C1(n21751), .C2(n19929), .A(n19913), .B(n19912), .ZN(
        P2_U3057) );
  AOI22_X1 U22959 ( .A1(n19925), .A2(n20410), .B1(n20409), .B2(n19924), .ZN(
        n19915) );
  AOI22_X1 U22960 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20411), .ZN(n19914) );
  OAI211_X1 U22961 ( .C1(n20414), .C2(n19929), .A(n19915), .B(n19914), .ZN(
        P2_U3058) );
  AOI22_X1 U22962 ( .A1(n19925), .A2(n20416), .B1(n20415), .B2(n19924), .ZN(
        n19917) );
  AOI22_X1 U22963 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20417), .ZN(n19916) );
  OAI211_X1 U22964 ( .C1(n20420), .C2(n19929), .A(n19917), .B(n19916), .ZN(
        P2_U3059) );
  AOI22_X1 U22965 ( .A1(n19925), .A2(n20422), .B1(n20421), .B2(n19924), .ZN(
        n19919) );
  AOI22_X1 U22966 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20423), .ZN(n19918) );
  OAI211_X1 U22967 ( .C1(n20426), .C2(n19929), .A(n19919), .B(n19918), .ZN(
        P2_U3060) );
  AOI22_X1 U22968 ( .A1(n19925), .A2(n20428), .B1(n20427), .B2(n19924), .ZN(
        n19921) );
  AOI22_X1 U22969 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20429), .ZN(n19920) );
  OAI211_X1 U22970 ( .C1(n20432), .C2(n19929), .A(n19921), .B(n19920), .ZN(
        P2_U3061) );
  AOI22_X1 U22971 ( .A1(n19925), .A2(n20434), .B1(n20433), .B2(n19924), .ZN(
        n19923) );
  AOI22_X1 U22972 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20435), .ZN(n19922) );
  OAI211_X1 U22973 ( .C1(n20438), .C2(n19929), .A(n19923), .B(n19922), .ZN(
        P2_U3062) );
  AOI22_X1 U22974 ( .A1(n19925), .A2(n20440), .B1(n20439), .B2(n19924), .ZN(
        n19928) );
  AOI22_X1 U22975 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19926), .B1(
        n19956), .B2(n20441), .ZN(n19927) );
  OAI211_X1 U22976 ( .C1(n20444), .C2(n19929), .A(n19928), .B(n19927), .ZN(
        P2_U3063) );
  NOR2_X1 U22977 ( .A1(n20197), .A2(n19960), .ZN(n19934) );
  AOI221_X1 U22978 ( .B1(n19989), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19956), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19934), .ZN(n19932) );
  INV_X1 U22979 ( .A(n11283), .ZN(n19933) );
  NOR2_X1 U22980 ( .A1(n20195), .A2(n19960), .ZN(n19954) );
  AOI211_X1 U22981 ( .C1(n19933), .C2(n20300), .A(n20528), .B(n19954), .ZN(
        n19931) );
  INV_X1 U22982 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n19939) );
  OAI21_X1 U22983 ( .B1(n19933), .B2(n19954), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19936) );
  INV_X1 U22984 ( .A(n19934), .ZN(n19935) );
  NAND2_X1 U22985 ( .A1(n19936), .A2(n19935), .ZN(n19955) );
  AOI22_X1 U22986 ( .A1(n19955), .A2(n20395), .B1(n19954), .B2(n9869), .ZN(
        n19938) );
  AOI22_X1 U22987 ( .A1(n19989), .A2(n20405), .B1(n19956), .B2(n20238), .ZN(
        n19937) );
  OAI211_X1 U22988 ( .C1(n19959), .C2(n19939), .A(n19938), .B(n19937), .ZN(
        P2_U3064) );
  AOI22_X1 U22989 ( .A1(n19955), .A2(n21743), .B1(n19954), .B2(n21741), .ZN(
        n19941) );
  AOI22_X1 U22990 ( .A1(n19956), .A2(n20310), .B1(n19989), .B2(n21745), .ZN(
        n19940) );
  OAI211_X1 U22991 ( .C1(n19959), .C2(n11196), .A(n19941), .B(n19940), .ZN(
        P2_U3065) );
  INV_X1 U22992 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19944) );
  AOI22_X1 U22993 ( .A1(n19955), .A2(n20410), .B1(n19954), .B2(n20409), .ZN(
        n19943) );
  AOI22_X1 U22994 ( .A1(n19989), .A2(n20411), .B1(n19956), .B2(n20313), .ZN(
        n19942) );
  OAI211_X1 U22995 ( .C1(n19959), .C2(n19944), .A(n19943), .B(n19942), .ZN(
        P2_U3066) );
  AOI22_X1 U22996 ( .A1(n19955), .A2(n20416), .B1(n19954), .B2(n20415), .ZN(
        n19946) );
  AOI22_X1 U22997 ( .A1(n19989), .A2(n20417), .B1(n19956), .B2(n20316), .ZN(
        n19945) );
  OAI211_X1 U22998 ( .C1(n19959), .C2(n11171), .A(n19946), .B(n19945), .ZN(
        P2_U3067) );
  INV_X1 U22999 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U23000 ( .A1(n19955), .A2(n20422), .B1(n19954), .B2(n20421), .ZN(
        n19948) );
  AOI22_X1 U23001 ( .A1(n19989), .A2(n20423), .B1(n19956), .B2(n20248), .ZN(
        n19947) );
  OAI211_X1 U23002 ( .C1(n19959), .C2(n19949), .A(n19948), .B(n19947), .ZN(
        P2_U3068) );
  AOI22_X1 U23003 ( .A1(n19955), .A2(n20428), .B1(n19954), .B2(n20427), .ZN(
        n19951) );
  AOI22_X1 U23004 ( .A1(n19989), .A2(n20429), .B1(n19956), .B2(n20322), .ZN(
        n19950) );
  OAI211_X1 U23005 ( .C1(n19959), .C2(n11285), .A(n19951), .B(n19950), .ZN(
        P2_U3069) );
  AOI22_X1 U23006 ( .A1(n19955), .A2(n20434), .B1(n19954), .B2(n20433), .ZN(
        n19953) );
  AOI22_X1 U23007 ( .A1(n19956), .A2(n20325), .B1(n19989), .B2(n20435), .ZN(
        n19952) );
  OAI211_X1 U23008 ( .C1(n19959), .C2(n11320), .A(n19953), .B(n19952), .ZN(
        P2_U3070) );
  AOI22_X1 U23009 ( .A1(n19955), .A2(n20440), .B1(n19954), .B2(n20439), .ZN(
        n19958) );
  AOI22_X1 U23010 ( .A1(n19989), .A2(n20441), .B1(n19956), .B2(n20331), .ZN(
        n19957) );
  OAI211_X1 U23011 ( .C1(n19959), .C2(n11361), .A(n19958), .B(n19957), .ZN(
        P2_U3071) );
  NOR2_X1 U23012 ( .A1(n20227), .A2(n19960), .ZN(n19988) );
  AOI22_X1 U23013 ( .A1(n20405), .A2(n20019), .B1(n19988), .B2(n9869), .ZN(
        n19971) );
  OAI21_X1 U23014 ( .B1(n20090), .B2(n19961), .A(n20528), .ZN(n19969) );
  AND2_X1 U23015 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19962), .ZN(
        n19964) );
  INV_X1 U23016 ( .A(n19988), .ZN(n19979) );
  OAI211_X1 U23017 ( .C1(n19965), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20343), 
        .B(n19979), .ZN(n19963) );
  OAI211_X1 U23018 ( .C1(n19969), .C2(n19964), .A(n20403), .B(n19963), .ZN(
        n19991) );
  INV_X1 U23019 ( .A(n19964), .ZN(n19968) );
  INV_X1 U23020 ( .A(n19965), .ZN(n19966) );
  OAI21_X1 U23021 ( .B1(n19966), .B2(n19988), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19967) );
  AOI22_X1 U23022 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19991), .B1(
        n20395), .B2(n19990), .ZN(n19970) );
  OAI211_X1 U23023 ( .C1(n20408), .C2(n19987), .A(n19971), .B(n19970), .ZN(
        P2_U3072) );
  AOI22_X1 U23024 ( .A1(n19989), .A2(n20310), .B1(n19988), .B2(n21741), .ZN(
        n19973) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19991), .B1(
        n21743), .B2(n19990), .ZN(n19972) );
  OAI211_X1 U23026 ( .C1(n20356), .C2(n20010), .A(n19973), .B(n19972), .ZN(
        P2_U3073) );
  AOI22_X1 U23027 ( .A1(n19989), .A2(n20313), .B1(n19988), .B2(n20409), .ZN(
        n19975) );
  AOI22_X1 U23028 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19991), .B1(
        n20410), .B2(n19990), .ZN(n19974) );
  OAI211_X1 U23029 ( .C1(n20361), .C2(n20010), .A(n19975), .B(n19974), .ZN(
        P2_U3074) );
  NOR2_X1 U23030 ( .A1(n20362), .A2(n19979), .ZN(n19976) );
  AOI21_X1 U23031 ( .B1(n20019), .B2(n20417), .A(n19976), .ZN(n19978) );
  AOI22_X1 U23032 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19991), .B1(
        n20416), .B2(n19990), .ZN(n19977) );
  OAI211_X1 U23033 ( .C1(n20420), .C2(n19987), .A(n19978), .B(n19977), .ZN(
        P2_U3075) );
  NOR2_X1 U23034 ( .A1(n20367), .A2(n19979), .ZN(n19980) );
  AOI21_X1 U23035 ( .B1(n20019), .B2(n20423), .A(n19980), .ZN(n19982) );
  AOI22_X1 U23036 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19991), .B1(
        n20422), .B2(n19990), .ZN(n19981) );
  OAI211_X1 U23037 ( .C1(n20426), .C2(n19987), .A(n19982), .B(n19981), .ZN(
        P2_U3076) );
  AOI22_X1 U23038 ( .A1(n20019), .A2(n20429), .B1(n19988), .B2(n20427), .ZN(
        n19984) );
  AOI22_X1 U23039 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19991), .B1(
        n20428), .B2(n19990), .ZN(n19983) );
  OAI211_X1 U23040 ( .C1(n20432), .C2(n19987), .A(n19984), .B(n19983), .ZN(
        P2_U3077) );
  AOI22_X1 U23041 ( .A1(n20435), .A2(n20019), .B1(n19988), .B2(n20433), .ZN(
        n19986) );
  AOI22_X1 U23042 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19991), .B1(
        n20434), .B2(n19990), .ZN(n19985) );
  OAI211_X1 U23043 ( .C1(n20438), .C2(n19987), .A(n19986), .B(n19985), .ZN(
        P2_U3078) );
  AOI22_X1 U23044 ( .A1(n20331), .A2(n19989), .B1(n19988), .B2(n20439), .ZN(
        n19993) );
  AOI22_X1 U23045 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19991), .B1(
        n20440), .B2(n19990), .ZN(n19992) );
  OAI211_X1 U23046 ( .C1(n20383), .C2(n20010), .A(n19993), .B(n19992), .ZN(
        P2_U3079) );
  INV_X1 U23047 ( .A(n20342), .ZN(n20265) );
  NAND2_X1 U23048 ( .A1(n20265), .A2(n19994), .ZN(n20273) );
  OR2_X1 U23049 ( .A1(n20273), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19999) );
  INV_X1 U23050 ( .A(n19997), .ZN(n19995) );
  NAND2_X1 U23051 ( .A1(n20533), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20085) );
  NOR2_X1 U23052 ( .A1(n20085), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20026) );
  INV_X1 U23053 ( .A(n20026), .ZN(n20029) );
  NOR2_X1 U23054 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20029), .ZN(
        n20017) );
  OAI21_X1 U23055 ( .B1(n19995), .B2(n20017), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19996) );
  AOI22_X1 U23056 ( .A1(n20018), .A2(n20395), .B1(n9869), .B2(n20017), .ZN(
        n20003) );
  AOI21_X1 U23057 ( .B1(n19997), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20001) );
  OAI221_X1 U23058 ( .B1(n20198), .B2(n20010), .C1(n20198), .C2(n20049), .A(
        n19999), .ZN(n20000) );
  OAI211_X1 U23059 ( .C1(n20001), .C2(n20017), .A(n20403), .B(n20000), .ZN(
        n20020) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20020), .B1(
        n20051), .B2(n20405), .ZN(n20002) );
  OAI211_X1 U23061 ( .C1(n20408), .C2(n20010), .A(n20003), .B(n20002), .ZN(
        P2_U3080) );
  AOI22_X1 U23062 ( .A1(n20018), .A2(n21743), .B1(n21741), .B2(n20017), .ZN(
        n20005) );
  AOI22_X1 U23063 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20020), .B1(
        n20019), .B2(n20310), .ZN(n20004) );
  OAI211_X1 U23064 ( .C1(n20356), .C2(n20049), .A(n20005), .B(n20004), .ZN(
        P2_U3081) );
  AOI22_X1 U23065 ( .A1(n20018), .A2(n20410), .B1(n20409), .B2(n20017), .ZN(
        n20007) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20020), .B1(
        n20051), .B2(n20411), .ZN(n20006) );
  OAI211_X1 U23067 ( .C1(n20414), .C2(n20010), .A(n20007), .B(n20006), .ZN(
        P2_U3082) );
  AOI22_X1 U23068 ( .A1(n20018), .A2(n20416), .B1(n20415), .B2(n20017), .ZN(
        n20009) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20020), .B1(
        n20051), .B2(n20417), .ZN(n20008) );
  OAI211_X1 U23070 ( .C1(n20420), .C2(n20010), .A(n20009), .B(n20008), .ZN(
        P2_U3083) );
  AOI22_X1 U23071 ( .A1(n20018), .A2(n20422), .B1(n20421), .B2(n20017), .ZN(
        n20012) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20020), .B1(
        n20019), .B2(n20248), .ZN(n20011) );
  OAI211_X1 U23073 ( .C1(n20371), .C2(n20049), .A(n20012), .B(n20011), .ZN(
        P2_U3084) );
  AOI22_X1 U23074 ( .A1(n20018), .A2(n20428), .B1(n20427), .B2(n20017), .ZN(
        n20014) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20020), .B1(
        n20019), .B2(n20322), .ZN(n20013) );
  OAI211_X1 U23076 ( .C1(n20376), .C2(n20049), .A(n20014), .B(n20013), .ZN(
        P2_U3085) );
  AOI22_X1 U23077 ( .A1(n20018), .A2(n20434), .B1(n20433), .B2(n20017), .ZN(
        n20016) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20020), .B1(
        n20019), .B2(n20325), .ZN(n20015) );
  OAI211_X1 U23079 ( .C1(n20328), .C2(n20049), .A(n20016), .B(n20015), .ZN(
        P2_U3086) );
  AOI22_X1 U23080 ( .A1(n20018), .A2(n20440), .B1(n20439), .B2(n20017), .ZN(
        n20022) );
  AOI22_X1 U23081 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20020), .B1(
        n20019), .B2(n20331), .ZN(n20021) );
  OAI211_X1 U23082 ( .C1(n20383), .C2(n20049), .A(n20022), .B(n20021), .ZN(
        P2_U3087) );
  OR2_X1 U23083 ( .A1(n20297), .A2(n20085), .ZN(n20061) );
  INV_X1 U23084 ( .A(n20061), .ZN(n20050) );
  AOI22_X1 U23085 ( .A1(n20405), .A2(n20081), .B1(n20050), .B2(n9869), .ZN(
        n20032) );
  OAI21_X1 U23086 ( .B1(n20269), .B2(n20090), .A(n20528), .ZN(n20030) );
  OAI211_X1 U23087 ( .C1(n20024), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20343), 
        .B(n20061), .ZN(n20025) );
  OAI211_X1 U23088 ( .C1(n20030), .C2(n20026), .A(n20403), .B(n20025), .ZN(
        n20053) );
  OAI21_X1 U23089 ( .B1(n20027), .B2(n20050), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20028) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20053), .B1(
        n20395), .B2(n20052), .ZN(n20031) );
  OAI211_X1 U23091 ( .C1(n20408), .C2(n20049), .A(n20032), .B(n20031), .ZN(
        P2_U3088) );
  OAI22_X1 U23092 ( .A1(n20074), .A2(n20356), .B1(n20061), .B2(n20352), .ZN(
        n20033) );
  INV_X1 U23093 ( .A(n20033), .ZN(n20035) );
  AOI22_X1 U23094 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20053), .B1(
        n21743), .B2(n20052), .ZN(n20034) );
  OAI211_X1 U23095 ( .C1(n21751), .C2(n20049), .A(n20035), .B(n20034), .ZN(
        P2_U3089) );
  AOI22_X1 U23096 ( .A1(n20051), .A2(n20313), .B1(n20050), .B2(n20409), .ZN(
        n20037) );
  AOI22_X1 U23097 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20053), .B1(
        n20410), .B2(n20052), .ZN(n20036) );
  OAI211_X1 U23098 ( .C1(n20361), .C2(n20074), .A(n20037), .B(n20036), .ZN(
        P2_U3090) );
  OAI22_X1 U23099 ( .A1(n20074), .A2(n20363), .B1(n20061), .B2(n20362), .ZN(
        n20038) );
  INV_X1 U23100 ( .A(n20038), .ZN(n20040) );
  AOI22_X1 U23101 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20053), .B1(
        n20416), .B2(n20052), .ZN(n20039) );
  OAI211_X1 U23102 ( .C1(n20420), .C2(n20049), .A(n20040), .B(n20039), .ZN(
        P2_U3091) );
  OAI22_X1 U23103 ( .A1(n20074), .A2(n20371), .B1(n20061), .B2(n20367), .ZN(
        n20041) );
  INV_X1 U23104 ( .A(n20041), .ZN(n20043) );
  AOI22_X1 U23105 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20053), .B1(
        n20422), .B2(n20052), .ZN(n20042) );
  OAI211_X1 U23106 ( .C1(n20426), .C2(n20049), .A(n20043), .B(n20042), .ZN(
        P2_U3092) );
  OAI22_X1 U23107 ( .A1(n20074), .A2(n20376), .B1(n20061), .B2(n20372), .ZN(
        n20044) );
  INV_X1 U23108 ( .A(n20044), .ZN(n20046) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20053), .B1(
        n20428), .B2(n20052), .ZN(n20045) );
  OAI211_X1 U23110 ( .C1(n20432), .C2(n20049), .A(n20046), .B(n20045), .ZN(
        P2_U3093) );
  AOI22_X1 U23111 ( .A1(n20435), .A2(n20081), .B1(n20050), .B2(n20433), .ZN(
        n20048) );
  AOI22_X1 U23112 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20053), .B1(
        n20434), .B2(n20052), .ZN(n20047) );
  OAI211_X1 U23113 ( .C1(n20438), .C2(n20049), .A(n20048), .B(n20047), .ZN(
        P2_U3094) );
  AOI22_X1 U23114 ( .A1(n20331), .A2(n20051), .B1(n20050), .B2(n20439), .ZN(
        n20055) );
  AOI22_X1 U23115 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20053), .B1(
        n20440), .B2(n20052), .ZN(n20054) );
  OAI211_X1 U23116 ( .C1(n20383), .C2(n20074), .A(n20055), .B(n20054), .ZN(
        P2_U3095) );
  NOR2_X1 U23117 ( .A1(n20195), .A2(n20085), .ZN(n20079) );
  OAI21_X1 U23118 ( .B1(n20059), .B2(n20079), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20056) );
  OAI21_X1 U23119 ( .B1(n20085), .B2(n20197), .A(n20056), .ZN(n20080) );
  AOI22_X1 U23120 ( .A1(n20080), .A2(n20395), .B1(n20079), .B2(n9869), .ZN(
        n20065) );
  INV_X1 U23121 ( .A(n20057), .ZN(n20058) );
  OAI21_X1 U23122 ( .B1(n20081), .B2(n20108), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20062) );
  OAI21_X1 U23123 ( .B1(n20059), .B2(n20393), .A(n20300), .ZN(n20060) );
  AOI21_X1 U23124 ( .B1(n20062), .B2(n20061), .A(n20060), .ZN(n20063) );
  AOI22_X1 U23125 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20082), .B1(
        n20108), .B2(n20405), .ZN(n20064) );
  OAI211_X1 U23126 ( .C1(n20408), .C2(n20074), .A(n20065), .B(n20064), .ZN(
        P2_U3096) );
  AOI22_X1 U23127 ( .A1(n20080), .A2(n21743), .B1(n21741), .B2(n20079), .ZN(
        n20067) );
  AOI22_X1 U23128 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20082), .B1(
        n20108), .B2(n21745), .ZN(n20066) );
  OAI211_X1 U23129 ( .C1(n21751), .C2(n20074), .A(n20067), .B(n20066), .ZN(
        P2_U3097) );
  AOI22_X1 U23130 ( .A1(n20080), .A2(n20410), .B1(n20079), .B2(n20409), .ZN(
        n20069) );
  AOI22_X1 U23131 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20082), .B1(
        n20108), .B2(n20411), .ZN(n20068) );
  OAI211_X1 U23132 ( .C1(n20414), .C2(n20074), .A(n20069), .B(n20068), .ZN(
        P2_U3098) );
  AOI22_X1 U23133 ( .A1(n20080), .A2(n20416), .B1(n20415), .B2(n20079), .ZN(
        n20071) );
  AOI22_X1 U23134 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20082), .B1(
        n20108), .B2(n20417), .ZN(n20070) );
  OAI211_X1 U23135 ( .C1(n20420), .C2(n20074), .A(n20071), .B(n20070), .ZN(
        P2_U3099) );
  AOI22_X1 U23136 ( .A1(n20080), .A2(n20422), .B1(n20079), .B2(n20421), .ZN(
        n20073) );
  AOI22_X1 U23137 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20082), .B1(
        n20108), .B2(n20423), .ZN(n20072) );
  OAI211_X1 U23138 ( .C1(n20426), .C2(n20074), .A(n20073), .B(n20072), .ZN(
        P2_U3100) );
  AOI22_X1 U23139 ( .A1(n20080), .A2(n20428), .B1(n20079), .B2(n20427), .ZN(
        n20076) );
  AOI22_X1 U23140 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20322), .ZN(n20075) );
  OAI211_X1 U23141 ( .C1(n20376), .C2(n20115), .A(n20076), .B(n20075), .ZN(
        P2_U3101) );
  AOI22_X1 U23142 ( .A1(n20080), .A2(n20434), .B1(n20079), .B2(n20433), .ZN(
        n20078) );
  AOI22_X1 U23143 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20325), .ZN(n20077) );
  OAI211_X1 U23144 ( .C1(n20328), .C2(n20115), .A(n20078), .B(n20077), .ZN(
        P2_U3102) );
  AOI22_X1 U23145 ( .A1(n20080), .A2(n20440), .B1(n20079), .B2(n20439), .ZN(
        n20084) );
  AOI22_X1 U23146 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20331), .ZN(n20083) );
  OAI211_X1 U23147 ( .C1(n20383), .C2(n20115), .A(n20084), .B(n20083), .ZN(
        P2_U3103) );
  INV_X1 U23148 ( .A(n20085), .ZN(n20091) );
  NAND3_X1 U23149 ( .A1(n20300), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n20091), .ZN(n20089) );
  NOR2_X1 U23150 ( .A1(n20227), .A2(n20085), .ZN(n20121) );
  NOR2_X1 U23151 ( .A1(n20121), .A2(n20393), .ZN(n20086) );
  NAND2_X1 U23152 ( .A1(n20087), .A2(n20086), .ZN(n20092) );
  INV_X1 U23153 ( .A(n20092), .ZN(n20088) );
  AOI22_X1 U23154 ( .A1(n20111), .A2(n20395), .B1(n20121), .B2(n9869), .ZN(
        n20097) );
  NOR2_X1 U23155 ( .A1(n20090), .A2(n20398), .ZN(n20527) );
  AOI21_X1 U23156 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20091), .A(
        n20527), .ZN(n20094) );
  OAI211_X1 U23157 ( .C1(n20121), .C2(n20300), .A(n20092), .B(n20403), .ZN(
        n20093) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20112), .B1(
        n20117), .B2(n20405), .ZN(n20096) );
  OAI211_X1 U23159 ( .C1(n20408), .C2(n20115), .A(n20097), .B(n20096), .ZN(
        P2_U3104) );
  AOI22_X1 U23160 ( .A1(n20111), .A2(n21743), .B1(n21741), .B2(n20121), .ZN(
        n20099) );
  AOI22_X1 U23161 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20112), .B1(
        n20117), .B2(n21745), .ZN(n20098) );
  OAI211_X1 U23162 ( .C1(n21751), .C2(n20115), .A(n20099), .B(n20098), .ZN(
        P2_U3105) );
  AOI22_X1 U23163 ( .A1(n20111), .A2(n20410), .B1(n20121), .B2(n20409), .ZN(
        n20101) );
  AOI22_X1 U23164 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20112), .B1(
        n20108), .B2(n20313), .ZN(n20100) );
  OAI211_X1 U23165 ( .C1(n20361), .C2(n20154), .A(n20101), .B(n20100), .ZN(
        P2_U3106) );
  AOI22_X1 U23166 ( .A1(n20111), .A2(n20416), .B1(n20415), .B2(n20121), .ZN(
        n20103) );
  AOI22_X1 U23167 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20112), .B1(
        n20108), .B2(n20316), .ZN(n20102) );
  OAI211_X1 U23168 ( .C1(n20363), .C2(n20154), .A(n20103), .B(n20102), .ZN(
        P2_U3107) );
  AOI22_X1 U23169 ( .A1(n20111), .A2(n20422), .B1(n20121), .B2(n20421), .ZN(
        n20105) );
  AOI22_X1 U23170 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20112), .B1(
        n20117), .B2(n20423), .ZN(n20104) );
  OAI211_X1 U23171 ( .C1(n20426), .C2(n20115), .A(n20105), .B(n20104), .ZN(
        P2_U3108) );
  AOI22_X1 U23172 ( .A1(n20111), .A2(n20428), .B1(n20121), .B2(n20427), .ZN(
        n20107) );
  AOI22_X1 U23173 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20112), .B1(
        n20108), .B2(n20322), .ZN(n20106) );
  OAI211_X1 U23174 ( .C1(n20376), .C2(n20154), .A(n20107), .B(n20106), .ZN(
        P2_U3109) );
  AOI22_X1 U23175 ( .A1(n20111), .A2(n20434), .B1(n20121), .B2(n20433), .ZN(
        n20110) );
  AOI22_X1 U23176 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20112), .B1(
        n20108), .B2(n20325), .ZN(n20109) );
  OAI211_X1 U23177 ( .C1(n20328), .C2(n20154), .A(n20110), .B(n20109), .ZN(
        P2_U3110) );
  AOI22_X1 U23178 ( .A1(n20111), .A2(n20440), .B1(n20121), .B2(n20439), .ZN(
        n20114) );
  AOI22_X1 U23179 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20112), .B1(
        n20117), .B2(n20441), .ZN(n20113) );
  OAI211_X1 U23180 ( .C1(n20444), .C2(n20115), .A(n20114), .B(n20113), .ZN(
        P2_U3111) );
  INV_X1 U23181 ( .A(n20194), .ZN(n20166) );
  NAND2_X1 U23182 ( .A1(n20542), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20225) );
  NOR2_X1 U23183 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20225), .ZN(
        n20161) );
  AND2_X1 U23184 ( .A1(n20161), .A2(n20338), .ZN(n20128) );
  AOI22_X1 U23185 ( .A1(n20405), .A2(n20166), .B1(n20128), .B2(n9869), .ZN(
        n20127) );
  OAI21_X1 U23186 ( .B1(n20166), .B2(n20117), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20118) );
  NAND2_X1 U23187 ( .A1(n20118), .A2(n20528), .ZN(n20125) );
  NOR2_X1 U23188 ( .A1(n20125), .A2(n20121), .ZN(n20119) );
  OAI21_X2 U23189 ( .B1(n20120), .B2(n20128), .A(n20403), .ZN(n20151) );
  NOR2_X1 U23190 ( .A1(n20128), .A2(n20121), .ZN(n20124) );
  OAI21_X1 U23191 ( .B1(n20122), .B2(n20128), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20123) );
  AOI22_X1 U23192 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20151), .B1(
        n20395), .B2(n20150), .ZN(n20126) );
  OAI211_X1 U23193 ( .C1(n20408), .C2(n20154), .A(n20127), .B(n20126), .ZN(
        P2_U3112) );
  INV_X1 U23194 ( .A(n20128), .ZN(n20148) );
  OAI22_X1 U23195 ( .A1(n20154), .A2(n21751), .B1(n20148), .B2(n20352), .ZN(
        n20129) );
  INV_X1 U23196 ( .A(n20129), .ZN(n20131) );
  AOI22_X1 U23197 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n21743), .ZN(n20130) );
  OAI211_X1 U23198 ( .C1(n20356), .C2(n20194), .A(n20131), .B(n20130), .ZN(
        P2_U3113) );
  OAI22_X1 U23199 ( .A1(n20194), .A2(n20361), .B1(n20148), .B2(n20357), .ZN(
        n20132) );
  INV_X1 U23200 ( .A(n20132), .ZN(n20134) );
  AOI22_X1 U23201 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n20410), .ZN(n20133) );
  OAI211_X1 U23202 ( .C1(n20414), .C2(n20154), .A(n20134), .B(n20133), .ZN(
        P2_U3114) );
  OAI22_X1 U23203 ( .A1(n20194), .A2(n20363), .B1(n20148), .B2(n20362), .ZN(
        n20135) );
  INV_X1 U23204 ( .A(n20135), .ZN(n20137) );
  AOI22_X1 U23205 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n20416), .ZN(n20136) );
  OAI211_X1 U23206 ( .C1(n20420), .C2(n20154), .A(n20137), .B(n20136), .ZN(
        P2_U3115) );
  OAI22_X1 U23207 ( .A1(n20194), .A2(n20371), .B1(n20148), .B2(n20367), .ZN(
        n20138) );
  INV_X1 U23208 ( .A(n20138), .ZN(n20140) );
  AOI22_X1 U23209 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n20422), .ZN(n20139) );
  OAI211_X1 U23210 ( .C1(n20426), .C2(n20154), .A(n20140), .B(n20139), .ZN(
        P2_U3116) );
  OAI22_X1 U23211 ( .A1(n20194), .A2(n20376), .B1(n20148), .B2(n20372), .ZN(
        n20141) );
  INV_X1 U23212 ( .A(n20141), .ZN(n20143) );
  AOI22_X1 U23213 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n20428), .ZN(n20142) );
  OAI211_X1 U23214 ( .C1(n20432), .C2(n20154), .A(n20143), .B(n20142), .ZN(
        P2_U3117) );
  OAI22_X1 U23215 ( .A1(n20154), .A2(n20438), .B1(n20148), .B2(n20144), .ZN(
        n20145) );
  INV_X1 U23216 ( .A(n20145), .ZN(n20147) );
  AOI22_X1 U23217 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n20434), .ZN(n20146) );
  OAI211_X1 U23218 ( .C1(n20328), .C2(n20194), .A(n20147), .B(n20146), .ZN(
        P2_U3118) );
  OAI22_X1 U23219 ( .A1(n20194), .A2(n20383), .B1(n20148), .B2(n20381), .ZN(
        n20149) );
  INV_X1 U23220 ( .A(n20149), .ZN(n20153) );
  AOI22_X1 U23221 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20151), .B1(
        n20150), .B2(n20440), .ZN(n20152) );
  OAI211_X1 U23222 ( .C1(n20444), .C2(n20154), .A(n20153), .B(n20152), .ZN(
        P2_U3119) );
  NOR2_X1 U23223 ( .A1(n20155), .A2(n20198), .ZN(n20396) );
  NAND2_X1 U23224 ( .A1(n20396), .A2(n20160), .ZN(n20162) );
  INV_X1 U23225 ( .A(n20161), .ZN(n20156) );
  NAND2_X1 U23226 ( .A1(n20162), .A2(n20156), .ZN(n20159) );
  NOR2_X1 U23227 ( .A1(n20297), .A2(n20225), .ZN(n20199) );
  INV_X1 U23228 ( .A(n20199), .ZN(n20188) );
  AND2_X1 U23229 ( .A1(n20157), .A2(n20403), .ZN(n20158) );
  INV_X1 U23230 ( .A(n20224), .ZN(n20216) );
  AOI22_X1 U23231 ( .A1(n20405), .A2(n20216), .B1(n20199), .B2(n9869), .ZN(
        n20168) );
  NAND3_X1 U23232 ( .A1(n20162), .A2(n20161), .A3(n20528), .ZN(n20165) );
  OAI21_X1 U23233 ( .B1(n20163), .B2(n20199), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20164) );
  AOI22_X1 U23234 ( .A1(n20395), .A2(n20190), .B1(n20166), .B2(n20238), .ZN(
        n20167) );
  OAI211_X1 U23235 ( .C1(n20171), .C2(n20169), .A(n20168), .B(n20167), .ZN(
        P2_U3120) );
  OAI22_X1 U23236 ( .A1(n20194), .A2(n21751), .B1(n20188), .B2(n20352), .ZN(
        n20170) );
  INV_X1 U23237 ( .A(n20170), .ZN(n20173) );
  AOI22_X1 U23238 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20191), .B1(
        n21743), .B2(n20190), .ZN(n20172) );
  OAI211_X1 U23239 ( .C1(n20356), .C2(n20224), .A(n20173), .B(n20172), .ZN(
        P2_U3121) );
  OAI22_X1 U23240 ( .A1(n20224), .A2(n20361), .B1(n20188), .B2(n20357), .ZN(
        n20174) );
  INV_X1 U23241 ( .A(n20174), .ZN(n20176) );
  AOI22_X1 U23242 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20191), .B1(
        n20410), .B2(n20190), .ZN(n20175) );
  OAI211_X1 U23243 ( .C1(n20414), .C2(n20194), .A(n20176), .B(n20175), .ZN(
        P2_U3122) );
  OAI22_X1 U23244 ( .A1(n20194), .A2(n20420), .B1(n20188), .B2(n20362), .ZN(
        n20177) );
  INV_X1 U23245 ( .A(n20177), .ZN(n20179) );
  AOI22_X1 U23246 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20191), .B1(
        n20416), .B2(n20190), .ZN(n20178) );
  OAI211_X1 U23247 ( .C1(n20363), .C2(n20224), .A(n20179), .B(n20178), .ZN(
        P2_U3123) );
  OAI22_X1 U23248 ( .A1(n20194), .A2(n20426), .B1(n20188), .B2(n20367), .ZN(
        n20180) );
  INV_X1 U23249 ( .A(n20180), .ZN(n20182) );
  AOI22_X1 U23250 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20191), .B1(
        n20422), .B2(n20190), .ZN(n20181) );
  OAI211_X1 U23251 ( .C1(n20371), .C2(n20224), .A(n20182), .B(n20181), .ZN(
        P2_U3124) );
  OAI22_X1 U23252 ( .A1(n20224), .A2(n20376), .B1(n20188), .B2(n20372), .ZN(
        n20183) );
  INV_X1 U23253 ( .A(n20183), .ZN(n20185) );
  AOI22_X1 U23254 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20191), .B1(
        n20428), .B2(n20190), .ZN(n20184) );
  OAI211_X1 U23255 ( .C1(n20432), .C2(n20194), .A(n20185), .B(n20184), .ZN(
        P2_U3125) );
  AOI22_X1 U23256 ( .A1(n20435), .A2(n20216), .B1(n20199), .B2(n20433), .ZN(
        n20187) );
  AOI22_X1 U23257 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20191), .B1(
        n20434), .B2(n20190), .ZN(n20186) );
  OAI211_X1 U23258 ( .C1(n20438), .C2(n20194), .A(n20187), .B(n20186), .ZN(
        P2_U3126) );
  OAI22_X1 U23259 ( .A1(n20224), .A2(n20383), .B1(n20188), .B2(n20381), .ZN(
        n20189) );
  INV_X1 U23260 ( .A(n20189), .ZN(n20193) );
  AOI22_X1 U23261 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20191), .B1(
        n20440), .B2(n20190), .ZN(n20192) );
  OAI211_X1 U23262 ( .C1(n20444), .C2(n20194), .A(n20193), .B(n20192), .ZN(
        P2_U3127) );
  NOR2_X1 U23263 ( .A1(n20195), .A2(n20225), .ZN(n20219) );
  OAI21_X1 U23264 ( .B1(n11328), .B2(n20219), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20196) );
  AOI22_X1 U23265 ( .A1(n20220), .A2(n20395), .B1(n20219), .B2(n9869), .ZN(
        n20205) );
  NAND2_X1 U23266 ( .A1(n20337), .A2(n20522), .ZN(n20263) );
  AOI21_X1 U23267 ( .B1(n20224), .B2(n20263), .A(n20198), .ZN(n20200) );
  NOR2_X1 U23268 ( .A1(n20200), .A2(n20199), .ZN(n20201) );
  AOI211_X1 U23269 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20202), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20201), .ZN(n20203) );
  AOI22_X1 U23270 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20221), .B1(
        n20253), .B2(n20405), .ZN(n20204) );
  OAI211_X1 U23271 ( .C1(n20408), .C2(n20224), .A(n20205), .B(n20204), .ZN(
        P2_U3128) );
  AOI22_X1 U23272 ( .A1(n20220), .A2(n21743), .B1(n21741), .B2(n20219), .ZN(
        n20207) );
  AOI22_X1 U23273 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20221), .B1(
        n20216), .B2(n20310), .ZN(n20206) );
  OAI211_X1 U23274 ( .C1(n20356), .C2(n20263), .A(n20207), .B(n20206), .ZN(
        P2_U3129) );
  AOI22_X1 U23275 ( .A1(n20220), .A2(n20410), .B1(n20219), .B2(n20409), .ZN(
        n20209) );
  AOI22_X1 U23276 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20221), .B1(
        n20253), .B2(n20411), .ZN(n20208) );
  OAI211_X1 U23277 ( .C1(n20414), .C2(n20224), .A(n20209), .B(n20208), .ZN(
        P2_U3130) );
  AOI22_X1 U23278 ( .A1(n20220), .A2(n20416), .B1(n20415), .B2(n20219), .ZN(
        n20211) );
  AOI22_X1 U23279 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20221), .B1(
        n20253), .B2(n20417), .ZN(n20210) );
  OAI211_X1 U23280 ( .C1(n20420), .C2(n20224), .A(n20211), .B(n20210), .ZN(
        P2_U3131) );
  AOI22_X1 U23281 ( .A1(n20220), .A2(n20422), .B1(n20219), .B2(n20421), .ZN(
        n20213) );
  AOI22_X1 U23282 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20221), .B1(
        n20253), .B2(n20423), .ZN(n20212) );
  OAI211_X1 U23283 ( .C1(n20426), .C2(n20224), .A(n20213), .B(n20212), .ZN(
        P2_U3132) );
  AOI22_X1 U23284 ( .A1(n20220), .A2(n20428), .B1(n20219), .B2(n20427), .ZN(
        n20215) );
  AOI22_X1 U23285 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20221), .B1(
        n20253), .B2(n20429), .ZN(n20214) );
  OAI211_X1 U23286 ( .C1(n20432), .C2(n20224), .A(n20215), .B(n20214), .ZN(
        P2_U3133) );
  AOI22_X1 U23287 ( .A1(n20220), .A2(n20434), .B1(n20219), .B2(n20433), .ZN(
        n20218) );
  AOI22_X1 U23288 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20221), .B1(
        n20216), .B2(n20325), .ZN(n20217) );
  OAI211_X1 U23289 ( .C1(n20328), .C2(n20263), .A(n20218), .B(n20217), .ZN(
        P2_U3134) );
  AOI22_X1 U23290 ( .A1(n20220), .A2(n20440), .B1(n20219), .B2(n20439), .ZN(
        n20223) );
  AOI22_X1 U23291 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20221), .B1(
        n20253), .B2(n20441), .ZN(n20222) );
  OAI211_X1 U23292 ( .C1(n20444), .C2(n20224), .A(n20223), .B(n20222), .ZN(
        P2_U3135) );
  NAND2_X1 U23293 ( .A1(n20396), .A2(n20522), .ZN(n20226) );
  INV_X1 U23294 ( .A(n20225), .ZN(n20228) );
  NAND2_X1 U23295 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20228), .ZN(
        n20235) );
  NAND2_X1 U23296 ( .A1(n20226), .A2(n20235), .ZN(n20234) );
  INV_X1 U23297 ( .A(n20227), .ZN(n20229) );
  NAND2_X1 U23298 ( .A1(n20229), .A2(n20228), .ZN(n20230) );
  INV_X1 U23299 ( .A(n20230), .ZN(n20258) );
  AND2_X1 U23300 ( .A1(n20230), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20231) );
  OAI211_X1 U23301 ( .C1(n20258), .C2(n20300), .A(n20237), .B(n20403), .ZN(
        n20232) );
  INV_X1 U23302 ( .A(n20232), .ZN(n20233) );
  OAI21_X1 U23303 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20235), .A(n20393), 
        .ZN(n20236) );
  AOI22_X1 U23304 ( .A1(n20259), .A2(n20395), .B1(n9869), .B2(n20258), .ZN(
        n20240) );
  AOI22_X1 U23305 ( .A1(n20271), .A2(n20405), .B1(n20253), .B2(n20238), .ZN(
        n20239) );
  OAI211_X1 U23306 ( .C1(n20252), .C2(n20241), .A(n20240), .B(n20239), .ZN(
        P2_U3136) );
  AOI22_X1 U23307 ( .A1(n20259), .A2(n21743), .B1(n21741), .B2(n20258), .ZN(
        n20243) );
  AOI22_X1 U23308 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20260), .B1(
        n20253), .B2(n20310), .ZN(n20242) );
  OAI211_X1 U23309 ( .C1(n20356), .C2(n20295), .A(n20243), .B(n20242), .ZN(
        P2_U3137) );
  AOI22_X1 U23310 ( .A1(n20259), .A2(n20410), .B1(n20409), .B2(n20258), .ZN(
        n20245) );
  AOI22_X1 U23311 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20260), .B1(
        n20253), .B2(n20313), .ZN(n20244) );
  OAI211_X1 U23312 ( .C1(n20361), .C2(n20295), .A(n20245), .B(n20244), .ZN(
        P2_U3138) );
  AOI22_X1 U23313 ( .A1(n20259), .A2(n20416), .B1(n20415), .B2(n20258), .ZN(
        n20247) );
  AOI22_X1 U23314 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20260), .B1(
        n20271), .B2(n20417), .ZN(n20246) );
  OAI211_X1 U23315 ( .C1(n20420), .C2(n20263), .A(n20247), .B(n20246), .ZN(
        P2_U3139) );
  INV_X1 U23316 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20251) );
  AOI22_X1 U23317 ( .A1(n20259), .A2(n20422), .B1(n20421), .B2(n20258), .ZN(
        n20250) );
  AOI22_X1 U23318 ( .A1(n20271), .A2(n20423), .B1(n20253), .B2(n20248), .ZN(
        n20249) );
  OAI211_X1 U23319 ( .C1(n20252), .C2(n20251), .A(n20250), .B(n20249), .ZN(
        P2_U3140) );
  AOI22_X1 U23320 ( .A1(n20259), .A2(n20428), .B1(n20427), .B2(n20258), .ZN(
        n20255) );
  AOI22_X1 U23321 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20260), .B1(
        n20253), .B2(n20322), .ZN(n20254) );
  OAI211_X1 U23322 ( .C1(n20376), .C2(n20295), .A(n20255), .B(n20254), .ZN(
        P2_U3141) );
  AOI22_X1 U23323 ( .A1(n20259), .A2(n20434), .B1(n20433), .B2(n20258), .ZN(
        n20257) );
  AOI22_X1 U23324 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20260), .B1(
        n20271), .B2(n20435), .ZN(n20256) );
  OAI211_X1 U23325 ( .C1(n20438), .C2(n20263), .A(n20257), .B(n20256), .ZN(
        P2_U3142) );
  AOI22_X1 U23326 ( .A1(n20259), .A2(n20440), .B1(n20439), .B2(n20258), .ZN(
        n20262) );
  AOI22_X1 U23327 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20260), .B1(
        n20271), .B2(n20441), .ZN(n20261) );
  OAI211_X1 U23328 ( .C1(n20444), .C2(n20263), .A(n20262), .B(n20261), .ZN(
        P2_U3143) );
  NOR3_X2 U23329 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20296), .ZN(n20290) );
  OAI21_X1 U23330 ( .B1(n20264), .B2(n20290), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20268) );
  NAND3_X1 U23331 ( .A1(n20266), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20265), .ZN(n20267) );
  NAND2_X1 U23332 ( .A1(n20268), .A2(n20267), .ZN(n20291) );
  AOI22_X1 U23333 ( .A1(n20291), .A2(n20395), .B1(n9869), .B2(n20290), .ZN(
        n20277) );
  INV_X1 U23334 ( .A(n20337), .ZN(n20270) );
  OAI21_X1 U23335 ( .B1(n20332), .B2(n20271), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20272) );
  OAI21_X1 U23336 ( .B1(n20533), .B2(n20273), .A(n20272), .ZN(n20275) );
  NAND3_X1 U23337 ( .A1(n20275), .A2(n20403), .A3(n20274), .ZN(n20292) );
  AOI22_X1 U23338 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20405), .ZN(n20276) );
  OAI211_X1 U23339 ( .C1(n20408), .C2(n20295), .A(n20277), .B(n20276), .ZN(
        P2_U3144) );
  AOI22_X1 U23340 ( .A1(n20291), .A2(n21743), .B1(n21741), .B2(n20290), .ZN(
        n20279) );
  AOI22_X1 U23341 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n21745), .ZN(n20278) );
  OAI211_X1 U23342 ( .C1(n21751), .C2(n20295), .A(n20279), .B(n20278), .ZN(
        P2_U3145) );
  AOI22_X1 U23343 ( .A1(n20291), .A2(n20410), .B1(n20409), .B2(n20290), .ZN(
        n20281) );
  AOI22_X1 U23344 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20411), .ZN(n20280) );
  OAI211_X1 U23345 ( .C1(n20414), .C2(n20295), .A(n20281), .B(n20280), .ZN(
        P2_U3146) );
  AOI22_X1 U23346 ( .A1(n20291), .A2(n20416), .B1(n20415), .B2(n20290), .ZN(
        n20283) );
  AOI22_X1 U23347 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20417), .ZN(n20282) );
  OAI211_X1 U23348 ( .C1(n20420), .C2(n20295), .A(n20283), .B(n20282), .ZN(
        P2_U3147) );
  AOI22_X1 U23349 ( .A1(n20291), .A2(n20422), .B1(n20421), .B2(n20290), .ZN(
        n20285) );
  AOI22_X1 U23350 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20423), .ZN(n20284) );
  OAI211_X1 U23351 ( .C1(n20426), .C2(n20295), .A(n20285), .B(n20284), .ZN(
        P2_U3148) );
  AOI22_X1 U23352 ( .A1(n20291), .A2(n20428), .B1(n20427), .B2(n20290), .ZN(
        n20287) );
  AOI22_X1 U23353 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20429), .ZN(n20286) );
  OAI211_X1 U23354 ( .C1(n20432), .C2(n20295), .A(n20287), .B(n20286), .ZN(
        P2_U3149) );
  AOI22_X1 U23355 ( .A1(n20291), .A2(n20434), .B1(n20433), .B2(n20290), .ZN(
        n20289) );
  AOI22_X1 U23356 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20435), .ZN(n20288) );
  OAI211_X1 U23357 ( .C1(n20438), .C2(n20295), .A(n20289), .B(n20288), .ZN(
        P2_U3150) );
  AOI22_X1 U23358 ( .A1(n20291), .A2(n20440), .B1(n20439), .B2(n20290), .ZN(
        n20294) );
  AOI22_X1 U23359 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20292), .B1(
        n20332), .B2(n20441), .ZN(n20293) );
  OAI211_X1 U23360 ( .C1(n20444), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        P2_U3151) );
  INV_X1 U23361 ( .A(n20332), .ZN(n20321) );
  OR2_X1 U23362 ( .A1(n20296), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20302) );
  NOR2_X1 U23363 ( .A1(n20297), .A2(n20296), .ZN(n20329) );
  AOI211_X2 U23364 ( .C1(n20302), .C2(n20393), .A(n20298), .B(n20299), .ZN(
        n20330) );
  AOI22_X1 U23365 ( .A1(n20330), .A2(n20395), .B1(n9869), .B2(n20329), .ZN(
        n20309) );
  INV_X1 U23366 ( .A(n20299), .ZN(n20305) );
  NAND3_X1 U23367 ( .A1(n20306), .A2(n20396), .A3(n20300), .ZN(n20301) );
  OAI21_X1 U23368 ( .B1(n20303), .B2(n20302), .A(n20301), .ZN(n20304) );
  NAND3_X1 U23369 ( .A1(n20305), .A2(n20403), .A3(n20304), .ZN(n20333) );
  AOI22_X1 U23370 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20333), .B1(
        n20339), .B2(n20405), .ZN(n20308) );
  OAI211_X1 U23371 ( .C1(n20408), .C2(n20321), .A(n20309), .B(n20308), .ZN(
        P2_U3152) );
  AOI22_X1 U23372 ( .A1(n20330), .A2(n21743), .B1(n21741), .B2(n20329), .ZN(
        n20312) );
  AOI22_X1 U23373 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20310), .ZN(n20311) );
  OAI211_X1 U23374 ( .C1(n20356), .C2(n20389), .A(n20312), .B(n20311), .ZN(
        P2_U3153) );
  AOI22_X1 U23375 ( .A1(n20330), .A2(n20410), .B1(n20409), .B2(n20329), .ZN(
        n20315) );
  AOI22_X1 U23376 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20313), .ZN(n20314) );
  OAI211_X1 U23377 ( .C1(n20361), .C2(n20389), .A(n20315), .B(n20314), .ZN(
        P2_U3154) );
  AOI22_X1 U23378 ( .A1(n20330), .A2(n20416), .B1(n20415), .B2(n20329), .ZN(
        n20318) );
  AOI22_X1 U23379 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20316), .ZN(n20317) );
  OAI211_X1 U23380 ( .C1(n20363), .C2(n20389), .A(n20318), .B(n20317), .ZN(
        P2_U3155) );
  AOI22_X1 U23381 ( .A1(n20330), .A2(n20422), .B1(n20421), .B2(n20329), .ZN(
        n20320) );
  AOI22_X1 U23382 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20333), .B1(
        n20339), .B2(n20423), .ZN(n20319) );
  OAI211_X1 U23383 ( .C1(n20426), .C2(n20321), .A(n20320), .B(n20319), .ZN(
        P2_U3156) );
  AOI22_X1 U23384 ( .A1(n20330), .A2(n20428), .B1(n20427), .B2(n20329), .ZN(
        n20324) );
  AOI22_X1 U23385 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20322), .ZN(n20323) );
  OAI211_X1 U23386 ( .C1(n20376), .C2(n20389), .A(n20324), .B(n20323), .ZN(
        P2_U3157) );
  AOI22_X1 U23387 ( .A1(n20330), .A2(n20434), .B1(n20433), .B2(n20329), .ZN(
        n20327) );
  AOI22_X1 U23388 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20325), .ZN(n20326) );
  OAI211_X1 U23389 ( .C1(n20328), .C2(n20389), .A(n20327), .B(n20326), .ZN(
        P2_U3158) );
  AOI22_X1 U23390 ( .A1(n20330), .A2(n20440), .B1(n20439), .B2(n20329), .ZN(
        n20335) );
  AOI22_X1 U23391 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20331), .ZN(n20334) );
  OAI211_X1 U23392 ( .C1(n20383), .C2(n20389), .A(n20335), .B(n20334), .ZN(
        P2_U3159) );
  INV_X1 U23393 ( .A(n21750), .ZN(n20378) );
  NAND2_X1 U23394 ( .A1(n20392), .A2(n20338), .ZN(n20382) );
  INV_X1 U23395 ( .A(n20382), .ZN(n20377) );
  AOI22_X1 U23396 ( .A1(n20405), .A2(n20378), .B1(n20377), .B2(n9869), .ZN(
        n20351) );
  OAI21_X1 U23397 ( .B1(n20378), .B2(n20339), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20340) );
  NAND2_X1 U23398 ( .A1(n20340), .A2(n20528), .ZN(n20349) );
  AND2_X1 U23399 ( .A1(n20342), .A2(n20341), .ZN(n20345) );
  OAI211_X1 U23400 ( .C1(n11289), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20343), 
        .B(n20382), .ZN(n20344) );
  OAI211_X1 U23401 ( .C1(n20349), .C2(n20345), .A(n20403), .B(n20344), .ZN(
        n20386) );
  INV_X1 U23402 ( .A(n20345), .ZN(n20348) );
  OAI21_X1 U23403 ( .B1(n20346), .B2(n20377), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20347) );
  AOI22_X1 U23404 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20386), .B1(
        n20395), .B2(n20385), .ZN(n20350) );
  OAI211_X1 U23405 ( .C1(n20408), .C2(n20389), .A(n20351), .B(n20350), .ZN(
        P2_U3160) );
  OAI22_X1 U23406 ( .A1(n20389), .A2(n21751), .B1(n20382), .B2(n20352), .ZN(
        n20353) );
  INV_X1 U23407 ( .A(n20353), .ZN(n20355) );
  AOI22_X1 U23408 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20386), .B1(
        n21743), .B2(n20385), .ZN(n20354) );
  OAI211_X1 U23409 ( .C1(n20356), .C2(n21750), .A(n20355), .B(n20354), .ZN(
        P2_U3161) );
  OAI22_X1 U23410 ( .A1(n20389), .A2(n20414), .B1(n20382), .B2(n20357), .ZN(
        n20358) );
  INV_X1 U23411 ( .A(n20358), .ZN(n20360) );
  AOI22_X1 U23412 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20386), .B1(
        n20410), .B2(n20385), .ZN(n20359) );
  OAI211_X1 U23413 ( .C1(n20361), .C2(n21750), .A(n20360), .B(n20359), .ZN(
        P2_U3162) );
  OAI22_X1 U23414 ( .A1(n21750), .A2(n20363), .B1(n20382), .B2(n20362), .ZN(
        n20364) );
  INV_X1 U23415 ( .A(n20364), .ZN(n20366) );
  AOI22_X1 U23416 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20386), .B1(
        n20416), .B2(n20385), .ZN(n20365) );
  OAI211_X1 U23417 ( .C1(n20420), .C2(n20389), .A(n20366), .B(n20365), .ZN(
        P2_U3163) );
  OAI22_X1 U23418 ( .A1(n20389), .A2(n20426), .B1(n20382), .B2(n20367), .ZN(
        n20368) );
  INV_X1 U23419 ( .A(n20368), .ZN(n20370) );
  AOI22_X1 U23420 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20386), .B1(
        n20422), .B2(n20385), .ZN(n20369) );
  OAI211_X1 U23421 ( .C1(n20371), .C2(n21750), .A(n20370), .B(n20369), .ZN(
        P2_U3164) );
  OAI22_X1 U23422 ( .A1(n20389), .A2(n20432), .B1(n20382), .B2(n20372), .ZN(
        n20373) );
  INV_X1 U23423 ( .A(n20373), .ZN(n20375) );
  AOI22_X1 U23424 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20386), .B1(
        n20428), .B2(n20385), .ZN(n20374) );
  OAI211_X1 U23425 ( .C1(n20376), .C2(n21750), .A(n20375), .B(n20374), .ZN(
        P2_U3165) );
  AOI22_X1 U23426 ( .A1(n20435), .A2(n20378), .B1(n20377), .B2(n20433), .ZN(
        n20380) );
  AOI22_X1 U23427 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20386), .B1(
        n20434), .B2(n20385), .ZN(n20379) );
  OAI211_X1 U23428 ( .C1(n20438), .C2(n20389), .A(n20380), .B(n20379), .ZN(
        P2_U3166) );
  OAI22_X1 U23429 ( .A1(n21750), .A2(n20383), .B1(n20382), .B2(n20381), .ZN(
        n20384) );
  INV_X1 U23430 ( .A(n20384), .ZN(n20388) );
  AOI22_X1 U23431 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20386), .B1(
        n20440), .B2(n20385), .ZN(n20387) );
  OAI211_X1 U23432 ( .C1(n20444), .C2(n20389), .A(n20388), .B(n20387), .ZN(
        P2_U3167) );
  AND2_X1 U23433 ( .A1(n20400), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20390) );
  NAND2_X1 U23434 ( .A1(n20391), .A2(n20390), .ZN(n20402) );
  INV_X1 U23435 ( .A(n20392), .ZN(n20397) );
  OAI21_X1 U23436 ( .B1(n20397), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20393), 
        .ZN(n20394) );
  INV_X1 U23437 ( .A(n20400), .ZN(n21742) );
  AOI22_X1 U23438 ( .A1(n21744), .A2(n20395), .B1(n21742), .B2(n9869), .ZN(
        n20407) );
  INV_X1 U23439 ( .A(n20396), .ZN(n20399) );
  OAI21_X1 U23440 ( .B1(n20399), .B2(n20398), .A(n20397), .ZN(n20404) );
  NAND2_X1 U23441 ( .A1(n20400), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20401) );
  NAND4_X1 U23442 ( .A1(n20404), .A2(n20403), .A3(n20402), .A4(n20401), .ZN(
        n21747) );
  AOI22_X1 U23443 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20405), .ZN(n20406) );
  OAI211_X1 U23444 ( .C1(n20408), .C2(n21750), .A(n20407), .B(n20406), .ZN(
        P2_U3168) );
  AOI22_X1 U23445 ( .A1(n21744), .A2(n20410), .B1(n21742), .B2(n20409), .ZN(
        n20413) );
  AOI22_X1 U23446 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20411), .ZN(n20412) );
  OAI211_X1 U23447 ( .C1(n20414), .C2(n21750), .A(n20413), .B(n20412), .ZN(
        P2_U3170) );
  AOI22_X1 U23448 ( .A1(n21744), .A2(n20416), .B1(n21742), .B2(n20415), .ZN(
        n20419) );
  AOI22_X1 U23449 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20417), .ZN(n20418) );
  OAI211_X1 U23450 ( .C1(n20420), .C2(n21750), .A(n20419), .B(n20418), .ZN(
        P2_U3171) );
  AOI22_X1 U23451 ( .A1(n21744), .A2(n20422), .B1(n21742), .B2(n20421), .ZN(
        n20425) );
  AOI22_X1 U23452 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20423), .ZN(n20424) );
  OAI211_X1 U23453 ( .C1(n20426), .C2(n21750), .A(n20425), .B(n20424), .ZN(
        P2_U3172) );
  AOI22_X1 U23454 ( .A1(n21744), .A2(n20428), .B1(n21742), .B2(n20427), .ZN(
        n20431) );
  AOI22_X1 U23455 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20429), .ZN(n20430) );
  OAI211_X1 U23456 ( .C1(n20432), .C2(n21750), .A(n20431), .B(n20430), .ZN(
        P2_U3173) );
  AOI22_X1 U23457 ( .A1(n21744), .A2(n20434), .B1(n21742), .B2(n20433), .ZN(
        n20437) );
  AOI22_X1 U23458 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20435), .ZN(n20436) );
  OAI211_X1 U23459 ( .C1(n20438), .C2(n21750), .A(n20437), .B(n20436), .ZN(
        P2_U3174) );
  AOI22_X1 U23460 ( .A1(n21744), .A2(n20440), .B1(n21742), .B2(n20439), .ZN(
        n20443) );
  AOI22_X1 U23461 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n20441), .ZN(n20442) );
  OAI211_X1 U23462 ( .C1(n20444), .C2(n21750), .A(n20443), .B(n20442), .ZN(
        P2_U3175) );
  AND2_X1 U23463 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20445), .ZN(
        P2_U3179) );
  AND2_X1 U23464 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20445), .ZN(
        P2_U3180) );
  AND2_X1 U23465 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20445), .ZN(
        P2_U3181) );
  AND2_X1 U23466 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20445), .ZN(
        P2_U3182) );
  AND2_X1 U23467 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20445), .ZN(
        P2_U3183) );
  AND2_X1 U23468 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20445), .ZN(
        P2_U3184) );
  AND2_X1 U23469 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20445), .ZN(
        P2_U3185) );
  AND2_X1 U23470 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20445), .ZN(
        P2_U3186) );
  AND2_X1 U23471 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20445), .ZN(
        P2_U3187) );
  AND2_X1 U23472 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20445), .ZN(
        P2_U3188) );
  AND2_X1 U23473 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20445), .ZN(
        P2_U3189) );
  AND2_X1 U23474 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20445), .ZN(
        P2_U3190) );
  AND2_X1 U23475 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20445), .ZN(
        P2_U3191) );
  AND2_X1 U23476 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20445), .ZN(
        P2_U3192) );
  AND2_X1 U23477 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20445), .ZN(
        P2_U3193) );
  AND2_X1 U23478 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20445), .ZN(
        P2_U3194) );
  AND2_X1 U23479 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20445), .ZN(
        P2_U3195) );
  AND2_X1 U23480 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20445), .ZN(
        P2_U3196) );
  AND2_X1 U23481 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20445), .ZN(
        P2_U3197) );
  AND2_X1 U23482 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20445), .ZN(
        P2_U3198) );
  AND2_X1 U23483 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20445), .ZN(
        P2_U3199) );
  AND2_X1 U23484 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20445), .ZN(
        P2_U3200) );
  AND2_X1 U23485 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20445), .ZN(P2_U3201) );
  AND2_X1 U23486 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20445), .ZN(P2_U3202) );
  AND2_X1 U23487 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20445), .ZN(P2_U3203) );
  AND2_X1 U23488 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20445), .ZN(P2_U3204) );
  AND2_X1 U23489 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20445), .ZN(P2_U3205) );
  AND2_X1 U23490 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20445), .ZN(P2_U3206) );
  AND2_X1 U23491 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20445), .ZN(P2_U3207) );
  AND2_X1 U23492 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20445), .ZN(P2_U3208) );
  NAND2_X1 U23493 ( .A1(n20456), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20458) );
  NAND3_X1 U23494 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20458), .ZN(n20448) );
  AOI211_X1 U23495 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21335), .A(
        n20446), .B(n20556), .ZN(n20447) );
  INV_X1 U23496 ( .A(NA), .ZN(n21340) );
  NOR3_X1 U23497 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21340), .ZN(n20463) );
  AOI211_X1 U23498 ( .C1(n20464), .C2(n20448), .A(n20447), .B(n20463), .ZN(
        n20449) );
  INV_X1 U23499 ( .A(n20449), .ZN(P2_U3209) );
  AOI21_X1 U23500 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21335), .A(n20464), 
        .ZN(n20455) );
  NOR2_X1 U23501 ( .A1(n19734), .A2(n20455), .ZN(n20451) );
  AOI21_X1 U23502 ( .B1(n20451), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n20450), .ZN(n20452) );
  OAI211_X1 U23503 ( .C1(n21335), .C2(n20453), .A(n20452), .B(n20458), .ZN(
        P2_U3210) );
  NOR2_X1 U23504 ( .A1(n20454), .A2(n20464), .ZN(n20457) );
  AOI21_X1 U23505 ( .B1(n20457), .B2(n20456), .A(n20455), .ZN(n20462) );
  OAI22_X1 U23506 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20459), .B1(NA), 
        .B2(n20458), .ZN(n20460) );
  OAI211_X1 U23507 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20460), .ZN(n20461) );
  OAI21_X1 U23508 ( .B1(n20463), .B2(n20462), .A(n20461), .ZN(P2_U3211) );
  NAND2_X2 U23509 ( .A1(n20556), .A2(n20464), .ZN(n20513) );
  NAND2_X2 U23510 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20556), .ZN(n20511) );
  OAI222_X1 U23511 ( .A1(n20513), .A2(n11130), .B1(n20466), .B2(n20556), .C1(
        n20465), .C2(n20511), .ZN(P2_U3212) );
  OAI222_X1 U23512 ( .A1(n20511), .A2(n11130), .B1(n20467), .B2(n20556), .C1(
        n16705), .C2(n20513), .ZN(P2_U3213) );
  OAI222_X1 U23513 ( .A1(n20511), .A2(n16705), .B1(n20468), .B2(n20556), .C1(
        n16691), .C2(n20513), .ZN(P2_U3214) );
  OAI222_X1 U23514 ( .A1(n20513), .A2(n16223), .B1(n20469), .B2(n20556), .C1(
        n16691), .C2(n20511), .ZN(P2_U3215) );
  OAI222_X1 U23515 ( .A1(n20513), .A2(n20471), .B1(n20470), .B2(n20556), .C1(
        n16223), .C2(n20511), .ZN(P2_U3216) );
  OAI222_X1 U23516 ( .A1(n20513), .A2(n16654), .B1(n20472), .B2(n20556), .C1(
        n20471), .C2(n20511), .ZN(P2_U3217) );
  OAI222_X1 U23517 ( .A1(n20513), .A2(n20474), .B1(n20473), .B2(n20556), .C1(
        n16654), .C2(n20511), .ZN(P2_U3218) );
  INV_X1 U23518 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20476) );
  OAI222_X1 U23519 ( .A1(n20513), .A2(n20476), .B1(n20475), .B2(n20556), .C1(
        n20474), .C2(n20511), .ZN(P2_U3219) );
  OAI222_X1 U23520 ( .A1(n20513), .A2(n20478), .B1(n20477), .B2(n20556), .C1(
        n20476), .C2(n20511), .ZN(P2_U3220) );
  OAI222_X1 U23521 ( .A1(n20513), .A2(n11558), .B1(n20479), .B2(n20556), .C1(
        n20478), .C2(n20511), .ZN(P2_U3221) );
  OAI222_X1 U23522 ( .A1(n20513), .A2(n20481), .B1(n20480), .B2(n20556), .C1(
        n11558), .C2(n20511), .ZN(P2_U3222) );
  OAI222_X1 U23523 ( .A1(n20513), .A2(n20483), .B1(n20482), .B2(n20556), .C1(
        n20481), .C2(n20511), .ZN(P2_U3223) );
  OAI222_X1 U23524 ( .A1(n20513), .A2(n20484), .B1(n21553), .B2(n20556), .C1(
        n20483), .C2(n20511), .ZN(P2_U3224) );
  OAI222_X1 U23525 ( .A1(n20513), .A2(n20485), .B1(n21680), .B2(n20556), .C1(
        n20484), .C2(n20511), .ZN(P2_U3225) );
  OAI222_X1 U23526 ( .A1(n20513), .A2(n20487), .B1(n20486), .B2(n20556), .C1(
        n20485), .C2(n20511), .ZN(P2_U3226) );
  OAI222_X1 U23527 ( .A1(n20513), .A2(n20488), .B1(n21569), .B2(n20556), .C1(
        n20487), .C2(n20511), .ZN(P2_U3227) );
  OAI222_X1 U23528 ( .A1(n20513), .A2(n20490), .B1(n20489), .B2(n20556), .C1(
        n20488), .C2(n20511), .ZN(P2_U3228) );
  OAI222_X1 U23529 ( .A1(n20513), .A2(n16079), .B1(n20491), .B2(n20556), .C1(
        n20490), .C2(n20511), .ZN(P2_U3229) );
  OAI222_X1 U23530 ( .A1(n20513), .A2(n20493), .B1(n20492), .B2(n20556), .C1(
        n16079), .C2(n20511), .ZN(P2_U3230) );
  OAI222_X1 U23531 ( .A1(n20513), .A2(n20495), .B1(n20494), .B2(n20556), .C1(
        n20493), .C2(n20511), .ZN(P2_U3231) );
  OAI222_X1 U23532 ( .A1(n20513), .A2(n20497), .B1(n20496), .B2(n20556), .C1(
        n20495), .C2(n20511), .ZN(P2_U3232) );
  OAI222_X1 U23533 ( .A1(n20513), .A2(n20499), .B1(n20498), .B2(n20556), .C1(
        n20497), .C2(n20511), .ZN(P2_U3233) );
  OAI222_X1 U23534 ( .A1(n20513), .A2(n20501), .B1(n20500), .B2(n20556), .C1(
        n20499), .C2(n20511), .ZN(P2_U3234) );
  OAI222_X1 U23535 ( .A1(n20513), .A2(n20503), .B1(n20502), .B2(n20556), .C1(
        n20501), .C2(n20511), .ZN(P2_U3235) );
  INV_X1 U23536 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20505) );
  OAI222_X1 U23537 ( .A1(n20513), .A2(n20505), .B1(n20504), .B2(n20556), .C1(
        n20503), .C2(n20511), .ZN(P2_U3236) );
  OAI222_X1 U23538 ( .A1(n20513), .A2(n16488), .B1(n20506), .B2(n20556), .C1(
        n20505), .C2(n20511), .ZN(P2_U3237) );
  OAI222_X1 U23539 ( .A1(n20511), .A2(n16488), .B1(n20507), .B2(n20556), .C1(
        n20508), .C2(n20513), .ZN(P2_U3238) );
  OAI222_X1 U23540 ( .A1(n20513), .A2(n15949), .B1(n20509), .B2(n20556), .C1(
        n20508), .C2(n20511), .ZN(P2_U3239) );
  OAI222_X1 U23541 ( .A1(n20513), .A2(n13652), .B1(n20510), .B2(n20556), .C1(
        n15949), .C2(n20511), .ZN(P2_U3240) );
  OAI222_X1 U23542 ( .A1(n20513), .A2(n13767), .B1(n20512), .B2(n20556), .C1(
        n13652), .C2(n20511), .ZN(P2_U3241) );
  OAI22_X1 U23543 ( .A1(n20557), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20556), .ZN(n20514) );
  INV_X1 U23544 ( .A(n20514), .ZN(P2_U3585) );
  MUX2_X1 U23545 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20557), .Z(P2_U3586) );
  OAI22_X1 U23546 ( .A1(n20557), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20556), .ZN(n20515) );
  INV_X1 U23547 ( .A(n20515), .ZN(P2_U3587) );
  OAI22_X1 U23548 ( .A1(n20557), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20556), .ZN(n20516) );
  INV_X1 U23549 ( .A(n20516), .ZN(P2_U3588) );
  OAI21_X1 U23550 ( .B1(n20520), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20518), 
        .ZN(n20517) );
  INV_X1 U23551 ( .A(n20517), .ZN(P2_U3591) );
  OAI21_X1 U23552 ( .B1(n20520), .B2(n20519), .A(n20518), .ZN(P2_U3592) );
  NAND2_X1 U23553 ( .A1(n20522), .A2(n20521), .ZN(n20539) );
  NAND3_X1 U23554 ( .A1(n20524), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20523), 
        .ZN(n20526) );
  NAND2_X1 U23555 ( .A1(n20526), .A2(n20525), .ZN(n20534) );
  NAND2_X1 U23556 ( .A1(n20539), .A2(n20534), .ZN(n20531) );
  AOI222_X1 U23557 ( .A1(n20531), .A2(n20530), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20529), .C1(n20528), .C2(n20527), .ZN(n20532) );
  AOI22_X1 U23558 ( .A1(n20543), .A2(n20533), .B1(n20532), .B2(n20540), .ZN(
        P2_U3602) );
  INV_X1 U23559 ( .A(n20534), .ZN(n20536) );
  AOI22_X1 U23560 ( .A1(n20537), .A2(n20536), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20535), .ZN(n20538) );
  AND2_X1 U23561 ( .A1(n20539), .A2(n20538), .ZN(n20541) );
  AOI22_X1 U23562 ( .A1(n20543), .A2(n20542), .B1(n20541), .B2(n20540), .ZN(
        P2_U3603) );
  INV_X1 U23563 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20544) );
  AOI22_X1 U23564 ( .A1(n20556), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20544), 
        .B2(n20557), .ZN(P2_U3608) );
  INV_X1 U23565 ( .A(n20545), .ZN(n20549) );
  INV_X1 U23566 ( .A(n20546), .ZN(n20548) );
  OAI22_X1 U23567 ( .A1(n20550), .A2(n20549), .B1(n20548), .B2(n20547), .ZN(
        n20551) );
  INV_X1 U23568 ( .A(n20551), .ZN(n20552) );
  NAND2_X1 U23569 ( .A1(n20553), .A2(n20552), .ZN(n20555) );
  MUX2_X1 U23570 ( .A(P2_MORE_REG_SCAN_IN), .B(n20555), .S(n20554), .Z(
        P2_U3609) );
  OAI22_X1 U23571 ( .A1(n20557), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20556), .ZN(n20558) );
  INV_X1 U23572 ( .A(n20558), .ZN(P2_U3611) );
  AOI21_X1 U23573 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21637), .A(n21332), 
        .ZN(n20566) );
  INV_X1 U23574 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20559) );
  NAND2_X2 U23575 ( .A1(n21332), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21380) );
  AOI21_X1 U23576 ( .B1(n20566), .B2(n20559), .A(n21392), .ZN(P1_U2802) );
  INV_X1 U23577 ( .A(n20560), .ZN(n20562) );
  OAI21_X1 U23578 ( .B1(n20562), .B2(n20561), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20563) );
  OAI21_X1 U23579 ( .B1(n20564), .B2(n17176), .A(n20563), .ZN(P1_U2803) );
  NOR2_X1 U23580 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20567) );
  OAI21_X1 U23581 ( .B1(n20567), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21380), .ZN(
        n20565) );
  OAI21_X1 U23582 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21380), .A(n20565), 
        .ZN(P1_U2804) );
  OAI21_X1 U23583 ( .B1(BS16), .B2(n20567), .A(n21397), .ZN(n21395) );
  OAI21_X1 U23584 ( .B1(n21397), .B2(n21232), .A(n21395), .ZN(P1_U2805) );
  AOI21_X1 U23585 ( .B1(n20568), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20716), .ZN(
        n20569) );
  INV_X1 U23586 ( .A(n20569), .ZN(P1_U2806) );
  NOR4_X1 U23587 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20573) );
  NOR4_X1 U23588 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20572) );
  NOR4_X1 U23589 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20571) );
  NOR4_X1 U23590 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20570) );
  NAND4_X1 U23591 ( .A1(n20573), .A2(n20572), .A3(n20571), .A4(n20570), .ZN(
        n20579) );
  NOR4_X1 U23592 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20577) );
  AOI211_X1 U23593 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_6__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20576) );
  NOR4_X1 U23594 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20575) );
  NOR4_X1 U23595 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20574) );
  NAND4_X1 U23596 ( .A1(n20577), .A2(n20576), .A3(n20575), .A4(n20574), .ZN(
        n20578) );
  NOR2_X1 U23597 ( .A1(n20579), .A2(n20578), .ZN(n21402) );
  INV_X1 U23598 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20581) );
  NOR3_X1 U23599 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20582) );
  OAI21_X1 U23600 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20582), .A(n21402), .ZN(
        n20580) );
  OAI21_X1 U23601 ( .B1(n21402), .B2(n20581), .A(n20580), .ZN(P1_U2807) );
  INV_X1 U23602 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21396) );
  AOI21_X1 U23603 ( .B1(n21398), .B2(n21396), .A(n20582), .ZN(n20583) );
  INV_X1 U23604 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21604) );
  INV_X1 U23605 ( .A(n21402), .ZN(n21405) );
  AOI22_X1 U23606 ( .A1(n21402), .A2(n20583), .B1(n21604), .B2(n21405), .ZN(
        P1_U2808) );
  NAND2_X1 U23607 ( .A1(n20585), .A2(n20584), .ZN(n20604) );
  NOR2_X1 U23608 ( .A1(n20637), .A2(n20586), .ZN(n20591) );
  AOI21_X1 U23609 ( .B1(n20608), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20607), .ZN(n20588) );
  NAND2_X1 U23610 ( .A1(n20641), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n20587) );
  OAI211_X1 U23611 ( .C1(n20648), .C2(n20589), .A(n20588), .B(n20587), .ZN(
        n20590) );
  AOI211_X1 U23612 ( .C1(n20592), .C2(n20601), .A(n20591), .B(n20590), .ZN(
        n20593) );
  OAI221_X1 U23613 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20594), .C1(n15662), 
        .C2(n20604), .A(n20593), .ZN(P1_U2833) );
  NAND2_X1 U23614 ( .A1(n20606), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n20605) );
  INV_X1 U23615 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21355) );
  NOR2_X1 U23616 ( .A1(n20637), .A2(n20595), .ZN(n20600) );
  AOI21_X1 U23617 ( .B1(n20608), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20607), .ZN(n20597) );
  NAND2_X1 U23618 ( .A1(n20641), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n20596) );
  OAI211_X1 U23619 ( .C1(n20648), .C2(n20598), .A(n20597), .B(n20596), .ZN(
        n20599) );
  AOI211_X1 U23620 ( .C1(n20602), .C2(n20601), .A(n20600), .B(n20599), .ZN(
        n20603) );
  OAI221_X1 U23621 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20605), .C1(n21355), 
        .C2(n20604), .A(n20603), .ZN(P1_U2834) );
  INV_X1 U23622 ( .A(n20606), .ZN(n20619) );
  AOI21_X1 U23623 ( .B1(n20608), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20607), .ZN(n20609) );
  INV_X1 U23624 ( .A(n20609), .ZN(n20613) );
  INV_X1 U23625 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20654) );
  OAI22_X1 U23626 ( .A1(n20637), .A2(n20611), .B1(n20654), .B2(n20610), .ZN(
        n20612) );
  AOI211_X1 U23627 ( .C1(n20627), .C2(n20649), .A(n20613), .B(n20612), .ZN(
        n20618) );
  OR2_X1 U23628 ( .A1(n20615), .A2(n20614), .ZN(n20633) );
  INV_X1 U23629 ( .A(n20633), .ZN(n20616) );
  AOI22_X1 U23630 ( .A1(n20652), .A2(n20635), .B1(n20616), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20617) );
  OAI211_X1 U23631 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20619), .A(n20618), .B(
        n20617), .ZN(P1_U2835) );
  INV_X1 U23632 ( .A(n20620), .ZN(n20714) );
  NOR2_X1 U23633 ( .A1(n20621), .A2(n20639), .ZN(n20626) );
  NAND2_X1 U23634 ( .A1(n20641), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n20623) );
  OAI211_X1 U23635 ( .C1(n20636), .C2(n20624), .A(n20623), .B(n20622), .ZN(
        n20625) );
  AOI211_X1 U23636 ( .C1(n20628), .C2(n20627), .A(n20626), .B(n20625), .ZN(
        n20629) );
  OAI21_X1 U23637 ( .B1(n20637), .B2(n20719), .A(n20629), .ZN(n20630) );
  AOI21_X1 U23638 ( .B1(n20714), .B2(n20635), .A(n20630), .ZN(n20631) );
  OAI221_X1 U23639 ( .B1(n20633), .B2(n21353), .C1(n20633), .C2(n20632), .A(
        n20631), .ZN(P1_U2836) );
  NAND2_X1 U23640 ( .A1(n20635), .A2(n20634), .ZN(n20644) );
  MUX2_X1 U23641 ( .A(n20637), .B(n20636), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n20643) );
  OAI22_X1 U23642 ( .A1(n20639), .A2(n21153), .B1(n20638), .B2(n21398), .ZN(
        n20640) );
  AOI21_X1 U23643 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(n20641), .A(n20640), .ZN(
        n20642) );
  AND3_X1 U23644 ( .A1(n20644), .A2(n20643), .A3(n20642), .ZN(n20647) );
  OR2_X1 U23645 ( .A1(n20645), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20646) );
  OAI211_X1 U23646 ( .C1(n20763), .C2(n20648), .A(n20647), .B(n20646), .ZN(
        P1_U2839) );
  AOI22_X1 U23647 ( .A1(n20652), .A2(n20651), .B1(n20650), .B2(n20649), .ZN(
        n20653) );
  OAI21_X1 U23648 ( .B1(n20655), .B2(n20654), .A(n20653), .ZN(P1_U2867) );
  OAI222_X1 U23649 ( .A1(n20680), .A2(n20657), .B1(n20686), .B2(n20656), .C1(
        n21633), .C2(n20678), .ZN(P1_U2921) );
  INV_X1 U23650 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20659) );
  AOI22_X1 U23651 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20658) );
  OAI21_X1 U23652 ( .B1(n20659), .B2(n20686), .A(n20658), .ZN(P1_U2922) );
  AOI22_X1 U23653 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20660) );
  OAI21_X1 U23654 ( .B1(n15410), .B2(n20686), .A(n20660), .ZN(P1_U2923) );
  AOI22_X1 U23655 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20661) );
  OAI21_X1 U23656 ( .B1(n15412), .B2(n20686), .A(n20661), .ZN(P1_U2924) );
  INV_X1 U23657 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n21526) );
  AOI22_X1 U23658 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n20671), .B1(n20683), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20662) );
  OAI21_X1 U23659 ( .B1(n21526), .B2(n20680), .A(n20662), .ZN(P1_U2925) );
  AOI222_X1 U23660 ( .A1(n20684), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20671), 
        .B2(P1_EAX_REG_10__SCAN_IN), .C1(P1_DATAO_REG_10__SCAN_IN), .C2(n20683), .ZN(n20663) );
  INV_X1 U23661 ( .A(n20663), .ZN(P1_U2926) );
  AOI22_X1 U23662 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20664) );
  OAI21_X1 U23663 ( .B1(n20665), .B2(n20686), .A(n20664), .ZN(P1_U2927) );
  AOI22_X1 U23664 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20666) );
  OAI21_X1 U23665 ( .B1(n21625), .B2(n20686), .A(n20666), .ZN(P1_U2928) );
  AOI22_X1 U23666 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20667) );
  OAI21_X1 U23667 ( .B1(n20668), .B2(n20686), .A(n20667), .ZN(P1_U2929) );
  AOI22_X1 U23668 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20669) );
  OAI21_X1 U23669 ( .B1(n20670), .B2(n20686), .A(n20669), .ZN(P1_U2930) );
  AOI222_X1 U23670 ( .A1(n20684), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20671), 
        .B2(P1_EAX_REG_5__SCAN_IN), .C1(P1_DATAO_REG_5__SCAN_IN), .C2(n20683), 
        .ZN(n20672) );
  INV_X1 U23671 ( .A(n20672), .ZN(P1_U2931) );
  INV_X1 U23672 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n21670) );
  OAI222_X1 U23673 ( .A1(n20680), .A2(n21670), .B1(n20686), .B2(n20674), .C1(
        n20678), .C2(n20673), .ZN(P1_U2932) );
  INV_X1 U23674 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n21592) );
  OAI222_X1 U23675 ( .A1(n20680), .A2(n21592), .B1(n20686), .B2(n20676), .C1(
        n20678), .C2(n20675), .ZN(P1_U2933) );
  INV_X1 U23676 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n21500) );
  OAI222_X1 U23677 ( .A1(n20680), .A2(n21500), .B1(n20686), .B2(n20679), .C1(
        n20678), .C2(n20677), .ZN(P1_U2934) );
  AOI22_X1 U23678 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20681) );
  OAI21_X1 U23679 ( .B1(n20682), .B2(n20686), .A(n20681), .ZN(P1_U2935) );
  AOI22_X1 U23680 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20684), .B1(n20683), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20685) );
  OAI21_X1 U23681 ( .B1(n20687), .B2(n20686), .A(n20685), .ZN(P1_U2936) );
  AOI22_X1 U23682 ( .A1(n14429), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20706), .ZN(n20690) );
  INV_X1 U23683 ( .A(n20688), .ZN(n20689) );
  NAND2_X1 U23684 ( .A1(n20698), .A2(n20689), .ZN(n20700) );
  NAND2_X1 U23685 ( .A1(n20690), .A2(n20700), .ZN(P1_U2948) );
  AOI22_X1 U23686 ( .A1(n14429), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20693) );
  INV_X1 U23687 ( .A(n20691), .ZN(n20692) );
  NAND2_X1 U23688 ( .A1(n20698), .A2(n20692), .ZN(n20702) );
  NAND2_X1 U23689 ( .A1(n20693), .A2(n20702), .ZN(P1_U2949) );
  AOI22_X1 U23690 ( .A1(n14429), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20696) );
  INV_X1 U23691 ( .A(n20694), .ZN(n20695) );
  NAND2_X1 U23692 ( .A1(n20698), .A2(n20695), .ZN(n20704) );
  NAND2_X1 U23693 ( .A1(n20696), .A2(n20704), .ZN(P1_U2950) );
  AOI22_X1 U23694 ( .A1(n14429), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20706), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20699) );
  NAND2_X1 U23695 ( .A1(n20698), .A2(n20697), .ZN(n20707) );
  NAND2_X1 U23696 ( .A1(n20699), .A2(n20707), .ZN(P1_U2951) );
  AOI22_X1 U23697 ( .A1(n14429), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20706), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20701) );
  NAND2_X1 U23698 ( .A1(n20701), .A2(n20700), .ZN(P1_U2963) );
  AOI22_X1 U23699 ( .A1(n14429), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20706), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20703) );
  NAND2_X1 U23700 ( .A1(n20703), .A2(n20702), .ZN(P1_U2964) );
  AOI22_X1 U23701 ( .A1(n14429), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20706), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20705) );
  NAND2_X1 U23702 ( .A1(n20705), .A2(n20704), .ZN(P1_U2965) );
  AOI22_X1 U23703 ( .A1(n14429), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20706), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20708) );
  NAND2_X1 U23704 ( .A1(n20708), .A2(n20707), .ZN(P1_U2966) );
  AOI22_X1 U23705 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20727), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20718) );
  AOI21_X1 U23706 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14625), .A(
        n20710), .ZN(n20713) );
  XNOR2_X1 U23707 ( .A(n20711), .B(n20733), .ZN(n20712) );
  XNOR2_X1 U23708 ( .A(n20713), .B(n20712), .ZN(n20731) );
  AOI22_X1 U23709 ( .A1(n20731), .A2(n20716), .B1(n20715), .B2(n20714), .ZN(
        n20717) );
  OAI211_X1 U23710 ( .C1(n20720), .C2(n20719), .A(n20718), .B(n20717), .ZN(
        P1_U2995) );
  NOR2_X1 U23711 ( .A1(n20722), .A2(n20721), .ZN(n20750) );
  OAI21_X1 U23712 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20723), .A(
        n20772), .ZN(n20743) );
  AOI211_X1 U23713 ( .C1(n20754), .C2(n20724), .A(n20750), .B(n20743), .ZN(
        n20742) );
  AOI211_X1 U23714 ( .C1(n20733), .C2(n9919), .A(n20725), .B(n20737), .ZN(
        n20726) );
  AOI21_X1 U23715 ( .B1(n20727), .B2(P1_REIP_REG_4__SCAN_IN), .A(n20726), .ZN(
        n20728) );
  OAI21_X1 U23716 ( .B1(n20774), .B2(n20729), .A(n20728), .ZN(n20730) );
  AOI21_X1 U23717 ( .B1(n20731), .B2(n20757), .A(n20730), .ZN(n20732) );
  OAI21_X1 U23718 ( .B1(n20742), .B2(n20733), .A(n20732), .ZN(P1_U3027) );
  AOI21_X1 U23719 ( .B1(n20736), .B2(n20735), .A(n20734), .ZN(n20741) );
  INV_X1 U23720 ( .A(n20737), .ZN(n20738) );
  AOI22_X1 U23721 ( .A1(n20739), .A2(n20757), .B1(n20738), .B2(n9919), .ZN(
        n20740) );
  OAI211_X1 U23722 ( .C1(n20742), .C2(n9919), .A(n20741), .B(n20740), .ZN(
        P1_U3028) );
  NOR2_X1 U23723 ( .A1(n20770), .A2(n20768), .ZN(n20744) );
  AOI21_X1 U23724 ( .B1(n20756), .B2(n20744), .A(n20743), .ZN(n20753) );
  AND3_X1 U23725 ( .A1(n20746), .A2(n20745), .A3(n20757), .ZN(n20751) );
  INV_X1 U23726 ( .A(n20747), .ZN(n20748) );
  OAI22_X1 U23727 ( .A1(n20774), .A2(n20748), .B1(n21350), .B2(n20781), .ZN(
        n20749) );
  NOR3_X1 U23728 ( .A1(n20751), .A2(n20750), .A3(n20749), .ZN(n20752) );
  OAI221_X1 U23729 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20755), .C1(
        n20754), .C2(n20753), .A(n20752), .ZN(P1_U3029) );
  NAND2_X1 U23730 ( .A1(n20756), .A2(n20770), .ZN(n20779) );
  AND3_X1 U23731 ( .A1(n20759), .A2(n20758), .A3(n20757), .ZN(n20766) );
  NOR3_X1 U23732 ( .A1(n20761), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20760), .ZN(n20765) );
  OAI21_X1 U23733 ( .B1(n20774), .B2(n20763), .A(n20762), .ZN(n20764) );
  NOR3_X1 U23734 ( .A1(n20766), .A2(n20765), .A3(n20764), .ZN(n20767) );
  OAI221_X1 U23735 ( .B1(n20768), .B2(n20772), .C1(n20768), .C2(n20779), .A(
        n20767), .ZN(P1_U3030) );
  INV_X1 U23736 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21404) );
  AOI22_X1 U23737 ( .A1(n20772), .A2(n20771), .B1(n20770), .B2(n20769), .ZN(
        n20778) );
  OAI22_X1 U23738 ( .A1(n20776), .A2(n20775), .B1(n20774), .B2(n20773), .ZN(
        n20777) );
  NOR2_X1 U23739 ( .A1(n20778), .A2(n20777), .ZN(n20780) );
  OAI211_X1 U23740 ( .C1(n21404), .C2(n20781), .A(n20780), .B(n20779), .ZN(
        P1_U3031) );
  NOR2_X1 U23741 ( .A1(n20783), .A2(n20782), .ZN(P1_U3032) );
  AOI21_X1 U23742 ( .B1(n20785), .B2(n21326), .A(n21232), .ZN(n20786) );
  NOR2_X1 U23743 ( .A1(n20786), .A2(n21266), .ZN(n20795) );
  NOR2_X1 U23744 ( .A1(n20854), .A2(n14513), .ZN(n20793) );
  INV_X1 U23745 ( .A(n20787), .ZN(n20792) );
  NAND2_X1 U23746 ( .A1(n20792), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21034) );
  INV_X1 U23747 ( .A(n21034), .ZN(n21089) );
  INV_X1 U23748 ( .A(n21032), .ZN(n20788) );
  NAND2_X1 U23749 ( .A1(n20788), .A2(n21087), .ZN(n20915) );
  INV_X1 U23750 ( .A(n20915), .ZN(n20789) );
  NOR2_X1 U23751 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20791), .ZN(
        n20828) );
  AOI22_X1 U23752 ( .A1(n21263), .A2(n20828), .B1(n21288), .B2(n21163), .ZN(
        n20799) );
  NOR2_X1 U23753 ( .A1(n20792), .A2(n21201), .ZN(n21154) );
  INV_X1 U23754 ( .A(n20793), .ZN(n20794) );
  AOI22_X1 U23755 ( .A1(n20795), .A2(n20794), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20915), .ZN(n20796) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21275), .ZN(n20798) );
  OAI211_X1 U23757 ( .C1(n20833), .C2(n21166), .A(n20799), .B(n20798), .ZN(
        P1_U3033) );
  AOI22_X1 U23758 ( .A1(n21279), .A2(n20828), .B1(n21288), .B2(n21167), .ZN(
        n20802) );
  INV_X1 U23759 ( .A(n20894), .ZN(n21281) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21281), .ZN(n20801) );
  OAI211_X1 U23761 ( .C1(n20833), .C2(n21170), .A(n20802), .B(n20801), .ZN(
        P1_U3034) );
  INV_X1 U23762 ( .A(n21286), .ZN(n21174) );
  NOR2_X2 U23763 ( .A1(n20827), .A2(n20804), .ZN(n21285) );
  AOI22_X1 U23764 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20829), .B1(DATAI_26_), 
        .B2(n14553), .ZN(n21292) );
  INV_X1 U23765 ( .A(n21292), .ZN(n21171) );
  AOI22_X1 U23766 ( .A1(n21285), .A2(n20828), .B1(n21288), .B2(n21171), .ZN(
        n20806) );
  AOI22_X1 U23767 ( .A1(DATAI_18_), .A2(n14553), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20829), .ZN(n20897) );
  INV_X1 U23768 ( .A(n20897), .ZN(n21287) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21287), .ZN(n20805) );
  OAI211_X1 U23770 ( .C1(n20833), .C2(n21174), .A(n20806), .B(n20805), .ZN(
        P1_U3035) );
  NOR2_X2 U23771 ( .A1(n20827), .A2(n12648), .ZN(n21293) );
  AOI22_X1 U23772 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20829), .B1(DATAI_27_), 
        .B2(n14553), .ZN(n20808) );
  AOI22_X1 U23773 ( .A1(n21293), .A2(n20828), .B1(n21288), .B2(n21295), .ZN(
        n20810) );
  AOI22_X2 U23774 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20829), .B1(DATAI_19_), 
        .B2(n14553), .ZN(n21298) );
  INV_X1 U23775 ( .A(n21298), .ZN(n21175) );
  AOI22_X1 U23776 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21175), .ZN(n20809) );
  OAI211_X1 U23777 ( .C1(n20833), .C2(n21178), .A(n20810), .B(n20809), .ZN(
        P1_U3036) );
  INV_X1 U23778 ( .A(n21300), .ZN(n21182) );
  NOR2_X2 U23779 ( .A1(n20827), .A2(n20812), .ZN(n21299) );
  AOI22_X1 U23780 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20829), .B1(DATAI_28_), 
        .B2(n14553), .ZN(n20813) );
  AOI22_X1 U23781 ( .A1(n21299), .A2(n20828), .B1(n21288), .B2(n21301), .ZN(
        n20815) );
  AOI22_X2 U23782 ( .A1(DATAI_20_), .A2(n14553), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20829), .ZN(n21304) );
  INV_X1 U23783 ( .A(n21304), .ZN(n21179) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21179), .ZN(n20814) );
  OAI211_X1 U23785 ( .C1(n20833), .C2(n21182), .A(n20815), .B(n20814), .ZN(
        P1_U3037) );
  INV_X1 U23786 ( .A(n21306), .ZN(n21186) );
  NOR2_X2 U23787 ( .A1(n20827), .A2(n12658), .ZN(n21305) );
  AOI22_X1 U23788 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20829), .B1(DATAI_29_), 
        .B2(n14553), .ZN(n20817) );
  AOI22_X1 U23789 ( .A1(n21305), .A2(n20828), .B1(n21288), .B2(n21307), .ZN(
        n20819) );
  INV_X1 U23790 ( .A(n21310), .ZN(n21183) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21183), .ZN(n20818) );
  OAI211_X1 U23792 ( .C1(n20833), .C2(n21186), .A(n20819), .B(n20818), .ZN(
        P1_U3038) );
  INV_X1 U23793 ( .A(n21312), .ZN(n21190) );
  NOR2_X2 U23794 ( .A1(n20827), .A2(n12630), .ZN(n21311) );
  AOI22_X1 U23795 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20829), .B1(DATAI_30_), 
        .B2(n14553), .ZN(n20821) );
  AOI22_X1 U23796 ( .A1(n21311), .A2(n20828), .B1(n21288), .B2(n21313), .ZN(
        n20823) );
  AOI22_X2 U23797 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20829), .B1(DATAI_22_), 
        .B2(n14553), .ZN(n21316) );
  INV_X1 U23798 ( .A(n21316), .ZN(n21187) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21187), .ZN(n20822) );
  OAI211_X1 U23800 ( .C1(n20833), .C2(n21190), .A(n20823), .B(n20822), .ZN(
        P1_U3039) );
  NOR2_X2 U23801 ( .A1(n20827), .A2(n20826), .ZN(n21320) );
  AOI22_X1 U23802 ( .A1(DATAI_31_), .A2(n14553), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20829), .ZN(n21030) );
  INV_X1 U23803 ( .A(n21030), .ZN(n21321) );
  AOI22_X1 U23804 ( .A1(n21320), .A2(n20828), .B1(n21288), .B2(n21321), .ZN(
        n20832) );
  AOI22_X1 U23805 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20829), .B1(DATAI_23_), 
        .B2(n14553), .ZN(n21327) );
  INV_X1 U23806 ( .A(n21327), .ZN(n21191) );
  AOI22_X1 U23807 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20830), .B1(
        n20848), .B2(n21191), .ZN(n20831) );
  OAI211_X1 U23808 ( .C1(n20833), .C2(n21197), .A(n20832), .B(n20831), .ZN(
        P1_U3040) );
  INV_X1 U23809 ( .A(n20834), .ZN(n20846) );
  AOI22_X1 U23810 ( .A1(n21286), .A2(n20846), .B1(n21285), .B2(n20847), .ZN(
        n20836) );
  AOI22_X1 U23811 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20849), .B1(
        n20848), .B2(n21171), .ZN(n20835) );
  OAI211_X1 U23812 ( .C1(n20897), .C2(n20866), .A(n20836), .B(n20835), .ZN(
        P1_U3043) );
  AOI22_X1 U23813 ( .A1(n21294), .A2(n20846), .B1(n21293), .B2(n20847), .ZN(
        n20838) );
  AOI22_X1 U23814 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20849), .B1(
        n20848), .B2(n21295), .ZN(n20837) );
  OAI211_X1 U23815 ( .C1(n21298), .C2(n20866), .A(n20838), .B(n20837), .ZN(
        P1_U3044) );
  AOI22_X1 U23816 ( .A1(n21300), .A2(n20846), .B1(n21299), .B2(n20847), .ZN(
        n20840) );
  AOI22_X1 U23817 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20849), .B1(
        n20848), .B2(n21301), .ZN(n20839) );
  OAI211_X1 U23818 ( .C1(n21304), .C2(n20866), .A(n20840), .B(n20839), .ZN(
        P1_U3045) );
  INV_X1 U23819 ( .A(n20849), .ZN(n20843) );
  INV_X1 U23820 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n21473) );
  AOI22_X1 U23821 ( .A1(n21306), .A2(n20846), .B1(n21305), .B2(n20847), .ZN(
        n20842) );
  AOI22_X1 U23822 ( .A1(n20875), .A2(n21183), .B1(n20848), .B2(n21307), .ZN(
        n20841) );
  OAI211_X1 U23823 ( .C1(n20843), .C2(n21473), .A(n20842), .B(n20841), .ZN(
        P1_U3046) );
  AOI22_X1 U23824 ( .A1(n21312), .A2(n20846), .B1(n21311), .B2(n20847), .ZN(
        n20845) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20849), .B1(
        n20848), .B2(n21313), .ZN(n20844) );
  OAI211_X1 U23826 ( .C1(n21316), .C2(n20866), .A(n20845), .B(n20844), .ZN(
        P1_U3047) );
  AOI22_X1 U23827 ( .A1(n21320), .A2(n20847), .B1(n21318), .B2(n20846), .ZN(
        n20851) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20849), .B1(
        n20848), .B2(n21321), .ZN(n20850) );
  OAI211_X1 U23829 ( .C1(n21327), .C2(n20866), .A(n20851), .B(n20850), .ZN(
        P1_U3048) );
  NAND3_X1 U23830 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21156), .A3(
        n21157), .ZN(n20887) );
  NOR2_X1 U23831 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20887), .ZN(
        n20876) );
  NAND2_X1 U23832 ( .A1(n9707), .A2(n13816), .ZN(n21231) );
  AOI22_X1 U23833 ( .A1(n21263), .A2(n20876), .B1(n20904), .B2(n21275), .ZN(
        n20861) );
  AOI21_X1 U23834 ( .B1(n20866), .B2(n20912), .A(n21232), .ZN(n20853) );
  NOR2_X1 U23835 ( .A1(n20853), .A2(n21266), .ZN(n20857) );
  INV_X1 U23836 ( .A(n20854), .ZN(n20884) );
  NAND2_X1 U23837 ( .A1(n20884), .A2(n14513), .ZN(n20858) );
  INV_X1 U23838 ( .A(n20876), .ZN(n20855) );
  AOI22_X1 U23839 ( .A1(n20857), .A2(n20858), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20855), .ZN(n20856) );
  OAI21_X1 U23840 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21087), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20980) );
  NAND3_X1 U23841 ( .A1(n21096), .A2(n20856), .A3(n20980), .ZN(n20878) );
  INV_X1 U23842 ( .A(n20857), .ZN(n20859) );
  OR2_X1 U23843 ( .A1(n21087), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20974) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20878), .B1(
        n21264), .B2(n20877), .ZN(n20860) );
  OAI211_X1 U23845 ( .C1(n21278), .C2(n20866), .A(n20861), .B(n20860), .ZN(
        P1_U3049) );
  AOI22_X1 U23846 ( .A1(n21279), .A2(n20876), .B1(n20904), .B2(n21281), .ZN(
        n20863) );
  AOI22_X1 U23847 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20878), .B1(
        n21280), .B2(n20877), .ZN(n20862) );
  OAI211_X1 U23848 ( .C1(n21284), .C2(n20866), .A(n20863), .B(n20862), .ZN(
        P1_U3050) );
  AOI22_X1 U23849 ( .A1(n21285), .A2(n20876), .B1(n20904), .B2(n21287), .ZN(
        n20865) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20878), .B1(
        n21286), .B2(n20877), .ZN(n20864) );
  OAI211_X1 U23851 ( .C1(n21292), .C2(n20866), .A(n20865), .B(n20864), .ZN(
        P1_U3051) );
  AOI22_X1 U23852 ( .A1(n21293), .A2(n20876), .B1(n20875), .B2(n21295), .ZN(
        n20868) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20878), .B1(
        n21294), .B2(n20877), .ZN(n20867) );
  OAI211_X1 U23854 ( .C1(n21298), .C2(n20912), .A(n20868), .B(n20867), .ZN(
        P1_U3052) );
  AOI22_X1 U23855 ( .A1(n21299), .A2(n20876), .B1(n20875), .B2(n21301), .ZN(
        n20870) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20878), .B1(
        n21300), .B2(n20877), .ZN(n20869) );
  OAI211_X1 U23857 ( .C1(n21304), .C2(n20912), .A(n20870), .B(n20869), .ZN(
        P1_U3053) );
  AOI22_X1 U23858 ( .A1(n21305), .A2(n20876), .B1(n20875), .B2(n21307), .ZN(
        n20872) );
  AOI22_X1 U23859 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20878), .B1(
        n21306), .B2(n20877), .ZN(n20871) );
  OAI211_X1 U23860 ( .C1(n21310), .C2(n20912), .A(n20872), .B(n20871), .ZN(
        P1_U3054) );
  AOI22_X1 U23861 ( .A1(n21311), .A2(n20876), .B1(n20875), .B2(n21313), .ZN(
        n20874) );
  AOI22_X1 U23862 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20878), .B1(
        n21312), .B2(n20877), .ZN(n20873) );
  OAI211_X1 U23863 ( .C1(n21316), .C2(n20912), .A(n20874), .B(n20873), .ZN(
        P1_U3055) );
  AOI22_X1 U23864 ( .A1(n21320), .A2(n20876), .B1(n20875), .B2(n21321), .ZN(
        n20880) );
  AOI22_X1 U23865 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20878), .B1(
        n21318), .B2(n20877), .ZN(n20879) );
  OAI211_X1 U23866 ( .C1(n21327), .C2(n20912), .A(n20880), .B(n20879), .ZN(
        P1_U3056) );
  NOR2_X1 U23867 ( .A1(n21117), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20907) );
  AOI22_X1 U23868 ( .A1(n21263), .A2(n20907), .B1(n20938), .B2(n21275), .ZN(
        n20891) );
  AOI21_X1 U23869 ( .B1(n20881), .B2(n21273), .A(n21270), .ZN(n20888) );
  AND2_X1 U23870 ( .A1(n20883), .A2(n20882), .ZN(n21260) );
  AOI21_X1 U23871 ( .B1(n20884), .B2(n21260), .A(n20907), .ZN(n20889) );
  INV_X1 U23872 ( .A(n20889), .ZN(n20886) );
  NAND2_X1 U23873 ( .A1(n21266), .A2(n20887), .ZN(n20885) );
  OAI211_X1 U23874 ( .C1(n20888), .C2(n20886), .A(n21272), .B(n20885), .ZN(
        n20909) );
  OAI22_X1 U23875 ( .A1(n20889), .A2(n20888), .B1(n21201), .B2(n20887), .ZN(
        n20908) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20909), .B1(
        n21264), .B2(n20908), .ZN(n20890) );
  OAI211_X1 U23877 ( .C1(n21278), .C2(n20912), .A(n20891), .B(n20890), .ZN(
        P1_U3057) );
  AOI22_X1 U23878 ( .A1(n21279), .A2(n20907), .B1(n20904), .B2(n21167), .ZN(
        n20893) );
  AOI22_X1 U23879 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20909), .B1(
        n21280), .B2(n20908), .ZN(n20892) );
  OAI211_X1 U23880 ( .C1(n20894), .C2(n20927), .A(n20893), .B(n20892), .ZN(
        P1_U3058) );
  AOI22_X1 U23881 ( .A1(n21285), .A2(n20907), .B1(n20904), .B2(n21171), .ZN(
        n20896) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20909), .B1(
        n21286), .B2(n20908), .ZN(n20895) );
  OAI211_X1 U23883 ( .C1(n20897), .C2(n20927), .A(n20896), .B(n20895), .ZN(
        P1_U3059) );
  AOI22_X1 U23884 ( .A1(n21293), .A2(n20907), .B1(n20904), .B2(n21295), .ZN(
        n20899) );
  AOI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20909), .B1(
        n21294), .B2(n20908), .ZN(n20898) );
  OAI211_X1 U23886 ( .C1(n21298), .C2(n20927), .A(n20899), .B(n20898), .ZN(
        P1_U3060) );
  AOI22_X1 U23887 ( .A1(n21299), .A2(n20907), .B1(n20904), .B2(n21301), .ZN(
        n20901) );
  AOI22_X1 U23888 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20909), .B1(
        n21300), .B2(n20908), .ZN(n20900) );
  OAI211_X1 U23889 ( .C1(n21304), .C2(n20927), .A(n20901), .B(n20900), .ZN(
        P1_U3061) );
  AOI22_X1 U23890 ( .A1(n21305), .A2(n20907), .B1(n20904), .B2(n21307), .ZN(
        n20903) );
  AOI22_X1 U23891 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20909), .B1(
        n21306), .B2(n20908), .ZN(n20902) );
  OAI211_X1 U23892 ( .C1(n21310), .C2(n20927), .A(n20903), .B(n20902), .ZN(
        P1_U3062) );
  AOI22_X1 U23893 ( .A1(n21311), .A2(n20907), .B1(n20904), .B2(n21313), .ZN(
        n20906) );
  AOI22_X1 U23894 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20909), .B1(
        n21312), .B2(n20908), .ZN(n20905) );
  OAI211_X1 U23895 ( .C1(n21316), .C2(n20927), .A(n20906), .B(n20905), .ZN(
        P1_U3063) );
  AOI22_X1 U23896 ( .A1(n21320), .A2(n20907), .B1(n20938), .B2(n21191), .ZN(
        n20911) );
  AOI22_X1 U23897 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20909), .B1(
        n21318), .B2(n20908), .ZN(n20910) );
  OAI211_X1 U23898 ( .C1(n21030), .C2(n20912), .A(n20911), .B(n20910), .ZN(
        P1_U3064) );
  INV_X1 U23899 ( .A(n21154), .ZN(n21230) );
  NOR2_X1 U23900 ( .A1(n21152), .A2(n20913), .ZN(n21003) );
  NAND3_X1 U23901 ( .A1(n21003), .A2(n21273), .A3(n21153), .ZN(n20914) );
  OAI21_X1 U23902 ( .B1(n20915), .B2(n21230), .A(n20914), .ZN(n20936) );
  NOR3_X1 U23903 ( .A1(n21157), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20945) );
  INV_X1 U23904 ( .A(n20945), .ZN(n20946) );
  NOR2_X1 U23905 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20946), .ZN(
        n20937) );
  AOI22_X1 U23906 ( .A1(n21264), .A2(n20936), .B1(n21263), .B2(n20937), .ZN(
        n20922) );
  INV_X1 U23907 ( .A(n21148), .ZN(n20916) );
  AOI21_X1 U23908 ( .B1(n20927), .B2(n20970), .A(n21232), .ZN(n20917) );
  AOI21_X1 U23909 ( .B1(n21003), .B2(n21153), .A(n20917), .ZN(n20918) );
  NOR2_X1 U23910 ( .A1(n20918), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20920) );
  AOI22_X1 U23911 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20939), .B1(
        n20962), .B2(n21275), .ZN(n20921) );
  OAI211_X1 U23912 ( .C1(n21278), .C2(n20927), .A(n20922), .B(n20921), .ZN(
        P1_U3065) );
  AOI22_X1 U23913 ( .A1(n21280), .A2(n20936), .B1(n21279), .B2(n20937), .ZN(
        n20924) );
  AOI22_X1 U23914 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20939), .B1(
        n20962), .B2(n21281), .ZN(n20923) );
  OAI211_X1 U23915 ( .C1(n21284), .C2(n20927), .A(n20924), .B(n20923), .ZN(
        P1_U3066) );
  AOI22_X1 U23916 ( .A1(n21286), .A2(n20936), .B1(n21285), .B2(n20937), .ZN(
        n20926) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20939), .B1(
        n20962), .B2(n21287), .ZN(n20925) );
  OAI211_X1 U23918 ( .C1(n21292), .C2(n20927), .A(n20926), .B(n20925), .ZN(
        P1_U3067) );
  AOI22_X1 U23919 ( .A1(n21294), .A2(n20936), .B1(n21293), .B2(n20937), .ZN(
        n20929) );
  AOI22_X1 U23920 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n21295), .ZN(n20928) );
  OAI211_X1 U23921 ( .C1(n21298), .C2(n20970), .A(n20929), .B(n20928), .ZN(
        P1_U3068) );
  AOI22_X1 U23922 ( .A1(n21300), .A2(n20936), .B1(n21299), .B2(n20937), .ZN(
        n20931) );
  AOI22_X1 U23923 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n21301), .ZN(n20930) );
  OAI211_X1 U23924 ( .C1(n21304), .C2(n20970), .A(n20931), .B(n20930), .ZN(
        P1_U3069) );
  AOI22_X1 U23925 ( .A1(n21306), .A2(n20936), .B1(n21305), .B2(n20937), .ZN(
        n20933) );
  AOI22_X1 U23926 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n21307), .ZN(n20932) );
  OAI211_X1 U23927 ( .C1(n21310), .C2(n20970), .A(n20933), .B(n20932), .ZN(
        P1_U3070) );
  AOI22_X1 U23928 ( .A1(n21312), .A2(n20936), .B1(n21311), .B2(n20937), .ZN(
        n20935) );
  AOI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n21313), .ZN(n20934) );
  OAI211_X1 U23930 ( .C1(n21316), .C2(n20970), .A(n20935), .B(n20934), .ZN(
        P1_U3071) );
  AOI22_X1 U23931 ( .A1(n21320), .A2(n20937), .B1(n21318), .B2(n20936), .ZN(
        n20941) );
  AOI22_X1 U23932 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n21321), .ZN(n20940) );
  OAI211_X1 U23933 ( .C1(n21327), .C2(n20970), .A(n20941), .B(n20940), .ZN(
        P1_U3072) );
  OAI21_X1 U23934 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21266), .A(n21008), 
        .ZN(n20943) );
  INV_X1 U23935 ( .A(n20942), .ZN(n21200) );
  NOR2_X1 U23936 ( .A1(n21199), .A2(n20946), .ZN(n20966) );
  AOI21_X1 U23937 ( .B1(n21003), .B2(n21200), .A(n20966), .ZN(n20947) );
  NAND2_X1 U23938 ( .A1(n20943), .A2(n20947), .ZN(n20944) );
  OAI211_X1 U23939 ( .C1(n21273), .C2(n20945), .A(n20944), .B(n21272), .ZN(
        n20967) );
  INV_X1 U23940 ( .A(n20967), .ZN(n20951) );
  INV_X1 U23941 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n21725) );
  OAI22_X1 U23942 ( .A1(n20947), .A2(n21266), .B1(n20946), .B2(n21201), .ZN(
        n20965) );
  AOI22_X1 U23943 ( .A1(n21264), .A2(n20965), .B1(n21263), .B2(n20966), .ZN(
        n20950) );
  INV_X1 U23944 ( .A(n21206), .ZN(n20948) );
  AOI22_X1 U23945 ( .A1(n20996), .A2(n21275), .B1(n20962), .B2(n21163), .ZN(
        n20949) );
  OAI211_X1 U23946 ( .C1(n20951), .C2(n21725), .A(n20950), .B(n20949), .ZN(
        P1_U3073) );
  AOI22_X1 U23947 ( .A1(n21280), .A2(n20965), .B1(n21279), .B2(n20966), .ZN(
        n20953) );
  AOI22_X1 U23948 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20967), .B1(
        n20996), .B2(n21281), .ZN(n20952) );
  OAI211_X1 U23949 ( .C1(n21284), .C2(n20970), .A(n20953), .B(n20952), .ZN(
        P1_U3074) );
  AOI22_X1 U23950 ( .A1(n21286), .A2(n20965), .B1(n21285), .B2(n20966), .ZN(
        n20955) );
  AOI22_X1 U23951 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20967), .B1(
        n20996), .B2(n21287), .ZN(n20954) );
  OAI211_X1 U23952 ( .C1(n21292), .C2(n20970), .A(n20955), .B(n20954), .ZN(
        P1_U3075) );
  AOI22_X1 U23953 ( .A1(n21294), .A2(n20965), .B1(n21293), .B2(n20966), .ZN(
        n20957) );
  AOI22_X1 U23954 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20967), .B1(
        n20962), .B2(n21295), .ZN(n20956) );
  OAI211_X1 U23955 ( .C1(n21298), .C2(n20972), .A(n20957), .B(n20956), .ZN(
        P1_U3076) );
  AOI22_X1 U23956 ( .A1(n21300), .A2(n20965), .B1(n21299), .B2(n20966), .ZN(
        n20959) );
  AOI22_X1 U23957 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20967), .B1(
        n20962), .B2(n21301), .ZN(n20958) );
  OAI211_X1 U23958 ( .C1(n21304), .C2(n20972), .A(n20959), .B(n20958), .ZN(
        P1_U3077) );
  AOI22_X1 U23959 ( .A1(n21306), .A2(n20965), .B1(n21305), .B2(n20966), .ZN(
        n20961) );
  AOI22_X1 U23960 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20967), .B1(
        n20962), .B2(n21307), .ZN(n20960) );
  OAI211_X1 U23961 ( .C1(n21310), .C2(n20972), .A(n20961), .B(n20960), .ZN(
        P1_U3078) );
  AOI22_X1 U23962 ( .A1(n21312), .A2(n20965), .B1(n21311), .B2(n20966), .ZN(
        n20964) );
  AOI22_X1 U23963 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20967), .B1(
        n20962), .B2(n21313), .ZN(n20963) );
  OAI211_X1 U23964 ( .C1(n21316), .C2(n20972), .A(n20964), .B(n20963), .ZN(
        P1_U3079) );
  AOI22_X1 U23965 ( .A1(n21320), .A2(n20966), .B1(n21318), .B2(n20965), .ZN(
        n20969) );
  AOI22_X1 U23966 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20967), .B1(
        n20996), .B2(n21191), .ZN(n20968) );
  OAI211_X1 U23967 ( .C1(n21030), .C2(n20970), .A(n20969), .B(n20968), .ZN(
        P1_U3080) );
  INV_X1 U23968 ( .A(n21231), .ZN(n20971) );
  NAND2_X1 U23969 ( .A1(n21029), .A2(n20972), .ZN(n20973) );
  AOI21_X1 U23970 ( .B1(n20973), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21266), 
        .ZN(n20979) );
  NAND2_X1 U23971 ( .A1(n21003), .A2(n14513), .ZN(n20978) );
  INV_X1 U23972 ( .A(n20978), .ZN(n20976) );
  INV_X1 U23973 ( .A(n20974), .ZN(n20975) );
  NAND2_X1 U23974 ( .A1(n21199), .A2(n12779), .ZN(n20977) );
  INV_X1 U23975 ( .A(n20977), .ZN(n20997) );
  AOI22_X1 U23976 ( .A1(n21263), .A2(n20997), .B1(n20996), .B2(n21163), .ZN(
        n20983) );
  AOI22_X1 U23977 ( .A1(n20979), .A2(n20978), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20977), .ZN(n20981) );
  NAND3_X1 U23978 ( .A1(n21236), .A2(n20981), .A3(n20980), .ZN(n20998) );
  AOI22_X1 U23979 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20998), .B1(
        n21021), .B2(n21275), .ZN(n20982) );
  OAI211_X1 U23980 ( .C1(n21001), .C2(n21166), .A(n20983), .B(n20982), .ZN(
        P1_U3081) );
  AOI22_X1 U23981 ( .A1(n21279), .A2(n20997), .B1(n20996), .B2(n21167), .ZN(
        n20985) );
  AOI22_X1 U23982 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20998), .B1(
        n21021), .B2(n21281), .ZN(n20984) );
  OAI211_X1 U23983 ( .C1(n21001), .C2(n21170), .A(n20985), .B(n20984), .ZN(
        P1_U3082) );
  AOI22_X1 U23984 ( .A1(n21285), .A2(n20997), .B1(n20996), .B2(n21171), .ZN(
        n20987) );
  AOI22_X1 U23985 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20998), .B1(
        n21021), .B2(n21287), .ZN(n20986) );
  OAI211_X1 U23986 ( .C1(n21001), .C2(n21174), .A(n20987), .B(n20986), .ZN(
        P1_U3083) );
  AOI22_X1 U23987 ( .A1(n21293), .A2(n20997), .B1(n20996), .B2(n21295), .ZN(
        n20989) );
  AOI22_X1 U23988 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20998), .B1(
        n21021), .B2(n21175), .ZN(n20988) );
  OAI211_X1 U23989 ( .C1(n21001), .C2(n21178), .A(n20989), .B(n20988), .ZN(
        P1_U3084) );
  AOI22_X1 U23990 ( .A1(n21299), .A2(n20997), .B1(n21021), .B2(n21179), .ZN(
        n20991) );
  AOI22_X1 U23991 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20998), .B1(
        n20996), .B2(n21301), .ZN(n20990) );
  OAI211_X1 U23992 ( .C1(n21001), .C2(n21182), .A(n20991), .B(n20990), .ZN(
        P1_U3085) );
  AOI22_X1 U23993 ( .A1(n21305), .A2(n20997), .B1(n21021), .B2(n21183), .ZN(
        n20993) );
  AOI22_X1 U23994 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20998), .B1(
        n20996), .B2(n21307), .ZN(n20992) );
  OAI211_X1 U23995 ( .C1(n21001), .C2(n21186), .A(n20993), .B(n20992), .ZN(
        P1_U3086) );
  AOI22_X1 U23996 ( .A1(n21311), .A2(n20997), .B1(n20996), .B2(n21313), .ZN(
        n20995) );
  AOI22_X1 U23997 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20998), .B1(
        n21021), .B2(n21187), .ZN(n20994) );
  OAI211_X1 U23998 ( .C1(n21001), .C2(n21190), .A(n20995), .B(n20994), .ZN(
        P1_U3087) );
  AOI22_X1 U23999 ( .A1(n21320), .A2(n20997), .B1(n20996), .B2(n21321), .ZN(
        n21000) );
  AOI22_X1 U24000 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20998), .B1(
        n21021), .B2(n21191), .ZN(n20999) );
  OAI211_X1 U24001 ( .C1(n21001), .C2(n21197), .A(n21000), .B(n20999), .ZN(
        P1_U3088) );
  INV_X1 U24002 ( .A(n21002), .ZN(n21025) );
  AOI21_X1 U24003 ( .B1(n21003), .B2(n21260), .A(n21025), .ZN(n21005) );
  OAI22_X1 U24004 ( .A1(n21005), .A2(n21266), .B1(n21004), .B2(n21201), .ZN(
        n21024) );
  AOI22_X1 U24005 ( .A1(n21264), .A2(n21024), .B1(n21025), .B2(n21263), .ZN(
        n21010) );
  INV_X1 U24006 ( .A(n21125), .ZN(n21007) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21026), .B1(
        n21055), .B2(n21275), .ZN(n21009) );
  OAI211_X1 U24008 ( .C1(n21278), .C2(n21029), .A(n21010), .B(n21009), .ZN(
        P1_U3089) );
  AOI22_X1 U24009 ( .A1(n21280), .A2(n21024), .B1(n21025), .B2(n21279), .ZN(
        n21012) );
  AOI22_X1 U24010 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21026), .B1(
        n21055), .B2(n21281), .ZN(n21011) );
  OAI211_X1 U24011 ( .C1(n21284), .C2(n21029), .A(n21012), .B(n21011), .ZN(
        P1_U3090) );
  AOI22_X1 U24012 ( .A1(n21286), .A2(n21024), .B1(n21025), .B2(n21285), .ZN(
        n21014) );
  AOI22_X1 U24013 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21026), .B1(
        n21055), .B2(n21287), .ZN(n21013) );
  OAI211_X1 U24014 ( .C1(n21292), .C2(n21029), .A(n21014), .B(n21013), .ZN(
        P1_U3091) );
  AOI22_X1 U24015 ( .A1(n21294), .A2(n21024), .B1(n21025), .B2(n21293), .ZN(
        n21016) );
  AOI22_X1 U24016 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21026), .B1(
        n21021), .B2(n21295), .ZN(n21015) );
  OAI211_X1 U24017 ( .C1(n21298), .C2(n21044), .A(n21016), .B(n21015), .ZN(
        P1_U3092) );
  AOI22_X1 U24018 ( .A1(n21300), .A2(n21024), .B1(n21025), .B2(n21299), .ZN(
        n21018) );
  AOI22_X1 U24019 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21026), .B1(
        n21021), .B2(n21301), .ZN(n21017) );
  OAI211_X1 U24020 ( .C1(n21304), .C2(n21044), .A(n21018), .B(n21017), .ZN(
        P1_U3093) );
  AOI22_X1 U24021 ( .A1(n21306), .A2(n21024), .B1(n21025), .B2(n21305), .ZN(
        n21020) );
  AOI22_X1 U24022 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21026), .B1(
        n21021), .B2(n21307), .ZN(n21019) );
  OAI211_X1 U24023 ( .C1(n21310), .C2(n21044), .A(n21020), .B(n21019), .ZN(
        P1_U3094) );
  AOI22_X1 U24024 ( .A1(n21312), .A2(n21024), .B1(n21025), .B2(n21311), .ZN(
        n21023) );
  AOI22_X1 U24025 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21026), .B1(
        n21021), .B2(n21313), .ZN(n21022) );
  OAI211_X1 U24026 ( .C1(n21316), .C2(n21044), .A(n21023), .B(n21022), .ZN(
        P1_U3095) );
  AOI22_X1 U24027 ( .A1(n21320), .A2(n21025), .B1(n21318), .B2(n21024), .ZN(
        n21028) );
  AOI22_X1 U24028 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21026), .B1(
        n21055), .B2(n21191), .ZN(n21027) );
  OAI211_X1 U24029 ( .C1(n21030), .C2(n21029), .A(n21028), .B(n21027), .ZN(
        P1_U3096) );
  NAND2_X1 U24030 ( .A1(n21031), .A2(n21152), .ZN(n21086) );
  INV_X1 U24031 ( .A(n21086), .ZN(n21118) );
  NOR3_X1 U24032 ( .A1(n21156), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21062) );
  INV_X1 U24033 ( .A(n21062), .ZN(n21059) );
  NOR2_X1 U24034 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21059), .ZN(
        n21054) );
  AOI21_X1 U24035 ( .B1(n21118), .B2(n21153), .A(n21054), .ZN(n21035) );
  AND2_X1 U24036 ( .A1(n21032), .A2(n21087), .ZN(n21162) );
  INV_X1 U24037 ( .A(n21162), .ZN(n21033) );
  OAI22_X1 U24038 ( .A1(n21035), .A2(n21266), .B1(n21034), .B2(n21033), .ZN(
        n21053) );
  AOI22_X1 U24039 ( .A1(n21264), .A2(n21053), .B1(n21263), .B2(n21054), .ZN(
        n21039) );
  OAI21_X1 U24040 ( .B1(n21080), .B2(n21055), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21036) );
  NAND2_X1 U24041 ( .A1(n21036), .A2(n21035), .ZN(n21037) );
  AOI22_X1 U24042 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21056), .B1(
        n21080), .B2(n21275), .ZN(n21038) );
  OAI211_X1 U24043 ( .C1(n21278), .C2(n21044), .A(n21039), .B(n21038), .ZN(
        P1_U3097) );
  AOI22_X1 U24044 ( .A1(n21280), .A2(n21053), .B1(n21279), .B2(n21054), .ZN(
        n21041) );
  AOI22_X1 U24045 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21056), .B1(
        n21080), .B2(n21281), .ZN(n21040) );
  OAI211_X1 U24046 ( .C1(n21284), .C2(n21044), .A(n21041), .B(n21040), .ZN(
        P1_U3098) );
  AOI22_X1 U24047 ( .A1(n21286), .A2(n21053), .B1(n21285), .B2(n21054), .ZN(
        n21043) );
  AOI22_X1 U24048 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21056), .B1(
        n21080), .B2(n21287), .ZN(n21042) );
  OAI211_X1 U24049 ( .C1(n21292), .C2(n21044), .A(n21043), .B(n21042), .ZN(
        P1_U3099) );
  AOI22_X1 U24050 ( .A1(n21294), .A2(n21053), .B1(n21293), .B2(n21054), .ZN(
        n21046) );
  AOI22_X1 U24051 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21056), .B1(
        n21055), .B2(n21295), .ZN(n21045) );
  OAI211_X1 U24052 ( .C1(n21298), .C2(n21069), .A(n21046), .B(n21045), .ZN(
        P1_U3100) );
  AOI22_X1 U24053 ( .A1(n21300), .A2(n21053), .B1(n21299), .B2(n21054), .ZN(
        n21048) );
  AOI22_X1 U24054 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21056), .B1(
        n21055), .B2(n21301), .ZN(n21047) );
  OAI211_X1 U24055 ( .C1(n21304), .C2(n21069), .A(n21048), .B(n21047), .ZN(
        P1_U3101) );
  AOI22_X1 U24056 ( .A1(n21306), .A2(n21053), .B1(n21305), .B2(n21054), .ZN(
        n21050) );
  AOI22_X1 U24057 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21056), .B1(
        n21055), .B2(n21307), .ZN(n21049) );
  OAI211_X1 U24058 ( .C1(n21310), .C2(n21069), .A(n21050), .B(n21049), .ZN(
        P1_U3102) );
  AOI22_X1 U24059 ( .A1(n21312), .A2(n21053), .B1(n21311), .B2(n21054), .ZN(
        n21052) );
  AOI22_X1 U24060 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21056), .B1(
        n21055), .B2(n21313), .ZN(n21051) );
  OAI211_X1 U24061 ( .C1(n21316), .C2(n21069), .A(n21052), .B(n21051), .ZN(
        P1_U3103) );
  AOI22_X1 U24062 ( .A1(n21320), .A2(n21054), .B1(n21318), .B2(n21053), .ZN(
        n21058) );
  AOI22_X1 U24063 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21056), .B1(
        n21055), .B2(n21321), .ZN(n21057) );
  OAI211_X1 U24064 ( .C1(n21327), .C2(n21069), .A(n21058), .B(n21057), .ZN(
        P1_U3104) );
  NOR2_X1 U24065 ( .A1(n21199), .A2(n21059), .ZN(n21079) );
  AOI21_X1 U24066 ( .B1(n21118), .B2(n21200), .A(n21079), .ZN(n21060) );
  OAI22_X1 U24067 ( .A1(n21060), .A2(n21266), .B1(n21059), .B2(n21201), .ZN(
        n21078) );
  AOI22_X1 U24068 ( .A1(n21264), .A2(n21078), .B1(n21263), .B2(n21079), .ZN(
        n21064) );
  OAI211_X1 U24069 ( .C1(n21126), .C2(n21232), .A(n21273), .B(n21060), .ZN(
        n21061) );
  OAI211_X1 U24070 ( .C1(n21273), .C2(n21062), .A(n21272), .B(n21061), .ZN(
        n21081) );
  AOI22_X1 U24071 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21081), .B1(
        n21111), .B2(n21275), .ZN(n21063) );
  OAI211_X1 U24072 ( .C1(n21278), .C2(n21069), .A(n21064), .B(n21063), .ZN(
        P1_U3105) );
  AOI22_X1 U24073 ( .A1(n21280), .A2(n21078), .B1(n21279), .B2(n21079), .ZN(
        n21066) );
  AOI22_X1 U24074 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21081), .B1(
        n21111), .B2(n21281), .ZN(n21065) );
  OAI211_X1 U24075 ( .C1(n21284), .C2(n21069), .A(n21066), .B(n21065), .ZN(
        P1_U3106) );
  AOI22_X1 U24076 ( .A1(n21286), .A2(n21078), .B1(n21285), .B2(n21079), .ZN(
        n21068) );
  AOI22_X1 U24077 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21081), .B1(
        n21111), .B2(n21287), .ZN(n21067) );
  OAI211_X1 U24078 ( .C1(n21292), .C2(n21069), .A(n21068), .B(n21067), .ZN(
        P1_U3107) );
  AOI22_X1 U24079 ( .A1(n21294), .A2(n21078), .B1(n21293), .B2(n21079), .ZN(
        n21071) );
  AOI22_X1 U24080 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21081), .B1(
        n21080), .B2(n21295), .ZN(n21070) );
  OAI211_X1 U24081 ( .C1(n21298), .C2(n21084), .A(n21071), .B(n21070), .ZN(
        P1_U3108) );
  AOI22_X1 U24082 ( .A1(n21300), .A2(n21078), .B1(n21299), .B2(n21079), .ZN(
        n21073) );
  AOI22_X1 U24083 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21081), .B1(
        n21080), .B2(n21301), .ZN(n21072) );
  OAI211_X1 U24084 ( .C1(n21304), .C2(n21084), .A(n21073), .B(n21072), .ZN(
        P1_U3109) );
  AOI22_X1 U24085 ( .A1(n21306), .A2(n21078), .B1(n21305), .B2(n21079), .ZN(
        n21075) );
  AOI22_X1 U24086 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21081), .B1(
        n21080), .B2(n21307), .ZN(n21074) );
  OAI211_X1 U24087 ( .C1(n21310), .C2(n21084), .A(n21075), .B(n21074), .ZN(
        P1_U3110) );
  AOI22_X1 U24088 ( .A1(n21312), .A2(n21078), .B1(n21311), .B2(n21079), .ZN(
        n21077) );
  AOI22_X1 U24089 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21081), .B1(
        n21080), .B2(n21313), .ZN(n21076) );
  OAI211_X1 U24090 ( .C1(n21316), .C2(n21084), .A(n21077), .B(n21076), .ZN(
        P1_U3111) );
  AOI22_X1 U24091 ( .A1(n21320), .A2(n21079), .B1(n21318), .B2(n21078), .ZN(
        n21083) );
  AOI22_X1 U24092 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21081), .B1(
        n21080), .B2(n21321), .ZN(n21082) );
  OAI211_X1 U24093 ( .C1(n21327), .C2(n21084), .A(n21083), .B(n21082), .ZN(
        P1_U3112) );
  NAND2_X1 U24094 ( .A1(n21133), .A2(n21084), .ZN(n21085) );
  AOI21_X1 U24095 ( .B1(n21085), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21266), 
        .ZN(n21094) );
  OR2_X1 U24096 ( .A1(n21086), .A2(n21153), .ZN(n21093) );
  INV_X1 U24097 ( .A(n21093), .ZN(n21090) );
  OR2_X1 U24098 ( .A1(n21087), .A2(n21156), .ZN(n21229) );
  INV_X1 U24099 ( .A(n21229), .ZN(n21088) );
  NOR3_X1 U24100 ( .A1(n21156), .A2(n13362), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21124) );
  INV_X1 U24101 ( .A(n21124), .ZN(n21119) );
  NOR2_X1 U24102 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21119), .ZN(
        n21112) );
  AOI22_X1 U24103 ( .A1(n21263), .A2(n21112), .B1(n21111), .B2(n21163), .ZN(
        n21098) );
  NOR2_X1 U24104 ( .A1(n21112), .A2(n21091), .ZN(n21092) );
  AOI21_X1 U24105 ( .B1(n21094), .B2(n21093), .A(n21092), .ZN(n21095) );
  NAND2_X1 U24106 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21229), .ZN(n21235) );
  NAND3_X1 U24107 ( .A1(n21096), .A2(n21095), .A3(n21235), .ZN(n21113) );
  AOI22_X1 U24108 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21113), .B1(
        n21144), .B2(n21275), .ZN(n21097) );
  OAI211_X1 U24109 ( .C1(n21116), .C2(n21166), .A(n21098), .B(n21097), .ZN(
        P1_U3113) );
  AOI22_X1 U24110 ( .A1(n21279), .A2(n21112), .B1(n21144), .B2(n21281), .ZN(
        n21100) );
  AOI22_X1 U24111 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21113), .B1(
        n21111), .B2(n21167), .ZN(n21099) );
  OAI211_X1 U24112 ( .C1(n21116), .C2(n21170), .A(n21100), .B(n21099), .ZN(
        P1_U3114) );
  AOI22_X1 U24113 ( .A1(n21285), .A2(n21112), .B1(n21111), .B2(n21171), .ZN(
        n21102) );
  AOI22_X1 U24114 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21113), .B1(
        n21144), .B2(n21287), .ZN(n21101) );
  OAI211_X1 U24115 ( .C1(n21116), .C2(n21174), .A(n21102), .B(n21101), .ZN(
        P1_U3115) );
  AOI22_X1 U24116 ( .A1(n21293), .A2(n21112), .B1(n21144), .B2(n21175), .ZN(
        n21104) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21113), .B1(
        n21111), .B2(n21295), .ZN(n21103) );
  OAI211_X1 U24118 ( .C1(n21116), .C2(n21178), .A(n21104), .B(n21103), .ZN(
        P1_U3116) );
  AOI22_X1 U24119 ( .A1(n21299), .A2(n21112), .B1(n21144), .B2(n21179), .ZN(
        n21106) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21113), .B1(
        n21111), .B2(n21301), .ZN(n21105) );
  OAI211_X1 U24121 ( .C1(n21116), .C2(n21182), .A(n21106), .B(n21105), .ZN(
        P1_U3117) );
  AOI22_X1 U24122 ( .A1(n21305), .A2(n21112), .B1(n21144), .B2(n21183), .ZN(
        n21108) );
  AOI22_X1 U24123 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21113), .B1(
        n21111), .B2(n21307), .ZN(n21107) );
  OAI211_X1 U24124 ( .C1(n21116), .C2(n21186), .A(n21108), .B(n21107), .ZN(
        P1_U3118) );
  AOI22_X1 U24125 ( .A1(n21311), .A2(n21112), .B1(n21144), .B2(n21187), .ZN(
        n21110) );
  AOI22_X1 U24126 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21113), .B1(
        n21111), .B2(n21313), .ZN(n21109) );
  OAI211_X1 U24127 ( .C1(n21116), .C2(n21190), .A(n21110), .B(n21109), .ZN(
        P1_U3119) );
  AOI22_X1 U24128 ( .A1(n21320), .A2(n21112), .B1(n21111), .B2(n21321), .ZN(
        n21115) );
  AOI22_X1 U24129 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21113), .B1(
        n21144), .B2(n21191), .ZN(n21114) );
  OAI211_X1 U24130 ( .C1(n21116), .C2(n21197), .A(n21115), .B(n21114), .ZN(
        P1_U3120) );
  NOR2_X1 U24131 ( .A1(n21117), .A2(n21156), .ZN(n21143) );
  AOI21_X1 U24132 ( .B1(n21118), .B2(n21260), .A(n21143), .ZN(n21121) );
  OAI22_X1 U24133 ( .A1(n21121), .A2(n21266), .B1(n21119), .B2(n21201), .ZN(
        n21142) );
  AOI22_X1 U24134 ( .A1(n21264), .A2(n21142), .B1(n21263), .B2(n21143), .ZN(
        n21128) );
  INV_X1 U24135 ( .A(n21126), .ZN(n21120) );
  NOR2_X1 U24136 ( .A1(n21120), .A2(n21266), .ZN(n21122) );
  OAI21_X1 U24137 ( .B1(n21270), .B2(n21122), .A(n21121), .ZN(n21123) );
  OAI211_X1 U24138 ( .C1(n21273), .C2(n21124), .A(n21272), .B(n21123), .ZN(
        n21145) );
  AOI22_X1 U24139 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21145), .B1(
        n21193), .B2(n21275), .ZN(n21127) );
  OAI211_X1 U24140 ( .C1(n21278), .C2(n21133), .A(n21128), .B(n21127), .ZN(
        P1_U3121) );
  AOI22_X1 U24141 ( .A1(n21280), .A2(n21142), .B1(n21279), .B2(n21143), .ZN(
        n21130) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21145), .B1(
        n21193), .B2(n21281), .ZN(n21129) );
  OAI211_X1 U24143 ( .C1(n21284), .C2(n21133), .A(n21130), .B(n21129), .ZN(
        P1_U3122) );
  AOI22_X1 U24144 ( .A1(n21286), .A2(n21142), .B1(n21285), .B2(n21143), .ZN(
        n21132) );
  AOI22_X1 U24145 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21145), .B1(
        n21193), .B2(n21287), .ZN(n21131) );
  OAI211_X1 U24146 ( .C1(n21292), .C2(n21133), .A(n21132), .B(n21131), .ZN(
        P1_U3123) );
  AOI22_X1 U24147 ( .A1(n21294), .A2(n21142), .B1(n21293), .B2(n21143), .ZN(
        n21135) );
  AOI22_X1 U24148 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n21295), .ZN(n21134) );
  OAI211_X1 U24149 ( .C1(n21298), .C2(n21149), .A(n21135), .B(n21134), .ZN(
        P1_U3124) );
  AOI22_X1 U24150 ( .A1(n21300), .A2(n21142), .B1(n21299), .B2(n21143), .ZN(
        n21137) );
  AOI22_X1 U24151 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n21301), .ZN(n21136) );
  OAI211_X1 U24152 ( .C1(n21304), .C2(n21149), .A(n21137), .B(n21136), .ZN(
        P1_U3125) );
  AOI22_X1 U24153 ( .A1(n21306), .A2(n21142), .B1(n21305), .B2(n21143), .ZN(
        n21139) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n21307), .ZN(n21138) );
  OAI211_X1 U24155 ( .C1(n21310), .C2(n21149), .A(n21139), .B(n21138), .ZN(
        P1_U3126) );
  AOI22_X1 U24156 ( .A1(n21312), .A2(n21142), .B1(n21311), .B2(n21143), .ZN(
        n21141) );
  AOI22_X1 U24157 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n21313), .ZN(n21140) );
  OAI211_X1 U24158 ( .C1(n21316), .C2(n21149), .A(n21141), .B(n21140), .ZN(
        P1_U3127) );
  AOI22_X1 U24159 ( .A1(n21320), .A2(n21143), .B1(n21318), .B2(n21142), .ZN(
        n21147) );
  AOI22_X1 U24160 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n21321), .ZN(n21146) );
  OAI211_X1 U24161 ( .C1(n21327), .C2(n21149), .A(n21147), .B(n21146), .ZN(
        P1_U3128) );
  NAND2_X1 U24162 ( .A1(n21149), .A2(n21213), .ZN(n21150) );
  AOI21_X1 U24163 ( .B1(n21150), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21266), 
        .ZN(n21160) );
  NAND2_X1 U24164 ( .A1(n21261), .A2(n21153), .ZN(n21159) );
  INV_X1 U24165 ( .A(n21159), .ZN(n21155) );
  NOR3_X1 U24166 ( .A1(n21157), .A2(n21156), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21205) );
  NAND2_X1 U24167 ( .A1(n21199), .A2(n21205), .ZN(n21158) );
  INV_X1 U24168 ( .A(n21158), .ZN(n21192) );
  AOI22_X1 U24169 ( .A1(n21263), .A2(n21192), .B1(n21224), .B2(n21275), .ZN(
        n21165) );
  AOI22_X1 U24170 ( .A1(n21160), .A2(n21159), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21158), .ZN(n21161) );
  AOI22_X1 U24171 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21163), .ZN(n21164) );
  OAI211_X1 U24172 ( .C1(n21198), .C2(n21166), .A(n21165), .B(n21164), .ZN(
        P1_U3129) );
  AOI22_X1 U24173 ( .A1(n21279), .A2(n21192), .B1(n21224), .B2(n21281), .ZN(
        n21169) );
  AOI22_X1 U24174 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21167), .ZN(n21168) );
  OAI211_X1 U24175 ( .C1(n21198), .C2(n21170), .A(n21169), .B(n21168), .ZN(
        P1_U3130) );
  AOI22_X1 U24176 ( .A1(n21285), .A2(n21192), .B1(n21224), .B2(n21287), .ZN(
        n21173) );
  AOI22_X1 U24177 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21171), .ZN(n21172) );
  OAI211_X1 U24178 ( .C1(n21198), .C2(n21174), .A(n21173), .B(n21172), .ZN(
        P1_U3131) );
  AOI22_X1 U24179 ( .A1(n21293), .A2(n21192), .B1(n21224), .B2(n21175), .ZN(
        n21177) );
  AOI22_X1 U24180 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21295), .ZN(n21176) );
  OAI211_X1 U24181 ( .C1(n21198), .C2(n21178), .A(n21177), .B(n21176), .ZN(
        P1_U3132) );
  AOI22_X1 U24182 ( .A1(n21299), .A2(n21192), .B1(n21224), .B2(n21179), .ZN(
        n21181) );
  AOI22_X1 U24183 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21301), .ZN(n21180) );
  OAI211_X1 U24184 ( .C1(n21198), .C2(n21182), .A(n21181), .B(n21180), .ZN(
        P1_U3133) );
  AOI22_X1 U24185 ( .A1(n21305), .A2(n21192), .B1(n21224), .B2(n21183), .ZN(
        n21185) );
  AOI22_X1 U24186 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21307), .ZN(n21184) );
  OAI211_X1 U24187 ( .C1(n21198), .C2(n21186), .A(n21185), .B(n21184), .ZN(
        P1_U3134) );
  AOI22_X1 U24188 ( .A1(n21311), .A2(n21192), .B1(n21224), .B2(n21187), .ZN(
        n21189) );
  AOI22_X1 U24189 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21313), .ZN(n21188) );
  OAI211_X1 U24190 ( .C1(n21198), .C2(n21190), .A(n21189), .B(n21188), .ZN(
        P1_U3135) );
  AOI22_X1 U24191 ( .A1(n21320), .A2(n21192), .B1(n21224), .B2(n21191), .ZN(
        n21196) );
  AOI22_X1 U24192 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21194), .B1(
        n21193), .B2(n21321), .ZN(n21195) );
  OAI211_X1 U24193 ( .C1(n21198), .C2(n21197), .A(n21196), .B(n21195), .ZN(
        P1_U3136) );
  INV_X1 U24194 ( .A(n21205), .ZN(n21202) );
  NOR2_X1 U24195 ( .A1(n21199), .A2(n21202), .ZN(n21223) );
  AOI21_X1 U24196 ( .B1(n21261), .B2(n21200), .A(n21223), .ZN(n21203) );
  OAI22_X1 U24197 ( .A1(n21203), .A2(n21266), .B1(n21202), .B2(n21201), .ZN(
        n21222) );
  AOI22_X1 U24198 ( .A1(n21264), .A2(n21222), .B1(n21263), .B2(n21223), .ZN(
        n21208) );
  OAI211_X1 U24199 ( .C1(n21265), .C2(n21232), .A(n21273), .B(n21203), .ZN(
        n21204) );
  OAI211_X1 U24200 ( .C1(n21273), .C2(n21205), .A(n21272), .B(n21204), .ZN(
        n21225) );
  AOI22_X1 U24201 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21225), .B1(
        n21255), .B2(n21275), .ZN(n21207) );
  OAI211_X1 U24202 ( .C1(n21278), .C2(n21213), .A(n21208), .B(n21207), .ZN(
        P1_U3137) );
  AOI22_X1 U24203 ( .A1(n21280), .A2(n21222), .B1(n21279), .B2(n21223), .ZN(
        n21210) );
  AOI22_X1 U24204 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21225), .B1(
        n21255), .B2(n21281), .ZN(n21209) );
  OAI211_X1 U24205 ( .C1(n21284), .C2(n21213), .A(n21210), .B(n21209), .ZN(
        P1_U3138) );
  AOI22_X1 U24206 ( .A1(n21286), .A2(n21222), .B1(n21285), .B2(n21223), .ZN(
        n21212) );
  AOI22_X1 U24207 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21225), .B1(
        n21255), .B2(n21287), .ZN(n21211) );
  OAI211_X1 U24208 ( .C1(n21292), .C2(n21213), .A(n21212), .B(n21211), .ZN(
        P1_U3139) );
  AOI22_X1 U24209 ( .A1(n21294), .A2(n21222), .B1(n21293), .B2(n21223), .ZN(
        n21215) );
  AOI22_X1 U24210 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21295), .ZN(n21214) );
  OAI211_X1 U24211 ( .C1(n21298), .C2(n21244), .A(n21215), .B(n21214), .ZN(
        P1_U3140) );
  AOI22_X1 U24212 ( .A1(n21300), .A2(n21222), .B1(n21299), .B2(n21223), .ZN(
        n21217) );
  AOI22_X1 U24213 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21301), .ZN(n21216) );
  OAI211_X1 U24214 ( .C1(n21304), .C2(n21244), .A(n21217), .B(n21216), .ZN(
        P1_U3141) );
  AOI22_X1 U24215 ( .A1(n21306), .A2(n21222), .B1(n21305), .B2(n21223), .ZN(
        n21219) );
  AOI22_X1 U24216 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21307), .ZN(n21218) );
  OAI211_X1 U24217 ( .C1(n21310), .C2(n21244), .A(n21219), .B(n21218), .ZN(
        P1_U3142) );
  AOI22_X1 U24218 ( .A1(n21312), .A2(n21222), .B1(n21311), .B2(n21223), .ZN(
        n21221) );
  AOI22_X1 U24219 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21313), .ZN(n21220) );
  OAI211_X1 U24220 ( .C1(n21316), .C2(n21244), .A(n21221), .B(n21220), .ZN(
        P1_U3143) );
  AOI22_X1 U24221 ( .A1(n21320), .A2(n21223), .B1(n21318), .B2(n21222), .ZN(
        n21227) );
  AOI22_X1 U24222 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21321), .ZN(n21226) );
  OAI211_X1 U24223 ( .C1(n21327), .C2(n21244), .A(n21227), .B(n21226), .ZN(
        P1_U3144) );
  NAND3_X1 U24224 ( .A1(n21261), .A2(n14513), .A3(n21273), .ZN(n21228) );
  OAI21_X1 U24225 ( .B1(n21230), .B2(n21229), .A(n21228), .ZN(n21253) );
  INV_X1 U24226 ( .A(n21274), .ZN(n21262) );
  NOR2_X1 U24227 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21262), .ZN(
        n21254) );
  AOI22_X1 U24228 ( .A1(n21264), .A2(n21253), .B1(n21263), .B2(n21254), .ZN(
        n21239) );
  AOI21_X1 U24229 ( .B1(n21291), .B2(n21244), .A(n21232), .ZN(n21233) );
  AOI21_X1 U24230 ( .B1(n21261), .B2(n14513), .A(n21233), .ZN(n21234) );
  NOR2_X1 U24231 ( .A1(n21234), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21237) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21256), .B1(
        n21322), .B2(n21275), .ZN(n21238) );
  OAI211_X1 U24233 ( .C1(n21278), .C2(n21244), .A(n21239), .B(n21238), .ZN(
        P1_U3145) );
  AOI22_X1 U24234 ( .A1(n21280), .A2(n21253), .B1(n21279), .B2(n21254), .ZN(
        n21241) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21256), .B1(
        n21322), .B2(n21281), .ZN(n21240) );
  OAI211_X1 U24236 ( .C1(n21284), .C2(n21244), .A(n21241), .B(n21240), .ZN(
        P1_U3146) );
  AOI22_X1 U24237 ( .A1(n21286), .A2(n21253), .B1(n21285), .B2(n21254), .ZN(
        n21243) );
  AOI22_X1 U24238 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21256), .B1(
        n21322), .B2(n21287), .ZN(n21242) );
  OAI211_X1 U24239 ( .C1(n21292), .C2(n21244), .A(n21243), .B(n21242), .ZN(
        P1_U3147) );
  AOI22_X1 U24240 ( .A1(n21294), .A2(n21253), .B1(n21293), .B2(n21254), .ZN(
        n21246) );
  AOI22_X1 U24241 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21256), .B1(
        n21255), .B2(n21295), .ZN(n21245) );
  OAI211_X1 U24242 ( .C1(n21298), .C2(n21291), .A(n21246), .B(n21245), .ZN(
        P1_U3148) );
  AOI22_X1 U24243 ( .A1(n21300), .A2(n21253), .B1(n21299), .B2(n21254), .ZN(
        n21248) );
  AOI22_X1 U24244 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21256), .B1(
        n21255), .B2(n21301), .ZN(n21247) );
  OAI211_X1 U24245 ( .C1(n21304), .C2(n21291), .A(n21248), .B(n21247), .ZN(
        P1_U3149) );
  AOI22_X1 U24246 ( .A1(n21306), .A2(n21253), .B1(n21305), .B2(n21254), .ZN(
        n21250) );
  AOI22_X1 U24247 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21256), .B1(
        n21255), .B2(n21307), .ZN(n21249) );
  OAI211_X1 U24248 ( .C1(n21310), .C2(n21291), .A(n21250), .B(n21249), .ZN(
        P1_U3150) );
  AOI22_X1 U24249 ( .A1(n21312), .A2(n21253), .B1(n21311), .B2(n21254), .ZN(
        n21252) );
  AOI22_X1 U24250 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21256), .B1(
        n21255), .B2(n21313), .ZN(n21251) );
  OAI211_X1 U24251 ( .C1(n21316), .C2(n21291), .A(n21252), .B(n21251), .ZN(
        P1_U3151) );
  AOI22_X1 U24252 ( .A1(n21320), .A2(n21254), .B1(n21318), .B2(n21253), .ZN(
        n21258) );
  AOI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21256), .B1(
        n21255), .B2(n21321), .ZN(n21257) );
  OAI211_X1 U24254 ( .C1(n21327), .C2(n21291), .A(n21258), .B(n21257), .ZN(
        P1_U3152) );
  INV_X1 U24255 ( .A(n21259), .ZN(n21319) );
  AOI21_X1 U24256 ( .B1(n21261), .B2(n21260), .A(n21319), .ZN(n21268) );
  OAI22_X1 U24257 ( .A1(n21268), .A2(n21266), .B1(n21201), .B2(n21262), .ZN(
        n21317) );
  AOI22_X1 U24258 ( .A1(n21264), .A2(n21317), .B1(n21319), .B2(n21263), .ZN(
        n21277) );
  INV_X1 U24259 ( .A(n21265), .ZN(n21267) );
  NOR2_X1 U24260 ( .A1(n21267), .A2(n21266), .ZN(n21269) );
  OAI21_X1 U24261 ( .B1(n21270), .B2(n21269), .A(n21268), .ZN(n21271) );
  OAI211_X1 U24262 ( .C1(n21274), .C2(n21273), .A(n21272), .B(n21271), .ZN(
        n21323) );
  AOI22_X1 U24263 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21323), .B1(
        n21288), .B2(n21275), .ZN(n21276) );
  OAI211_X1 U24264 ( .C1(n21278), .C2(n21291), .A(n21277), .B(n21276), .ZN(
        P1_U3153) );
  AOI22_X1 U24265 ( .A1(n21280), .A2(n21317), .B1(n21319), .B2(n21279), .ZN(
        n21283) );
  AOI22_X1 U24266 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21323), .B1(
        n21288), .B2(n21281), .ZN(n21282) );
  OAI211_X1 U24267 ( .C1(n21284), .C2(n21291), .A(n21283), .B(n21282), .ZN(
        P1_U3154) );
  AOI22_X1 U24268 ( .A1(n21286), .A2(n21317), .B1(n21319), .B2(n21285), .ZN(
        n21290) );
  AOI22_X1 U24269 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21323), .B1(
        n21288), .B2(n21287), .ZN(n21289) );
  OAI211_X1 U24270 ( .C1(n21292), .C2(n21291), .A(n21290), .B(n21289), .ZN(
        P1_U3155) );
  AOI22_X1 U24271 ( .A1(n21294), .A2(n21317), .B1(n21319), .B2(n21293), .ZN(
        n21297) );
  AOI22_X1 U24272 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21323), .B1(
        n21322), .B2(n21295), .ZN(n21296) );
  OAI211_X1 U24273 ( .C1(n21298), .C2(n21326), .A(n21297), .B(n21296), .ZN(
        P1_U3156) );
  AOI22_X1 U24274 ( .A1(n21300), .A2(n21317), .B1(n21319), .B2(n21299), .ZN(
        n21303) );
  AOI22_X1 U24275 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21323), .B1(
        n21322), .B2(n21301), .ZN(n21302) );
  OAI211_X1 U24276 ( .C1(n21304), .C2(n21326), .A(n21303), .B(n21302), .ZN(
        P1_U3157) );
  AOI22_X1 U24277 ( .A1(n21306), .A2(n21317), .B1(n21319), .B2(n21305), .ZN(
        n21309) );
  AOI22_X1 U24278 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21323), .B1(
        n21322), .B2(n21307), .ZN(n21308) );
  OAI211_X1 U24279 ( .C1(n21310), .C2(n21326), .A(n21309), .B(n21308), .ZN(
        P1_U3158) );
  AOI22_X1 U24280 ( .A1(n21312), .A2(n21317), .B1(n21319), .B2(n21311), .ZN(
        n21315) );
  AOI22_X1 U24281 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21323), .B1(
        n21322), .B2(n21313), .ZN(n21314) );
  OAI211_X1 U24282 ( .C1(n21316), .C2(n21326), .A(n21315), .B(n21314), .ZN(
        P1_U3159) );
  AOI22_X1 U24283 ( .A1(n21320), .A2(n21319), .B1(n21318), .B2(n21317), .ZN(
        n21325) );
  AOI22_X1 U24284 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21323), .B1(
        n21322), .B2(n21321), .ZN(n21324) );
  OAI211_X1 U24285 ( .C1(n21327), .C2(n21326), .A(n21325), .B(n21324), .ZN(
        P1_U3160) );
  AOI21_X1 U24286 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n17176), .A(n21328), 
        .ZN(n21330) );
  NAND2_X1 U24287 ( .A1(n21330), .A2(n21329), .ZN(P1_U3163) );
  AND2_X1 U24288 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21331), .ZN(
        P1_U3164) );
  AND2_X1 U24289 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21331), .ZN(
        P1_U3165) );
  AND2_X1 U24290 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21331), .ZN(
        P1_U3166) );
  AND2_X1 U24291 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21331), .ZN(
        P1_U3167) );
  AND2_X1 U24292 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21331), .ZN(
        P1_U3168) );
  AND2_X1 U24293 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21331), .ZN(
        P1_U3169) );
  AND2_X1 U24294 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21331), .ZN(
        P1_U3170) );
  AND2_X1 U24295 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21331), .ZN(
        P1_U3171) );
  AND2_X1 U24296 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21331), .ZN(
        P1_U3172) );
  AND2_X1 U24297 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21331), .ZN(
        P1_U3173) );
  AND2_X1 U24298 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21331), .ZN(
        P1_U3174) );
  AND2_X1 U24299 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21331), .ZN(
        P1_U3175) );
  AND2_X1 U24300 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21331), .ZN(
        P1_U3176) );
  AND2_X1 U24301 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21331), .ZN(
        P1_U3177) );
  AND2_X1 U24302 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21331), .ZN(
        P1_U3178) );
  AND2_X1 U24303 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21331), .ZN(
        P1_U3179) );
  AND2_X1 U24304 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21331), .ZN(
        P1_U3180) );
  AND2_X1 U24305 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21331), .ZN(
        P1_U3181) );
  AND2_X1 U24306 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21331), .ZN(
        P1_U3182) );
  AND2_X1 U24307 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21331), .ZN(
        P1_U3183) );
  AND2_X1 U24308 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21331), .ZN(
        P1_U3184) );
  AND2_X1 U24309 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21331), .ZN(
        P1_U3185) );
  AND2_X1 U24310 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21331), .ZN(P1_U3186) );
  AND2_X1 U24311 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21331), .ZN(P1_U3187) );
  AND2_X1 U24312 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21331), .ZN(P1_U3188) );
  INV_X1 U24313 ( .A(P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n21562) );
  NOR2_X1 U24314 ( .A1(n21397), .A2(n21562), .ZN(P1_U3189) );
  AND2_X1 U24315 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21331), .ZN(P1_U3190) );
  AND2_X1 U24316 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21331), .ZN(P1_U3191) );
  AND2_X1 U24317 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21331), .ZN(P1_U3192) );
  AND2_X1 U24318 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21331), .ZN(P1_U3193) );
  AOI21_X1 U24319 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21341), .A(n21332), 
        .ZN(n21338) );
  NOR2_X1 U24320 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21334) );
  NAND2_X1 U24321 ( .A1(n21332), .A2(NA), .ZN(n21333) );
  OAI211_X1 U24322 ( .C1(n21335), .C2(n21334), .A(n21333), .B(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21336) );
  INV_X1 U24323 ( .A(n21336), .ZN(n21337) );
  OAI22_X1 U24324 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21338), .B1(n21392), 
        .B2(n21337), .ZN(P1_U3194) );
  NAND3_X1 U24325 ( .A1(n21341), .A2(P1_STATE_REG_1__SCAN_IN), .A3(n21340), 
        .ZN(n21346) );
  INV_X1 U24326 ( .A(n21338), .ZN(n21339) );
  OAI211_X1 U24327 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21340), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21339), .ZN(n21345) );
  NAND2_X1 U24328 ( .A1(n21341), .A2(n21340), .ZN(n21342) );
  OAI221_X1 U24329 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n21342), .A(n21637), .ZN(n21343) );
  NAND3_X1 U24330 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n21343), .ZN(
        n21344) );
  OAI211_X1 U24331 ( .C1(n21347), .C2(n21346), .A(n21345), .B(n21344), .ZN(
        P1_U3196) );
  OR2_X1 U24332 ( .A1(n21380), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21389) );
  INV_X1 U24333 ( .A(n21389), .ZN(n21383) );
  NOR2_X1 U24334 ( .A1(n21637), .A2(n21380), .ZN(n21381) );
  AOI222_X1 U24335 ( .A1(n21383), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21387), .ZN(n21348) );
  INV_X1 U24336 ( .A(n21348), .ZN(P1_U3197) );
  AOI22_X1 U24337 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21380), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n21383), .ZN(n21349) );
  OAI21_X1 U24338 ( .B1(n21350), .B2(n21385), .A(n21349), .ZN(P1_U3198) );
  AOI222_X1 U24339 ( .A1(n21387), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21383), .ZN(n21351) );
  INV_X1 U24340 ( .A(n21351), .ZN(P1_U3199) );
  AOI22_X1 U24341 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n21380), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21383), .ZN(n21352) );
  OAI21_X1 U24342 ( .B1(n21353), .B2(n21385), .A(n21352), .ZN(P1_U3200) );
  AOI22_X1 U24343 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21380), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21387), .ZN(n21354) );
  OAI21_X1 U24344 ( .B1(n21355), .B2(n21389), .A(n21354), .ZN(P1_U3201) );
  AOI222_X1 U24345 ( .A1(n21383), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21387), .ZN(n21356) );
  INV_X1 U24346 ( .A(n21356), .ZN(P1_U3202) );
  AOI222_X1 U24347 ( .A1(n21381), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21383), .ZN(n21357) );
  INV_X1 U24348 ( .A(n21357), .ZN(P1_U3203) );
  AOI222_X1 U24349 ( .A1(n21383), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21387), .ZN(n21358) );
  INV_X1 U24350 ( .A(n21358), .ZN(P1_U3204) );
  AOI222_X1 U24351 ( .A1(n21381), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21383), .ZN(n21359) );
  INV_X1 U24352 ( .A(n21359), .ZN(P1_U3205) );
  AOI222_X1 U24353 ( .A1(n21383), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21387), .ZN(n21360) );
  INV_X1 U24354 ( .A(n21360), .ZN(P1_U3206) );
  AOI222_X1 U24355 ( .A1(n21381), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21383), .ZN(n21361) );
  INV_X1 U24356 ( .A(n21361), .ZN(P1_U3207) );
  AOI222_X1 U24357 ( .A1(n21381), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21383), .ZN(n21362) );
  INV_X1 U24358 ( .A(n21362), .ZN(P1_U3208) );
  AOI222_X1 U24359 ( .A1(n21381), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21383), .ZN(n21363) );
  INV_X1 U24360 ( .A(n21363), .ZN(P1_U3209) );
  AOI222_X1 U24361 ( .A1(n21383), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21387), .ZN(n21364) );
  INV_X1 U24362 ( .A(n21364), .ZN(P1_U3210) );
  AOI222_X1 U24363 ( .A1(n21387), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21383), .ZN(n21365) );
  INV_X1 U24364 ( .A(n21365), .ZN(P1_U3211) );
  INV_X1 U24365 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21716) );
  INV_X1 U24366 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21366) );
  OAI222_X1 U24367 ( .A1(n21385), .A2(n21367), .B1(n21716), .B2(n21392), .C1(
        n21366), .C2(n21389), .ZN(P1_U3212) );
  AOI222_X1 U24368 ( .A1(n21387), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n21383), .ZN(n21368) );
  INV_X1 U24369 ( .A(n21368), .ZN(P1_U3213) );
  INV_X1 U24370 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21719) );
  OAI222_X1 U24371 ( .A1(n21385), .A2(n21369), .B1(n21719), .B2(n21392), .C1(
        n21571), .C2(n21389), .ZN(P1_U3214) );
  AOI222_X1 U24372 ( .A1(n21383), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21387), .ZN(n21370) );
  INV_X1 U24373 ( .A(n21370), .ZN(P1_U3215) );
  AOI222_X1 U24374 ( .A1(n21387), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21383), .ZN(n21371) );
  INV_X1 U24375 ( .A(n21371), .ZN(P1_U3216) );
  AOI222_X1 U24376 ( .A1(n21387), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21383), .ZN(n21372) );
  INV_X1 U24377 ( .A(n21372), .ZN(P1_U3217) );
  INV_X1 U24378 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21706) );
  OAI222_X1 U24379 ( .A1(n21385), .A2(n21374), .B1(n21706), .B2(n21392), .C1(
        n21373), .C2(n21389), .ZN(P1_U3218) );
  AOI222_X1 U24380 ( .A1(n21383), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21387), .ZN(n21375) );
  INV_X1 U24381 ( .A(n21375), .ZN(P1_U3219) );
  AOI222_X1 U24382 ( .A1(n21387), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21383), .ZN(n21376) );
  INV_X1 U24383 ( .A(n21376), .ZN(P1_U3220) );
  AOI222_X1 U24384 ( .A1(n21387), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21383), .ZN(n21377) );
  INV_X1 U24385 ( .A(n21377), .ZN(P1_U3221) );
  AOI222_X1 U24386 ( .A1(n21381), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21383), .ZN(n21378) );
  INV_X1 U24387 ( .A(n21378), .ZN(P1_U3222) );
  AOI222_X1 U24388 ( .A1(n21381), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21383), .ZN(n21379) );
  INV_X1 U24389 ( .A(n21379), .ZN(P1_U3223) );
  AOI222_X1 U24390 ( .A1(n21381), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21380), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21383), .ZN(n21382) );
  INV_X1 U24391 ( .A(n21382), .ZN(P1_U3224) );
  AOI22_X1 U24392 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21383), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21380), .ZN(n21384) );
  OAI21_X1 U24393 ( .B1(n21386), .B2(n21385), .A(n21384), .ZN(P1_U3225) );
  AOI22_X1 U24394 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21387), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21380), .ZN(n21388) );
  OAI21_X1 U24395 ( .B1(n10683), .B2(n21389), .A(n21388), .ZN(P1_U3226) );
  INV_X1 U24396 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21493) );
  AOI22_X1 U24397 ( .A1(n21392), .A2(n21604), .B1(n21493), .B2(n21380), .ZN(
        P1_U3458) );
  OAI22_X1 U24398 ( .A1(n21380), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21392), .ZN(n21390) );
  INV_X1 U24399 ( .A(n21390), .ZN(P1_U3459) );
  OAI22_X1 U24400 ( .A1(n21380), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21392), .ZN(n21391) );
  INV_X1 U24401 ( .A(n21391), .ZN(P1_U3460) );
  OAI22_X1 U24402 ( .A1(n21380), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21392), .ZN(n21393) );
  INV_X1 U24403 ( .A(n21393), .ZN(P1_U3461) );
  OAI21_X1 U24404 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21397), .A(n21395), 
        .ZN(n21394) );
  INV_X1 U24405 ( .A(n21394), .ZN(P1_U3464) );
  OAI21_X1 U24406 ( .B1(n21397), .B2(n21396), .A(n21395), .ZN(P1_U3465) );
  AOI21_X1 U24407 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21399) );
  AOI22_X1 U24408 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21399), .B2(n21398), .ZN(n21401) );
  INV_X1 U24409 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21400) );
  AOI22_X1 U24410 ( .A1(n21402), .A2(n21401), .B1(n21400), .B2(n21405), .ZN(
        P1_U3481) );
  INV_X1 U24411 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21585) );
  NOR2_X1 U24412 ( .A1(n21405), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21403) );
  AOI22_X1 U24413 ( .A1(n21585), .A2(n21405), .B1(n21404), .B2(n21403), .ZN(
        P1_U3482) );
  AOI22_X1 U24414 ( .A1(n21392), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21406), 
        .B2(n21380), .ZN(P1_U3483) );
  AOI211_X1 U24415 ( .C1(n20684), .C2(n21409), .A(n21408), .B(n21407), .ZN(
        n21417) );
  INV_X1 U24416 ( .A(n21410), .ZN(n21411) );
  OAI211_X1 U24417 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21412), .A(n21411), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21414) );
  AOI21_X1 U24418 ( .B1(n21414), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21413), 
        .ZN(n21416) );
  NAND2_X1 U24419 ( .A1(n21417), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21415) );
  OAI21_X1 U24420 ( .B1(n21417), .B2(n21416), .A(n21415), .ZN(P1_U3485) );
  OAI22_X1 U24421 ( .A1(n21380), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n21392), .ZN(n21418) );
  INV_X1 U24422 ( .A(n21418), .ZN(P1_U3486) );
  INV_X1 U24423 ( .A(P3_LWORD_REG_12__SCAN_IN), .ZN(n21740) );
  NOR4_X1 U24424 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(P2_ADDRESS_REG_13__SCAN_IN), .A3(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A4(n21419), .ZN(n21420) );
  NAND3_X1 U24425 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n21420), .A3(
        n9919), .ZN(n21434) );
  NOR4_X1 U24426 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(n21691), .A4(n21688), .ZN(
        n21432) );
  NAND4_X1 U24427 ( .A1(n21421), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_8__SCAN_IN), .A4(n11241), .ZN(n21423) );
  NAND4_X1 U24428 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        P1_EAX_REG_10__SCAN_IN), .A3(P3_ADDRESS_REG_6__SCAN_IN), .A4(n21725), 
        .ZN(n21422) );
  NOR2_X1 U24429 ( .A1(n21423), .A2(n21422), .ZN(n21429) );
  NAND2_X1 U24430 ( .A1(n14680), .A2(n21424), .ZN(n21426) );
  NAND4_X1 U24431 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(n21715), .A4(n21673), .ZN(n21425) );
  NOR2_X1 U24432 ( .A1(n21426), .A2(n21425), .ZN(n21428) );
  AND4_X1 U24433 ( .A1(n21430), .A2(n21429), .A3(n21428), .A4(n21427), .ZN(
        n21431) );
  NAND2_X1 U24434 ( .A1(n21432), .A2(n21431), .ZN(n21433) );
  NOR4_X1 U24435 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(
        P1_LWORD_REG_4__SCAN_IN), .A3(n21434), .A4(n21433), .ZN(n21468) );
  NAND4_X1 U24436 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_2__SCAN_IN), .A3(P1_REIP_REG_19__SCAN_IN), .A4(
        BUF1_REG_18__SCAN_IN), .ZN(n21438) );
  NAND4_X1 U24437 ( .A1(BUF2_REG_31__SCAN_IN), .A2(P2_ADDRESS_REG_15__SCAN_IN), 
        .A3(n21568), .A4(n21562), .ZN(n21437) );
  NAND4_X1 U24438 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_31__SCAN_IN), .A3(P1_LWORD_REG_3__SCAN_IN), .A4(
        n21589), .ZN(n21436) );
  NAND4_X1 U24439 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n21587), .A3(n21584), 
        .A4(n21585), .ZN(n21435) );
  NOR4_X1 U24440 ( .A1(n21438), .A2(n21437), .A3(n21436), .A4(n21435), .ZN(
        n21467) );
  INV_X1 U24441 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n21542) );
  NAND4_X1 U24442 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(P3_LWORD_REG_3__SCAN_IN), 
        .A4(n21542), .ZN(n21442) );
  NAND4_X1 U24443 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(
        P3_LWORD_REG_8__SCAN_IN), .A3(P1_LWORD_REG_11__SCAN_IN), .A4(n21537), 
        .ZN(n21441) );
  NAND4_X1 U24444 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        P3_EBX_REG_26__SCAN_IN), .A3(P3_DATAO_REG_13__SCAN_IN), .A4(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n21440) );
  NAND4_X1 U24445 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n21546), .A3(n21552), 
        .A4(n21553), .ZN(n21439) );
  NOR4_X1 U24446 ( .A1(n21442), .A2(n21441), .A3(n21440), .A4(n21439), .ZN(
        n21466) );
  NOR4_X1 U24447 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A3(P3_REIP_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21446) );
  INV_X1 U24448 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n21602) );
  NOR4_X1 U24449 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n21602), .A4(n21612), .ZN(
        n21445) );
  NOR4_X1 U24450 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P2_DATAO_REG_20__SCAN_IN), 
        .A3(n21655), .A4(n21656), .ZN(n21444) );
  NOR4_X1 U24451 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P1_DATAO_REG_5__SCAN_IN), 
        .A3(n21659), .A4(n21650), .ZN(n21443) );
  NAND4_X1 U24452 ( .A1(n21446), .A2(n21445), .A3(n21444), .A4(n21443), .ZN(
        n21464) );
  NOR4_X1 U24453 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n21709), .A3(n21708), .A4(
        n21699), .ZN(n21450) );
  NOR4_X1 U24454 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(n21718), .A4(n21702), .ZN(n21449) );
  NOR4_X1 U24455 ( .A1(BUF2_REG_22__SCAN_IN), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .A3(n21625), .A4(n21627), .ZN(n21448) );
  NOR4_X1 U24456 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .A3(n21621), .A4(n21619), .ZN(n21447) );
  NAND4_X1 U24457 ( .A1(n21450), .A2(n21449), .A3(n21448), .A4(n21447), .ZN(
        n21463) );
  NOR4_X1 U24458 ( .A1(n11326), .A2(n21501), .A3(n21500), .A4(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21452) );
  NOR2_X1 U24459 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21451) );
  AND4_X1 U24460 ( .A1(n21452), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A3(
        n21451), .A4(n21508), .ZN(n21455) );
  NOR4_X1 U24461 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21517), .A3(
        n21516), .A4(n21523), .ZN(n21454) );
  INV_X1 U24462 ( .A(DATAI_3_), .ZN(n21503) );
  NOR4_X1 U24463 ( .A1(DATAI_29_), .A2(P2_LWORD_REG_5__SCAN_IN), .A3(n21506), 
        .A4(n21503), .ZN(n21453) );
  NAND3_X1 U24464 ( .A1(n21455), .A2(n21454), .A3(n21453), .ZN(n21462) );
  NOR2_X1 U24465 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21456) );
  NAND4_X1 U24466 ( .A1(n21456), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(n21471), .ZN(n21457) );
  NOR4_X1 U24467 ( .A1(n21470), .A2(n21487), .A3(n21640), .A4(n21457), .ZN(
        n21460) );
  NOR4_X1 U24468 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11287), .A3(
        n21476), .A4(n21474), .ZN(n21459) );
  NOR4_X1 U24469 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(
        P1_DATAO_REG_15__SCAN_IN), .A3(n21643), .A4(n21642), .ZN(n21458) );
  NAND3_X1 U24470 ( .A1(n21460), .A2(n21459), .A3(n21458), .ZN(n21461) );
  NOR4_X1 U24471 ( .A1(n21464), .A2(n21463), .A3(n21462), .A4(n21461), .ZN(
        n21465) );
  NAND4_X1 U24472 ( .A1(n21468), .A2(n21467), .A3(n21466), .A4(n21465), .ZN(
        n21739) );
  AOI22_X1 U24473 ( .A1(n21471), .A2(keyinput67), .B1(n21470), .B2(keyinput77), 
        .ZN(n21469) );
  OAI221_X1 U24474 ( .B1(n21471), .B2(keyinput67), .C1(n21470), .C2(keyinput77), .A(n21469), .ZN(n21483) );
  AOI22_X1 U24475 ( .A1(n21474), .A2(keyinput62), .B1(n21473), .B2(keyinput123), .ZN(n21472) );
  OAI221_X1 U24476 ( .B1(n21474), .B2(keyinput62), .C1(n21473), .C2(
        keyinput123), .A(n21472), .ZN(n21482) );
  AOI22_X1 U24477 ( .A1(n11287), .A2(keyinput122), .B1(keyinput79), .B2(n21476), .ZN(n21475) );
  OAI221_X1 U24478 ( .B1(n11287), .B2(keyinput122), .C1(n21476), .C2(
        keyinput79), .A(n21475), .ZN(n21481) );
  INV_X1 U24479 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21477) );
  XOR2_X1 U24480 ( .A(n21477), .B(keyinput24), .Z(n21479) );
  XNOR2_X1 U24481 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B(keyinput12), .ZN(
        n21478) );
  NAND2_X1 U24482 ( .A1(n21479), .A2(n21478), .ZN(n21480) );
  NOR4_X1 U24483 ( .A1(n21483), .A2(n21482), .A3(n21481), .A4(n21480), .ZN(
        n21534) );
  AOI22_X1 U24484 ( .A1(n21486), .A2(keyinput71), .B1(n21485), .B2(keyinput3), 
        .ZN(n21484) );
  OAI221_X1 U24485 ( .B1(n21486), .B2(keyinput71), .C1(n21485), .C2(keyinput3), 
        .A(n21484), .ZN(n21490) );
  XNOR2_X1 U24486 ( .A(n21487), .B(keyinput40), .ZN(n21489) );
  XNOR2_X1 U24487 ( .A(n12666), .B(keyinput110), .ZN(n21488) );
  OR3_X1 U24488 ( .A1(n21490), .A2(n21489), .A3(n21488), .ZN(n21498) );
  AOI22_X1 U24489 ( .A1(n21493), .A2(keyinput87), .B1(keyinput102), .B2(n21492), .ZN(n21491) );
  OAI221_X1 U24490 ( .B1(n21493), .B2(keyinput87), .C1(n21492), .C2(
        keyinput102), .A(n21491), .ZN(n21497) );
  AOI22_X1 U24491 ( .A1(n21495), .A2(keyinput104), .B1(n11326), .B2(keyinput69), .ZN(n21494) );
  OAI221_X1 U24492 ( .B1(n21495), .B2(keyinput104), .C1(n11326), .C2(
        keyinput69), .A(n21494), .ZN(n21496) );
  NOR3_X1 U24493 ( .A1(n21498), .A2(n21497), .A3(n21496), .ZN(n21533) );
  AOI22_X1 U24494 ( .A1(n21501), .A2(keyinput59), .B1(keyinput64), .B2(n21500), 
        .ZN(n21499) );
  OAI221_X1 U24495 ( .B1(n21501), .B2(keyinput59), .C1(n21500), .C2(keyinput64), .A(n21499), .ZN(n21514) );
  AOI22_X1 U24496 ( .A1(n21504), .A2(keyinput45), .B1(n21503), .B2(keyinput93), 
        .ZN(n21502) );
  OAI221_X1 U24497 ( .B1(n21504), .B2(keyinput45), .C1(n21503), .C2(keyinput93), .A(n21502), .ZN(n21513) );
  INV_X1 U24498 ( .A(DATAI_29_), .ZN(n21507) );
  AOI22_X1 U24499 ( .A1(n21507), .A2(keyinput46), .B1(n21506), .B2(keyinput22), 
        .ZN(n21505) );
  OAI221_X1 U24500 ( .B1(n21507), .B2(keyinput46), .C1(n21506), .C2(keyinput22), .A(n21505), .ZN(n21512) );
  XOR2_X1 U24501 ( .A(n21508), .B(keyinput48), .Z(n21510) );
  XNOR2_X1 U24502 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B(keyinput2), .ZN(
        n21509) );
  NAND2_X1 U24503 ( .A1(n21510), .A2(n21509), .ZN(n21511) );
  NOR4_X1 U24504 ( .A1(n21514), .A2(n21513), .A3(n21512), .A4(n21511), .ZN(
        n21532) );
  AOI22_X1 U24505 ( .A1(n21517), .A2(keyinput120), .B1(keyinput35), .B2(n21516), .ZN(n21515) );
  OAI221_X1 U24506 ( .B1(n21517), .B2(keyinput120), .C1(n21516), .C2(
        keyinput35), .A(n21515), .ZN(n21521) );
  XNOR2_X1 U24507 ( .A(n21518), .B(keyinput115), .ZN(n21520) );
  XOR2_X1 U24508 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B(keyinput90), .Z(
        n21519) );
  OR3_X1 U24509 ( .A1(n21521), .A2(n21520), .A3(n21519), .ZN(n21530) );
  INV_X1 U24510 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21524) );
  AOI22_X1 U24511 ( .A1(n21524), .A2(keyinput75), .B1(keyinput94), .B2(n21523), 
        .ZN(n21522) );
  OAI221_X1 U24512 ( .B1(n21524), .B2(keyinput75), .C1(n21523), .C2(keyinput94), .A(n21522), .ZN(n21529) );
  AOI22_X1 U24513 ( .A1(n21527), .A2(keyinput116), .B1(keyinput81), .B2(n21526), .ZN(n21525) );
  OAI221_X1 U24514 ( .B1(n21527), .B2(keyinput116), .C1(n21526), .C2(
        keyinput81), .A(n21525), .ZN(n21528) );
  NOR3_X1 U24515 ( .A1(n21530), .A2(n21529), .A3(n21528), .ZN(n21531) );
  NAND4_X1 U24516 ( .A1(n21534), .A2(n21533), .A3(n21532), .A4(n21531), .ZN(
        n21737) );
  AOI22_X1 U24517 ( .A1(n21537), .A2(keyinput100), .B1(keyinput78), .B2(n21536), .ZN(n21535) );
  OAI221_X1 U24518 ( .B1(n21537), .B2(keyinput100), .C1(n21536), .C2(
        keyinput78), .A(n21535), .ZN(n21550) );
  AOI22_X1 U24519 ( .A1(n21540), .A2(keyinput17), .B1(keyinput25), .B2(n21539), 
        .ZN(n21538) );
  OAI221_X1 U24520 ( .B1(n21540), .B2(keyinput17), .C1(n21539), .C2(keyinput25), .A(n21538), .ZN(n21549) );
  AOI22_X1 U24521 ( .A1(n21543), .A2(keyinput97), .B1(n21542), .B2(keyinput52), 
        .ZN(n21541) );
  OAI221_X1 U24522 ( .B1(n21543), .B2(keyinput97), .C1(n21542), .C2(keyinput52), .A(n21541), .ZN(n21548) );
  AOI22_X1 U24523 ( .A1(n21546), .A2(keyinput88), .B1(keyinput111), .B2(n21545), .ZN(n21544) );
  OAI221_X1 U24524 ( .B1(n21546), .B2(keyinput88), .C1(n21545), .C2(
        keyinput111), .A(n21544), .ZN(n21547) );
  NOR4_X1 U24525 ( .A1(n21550), .A2(n21549), .A3(n21548), .A4(n21547), .ZN(
        n21600) );
  AOI22_X1 U24526 ( .A1(n21553), .A2(keyinput47), .B1(n21552), .B2(keyinput33), 
        .ZN(n21551) );
  OAI221_X1 U24527 ( .B1(n21553), .B2(keyinput47), .C1(n21552), .C2(keyinput33), .A(n21551), .ZN(n21566) );
  AOI22_X1 U24528 ( .A1(n21556), .A2(keyinput0), .B1(keyinput61), .B2(n21555), 
        .ZN(n21554) );
  OAI221_X1 U24529 ( .B1(n21556), .B2(keyinput0), .C1(n21555), .C2(keyinput61), 
        .A(n21554), .ZN(n21565) );
  AOI22_X1 U24530 ( .A1(n21559), .A2(keyinput98), .B1(n21558), .B2(keyinput65), 
        .ZN(n21557) );
  OAI221_X1 U24531 ( .B1(n21559), .B2(keyinput98), .C1(n21558), .C2(keyinput65), .A(n21557), .ZN(n21564) );
  AOI22_X1 U24532 ( .A1(n21562), .A2(keyinput29), .B1(n21561), .B2(keyinput66), 
        .ZN(n21560) );
  OAI221_X1 U24533 ( .B1(n21562), .B2(keyinput29), .C1(n21561), .C2(keyinput66), .A(n21560), .ZN(n21563) );
  NOR4_X1 U24534 ( .A1(n21566), .A2(n21565), .A3(n21564), .A4(n21563), .ZN(
        n21599) );
  AOI22_X1 U24535 ( .A1(n21569), .A2(keyinput108), .B1(keyinput89), .B2(n21568), .ZN(n21567) );
  OAI221_X1 U24536 ( .B1(n21569), .B2(keyinput108), .C1(n21568), .C2(
        keyinput89), .A(n21567), .ZN(n21582) );
  INV_X1 U24537 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21572) );
  AOI22_X1 U24538 ( .A1(n21572), .A2(keyinput85), .B1(keyinput42), .B2(n21571), 
        .ZN(n21570) );
  OAI221_X1 U24539 ( .B1(n21572), .B2(keyinput85), .C1(n21571), .C2(keyinput42), .A(n21570), .ZN(n21581) );
  AOI22_X1 U24540 ( .A1(n21575), .A2(keyinput127), .B1(keyinput96), .B2(n21574), .ZN(n21573) );
  OAI221_X1 U24541 ( .B1(n21575), .B2(keyinput127), .C1(n21574), .C2(
        keyinput96), .A(n21573), .ZN(n21580) );
  AOI22_X1 U24542 ( .A1(n21578), .A2(keyinput27), .B1(keyinput101), .B2(n21577), .ZN(n21576) );
  OAI221_X1 U24543 ( .B1(n21578), .B2(keyinput27), .C1(n21577), .C2(
        keyinput101), .A(n21576), .ZN(n21579) );
  NOR4_X1 U24544 ( .A1(n21582), .A2(n21581), .A3(n21580), .A4(n21579), .ZN(
        n21598) );
  AOI22_X1 U24545 ( .A1(n21585), .A2(keyinput84), .B1(n21584), .B2(keyinput11), 
        .ZN(n21583) );
  OAI221_X1 U24546 ( .B1(n21585), .B2(keyinput84), .C1(n21584), .C2(keyinput11), .A(n21583), .ZN(n21596) );
  AOI22_X1 U24547 ( .A1(n21587), .A2(keyinput7), .B1(n11427), .B2(keyinput44), 
        .ZN(n21586) );
  OAI221_X1 U24548 ( .B1(n21587), .B2(keyinput7), .C1(n11427), .C2(keyinput44), 
        .A(n21586), .ZN(n21595) );
  AOI22_X1 U24549 ( .A1(n21590), .A2(keyinput26), .B1(n21589), .B2(keyinput95), 
        .ZN(n21588) );
  OAI221_X1 U24550 ( .B1(n21590), .B2(keyinput26), .C1(n21589), .C2(keyinput95), .A(n21588), .ZN(n21594) );
  AOI22_X1 U24551 ( .A1(n21592), .A2(keyinput32), .B1(n11241), .B2(keyinput82), 
        .ZN(n21591) );
  OAI221_X1 U24552 ( .B1(n21592), .B2(keyinput32), .C1(n11241), .C2(keyinput82), .A(n21591), .ZN(n21593) );
  NOR4_X1 U24553 ( .A1(n21596), .A2(n21595), .A3(n21594), .A4(n21593), .ZN(
        n21597) );
  NAND4_X1 U24554 ( .A1(n21600), .A2(n21599), .A3(n21598), .A4(n21597), .ZN(
        n21736) );
  AOI22_X1 U24555 ( .A1(n21603), .A2(keyinput37), .B1(keyinput28), .B2(n21602), 
        .ZN(n21601) );
  OAI221_X1 U24556 ( .B1(n21603), .B2(keyinput37), .C1(n21602), .C2(keyinput28), .A(n21601), .ZN(n21607) );
  XNOR2_X1 U24557 ( .A(n14680), .B(keyinput92), .ZN(n21606) );
  XNOR2_X1 U24558 ( .A(n21604), .B(keyinput4), .ZN(n21605) );
  OR3_X1 U24559 ( .A1(n21607), .A2(n21606), .A3(n21605), .ZN(n21616) );
  AOI22_X1 U24560 ( .A1(n21610), .A2(keyinput112), .B1(keyinput118), .B2(
        n21609), .ZN(n21608) );
  OAI221_X1 U24561 ( .B1(n21610), .B2(keyinput112), .C1(n21609), .C2(
        keyinput118), .A(n21608), .ZN(n21615) );
  AOI22_X1 U24562 ( .A1(n21613), .A2(keyinput126), .B1(keyinput56), .B2(n21612), .ZN(n21611) );
  OAI221_X1 U24563 ( .B1(n21613), .B2(keyinput126), .C1(n21612), .C2(
        keyinput56), .A(n21611), .ZN(n21614) );
  NOR3_X1 U24564 ( .A1(n21616), .A2(n21615), .A3(n21614), .ZN(n21667) );
  AOI22_X1 U24565 ( .A1(n21619), .A2(keyinput54), .B1(n21618), .B2(keyinput10), 
        .ZN(n21617) );
  OAI221_X1 U24566 ( .B1(n21619), .B2(keyinput54), .C1(n21618), .C2(keyinput10), .A(n21617), .ZN(n21631) );
  AOI22_X1 U24567 ( .A1(n21622), .A2(keyinput5), .B1(keyinput114), .B2(n21621), 
        .ZN(n21620) );
  OAI221_X1 U24568 ( .B1(n21622), .B2(keyinput5), .C1(n21621), .C2(keyinput114), .A(n21620), .ZN(n21630) );
  AOI22_X1 U24569 ( .A1(n21625), .A2(keyinput58), .B1(keyinput117), .B2(n21624), .ZN(n21623) );
  OAI221_X1 U24570 ( .B1(n21625), .B2(keyinput58), .C1(n21624), .C2(
        keyinput117), .A(n21623), .ZN(n21629) );
  AOI22_X1 U24571 ( .A1(n21627), .A2(keyinput103), .B1(keyinput16), .B2(n17354), .ZN(n21626) );
  OAI221_X1 U24572 ( .B1(n21627), .B2(keyinput103), .C1(n17354), .C2(
        keyinput16), .A(n21626), .ZN(n21628) );
  NOR4_X1 U24573 ( .A1(n21631), .A2(n21630), .A3(n21629), .A4(n21628), .ZN(
        n21666) );
  AOI22_X1 U24574 ( .A1(n21634), .A2(keyinput38), .B1(keyinput19), .B2(n21633), 
        .ZN(n21632) );
  OAI221_X1 U24575 ( .B1(n21634), .B2(keyinput38), .C1(n21633), .C2(keyinput19), .A(n21632), .ZN(n21647) );
  AOI22_X1 U24576 ( .A1(n21637), .A2(keyinput31), .B1(keyinput53), .B2(n21636), 
        .ZN(n21635) );
  OAI221_X1 U24577 ( .B1(n21637), .B2(keyinput31), .C1(n21636), .C2(keyinput53), .A(n21635), .ZN(n21646) );
  AOI22_X1 U24578 ( .A1(n21640), .A2(keyinput83), .B1(n21639), .B2(keyinput50), 
        .ZN(n21638) );
  OAI221_X1 U24579 ( .B1(n21640), .B2(keyinput83), .C1(n21639), .C2(keyinput50), .A(n21638), .ZN(n21645) );
  AOI22_X1 U24580 ( .A1(n21643), .A2(keyinput39), .B1(keyinput60), .B2(n21642), 
        .ZN(n21641) );
  OAI221_X1 U24581 ( .B1(n21643), .B2(keyinput39), .C1(n21642), .C2(keyinput60), .A(n21641), .ZN(n21644) );
  NOR4_X1 U24582 ( .A1(n21647), .A2(n21646), .A3(n21645), .A4(n21644), .ZN(
        n21665) );
  AOI22_X1 U24583 ( .A1(n21650), .A2(keyinput74), .B1(keyinput68), .B2(n21649), 
        .ZN(n21648) );
  OAI221_X1 U24584 ( .B1(n21650), .B2(keyinput74), .C1(n21649), .C2(keyinput68), .A(n21648), .ZN(n21663) );
  AOI22_X1 U24585 ( .A1(n21653), .A2(keyinput121), .B1(keyinput119), .B2(
        n21652), .ZN(n21651) );
  OAI221_X1 U24586 ( .B1(n21653), .B2(keyinput121), .C1(n21652), .C2(
        keyinput119), .A(n21651), .ZN(n21662) );
  AOI22_X1 U24587 ( .A1(n21656), .A2(keyinput1), .B1(n21655), .B2(keyinput18), 
        .ZN(n21654) );
  OAI221_X1 U24588 ( .B1(n21656), .B2(keyinput1), .C1(n21655), .C2(keyinput18), 
        .A(n21654), .ZN(n21661) );
  AOI22_X1 U24589 ( .A1(n21659), .A2(keyinput30), .B1(keyinput34), .B2(n21658), 
        .ZN(n21657) );
  OAI221_X1 U24590 ( .B1(n21659), .B2(keyinput30), .C1(n21658), .C2(keyinput34), .A(n21657), .ZN(n21660) );
  NOR4_X1 U24591 ( .A1(n21663), .A2(n21662), .A3(n21661), .A4(n21660), .ZN(
        n21664) );
  NAND4_X1 U24592 ( .A1(n21667), .A2(n21666), .A3(n21665), .A4(n21664), .ZN(
        n21735) );
  INV_X1 U24593 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21669) );
  AOI22_X1 U24594 ( .A1(n21670), .A2(keyinput106), .B1(n21669), .B2(
        keyinput107), .ZN(n21668) );
  OAI221_X1 U24595 ( .B1(n21670), .B2(keyinput106), .C1(n21669), .C2(
        keyinput107), .A(n21668), .ZN(n21677) );
  AOI22_X1 U24596 ( .A1(n21673), .A2(keyinput49), .B1(n21672), .B2(keyinput21), 
        .ZN(n21671) );
  OAI221_X1 U24597 ( .B1(n21673), .B2(keyinput49), .C1(n21672), .C2(keyinput21), .A(n21671), .ZN(n21676) );
  XNOR2_X1 U24598 ( .A(n21674), .B(keyinput91), .ZN(n21675) );
  OR3_X1 U24599 ( .A1(n21677), .A2(n21676), .A3(n21675), .ZN(n21683) );
  AOI22_X1 U24600 ( .A1(n9919), .A2(keyinput6), .B1(keyinput36), .B2(n21679), 
        .ZN(n21678) );
  OAI221_X1 U24601 ( .B1(n9919), .B2(keyinput6), .C1(n21679), .C2(keyinput36), 
        .A(n21678), .ZN(n21682) );
  XNOR2_X1 U24602 ( .A(n21680), .B(keyinput86), .ZN(n21681) );
  NOR3_X1 U24603 ( .A1(n21683), .A2(n21682), .A3(n21681), .ZN(n21733) );
  AOI22_X1 U24604 ( .A1(n21686), .A2(keyinput99), .B1(n21685), .B2(keyinput63), 
        .ZN(n21684) );
  OAI221_X1 U24605 ( .B1(n21686), .B2(keyinput99), .C1(n21685), .C2(keyinput63), .A(n21684), .ZN(n21697) );
  AOI22_X1 U24606 ( .A1(n21689), .A2(keyinput51), .B1(keyinput55), .B2(n21688), 
        .ZN(n21687) );
  OAI221_X1 U24607 ( .B1(n21689), .B2(keyinput51), .C1(n21688), .C2(keyinput55), .A(n21687), .ZN(n21696) );
  AOI22_X1 U24608 ( .A1(keyinput72), .A2(n21691), .B1(keyinput124), .B2(n21740), .ZN(n21690) );
  OAI21_X1 U24609 ( .B1(n21691), .B2(keyinput72), .A(n21690), .ZN(n21695) );
  XNOR2_X1 U24610 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B(keyinput8), .ZN(
        n21693) );
  XNOR2_X1 U24611 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B(keyinput43), 
        .ZN(n21692) );
  NAND2_X1 U24612 ( .A1(n21693), .A2(n21692), .ZN(n21694) );
  NOR4_X1 U24613 ( .A1(n21697), .A2(n21696), .A3(n21695), .A4(n21694), .ZN(
        n21732) );
  AOI22_X1 U24614 ( .A1(n21700), .A2(keyinput20), .B1(n21699), .B2(keyinput70), 
        .ZN(n21698) );
  OAI221_X1 U24615 ( .B1(n21700), .B2(keyinput20), .C1(n21699), .C2(keyinput70), .A(n21698), .ZN(n21713) );
  AOI22_X1 U24616 ( .A1(n21703), .A2(keyinput23), .B1(keyinput125), .B2(n21702), .ZN(n21701) );
  OAI221_X1 U24617 ( .B1(n21703), .B2(keyinput23), .C1(n21702), .C2(
        keyinput125), .A(n21701), .ZN(n21712) );
  AOI22_X1 U24618 ( .A1(n21706), .A2(keyinput15), .B1(keyinput57), .B2(n21705), 
        .ZN(n21704) );
  OAI221_X1 U24619 ( .B1(n21706), .B2(keyinput15), .C1(n21705), .C2(keyinput57), .A(n21704), .ZN(n21711) );
  AOI22_X1 U24620 ( .A1(n21709), .A2(keyinput109), .B1(n21708), .B2(keyinput76), .ZN(n21707) );
  OAI221_X1 U24621 ( .B1(n21709), .B2(keyinput109), .C1(n21708), .C2(
        keyinput76), .A(n21707), .ZN(n21710) );
  NOR4_X1 U24622 ( .A1(n21713), .A2(n21712), .A3(n21711), .A4(n21710), .ZN(
        n21731) );
  AOI22_X1 U24623 ( .A1(n21716), .A2(keyinput105), .B1(n21715), .B2(keyinput80), .ZN(n21714) );
  OAI221_X1 U24624 ( .B1(n21716), .B2(keyinput105), .C1(n21715), .C2(
        keyinput80), .A(n21714), .ZN(n21729) );
  AOI22_X1 U24625 ( .A1(n21719), .A2(keyinput73), .B1(n21718), .B2(keyinput13), 
        .ZN(n21717) );
  OAI221_X1 U24626 ( .B1(n21719), .B2(keyinput73), .C1(n21718), .C2(keyinput13), .A(n21717), .ZN(n21723) );
  XNOR2_X1 U24627 ( .A(n21720), .B(keyinput9), .ZN(n21722) );
  XOR2_X1 U24628 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B(keyinput41), .Z(
        n21721) );
  OR3_X1 U24629 ( .A1(n21723), .A2(n21722), .A3(n21721), .ZN(n21728) );
  AOI22_X1 U24630 ( .A1(n21726), .A2(keyinput14), .B1(n21725), .B2(keyinput113), .ZN(n21724) );
  OAI221_X1 U24631 ( .B1(n21726), .B2(keyinput14), .C1(n21725), .C2(
        keyinput113), .A(n21724), .ZN(n21727) );
  NOR3_X1 U24632 ( .A1(n21729), .A2(n21728), .A3(n21727), .ZN(n21730) );
  NAND4_X1 U24633 ( .A1(n21733), .A2(n21732), .A3(n21731), .A4(n21730), .ZN(
        n21734) );
  NOR4_X1 U24634 ( .A1(n21737), .A2(n21736), .A3(n21735), .A4(n21734), .ZN(
        n21738) );
  OAI221_X1 U24635 ( .B1(keyinput124), .B2(n21740), .C1(keyinput124), .C2(
        n21739), .A(n21738), .ZN(n21753) );
  AOI22_X1 U24636 ( .A1(n21744), .A2(n21743), .B1(n21742), .B2(n21741), .ZN(
        n21749) );
  AOI22_X1 U24637 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21747), .B1(
        n21746), .B2(n21745), .ZN(n21748) );
  OAI211_X1 U24638 ( .C1(n21751), .C2(n21750), .A(n21749), .B(n21748), .ZN(
        n21752) );
  XNOR2_X1 U24639 ( .A(n21753), .B(n21752), .ZN(P2_U3169) );
  NAND2_X1 U11233 ( .A1(n11828), .A2(n11076), .ZN(n11860) );
  INV_X1 U11604 ( .A(n18197), .ZN(n19105) );
  CLKBUF_X3 U11127 ( .A(n13880), .Z(n9689) );
  BUF_X2 U11192 ( .A(n11380), .Z(n16629) );
  AND2_X2 U11583 ( .A1(n9711), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11238) );
  CLKBUF_X3 U11143 ( .A(n11055), .Z(n11065) );
  CLKBUF_X2 U11154 ( .A(n12741), .Z(n12756) );
  CLKBUF_X1 U11162 ( .A(n11062), .Z(n11635) );
  CLKBUF_X1 U11172 ( .A(n12687), .Z(n12688) );
  CLKBUF_X2 U11177 ( .A(n11078), .Z(n11840) );
  CLKBUF_X1 U11181 ( .A(n11183), .Z(n9704) );
  CLKBUF_X1 U11182 ( .A(n13754), .Z(n9694) );
  AND2_X1 U11210 ( .A1(n13584), .A2(n13590), .ZN(n13777) );
  CLKBUF_X1 U11226 ( .A(n12677), .Z(n21412) );
  CLKBUF_X1 U11274 ( .A(n20852), .Z(n9707) );
  CLKBUF_X1 U11277 ( .A(n11518), .Z(n11516) );
  CLKBUF_X1 U11281 ( .A(n11099), .Z(n14264) );
  CLKBUF_X1 U11322 ( .A(n12482), .Z(n16036) );
  AND2_X1 U11522 ( .A1(n16802), .A2(n10738), .ZN(n10083) );
  CLKBUF_X1 U11971 ( .A(n16004), .Z(n16022) );
  CLKBUF_X1 U12593 ( .A(n13605), .Z(n15966) );
  NAND2_X2 U13603 ( .A1(n19548), .A2(n18949), .ZN(n19030) );
  CLKBUF_X1 U13637 ( .A(n11183), .Z(n9703) );
endmodule

