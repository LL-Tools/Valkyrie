

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558;

  CLKBUF_X2 U2256 ( .A(n2275), .Z(n2763) );
  INV_X1 U2257 ( .A(n2713), .ZN(n2318) );
  INV_X1 U2258 ( .A(n2689), .ZN(n2716) );
  INV_X2 U2259 ( .A(n2339), .ZN(n2611) );
  OR2_X1 U2260 ( .A1(n3341), .A2(n3617), .ZN(n2067) );
  INV_X1 U2261 ( .A(n2703), .ZN(n2014) );
  CLKBUF_X3 U2263 ( .A(n2301), .Z(n3586) );
  CLKBUF_X2 U2264 ( .A(n2322), .Z(n2915) );
  INV_X2 U2265 ( .A(n4453), .ZN(n4442) );
  NAND4_X2 U2266 ( .A1(n2712), .A2(n2711), .A3(n2710), .A4(n2709), .ZN(n3776)
         );
  OAI21_X2 U2267 ( .B1(n3782), .B2(n2836), .A(n2080), .ZN(n3765) );
  NAND2_X1 U2268 ( .A1(n3541), .A2(n3539), .ZN(n2844) );
  NAND2_X1 U2269 ( .A1(n3137), .A2(n3107), .ZN(n3539) );
  NAND2_X1 U2270 ( .A1(n2029), .A2(n2218), .ZN(n2438) );
  BUF_X1 U2271 ( .A(n4491), .Z(n2015) );
  AOI21_X1 U2272 ( .B1(n2876), .B2(n4534), .A(n2875), .ZN(n2894) );
  OAI22_X1 U2273 ( .A1(n3444), .A2(n2629), .B1(n2628), .B2(n2627), .ZN(n3407)
         );
  NAND2_X1 U2274 ( .A1(n2067), .A2(n2815), .ZN(n3353) );
  NOR2_X1 U2275 ( .A1(n2027), .A2(n3743), .ZN(n2120) );
  NAND2_X1 U2276 ( .A1(n2804), .A2(n2803), .ZN(n3235) );
  NAND2_X1 U2277 ( .A1(n2799), .A2(n2798), .ZN(n3118) );
  OR2_X1 U2278 ( .A1(n2680), .A2(n3510), .ZN(n2697) );
  NAND2_X1 U2279 ( .A1(n2325), .A2(n2324), .ZN(n3690) );
  INV_X1 U2280 ( .A(n3073), .ZN(n2270) );
  AND2_X1 U2281 ( .A1(n2769), .A2(n2742), .ZN(n3073) );
  AND4_X1 U2282 ( .A1(n2300), .A2(n2299), .A3(n2298), .A4(n2297), .ZN(n3137)
         );
  INV_X1 U2283 ( .A(n2797), .ZN(n3083) );
  AND2_X1 U2284 ( .A1(n2033), .A2(n2107), .ZN(n2109) );
  NAND2_X1 U2285 ( .A1(n2304), .A2(n2303), .ZN(n3107) );
  AND2_X1 U2286 ( .A1(n2838), .A2(n2751), .ZN(n4448) );
  NAND4_X1 U2287 ( .A1(n2281), .A2(n2280), .A3(n2279), .A4(n2278), .ZN(n2840)
         );
  XNOR2_X1 U2288 ( .A(n2251), .B(n2250), .ZN(n2769) );
  NAND2_X1 U2289 ( .A1(n3586), .A2(DATAI_2_), .ZN(n2303) );
  XNOR2_X1 U2290 ( .A(n2255), .B(n2221), .ZN(n2751) );
  OR2_X1 U2291 ( .A1(n3586), .A2(n2940), .ZN(n2304) );
  INV_X1 U2292 ( .A(n4421), .ZN(n4436) );
  NAND2_X1 U2293 ( .A1(n2254), .A2(IR_REG_31__SCAN_IN), .ZN(n2255) );
  NAND2_X1 U2294 ( .A1(n2269), .A2(IR_REG_31__SCAN_IN), .ZN(n2251) );
  OAI211_X1 U2295 ( .C1(n2925), .C2(IR_REG_27__SCAN_IN), .A(n2258), .B(n2259), 
        .ZN(n2301) );
  NAND2_X1 U2296 ( .A1(n2738), .A2(IR_REG_31__SCAN_IN), .ZN(n2243) );
  NAND2_X1 U2297 ( .A1(n2138), .A2(IR_REG_31__SCAN_IN), .ZN(n2925) );
  NOR2_X1 U2298 ( .A1(n2573), .A2(IR_REG_17__SCAN_IN), .ZN(n2586) );
  NOR2_X2 U2299 ( .A1(n2225), .A2(n2224), .ZN(n2241) );
  NOR2_X1 U2300 ( .A1(n2209), .A2(IR_REG_28__SCAN_IN), .ZN(n2208) );
  NOR2_X1 U2301 ( .A1(n2130), .A2(IR_REG_29__SCAN_IN), .ZN(n2129) );
  AND2_X1 U2302 ( .A1(n2266), .A2(n2250), .ZN(n2252) );
  AND2_X1 U2303 ( .A1(n2362), .A2(n2216), .ZN(n2218) );
  INV_X1 U2304 ( .A(IR_REG_0__SCAN_IN), .ZN(n4491) );
  INV_X1 U2305 ( .A(IR_REG_12__SCAN_IN), .ZN(n2504) );
  INV_X1 U2306 ( .A(IR_REG_14__SCAN_IN), .ZN(n2544) );
  INV_X1 U2307 ( .A(IR_REG_15__SCAN_IN), .ZN(n2558) );
  NOR2_X1 U2308 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2362)
         );
  INV_X1 U2309 ( .A(IR_REG_10__SCAN_IN), .ZN(n4107) );
  NOR2_X1 U2310 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2216)
         );
  INV_X1 U2311 ( .A(IR_REG_27__SCAN_IN), .ZN(n2924) );
  INV_X1 U2312 ( .A(IR_REG_24__SCAN_IN), .ZN(n2242) );
  INV_X1 U2313 ( .A(IR_REG_11__SCAN_IN), .ZN(n2503) );
  INV_X1 U2314 ( .A(IR_REG_20__SCAN_IN), .ZN(n2250) );
  INV_X1 U2315 ( .A(IR_REG_19__SCAN_IN), .ZN(n2266) );
  NOR2_X1 U2316 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2226)
         );
  OR2_X2 U2317 ( .A1(n2713), .A2(n4537), .ZN(n2703) );
  NAND3_X2 U2318 ( .A1(n2109), .A2(n2110), .A3(n2239), .ZN(n2790) );
  OAI21_X2 U2319 ( .B1(n3155), .B2(n2802), .A(n2801), .ZN(n3183) );
  OAI22_X2 U2320 ( .A1(n3118), .A2(n2800), .B1(n3127), .B2(n3688), .ZN(n3155)
         );
  XNOR2_X2 U2321 ( .A(n2231), .B(n2230), .ZN(n2238) );
  OAI21_X2 U2322 ( .B1(n3134), .B2(n2795), .A(n2794), .ZN(n3066) );
  NAND2_X2 U2323 ( .A1(n3099), .A2(n2793), .ZN(n3134) );
  OAI21_X2 U2324 ( .B1(n3235), .B2(n2806), .A(n2805), .ZN(n3208) );
  OAI22_X2 U2325 ( .A1(n3811), .A2(n2835), .B1(n3824), .B2(n3457), .ZN(n3782)
         );
  OAI21_X2 U2326 ( .B1(n3828), .B2(n2834), .A(n2833), .ZN(n3811) );
  AND2_X1 U2327 ( .A1(n2238), .A2(n2236), .ZN(n2322) );
  NAND2_X4 U2328 ( .A1(n4225), .A2(n2236), .ZN(n2319) );
  XNOR2_X2 U2329 ( .A(n2234), .B(n2233), .ZN(n2236) );
  INV_X1 U2330 ( .A(n3494), .ZN(n2176) );
  AND2_X1 U2331 ( .A1(n2171), .A2(n2173), .ZN(n2170) );
  INV_X1 U2332 ( .A(n3435), .ZN(n2171) );
  INV_X1 U2333 ( .A(n2064), .ZN(n2063) );
  AOI21_X1 U2334 ( .B1(n2181), .B2(n2185), .A(n2179), .ZN(n2178) );
  OAI21_X1 U2335 ( .B1(n2120), .B2(n3757), .A(n2117), .ZN(n2116) );
  NAND2_X1 U2336 ( .A1(n2120), .A2(n2118), .ZN(n2117) );
  NAND2_X1 U2337 ( .A1(n3742), .A2(n3756), .ZN(n2118) );
  NAND2_X1 U2338 ( .A1(n3136), .A2(n3545), .ZN(n3076) );
  INV_X1 U2339 ( .A(n2257), .ZN(n2099) );
  NAND2_X1 U2340 ( .A1(n2020), .A2(n2176), .ZN(n2173) );
  AND2_X1 U2341 ( .A1(n2271), .A2(n2270), .ZN(n2689) );
  AND2_X1 U2342 ( .A1(n2892), .A2(n2737), .ZN(n2774) );
  INV_X1 U2343 ( .A(n3788), .ZN(n3511) );
  NAND2_X1 U2344 ( .A1(n3779), .A2(n3513), .ZN(n2080) );
  NAND2_X1 U2345 ( .A1(n2069), .A2(n2019), .ZN(n3860) );
  NAND2_X1 U2346 ( .A1(n3904), .A2(n2070), .ZN(n2069) );
  NOR2_X1 U2347 ( .A1(n3594), .A2(n2042), .ZN(n2071) );
  NAND2_X1 U2348 ( .A1(n3957), .A2(n2818), .ZN(n2076) );
  OR2_X1 U2349 ( .A1(n3949), .A2(n3966), .ZN(n2818) );
  AND2_X1 U2350 ( .A1(n4234), .A2(n2920), .ZN(n4423) );
  OR2_X1 U2351 ( .A1(n4234), .A2(n2871), .ZN(n4426) );
  AND3_X1 U2352 ( .A1(n2110), .A2(n4421), .A3(n2239), .ZN(n2108) );
  INV_X1 U2353 ( .A(n3249), .ZN(n2184) );
  XNOR2_X1 U2354 ( .A(n2328), .B(n2716), .ZN(n2346) );
  NAND2_X1 U2355 ( .A1(n2327), .A2(n2326), .ZN(n2328) );
  NAND2_X1 U2356 ( .A1(n3690), .A2(n2611), .ZN(n2326) );
  OAI22_X1 U2357 ( .A1(n4319), .A2(n4317), .B1(n3724), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3725) );
  NOR2_X1 U2358 ( .A1(n3822), .A2(n3653), .ZN(n3801) );
  INV_X1 U2359 ( .A(n3576), .ZN(n2128) );
  NAND2_X1 U2360 ( .A1(n2857), .A2(n2856), .ZN(n3898) );
  INV_X1 U2361 ( .A(n2105), .ZN(n2104) );
  OAI21_X1 U2362 ( .B1(n2854), .B2(n2106), .A(n3368), .ZN(n2105) );
  INV_X1 U2363 ( .A(n3523), .ZN(n2106) );
  OAI21_X1 U2364 ( .B1(n2065), .B2(n2063), .A(n2812), .ZN(n2062) );
  OR2_X1 U2365 ( .A1(n2063), .A2(n2811), .ZN(n2059) );
  INV_X1 U2366 ( .A(n3551), .ZN(n2123) );
  NAND2_X1 U2367 ( .A1(n2846), .A2(n3133), .ZN(n3136) );
  NOR2_X1 U2368 ( .A1(n2528), .A2(IR_REG_13__SCAN_IN), .ZN(n2545) );
  NOR2_X1 U2369 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2085)
         );
  INV_X1 U2370 ( .A(n3473), .ZN(n2206) );
  AOI21_X1 U2371 ( .B1(n2193), .B2(n2195), .A(n2046), .ZN(n2191) );
  AOI21_X1 U2372 ( .B1(n2170), .B2(n2168), .A(n2045), .ZN(n2167) );
  INV_X1 U2373 ( .A(n2037), .ZN(n2168) );
  INV_X1 U2374 ( .A(n2170), .ZN(n2169) );
  OR2_X1 U2375 ( .A1(n3137), .A2(n2703), .ZN(n2308) );
  OAI21_X1 U2376 ( .B1(n3137), .B2(n2339), .A(n2305), .ZN(n2306) );
  OR2_X1 U2377 ( .A1(n2918), .A2(n2878), .ZN(n2986) );
  NAND2_X1 U2378 ( .A1(n2579), .A2(n2211), .ZN(n2175) );
  AND2_X1 U2379 ( .A1(n2774), .A2(n2773), .ZN(n3488) );
  OR2_X1 U2380 ( .A1(n2763), .A2(n3768), .ZN(n2700) );
  OR2_X1 U2381 ( .A1(n2763), .A2(n3833), .ZN(n2657) );
  AND2_X1 U2383 ( .A1(n2915), .A2(REG0_REG_3__SCAN_IN), .ZN(n2212) );
  NAND2_X1 U2384 ( .A1(n2972), .A2(n2090), .ZN(n2089) );
  NAND2_X1 U2385 ( .A1(n4232), .A2(REG2_REG_2__SCAN_IN), .ZN(n2090) );
  INV_X1 U2386 ( .A(n2145), .ZN(n2144) );
  OAI21_X1 U2387 ( .B1(n2944), .B2(n2147), .A(REG1_REG_3__SCAN_IN), .ZN(n2145)
         );
  OAI22_X1 U2388 ( .A1(n3009), .A2(n3008), .B1(n2147), .B2(n2088), .ZN(n3010)
         );
  INV_X1 U2389 ( .A(n2089), .ZN(n2088) );
  XNOR2_X1 U2390 ( .A(n3010), .B(n4231), .ZN(n3033) );
  NOR2_X1 U2391 ( .A1(n4247), .A2(n3001), .ZN(n3002) );
  AND2_X1 U2392 ( .A1(n3007), .A2(REG1_REG_5__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U2393 ( .A1(n2152), .A2(n2151), .ZN(n3692) );
  NAND2_X1 U2394 ( .A1(n2153), .A2(REG1_REG_7__SCAN_IN), .ZN(n2151) );
  OAI21_X1 U2395 ( .B1(n2153), .B2(REG1_REG_7__SCAN_IN), .A(n4230), .ZN(n2152)
         );
  XNOR2_X1 U2396 ( .A(n3713), .B(n4485), .ZN(n4267) );
  NAND2_X1 U2397 ( .A1(n3711), .A2(n2093), .ZN(n3713) );
  NAND2_X1 U2398 ( .A1(n4230), .A2(REG2_REG_7__SCAN_IN), .ZN(n2093) );
  NAND2_X1 U2399 ( .A1(n4267), .A2(REG2_REG_8__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U2400 ( .A1(n4278), .A2(n3715), .ZN(n3717) );
  XNOR2_X1 U2401 ( .A(n3721), .B(n4478), .ZN(n4309) );
  NAND2_X1 U2402 ( .A1(n4300), .A2(n3720), .ZN(n3721) );
  NAND2_X1 U2403 ( .A1(n3710), .A2(REG2_REG_11__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U2404 ( .A1(n4323), .A2(n2051), .ZN(n3702) );
  XNOR2_X1 U2405 ( .A(n3705), .B(n4470), .ZN(n4352) );
  NAND2_X1 U2406 ( .A1(n4349), .A2(n3729), .ZN(n4363) );
  NAND2_X1 U2407 ( .A1(n4363), .A2(n4365), .ZN(n4364) );
  NOR2_X1 U2408 ( .A1(n3760), .A2(n3761), .ZN(n3982) );
  INV_X1 U2409 ( .A(n3848), .ZN(n3807) );
  OR2_X1 U2410 ( .A1(n3848), .A2(n3474), .ZN(n2833) );
  NOR2_X1 U2411 ( .A1(n3807), .A2(n3832), .ZN(n2834) );
  AND2_X1 U2412 ( .A1(n3947), .A2(n2821), .ZN(n2822) );
  NAND2_X1 U2413 ( .A1(n3961), .A2(n3390), .ZN(n2077) );
  NAND2_X1 U2414 ( .A1(n3366), .A2(n3604), .ZN(n2078) );
  NAND2_X1 U2415 ( .A1(n2016), .A2(n2028), .ZN(n2064) );
  AND2_X1 U2416 ( .A1(n2016), .A2(n4387), .ZN(n2065) );
  NAND2_X1 U2417 ( .A1(n2850), .A2(n3560), .ZN(n3204) );
  OAI21_X1 U2418 ( .B1(n3120), .B2(n3119), .A(n3555), .ZN(n3150) );
  NAND2_X1 U2419 ( .A1(n3767), .A2(n2887), .ZN(n3760) );
  NAND2_X1 U2420 ( .A1(n4430), .A2(n4498), .ZN(n4534) );
  NAND2_X1 U2421 ( .A1(n2256), .A2(n2757), .ZN(n2918) );
  NAND2_X1 U2422 ( .A1(n3423), .A2(IR_REG_31__SCAN_IN), .ZN(n2231) );
  NAND2_X1 U2423 ( .A1(n2030), .A2(n2227), .ZN(n2209) );
  AND3_X1 U2424 ( .A1(n2240), .A2(n2241), .A3(n2226), .ZN(n2228) );
  NAND2_X1 U2425 ( .A1(n2099), .A2(n4108), .ZN(n2315) );
  NAND2_X1 U2426 ( .A1(n2015), .A2(n2084), .ZN(n2257) );
  INV_X1 U2427 ( .A(IR_REG_1__SCAN_IN), .ZN(n2084) );
  INV_X1 U2428 ( .A(n3301), .ZN(n3684) );
  XNOR2_X1 U2429 ( .A(n2089), .B(n2998), .ZN(n3009) );
  XNOR2_X1 U2430 ( .A(n3717), .B(n3716), .ZN(n4291) );
  NAND2_X1 U2431 ( .A1(n4301), .A2(n4302), .ZN(n4300) );
  XNOR2_X1 U2432 ( .A(n3702), .B(n4475), .ZN(n4335) );
  NAND2_X1 U2433 ( .A1(n4335), .A2(REG1_REG_14__SCAN_IN), .ZN(n4334) );
  OR2_X1 U2434 ( .A1(n4352), .A2(n2157), .ZN(n2154) );
  OR2_X1 U2435 ( .A1(n4368), .A2(REG1_REG_16__SCAN_IN), .ZN(n2157) );
  NAND2_X1 U2436 ( .A1(n3706), .A2(n2156), .ZN(n2155) );
  INV_X1 U2437 ( .A(n4368), .ZN(n2156) );
  INV_X1 U2438 ( .A(n4354), .ZN(n4380) );
  NAND2_X1 U2439 ( .A1(n3753), .A2(n3752), .ZN(n2079) );
  NAND2_X1 U2440 ( .A1(n2115), .A2(n4444), .ZN(n2113) );
  AOI21_X1 U2441 ( .B1(n2874), .B2(n4444), .A(n2873), .ZN(n3418) );
  AND2_X1 U2442 ( .A1(n4453), .A2(n3736), .ZN(n3954) );
  INV_X1 U2443 ( .A(n3905), .ZN(n3974) );
  OR2_X1 U2444 ( .A1(n2918), .A2(n2877), .ZN(n4457) );
  INV_X1 U2445 ( .A(n2194), .ZN(n2193) );
  OAI21_X1 U2446 ( .B1(n2196), .B2(n3398), .A(n3388), .ZN(n2194) );
  AND2_X1 U2447 ( .A1(n2196), .A2(n3398), .ZN(n2195) );
  NAND2_X1 U2448 ( .A1(n2925), .A2(IR_REG_28__SCAN_IN), .ZN(n2258) );
  AND2_X1 U2449 ( .A1(n2537), .A2(REG3_REG_15__SCAN_IN), .ZN(n2551) );
  AND2_X1 U2450 ( .A1(n2149), .A2(n2148), .ZN(n2999) );
  NAND2_X1 U2451 ( .A1(n4275), .A2(n3694), .ZN(n3695) );
  NAND2_X1 U2452 ( .A1(n4343), .A2(n2054), .ZN(n3705) );
  OR2_X1 U2453 ( .A1(n3585), .A2(n3637), .ZN(n3603) );
  OAI22_X1 U2454 ( .A1(n3898), .A2(n2125), .B1(n2126), .B2(n2865), .ZN(n3822)
         );
  AND2_X1 U2455 ( .A1(n2128), .A2(n3647), .ZN(n2126) );
  NAND2_X1 U2456 ( .A1(n3652), .A2(n2862), .ZN(n2125) );
  NAND2_X1 U2457 ( .A1(n2828), .A2(n2827), .ZN(n2832) );
  AND2_X1 U2458 ( .A1(n2074), .A2(n3593), .ZN(n2070) );
  NAND2_X1 U2459 ( .A1(n2551), .A2(REG3_REG_16__SCAN_IN), .ZN(n2568) );
  OR2_X1 U2460 ( .A1(n3268), .A2(n3530), .ZN(n3281) );
  NOR2_X1 U2461 ( .A1(n3831), .A2(n3812), .ZN(n2139) );
  NOR2_X1 U2462 ( .A1(n2886), .A2(n3486), .ZN(n2131) );
  AND2_X1 U2463 ( .A1(n4390), .A2(n3273), .ZN(n2137) );
  AND3_X1 U2464 ( .A1(n3145), .A2(n2133), .A3(n3157), .ZN(n3156) );
  AND2_X1 U2465 ( .A1(n3083), .A2(n3121), .ZN(n2133) );
  INV_X1 U2466 ( .A(IR_REG_9__SCAN_IN), .ZN(n2081) );
  INV_X1 U2467 ( .A(IR_REG_16__SCAN_IN), .ZN(n2082) );
  INV_X1 U2468 ( .A(IR_REG_13__SCAN_IN), .ZN(n2083) );
  OR2_X1 U2469 ( .A1(n2263), .A2(n2759), .ZN(n2740) );
  INV_X1 U2470 ( .A(IR_REG_23__SCAN_IN), .ZN(n2739) );
  OR2_X1 U2471 ( .A1(n2506), .A2(n2505), .ZN(n2528) );
  OR2_X1 U2472 ( .A1(n2506), .A2(IR_REG_10__SCAN_IN), .ZN(n2471) );
  OR2_X1 U2473 ( .A1(n2438), .A2(IR_REG_9__SCAN_IN), .ZN(n2506) );
  INV_X1 U2474 ( .A(IR_REG_2__SCAN_IN), .ZN(n4108) );
  NAND2_X1 U2475 ( .A1(n2373), .A2(n2188), .ZN(n2187) );
  NOR2_X1 U2476 ( .A1(n2189), .A2(n3090), .ZN(n2188) );
  INV_X1 U2477 ( .A(n2182), .ZN(n2181) );
  OAI21_X1 U2478 ( .B1(n2519), .B2(n2183), .A(n2518), .ZN(n2182) );
  NAND2_X1 U2479 ( .A1(n2184), .A2(n3250), .ZN(n2183) );
  NAND2_X1 U2480 ( .A1(n2186), .A2(n3250), .ZN(n2185) );
  INV_X1 U2481 ( .A(n2519), .ZN(n2186) );
  NOR2_X1 U2482 ( .A1(n3218), .A2(n2198), .ZN(n2197) );
  INV_X1 U2483 ( .A(n2200), .ZN(n2198) );
  NAND2_X1 U2484 ( .A1(n3194), .A2(n3195), .ZN(n2200) );
  NAND2_X1 U2485 ( .A1(n3197), .A2(n2201), .ZN(n2199) );
  NAND2_X1 U2486 ( .A1(n2203), .A2(n2202), .ZN(n2201) );
  INV_X1 U2487 ( .A(n3195), .ZN(n2202) );
  INV_X1 U2488 ( .A(n3194), .ZN(n2203) );
  AOI21_X1 U2489 ( .B1(n2167), .B2(n2169), .A(n2165), .ZN(n2164) );
  INV_X1 U2490 ( .A(n3482), .ZN(n2165) );
  AND2_X1 U2491 ( .A1(n2496), .A2(n2495), .ZN(n3329) );
  XNOR2_X1 U2492 ( .A(n2272), .B(n2689), .ZN(n2290) );
  OAI22_X1 U2493 ( .A1(n2993), .A2(n2339), .B1(n2713), .B2(n4436), .ZN(n2272)
         );
  INV_X1 U2494 ( .A(n3025), .ZN(n2312) );
  NAND2_X1 U2495 ( .A1(n2192), .A2(n2563), .ZN(n3396) );
  NAND2_X1 U2496 ( .A1(n2536), .A2(n2535), .ZN(n2192) );
  INV_X1 U2497 ( .A(n4464), .ZN(n2757) );
  AND4_X1 U2498 ( .A1(n2527), .A2(n2526), .A3(n2525), .A4(n2524), .ZN(n2813)
         );
  AND4_X1 U2499 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n3301)
         );
  NAND2_X1 U2500 ( .A1(n2295), .A2(REG1_REG_1__SCAN_IN), .ZN(n2110) );
  NAND2_X1 U2501 ( .A1(n2975), .A2(n2944), .ZN(n2143) );
  NOR2_X1 U2502 ( .A1(n4248), .A2(n2330), .ZN(n2162) );
  NOR2_X1 U2503 ( .A1(n2257), .A2(IR_REG_5__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U2504 ( .A1(n4251), .A2(n2043), .ZN(n3013) );
  OR2_X1 U2505 ( .A1(n4256), .A2(n3003), .ZN(n2153) );
  NAND2_X1 U2506 ( .A1(n4271), .A2(n3693), .ZN(n4276) );
  NAND2_X1 U2507 ( .A1(n4276), .A2(n4277), .ZN(n4275) );
  XNOR2_X1 U2508 ( .A(n3695), .B(n3716), .ZN(n4289) );
  NAND2_X1 U2509 ( .A1(n4289), .A2(REG1_REG_10__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U2510 ( .A1(n4297), .A2(n3697), .ZN(n3698) );
  OAI21_X1 U2511 ( .B1(n4330), .B2(n2095), .A(n2094), .ZN(n4339) );
  NAND2_X1 U2512 ( .A1(n2096), .A2(REG2_REG_14__SCAN_IN), .ZN(n2095) );
  NAND2_X1 U2513 ( .A1(n3726), .A2(n2096), .ZN(n2094) );
  INV_X1 U2514 ( .A(n4340), .ZN(n2096) );
  NOR2_X1 U2515 ( .A1(n4330), .A2(n4331), .ZN(n4329) );
  NAND2_X1 U2516 ( .A1(n4364), .A2(n2091), .ZN(n4374) );
  NAND2_X1 U2517 ( .A1(n4469), .A2(n3970), .ZN(n2091) );
  NOR2_X1 U2518 ( .A1(n2114), .A2(n4396), .ZN(n2112) );
  AND2_X1 U2519 ( .A1(n2036), .A2(n2116), .ZN(n2114) );
  NAND2_X1 U2520 ( .A1(n2116), .A2(n2119), .ZN(n2115) );
  NAND2_X1 U2521 ( .A1(n3744), .A2(n3757), .ZN(n2119) );
  INV_X1 U2522 ( .A(n2867), .ZN(n3775) );
  INV_X1 U2523 ( .A(n3603), .ZN(n3772) );
  AND2_X1 U2524 ( .A1(n3586), .A2(DATAI_25_), .ZN(n3812) );
  AND4_X1 U2525 ( .A1(n2644), .A2(n2643), .A3(n2642), .A4(n2641), .ZN(n3872)
         );
  NAND2_X1 U2526 ( .A1(n2654), .A2(REG3_REG_24__SCAN_IN), .ZN(n2669) );
  AND2_X1 U2527 ( .A1(n2639), .A2(REG3_REG_23__SCAN_IN), .ZN(n2654) );
  NOR2_X1 U2528 ( .A1(n2632), .A2(n2631), .ZN(n2639) );
  OR2_X1 U2529 ( .A1(n3898), .A2(n3650), .ZN(n2127) );
  AND4_X1 U2530 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n3896)
         );
  NAND2_X1 U2531 ( .A1(n2605), .A2(REG3_REG_20__SCAN_IN), .ZN(n2618) );
  NOR2_X1 U2532 ( .A1(n2593), .A2(n4083), .ZN(n2605) );
  NAND2_X1 U2533 ( .A1(n2581), .A2(REG3_REG_18__SCAN_IN), .ZN(n2593) );
  INV_X1 U2534 ( .A(n2568), .ZN(n2580) );
  AOI21_X1 U2535 ( .B1(n2104), .B2(n2106), .A(n2101), .ZN(n2100) );
  INV_X1 U2536 ( .A(n3645), .ZN(n2101) );
  OR2_X1 U2537 ( .A1(n3315), .A2(n3356), .ZN(n2816) );
  NAND2_X1 U2538 ( .A1(n3354), .A2(n2854), .ZN(n2103) );
  INV_X1 U2539 ( .A(n3604), .ZN(n3368) );
  NOR2_X1 U2540 ( .A1(n3295), .A2(n2884), .ZN(n3296) );
  AND2_X1 U2541 ( .A1(n2137), .A2(n2136), .ZN(n2135) );
  INV_X1 U2542 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2521) );
  NOR2_X1 U2543 ( .A1(n2522), .A2(n2521), .ZN(n2537) );
  OR2_X1 U2544 ( .A1(n2061), .A2(n2811), .ZN(n2057) );
  INV_X1 U2545 ( .A(n2062), .ZN(n2061) );
  NAND2_X1 U2546 ( .A1(n3296), .A2(n2135), .ZN(n3348) );
  INV_X1 U2547 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3336) );
  OR2_X1 U2548 ( .A1(n2484), .A2(n2483), .ZN(n2497) );
  OR2_X1 U2549 ( .A1(n2497), .A2(n3336), .ZN(n2522) );
  NAND2_X1 U2550 ( .A1(n2464), .A2(REG3_REG_11__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U2551 ( .A1(n3299), .A2(n3525), .ZN(n2851) );
  OAI21_X1 U2552 ( .B1(n3204), .B2(n3203), .A(n3567), .ZN(n3299) );
  NOR2_X1 U2553 ( .A1(n2431), .A2(n3219), .ZN(n2444) );
  AND2_X1 U2554 ( .A1(n2444), .A2(REG3_REG_10__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U2555 ( .A1(n2121), .A2(n3559), .ZN(n3236) );
  NOR2_X1 U2556 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
  INV_X1 U2557 ( .A(n2849), .ZN(n2124) );
  INV_X1 U2558 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2414) );
  OR2_X1 U2559 ( .A1(n2415), .A2(n2414), .ZN(n2431) );
  INV_X1 U2560 ( .A(n3686), .ZN(n3221) );
  NAND2_X1 U2561 ( .A1(n2848), .A2(n3551), .ZN(n3173) );
  INV_X1 U2562 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2375) );
  NOR2_X1 U2563 ( .A1(n2376), .A2(n2375), .ZN(n2397) );
  AND4_X1 U2564 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(n3151)
         );
  NAND2_X1 U2565 ( .A1(n2356), .A2(REG3_REG_5__SCAN_IN), .ZN(n2376) );
  OAI21_X1 U2566 ( .B1(n3076), .B2(n2847), .A(n3549), .ZN(n3120) );
  NAND2_X1 U2567 ( .A1(n3145), .A2(n3083), .ZN(n3126) );
  NAND2_X1 U2568 ( .A1(n2317), .A2(n2316), .ZN(n3544) );
  OR2_X1 U2569 ( .A1(n3586), .A2(n2147), .ZN(n2317) );
  NOR2_X1 U2570 ( .A1(n4504), .A2(n3544), .ZN(n3145) );
  NAND2_X1 U2571 ( .A1(n2097), .A2(n2844), .ZN(n3106) );
  NAND2_X1 U2572 ( .A1(n4420), .A2(n2842), .ZN(n2098) );
  INV_X1 U2573 ( .A(n4423), .ZN(n4447) );
  NOR2_X1 U2574 ( .A1(n3795), .A2(n3775), .ZN(n3767) );
  INV_X1 U2575 ( .A(n2139), .ZN(n3814) );
  NAND2_X1 U2576 ( .A1(n2139), .A2(n3513), .ZN(n3795) );
  AND2_X1 U2577 ( .A1(n3931), .A2(n2049), .ZN(n3851) );
  INV_X1 U2578 ( .A(n2886), .ZN(n3888) );
  NAND2_X1 U2579 ( .A1(n3931), .A2(n2131), .ZN(n3887) );
  NAND2_X1 U2580 ( .A1(n3931), .A2(n3907), .ZN(n3906) );
  NOR2_X1 U2581 ( .A1(n3965), .A2(n3946), .ZN(n3940) );
  AND2_X1 U2582 ( .A1(n3940), .A2(n3929), .ZN(n3931) );
  OR2_X1 U2583 ( .A1(n3964), .A2(n2885), .ZN(n3965) );
  NOR2_X1 U2584 ( .A1(n4171), .A2(n3400), .ZN(n3373) );
  NAND2_X1 U2585 ( .A1(n3296), .A2(n2137), .ZN(n3289) );
  AND2_X1 U2586 ( .A1(n3296), .A2(n4390), .ZN(n4400) );
  OR2_X1 U2587 ( .A1(n3234), .A2(n3209), .ZN(n3295) );
  OR2_X1 U2588 ( .A1(n4435), .A2(n3107), .ZN(n4504) );
  NOR2_X1 U2589 ( .A1(n2880), .A2(n3067), .ZN(n2893) );
  NAND2_X1 U2590 ( .A1(n2740), .A2(n2739), .ZN(n2738) );
  OAI21_X1 U2591 ( .B1(n2740), .B2(n2739), .A(n2738), .ZN(n2919) );
  NAND2_X1 U2592 ( .A1(n2265), .A2(n2264), .ZN(n2838) );
  NAND2_X1 U2593 ( .A1(n2382), .A2(n2099), .ZN(n2363) );
  AND4_X1 U2594 ( .A1(n2637), .A2(n2636), .A3(n2635), .A4(n2634), .ZN(n3880)
         );
  INV_X1 U2595 ( .A(n3426), .ZN(n3430) );
  NAND2_X1 U2596 ( .A1(n2295), .A2(REG1_REG_2__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2597 ( .A1(n2172), .A2(n2173), .ZN(n3436) );
  NAND2_X1 U2598 ( .A1(n2579), .A2(n2037), .ZN(n2172) );
  INV_X1 U2599 ( .A(n3685), .ZN(n3238) );
  XNOR2_X1 U2600 ( .A(n2290), .B(n2291), .ZN(n2984) );
  NAND2_X1 U2601 ( .A1(n3480), .A2(n3484), .ZN(n3444) );
  NAND2_X1 U2602 ( .A1(n3252), .A2(n3249), .ZN(n2180) );
  AOI21_X1 U2603 ( .B1(n2664), .B2(n2206), .A(n2205), .ZN(n2204) );
  AND2_X1 U2604 ( .A1(n2667), .A2(n2666), .ZN(n2205) );
  AND4_X1 U2605 ( .A1(n2338), .A2(n2337), .A3(n2336), .A4(n2335), .ZN(n2796)
         );
  OAI21_X1 U2606 ( .B1(n3426), .B2(n2667), .A(n2666), .ZN(n3471) );
  NAND2_X1 U2607 ( .A1(n3042), .A2(n2349), .ZN(n3053) );
  NAND2_X1 U2608 ( .A1(n2199), .A2(n2200), .ZN(n3217) );
  INV_X1 U2609 ( .A(n2882), .ZN(n4450) );
  INV_X1 U2610 ( .A(n4402), .ZN(n4390) );
  AND4_X1 U2611 ( .A1(n2572), .A2(n2571), .A3(n2570), .A4(n2569), .ZN(n3949)
         );
  INV_X1 U2612 ( .A(n2210), .ZN(n2174) );
  AND2_X1 U2613 ( .A1(n2774), .A2(n2762), .ZN(n3500) );
  AND4_X1 U2614 ( .A1(n2674), .A2(n2673), .A3(n2672), .A4(n2671), .ZN(n3824)
         );
  INV_X1 U2615 ( .A(n3487), .ZN(n3514) );
  INV_X1 U2616 ( .A(n3488), .ZN(n3515) );
  AOI21_X1 U2617 ( .B1(n3451), .B2(n3452), .A(n3454), .ZN(n3504) );
  INV_X1 U2618 ( .A(n3496), .ZN(n3520) );
  AND4_X1 U2619 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n3467)
         );
  INV_X1 U2620 ( .A(n3500), .ZN(n3512) );
  INV_X1 U2621 ( .A(n3503), .ZN(n3518) );
  NAND4_X1 U2622 ( .A1(n2702), .A2(n2701), .A3(n2700), .A4(n2699), .ZN(n3788)
         );
  NAND4_X1 U2623 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n3848)
         );
  NAND4_X1 U2624 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n3947)
         );
  INV_X1 U2625 ( .A(n4391), .ZN(n3683) );
  INV_X1 U2626 ( .A(n3151), .ZN(n3240) );
  INV_X1 U2627 ( .A(n2796), .ZN(n3123) );
  NOR2_X1 U2628 ( .A1(n2323), .A2(n2212), .ZN(n2324) );
  NAND2_X1 U2629 ( .A1(n2321), .A2(n2320), .ZN(n2323) );
  INV_X1 U2630 ( .A(n3137), .ZN(n4424) );
  OR2_X1 U2631 ( .A1(n2354), .A2(n2283), .ZN(n2279) );
  NOR2_X1 U2632 ( .A1(n2922), .A2(n2923), .ZN(n2974) );
  NAND2_X1 U2633 ( .A1(n2142), .A2(n2146), .ZN(n2945) );
  NAND2_X1 U2634 ( .A1(n2143), .A2(n2998), .ZN(n2142) );
  AND2_X1 U2635 ( .A1(n3032), .A2(REG1_REG_4__SCAN_IN), .ZN(n3038) );
  OAI22_X1 U2636 ( .A1(n3033), .A2(n3012), .B1(n3011), .B2(n3041), .ZN(n4252)
         );
  XNOR2_X1 U2637 ( .A(n3013), .B(n4264), .ZN(n4261) );
  XNOR2_X1 U2638 ( .A(n3002), .B(n4264), .ZN(n4257) );
  NOR2_X1 U2639 ( .A1(n4257), .A2(n2374), .ZN(n4256) );
  INV_X1 U2640 ( .A(n2153), .ZN(n3691) );
  XNOR2_X1 U2641 ( .A(n3692), .B(n4485), .ZN(n4272) );
  NAND2_X1 U2642 ( .A1(n4266), .A2(n3714), .ZN(n4279) );
  NAND2_X1 U2643 ( .A1(n4290), .A2(n3718), .ZN(n4301) );
  XNOR2_X1 U2644 ( .A(n3698), .B(n4478), .ZN(n4314) );
  NAND2_X1 U2645 ( .A1(n4308), .A2(n3723), .ZN(n4319) );
  NAND2_X1 U2646 ( .A1(n4334), .A2(n3703), .ZN(n4344) );
  NAND2_X1 U2647 ( .A1(n4344), .A2(n4345), .ZN(n4343) );
  NAND2_X1 U2648 ( .A1(n4350), .A2(n2553), .ZN(n4349) );
  AND3_X1 U2649 ( .A1(n2155), .A2(n2154), .A3(n2056), .ZN(n4381) );
  NAND2_X1 U2650 ( .A1(n2269), .A2(n2268), .ZN(n3736) );
  OR2_X1 U2651 ( .A1(n2698), .A2(n2705), .ZN(n3768) );
  AND2_X1 U2652 ( .A1(n2072), .A2(n2075), .ZN(n3885) );
  NAND2_X1 U2653 ( .A1(n3904), .A2(n3593), .ZN(n2072) );
  NAND2_X1 U2654 ( .A1(n3296), .A2(n2134), .ZN(n4171) );
  AND2_X1 U2655 ( .A1(n2135), .A2(n2814), .ZN(n2134) );
  NAND2_X1 U2656 ( .A1(n2060), .A2(n2064), .ZN(n3287) );
  NAND2_X1 U2657 ( .A1(n4386), .A2(n2065), .ZN(n2060) );
  AND2_X1 U2658 ( .A1(n2066), .A2(n2068), .ZN(n3272) );
  NAND2_X1 U2659 ( .A1(n4386), .A2(n4387), .ZN(n2066) );
  NAND2_X1 U2660 ( .A1(n3117), .A2(n3116), .ZN(n3905) );
  INV_X1 U2661 ( .A(n4558), .ZN(n4556) );
  AOI21_X1 U2662 ( .B1(n3991), .B2(n4537), .A(n3993), .ZN(n2140) );
  AND2_X2 U2663 ( .A1(n2893), .A2(n3069), .ZN(n4544) );
  INV_X1 U2664 ( .A(n2226), .ZN(n2130) );
  INV_X1 U2665 ( .A(n2209), .ZN(n2207) );
  XNOR2_X1 U2666 ( .A(n2247), .B(IR_REG_26__SCAN_IN), .ZN(n2912) );
  INV_X1 U2667 ( .A(n2838), .ZN(n3670) );
  NAND2_X1 U2668 ( .A1(n2257), .A2(IR_REG_31__SCAN_IN), .ZN(n2302) );
  OAI211_X1 U2669 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_1__SCAN_IN), .A(n2092), 
        .B(n2257), .ZN(n2938) );
  NAND2_X1 U2670 ( .A1(n2031), .A2(IR_REG_0__SCAN_IN), .ZN(n2092) );
  NAND2_X1 U2671 ( .A1(n2155), .A2(n2154), .ZN(n4369) );
  AOI211_X1 U2672 ( .C1(n4438), .C2(n2038), .A(n3420), .B(n3419), .ZN(n3421)
         );
  NAND2_X1 U2673 ( .A1(n2038), .A2(n2889), .ZN(n2890) );
  INV_X1 U2674 ( .A(n4168), .ZN(n2889) );
  NAND2_X1 U2675 ( .A1(n2038), .A2(n2896), .ZN(n2897) );
  OR2_X1 U2676 ( .A1(n2238), .A2(n2236), .ZN(n2275) );
  OAI21_X1 U2677 ( .B1(n3406), .B2(n2047), .A(n2204), .ZN(n3451) );
  NAND2_X1 U2678 ( .A1(n3683), .A2(n3267), .ZN(n2016) );
  OR2_X1 U2679 ( .A1(n3426), .A2(n2664), .ZN(n2017) );
  XNOR2_X1 U2680 ( .A(n2302), .B(IR_REG_2__SCAN_IN), .ZN(n4232) );
  AND2_X1 U2681 ( .A1(n3091), .A2(n2409), .ZN(n2018) );
  NAND4_X1 U2682 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(n3805)
         );
  INV_X1 U2683 ( .A(n3805), .ZN(n3779) );
  OR2_X1 U2684 ( .A1(n2071), .A2(n2824), .ZN(n2019) );
  AND2_X1 U2685 ( .A1(n3884), .A2(n3907), .ZN(n3650) );
  OR2_X1 U2686 ( .A1(n2210), .A2(n2048), .ZN(n2020) );
  OR2_X1 U2687 ( .A1(n3427), .A2(n3428), .ZN(n2021) );
  AND2_X1 U2688 ( .A1(n2131), .A2(n2825), .ZN(n2022) );
  NAND2_X2 U2689 ( .A1(n2256), .A2(n3073), .ZN(n2339) );
  OR2_X1 U2690 ( .A1(n2220), .A2(n2219), .ZN(n2023) );
  AND2_X1 U2691 ( .A1(n3000), .A2(n4231), .ZN(n2024) );
  NOR2_X1 U2692 ( .A1(n3407), .A2(n3408), .ZN(n3406) );
  AND2_X1 U2693 ( .A1(n3776), .A2(n2887), .ZN(n3742) );
  NAND2_X1 U2694 ( .A1(n2102), .A2(n2100), .ZN(n3915) );
  AND2_X1 U2695 ( .A1(n2127), .A2(n2128), .ZN(n2025) );
  AND2_X1 U2696 ( .A1(n4391), .A2(n3273), .ZN(n2026) );
  INV_X1 U2697 ( .A(n4248), .ZN(n2163) );
  AND2_X1 U2698 ( .A1(n3744), .A2(n3637), .ZN(n2027) );
  OR2_X1 U2699 ( .A1(n2810), .A2(n2026), .ZN(n2028) );
  AND4_X1 U2700 ( .A1(n2085), .A2(n2087), .A3(n2086), .A4(n4491), .ZN(n2029)
         );
  INV_X1 U2701 ( .A(n3706), .ZN(n2158) );
  AND2_X1 U2702 ( .A1(n2924), .A2(n2229), .ZN(n2030) );
  NAND2_X1 U2703 ( .A1(n2109), .A2(n2108), .ZN(n2843) );
  AND2_X1 U2704 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2031)
         );
  AND2_X1 U2705 ( .A1(n2944), .A2(n2147), .ZN(n2032) );
  OR2_X1 U2706 ( .A1(n2275), .A2(n2237), .ZN(n2033) );
  AND2_X1 U2707 ( .A1(n2159), .A2(n2158), .ZN(n2034) );
  AND2_X1 U2708 ( .A1(n2227), .A2(n2229), .ZN(n2035) );
  NAND2_X1 U2709 ( .A1(n2120), .A2(n3756), .ZN(n2036) );
  INV_X1 U2710 ( .A(IR_REG_29__SCAN_IN), .ZN(n2233) );
  NAND2_X1 U2711 ( .A1(n2180), .A2(n3250), .ZN(n3260) );
  NAND2_X2 U2712 ( .A1(n2270), .A2(n2256), .ZN(n2713) );
  AND3_X1 U2713 ( .A1(n2536), .A2(n2196), .A3(n2535), .ZN(n3387) );
  INV_X1 U2714 ( .A(n3310), .ZN(n2179) );
  NAND2_X1 U2715 ( .A1(n3931), .A2(n2022), .ZN(n2132) );
  AND2_X1 U2716 ( .A1(n2176), .A2(n2211), .ZN(n2037) );
  AND2_X1 U2717 ( .A1(n3760), .A2(n2888), .ZN(n2038) );
  NAND2_X1 U2718 ( .A1(n2076), .A2(n2215), .ZN(n3938) );
  AND2_X1 U2719 ( .A1(n2175), .A2(n2174), .ZN(n2039) );
  NAND2_X1 U2720 ( .A1(n2103), .A2(n3523), .ZN(n3367) );
  INV_X1 U2721 ( .A(IR_REG_25__SCAN_IN), .ZN(n2227) );
  AND2_X1 U2722 ( .A1(n2383), .A2(n2218), .ZN(n2386) );
  AND3_X1 U2723 ( .A1(n2749), .A2(n2750), .A3(n3496), .ZN(n2040) );
  NOR2_X1 U2724 ( .A1(n4329), .A2(n3726), .ZN(n2041) );
  AND2_X1 U2725 ( .A1(n3896), .A2(n3888), .ZN(n2042) );
  OR2_X1 U2726 ( .A1(n4489), .A2(n3129), .ZN(n2043) );
  INV_X1 U2727 ( .A(IR_REG_7__SCAN_IN), .ZN(n2087) );
  NAND2_X1 U2728 ( .A1(n2166), .A2(n2164), .ZN(n3480) );
  INV_X1 U2729 ( .A(n2824), .ZN(n2074) );
  INV_X1 U2730 ( .A(n3650), .ZN(n2862) );
  NOR2_X1 U2731 ( .A1(n2206), .A2(n2666), .ZN(n2044) );
  NOR2_X1 U2732 ( .A1(n2604), .A2(n2603), .ZN(n2045) );
  NAND2_X1 U2733 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  INV_X1 U2734 ( .A(IR_REG_5__SCAN_IN), .ZN(n2217) );
  AND2_X1 U2735 ( .A1(n2567), .A2(n2566), .ZN(n2046) );
  OR2_X1 U2736 ( .A1(n2021), .A2(n2044), .ZN(n2047) );
  XNOR2_X1 U2737 ( .A(n2243), .B(n2242), .ZN(n2721) );
  INV_X1 U2738 ( .A(n3288), .ZN(n2136) );
  INV_X1 U2739 ( .A(n2751), .ZN(n2742) );
  NAND2_X1 U2740 ( .A1(n2199), .A2(n2197), .ZN(n3215) );
  AND2_X1 U2741 ( .A1(n2592), .A2(n2591), .ZN(n2048) );
  NAND2_X1 U2742 ( .A1(n2187), .A2(n3091), .ZN(n3164) );
  AND2_X1 U2743 ( .A1(n3586), .A2(DATAI_22_), .ZN(n3873) );
  INV_X1 U2744 ( .A(n3847), .ZN(n3853) );
  AND2_X1 U2745 ( .A1(n3586), .A2(DATAI_23_), .ZN(n3847) );
  AND2_X1 U2746 ( .A1(n3853), .A2(n2022), .ZN(n2049) );
  INV_X1 U2747 ( .A(n3594), .ZN(n2075) );
  AND2_X1 U2748 ( .A1(n3156), .A2(n3174), .ZN(n3178) );
  AND2_X1 U2749 ( .A1(n3145), .A2(n2133), .ZN(n2050) );
  OR2_X1 U2750 ( .A1(n4477), .A2(n3700), .ZN(n2051) );
  AND2_X1 U2751 ( .A1(n4448), .A2(n2769), .ZN(n4537) );
  INV_X1 U2752 ( .A(n2790), .ZN(n2993) );
  OR2_X1 U2753 ( .A1(n4385), .A2(n4467), .ZN(n2052) );
  AND2_X1 U2754 ( .A1(n2870), .A2(n2869), .ZN(n4396) );
  NOR2_X1 U2755 ( .A1(n2024), .A2(n3038), .ZN(n2053) );
  OR2_X1 U2756 ( .A1(n4348), .A2(n3704), .ZN(n2054) );
  INV_X1 U2757 ( .A(n2810), .ZN(n2068) );
  AND2_X1 U2758 ( .A1(n2228), .A2(n2207), .ZN(n2055) );
  INV_X1 U2759 ( .A(n2998), .ZN(n2147) );
  OR2_X1 U2760 ( .A1(n3730), .A2(REG1_REG_17__SCAN_IN), .ZN(n2056) );
  INV_X1 U2761 ( .A(IR_REG_8__SCAN_IN), .ZN(n2086) );
  NAND2_X2 U2762 ( .A1(n2058), .A2(n2057), .ZN(n3341) );
  OR2_X2 U2763 ( .A1(n4386), .A2(n2059), .ZN(n2058) );
  NAND2_X2 U2764 ( .A1(n2073), .A2(n2831), .ZN(n3828) );
  OR2_X2 U2765 ( .A1(n3860), .A2(n2832), .ZN(n2073) );
  AOI21_X2 U2766 ( .B1(n3938), .B2(n3945), .A(n2819), .ZN(n3914) );
  AND2_X2 U2767 ( .A1(n2078), .A2(n2077), .ZN(n3957) );
  NAND2_X1 U2768 ( .A1(n2079), .A2(n3755), .ZN(n3758) );
  OAI22_X2 U2769 ( .A1(n3765), .A2(n2837), .B1(n3511), .B2(n2867), .ZN(n3753)
         );
  NAND4_X1 U2770 ( .A1(n2558), .A2(n2083), .A3(n2082), .A4(n2081), .ZN(n2219)
         );
  NAND2_X1 U2771 ( .A1(n2792), .A2(n2844), .ZN(n3099) );
  MUX2_X1 U2772 ( .A(n2941), .B(DATAI_1_), .S(n2301), .Z(n4421) );
  NAND3_X1 U2773 ( .A1(n4384), .A2(n4383), .A3(n2052), .ZN(U3258) );
  MUX2_X1 U2774 ( .A(REG2_REG_1__SCAN_IN), .B(n2235), .S(n2938), .Z(n2922) );
  XNOR2_X1 U2775 ( .A(n3725), .B(n4475), .ZN(n4330) );
  OAI21_X2 U2776 ( .B1(n3353), .B2(n2817), .A(n2816), .ZN(n3366) );
  OAI22_X2 U2777 ( .A1(n3208), .A2(n2807), .B1(n3238), .B2(n3220), .ZN(n3298)
         );
  NAND2_X1 U2778 ( .A1(n2252), .A2(n2221), .ZN(n2261) );
  NAND2_X1 U2779 ( .A1(n2841), .A2(n4429), .ZN(n4428) );
  NOR2_X4 U2780 ( .A1(n2438), .A2(n2023), .ZN(n2240) );
  NAND2_X1 U2781 ( .A1(n3994), .A2(n2140), .ZN(n4185) );
  NAND2_X1 U2782 ( .A1(n2098), .A2(n2843), .ZN(n2845) );
  OAI21_X1 U2783 ( .B1(n4420), .B2(n2842), .A(n2098), .ZN(n4433) );
  INV_X1 U2784 ( .A(n2845), .ZN(n2097) );
  NAND2_X1 U2785 ( .A1(n3354), .A2(n2104), .ZN(n2102) );
  OR2_X2 U2786 ( .A1(n2319), .A2(n2235), .ZN(n2107) );
  NAND2_X1 U2787 ( .A1(n3771), .A2(n2112), .ZN(n2111) );
  OAI211_X1 U2788 ( .C1(n3771), .C2(n2113), .A(n3750), .B(n2111), .ZN(n3993)
         );
  NAND2_X1 U2789 ( .A1(n3771), .A2(n2868), .ZN(n3745) );
  NAND2_X1 U2790 ( .A1(n2848), .A2(n2122), .ZN(n2121) );
  NAND4_X1 U2791 ( .A1(n2240), .A2(n2241), .A3(n2208), .A4(n2226), .ZN(n2232)
         );
  NAND4_X1 U2792 ( .A1(n2240), .A2(n2241), .A3(n2208), .A4(n2129), .ZN(n3423)
         );
  INV_X1 U2793 ( .A(n2132), .ZN(n3863) );
  NAND4_X1 U2794 ( .A1(n2240), .A2(n2241), .A3(n2035), .A4(n2226), .ZN(n2138)
         );
  NAND4_X1 U2795 ( .A1(n2240), .A2(n2241), .A3(n2226), .A4(n2227), .ZN(n2246)
         );
  INV_X1 U2796 ( .A(n2228), .ZN(n2244) );
  OR2_X1 U2797 ( .A1(n2975), .A2(n2147), .ZN(n2141) );
  NAND3_X1 U2798 ( .A1(n2146), .A2(n2144), .A3(n2141), .ZN(n2149) );
  NAND2_X1 U2799 ( .A1(n2975), .A2(n2032), .ZN(n2146) );
  NAND2_X1 U2800 ( .A1(n2975), .A2(n2944), .ZN(n2150) );
  INV_X1 U2801 ( .A(n2149), .ZN(n2997) );
  NAND2_X1 U2802 ( .A1(n2150), .A2(n2998), .ZN(n2148) );
  OR2_X1 U2803 ( .A1(n4352), .A2(REG1_REG_16__SCAN_IN), .ZN(n2159) );
  INV_X1 U2804 ( .A(n2159), .ZN(n4351) );
  NAND2_X1 U2805 ( .A1(n2024), .A2(n2163), .ZN(n2160) );
  NAND2_X1 U2806 ( .A1(n3032), .A2(n2162), .ZN(n2161) );
  NAND2_X1 U2807 ( .A1(n2161), .A2(n2160), .ZN(n4247) );
  OAI21_X1 U2808 ( .B1(n2579), .B2(n2169), .A(n2167), .ZN(n3481) );
  NAND2_X1 U2809 ( .A1(n2579), .A2(n2167), .ZN(n2166) );
  OAI21_X1 U2810 ( .B1(n3252), .B2(n2185), .A(n2181), .ZN(n3313) );
  NAND2_X1 U2811 ( .A1(n2177), .A2(n2178), .ZN(n2533) );
  NAND2_X1 U2812 ( .A1(n3252), .A2(n2181), .ZN(n2177) );
  NAND2_X1 U2813 ( .A1(n2187), .A2(n2018), .ZN(n3166) );
  NAND2_X1 U2814 ( .A1(n2373), .A2(n2372), .ZN(n3089) );
  INV_X1 U2815 ( .A(n2372), .ZN(n2189) );
  NAND2_X1 U2816 ( .A1(n2190), .A2(n2191), .ZN(n3463) );
  NAND3_X1 U2817 ( .A1(n2536), .A2(n2193), .A3(n2535), .ZN(n2190) );
  INV_X1 U2818 ( .A(n2563), .ZN(n2196) );
  NOR2_X1 U2819 ( .A1(n3406), .A2(n2021), .ZN(n3426) );
  NAND2_X1 U2820 ( .A1(n3538), .A2(n2843), .ZN(n2841) );
  NAND2_X1 U2821 ( .A1(n3023), .A2(n2314), .ZN(n3043) );
  OR2_X1 U2822 ( .A1(n2319), .A2(n2277), .ZN(n2278) );
  NAND2_X1 U2823 ( .A1(n2238), .A2(n4226), .ZN(n2354) );
  AND2_X1 U2824 ( .A1(n2578), .A2(n2214), .ZN(n2210) );
  OR2_X1 U2825 ( .A1(n2578), .A2(n2214), .ZN(n2211) );
  INV_X1 U2826 ( .A(n3464), .ZN(n2578) );
  AND2_X1 U2827 ( .A1(n3843), .A2(n2826), .ZN(n3868) );
  INV_X1 U2828 ( .A(n3868), .ZN(n2828) );
  INV_X1 U2829 ( .A(IR_REG_28__SCAN_IN), .ZN(n2760) );
  AND2_X1 U2830 ( .A1(n3731), .A2(REG2_REG_18__SCAN_IN), .ZN(n2213) );
  INV_X1 U2831 ( .A(n3756), .ZN(n3757) );
  INV_X1 U2832 ( .A(IR_REG_31__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U2833 ( .A1(n2577), .A2(n2576), .ZN(n2214) );
  INV_X1 U2834 ( .A(n3644), .ZN(n2856) );
  OR2_X1 U2835 ( .A1(n3679), .A2(n2885), .ZN(n2215) );
  INV_X1 U2836 ( .A(n3710), .ZN(n4480) );
  INV_X1 U2837 ( .A(n2565), .ZN(n2566) );
  INV_X1 U2838 ( .A(IR_REG_17__SCAN_IN), .ZN(n2223) );
  AND2_X1 U2839 ( .A1(n3282), .A2(n3280), .ZN(n3529) );
  INV_X1 U2840 ( .A(IR_REG_21__SCAN_IN), .ZN(n2221) );
  INV_X1 U2841 ( .A(n2829), .ZN(n2827) );
  NAND2_X1 U2842 ( .A1(n3586), .A2(DATAI_3_), .ZN(n2316) );
  INV_X1 U2843 ( .A(n4287), .ZN(n3716) );
  INV_X1 U2844 ( .A(n2830), .ZN(n2831) );
  AND2_X1 U2845 ( .A1(n3677), .A2(n2825), .ZN(n2863) );
  OR2_X1 U2846 ( .A1(n3467), .A2(n3390), .ZN(n3645) );
  NAND2_X1 U2847 ( .A1(n3776), .A2(n3754), .ZN(n3755) );
  INV_X1 U2848 ( .A(IR_REG_26__SCAN_IN), .ZN(n2229) );
  INV_X1 U2849 ( .A(n3165), .ZN(n2409) );
  INV_X1 U2850 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2483) );
  NOR2_X1 U2851 ( .A1(n2697), .A2(n4076), .ZN(n2705) );
  OR2_X1 U2852 ( .A1(n2669), .A2(n3456), .ZN(n2680) );
  OR2_X1 U2853 ( .A1(n2618), .A2(n3445), .ZN(n2632) );
  AND2_X1 U2854 ( .A1(n3959), .A2(n3498), .ZN(n2819) );
  OR2_X1 U2855 ( .A1(n3681), .A2(n3347), .ZN(n2815) );
  INV_X1 U2856 ( .A(n4537), .ZN(n3992) );
  INV_X1 U2857 ( .A(n2844), .ZN(n3105) );
  INV_X1 U2858 ( .A(IR_REG_30__SCAN_IN), .ZN(n2230) );
  INV_X1 U2859 ( .A(n3180), .ZN(n3174) );
  INV_X1 U2860 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4083) );
  INV_X1 U2861 ( .A(n3107), .ZN(n3027) );
  OR2_X1 U2862 ( .A1(n2763), .A2(n3815), .ZN(n2672) );
  NAND2_X1 U2863 ( .A1(n2248), .A2(n2912), .ZN(n2256) );
  INV_X1 U2864 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3219) );
  NOR2_X1 U2865 ( .A1(n4375), .A2(n4374), .ZN(n4373) );
  INV_X1 U2866 ( .A(n3828), .ZN(n3830) );
  AND2_X1 U2867 ( .A1(n3534), .A2(n3522), .ZN(n3617) );
  INV_X1 U2868 ( .A(n4438), .ZN(n3968) );
  AND2_X1 U2869 ( .A1(n2724), .A2(n2721), .ZN(n2725) );
  INV_X1 U2870 ( .A(n3513), .ZN(n3793) );
  AND2_X1 U2871 ( .A1(n3586), .A2(DATAI_21_), .ZN(n2886) );
  INV_X1 U2872 ( .A(n3390), .ZN(n3372) );
  OR2_X1 U2873 ( .A1(n2879), .A2(n2986), .ZN(n3067) );
  NAND2_X1 U2874 ( .A1(n2397), .A2(REG3_REG_7__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U2875 ( .A1(n3215), .A2(n2459), .ZN(n3228) );
  AND2_X1 U2876 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2356) );
  AND2_X1 U2877 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2580), .ZN(n2581) );
  AND2_X1 U2878 ( .A1(n2774), .A2(n2745), .ZN(n3496) );
  OR2_X1 U2879 ( .A1(n2763), .A2(n3416), .ZN(n2710) );
  OR2_X1 U2880 ( .A1(n2763), .A2(n3509), .ZN(n2684) );
  AND4_X1 U2881 ( .A1(n2585), .A2(n2584), .A3(n2583), .A4(n2582), .ZN(n3959)
         );
  AND4_X1 U2882 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n4391)
         );
  NAND2_X1 U2883 ( .A1(n4314), .A2(REG1_REG_12__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U2884 ( .A1(n4381), .A2(n4382), .ZN(n4379) );
  INV_X1 U2885 ( .A(n4389), .ZN(n4422) );
  INV_X1 U2886 ( .A(n4426), .ZN(n4394) );
  INV_X1 U2887 ( .A(n4430), .ZN(n4445) );
  AND2_X1 U2888 ( .A1(n3954), .A2(n4537), .ZN(n4438) );
  INV_X1 U2889 ( .A(n4396), .ZN(n4444) );
  AOI21_X1 U2890 ( .B1(n2726), .B2(n3415), .A(n2725), .ZN(n2892) );
  INV_X1 U2891 ( .A(n4221), .ZN(n2896) );
  NAND2_X1 U2892 ( .A1(n3586), .A2(DATAI_20_), .ZN(n3907) );
  INV_X1 U2893 ( .A(n3198), .ZN(n3237) );
  AND2_X1 U2894 ( .A1(n4451), .A2(n2838), .ZN(n4538) );
  NAND2_X1 U2895 ( .A1(n2723), .A2(n2912), .ZN(n2910) );
  AND2_X1 U2896 ( .A1(n2474), .A2(n2491), .ZN(n3710) );
  INV_X1 U2897 ( .A(n4264), .ZN(n4486) );
  AND2_X1 U2898 ( .A1(n2935), .A2(n2934), .ZN(n4378) );
  NAND2_X1 U2899 ( .A1(n2756), .A2(STATE_REG_SCAN_IN), .ZN(n3503) );
  NAND4_X1 U2900 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n3884)
         );
  INV_X1 U2901 ( .A(n2813), .ZN(n3681) );
  OR2_X1 U2902 ( .A1(n2256), .A2(n4464), .ZN(n3689) );
  OR2_X1 U2903 ( .A1(n4245), .A2(n2963), .ZN(n4385) );
  OR2_X1 U2904 ( .A1(n4245), .A2(n4242), .ZN(n4354) );
  NAND2_X1 U2905 ( .A1(n4558), .A2(n4537), .ZN(n4168) );
  AND2_X2 U2906 ( .A1(n2893), .A2(n2892), .ZN(n4558) );
  NAND2_X1 U2907 ( .A1(n4544), .A2(n4537), .ZN(n4221) );
  INV_X1 U2908 ( .A(n4544), .ZN(n4542) );
  NAND2_X1 U2909 ( .A1(n2911), .A2(n2910), .ZN(n4460) );
  INV_X1 U2910 ( .A(n3736), .ZN(n4229) );
  INV_X1 U2911 ( .A(n3722), .ZN(n4478) );
  AND2_X1 U2912 ( .A1(n2405), .A2(n2423), .ZN(n4230) );
  INV_X1 U2913 ( .A(n3689), .ZN(U4043) );
  INV_X2 U2914 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND4_X1 U2915 ( .A1(n2503), .A2(n2504), .A3(n4107), .A4(n2544), .ZN(n2220)
         );
  INV_X1 U2916 ( .A(n2261), .ZN(n2222) );
  NAND2_X1 U2917 ( .A1(n2222), .A2(n4024), .ZN(n2225) );
  INV_X1 U2918 ( .A(IR_REG_18__SCAN_IN), .ZN(n2249) );
  NAND2_X1 U2919 ( .A1(n2223), .A2(n2249), .ZN(n2224) );
  INV_X1 U2920 ( .A(n2238), .ZN(n4225) );
  NAND2_X1 U2921 ( .A1(n2232), .A2(IR_REG_31__SCAN_IN), .ZN(n2234) );
  INV_X1 U2922 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2235) );
  INV_X1 U2923 ( .A(n2236), .ZN(n4226) );
  INV_X1 U2924 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2237) );
  NAND2_X1 U2925 ( .A1(n2322), .A2(REG0_REG_1__SCAN_IN), .ZN(n2239) );
  AND2_X1 U2926 ( .A1(n2240), .A2(n2241), .ZN(n2263) );
  NAND2_X1 U2927 ( .A1(n2244), .A2(IR_REG_31__SCAN_IN), .ZN(n2245) );
  XNOR2_X1 U2928 ( .A(n2245), .B(n2227), .ZN(n2913) );
  NOR2_X1 U2929 ( .A1(n2721), .A2(n2913), .ZN(n2248) );
  NAND2_X1 U2930 ( .A1(n2246), .A2(IR_REG_31__SCAN_IN), .ZN(n2247) );
  INV_X1 U2931 ( .A(n2240), .ZN(n2573) );
  NAND2_X1 U2932 ( .A1(n2586), .A2(n2249), .ZN(n2260) );
  NAND2_X1 U2933 ( .A1(n2260), .A2(IR_REG_31__SCAN_IN), .ZN(n2267) );
  NAND2_X1 U2934 ( .A1(n2267), .A2(n2266), .ZN(n2269) );
  INV_X1 U2935 ( .A(n2260), .ZN(n2253) );
  NAND2_X1 U2936 ( .A1(n2253), .A2(n2252), .ZN(n2254) );
  INV_X1 U2937 ( .A(n2938), .ZN(n2941) );
  NAND2_X1 U2938 ( .A1(n2760), .A2(IR_REG_27__SCAN_IN), .ZN(n2259) );
  OAI21_X1 U2939 ( .B1(n2261), .B2(n2260), .A(IR_REG_31__SCAN_IN), .ZN(n2262)
         );
  MUX2_X1 U2940 ( .A(IR_REG_31__SCAN_IN), .B(n2262), .S(IR_REG_22__SCAN_IN), 
        .Z(n2265) );
  INV_X1 U2941 ( .A(n2263), .ZN(n2264) );
  OR2_X1 U2942 ( .A1(n2267), .A2(n2266), .ZN(n2268) );
  NAND2_X1 U2943 ( .A1(n3670), .A2(n3736), .ZN(n2271) );
  NAND2_X1 U2944 ( .A1(n2014), .A2(n2790), .ZN(n2274) );
  NAND2_X1 U2945 ( .A1(n4421), .A2(n2611), .ZN(n2273) );
  NAND2_X1 U2946 ( .A1(n2274), .A2(n2273), .ZN(n2291) );
  INV_X1 U2947 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2283) );
  NAND2_X1 U2948 ( .A1(n2322), .A2(REG0_REG_0__SCAN_IN), .ZN(n2281) );
  INV_X1 U2949 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2276) );
  OR2_X1 U2950 ( .A1(n2275), .A2(n2276), .ZN(n2280) );
  INV_X1 U2951 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2277) );
  NAND2_X1 U2952 ( .A1(n2840), .A2(n2611), .ZN(n2282) );
  MUX2_X1 U2953 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2301), .Z(n2882) );
  NAND2_X1 U2954 ( .A1(n2882), .A2(n2318), .ZN(n2287) );
  OAI211_X1 U2955 ( .C1(n2256), .C2(n2283), .A(n2282), .B(n2287), .ZN(n2961)
         );
  NAND2_X1 U2956 ( .A1(n2840), .A2(n2014), .ZN(n2286) );
  NOR2_X1 U2957 ( .A1(n2256), .A2(n2015), .ZN(n2284) );
  AOI21_X1 U2958 ( .B1(n2882), .B2(n2611), .A(n2284), .ZN(n2285) );
  NAND2_X1 U2959 ( .A1(n2286), .A2(n2285), .ZN(n2962) );
  NAND2_X1 U2960 ( .A1(n2961), .A2(n2962), .ZN(n2289) );
  NAND2_X1 U2961 ( .A1(n2287), .A2(n2689), .ZN(n2288) );
  NAND2_X1 U2962 ( .A1(n2289), .A2(n2288), .ZN(n2985) );
  NAND2_X1 U2963 ( .A1(n2984), .A2(n2985), .ZN(n2294) );
  INV_X1 U2964 ( .A(n2290), .ZN(n2292) );
  NAND2_X1 U2965 ( .A1(n2292), .A2(n2291), .ZN(n2293) );
  NAND2_X1 U2966 ( .A1(n2294), .A2(n2293), .ZN(n3022) );
  INV_X1 U2967 ( .A(n3022), .ZN(n2313) );
  NAND2_X1 U2968 ( .A1(n2322), .A2(REG0_REG_2__SCAN_IN), .ZN(n2300) );
  INV_X1 U2969 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3103) );
  OR2_X1 U2970 ( .A1(n2275), .A2(n3103), .ZN(n2299) );
  INV_X1 U2971 ( .A(n2354), .ZN(n2295) );
  INV_X1 U2972 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2296) );
  OR2_X1 U2973 ( .A1(n2319), .A2(n2296), .ZN(n2297) );
  NAND2_X1 U2974 ( .A1(n2318), .A2(n3107), .ZN(n2305) );
  XNOR2_X1 U2975 ( .A(n2306), .B(n2689), .ZN(n2310) );
  NAND2_X1 U2976 ( .A1(n3107), .A2(n2611), .ZN(n2307) );
  AND2_X1 U2977 ( .A1(n2308), .A2(n2307), .ZN(n2309) );
  OR2_X1 U2978 ( .A1(n2310), .A2(n2309), .ZN(n2311) );
  NAND2_X1 U2979 ( .A1(n2310), .A2(n2309), .ZN(n2314) );
  NAND2_X1 U2980 ( .A1(n2311), .A2(n2314), .ZN(n3025) );
  NAND2_X1 U2981 ( .A1(n2313), .A2(n2312), .ZN(n3023) );
  NAND2_X1 U2982 ( .A1(n2315), .A2(IR_REG_31__SCAN_IN), .ZN(n2340) );
  XNOR2_X1 U2983 ( .A(n2340), .B(IR_REG_3__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U2984 ( .A1(n3544), .A2(n2318), .ZN(n2327) );
  INV_X1 U2985 ( .A(n2319), .ZN(n2916) );
  INV_X1 U2986 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3008) );
  OR2_X1 U2987 ( .A1(n2319), .A2(n3008), .ZN(n2325) );
  OR2_X1 U2988 ( .A1(n2354), .A2(n4550), .ZN(n2321) );
  OR2_X1 U2989 ( .A1(n2275), .A2(REG3_REG_3__SCAN_IN), .ZN(n2320) );
  AND2_X1 U2990 ( .A1(n3544), .A2(n2611), .ZN(n2329) );
  AOI21_X1 U2991 ( .B1(n3690), .B2(n2014), .A(n2329), .ZN(n2347) );
  XNOR2_X1 U2992 ( .A(n2346), .B(n2347), .ZN(n3044) );
  NAND2_X1 U2993 ( .A1(n3043), .A2(n3044), .ZN(n3042) );
  NAND2_X1 U2994 ( .A1(n2915), .A2(REG0_REG_4__SCAN_IN), .ZN(n2338) );
  INV_X1 U2995 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2330) );
  OR2_X1 U2996 ( .A1(n2354), .A2(n2330), .ZN(n2337) );
  INV_X1 U2997 ( .A(n2356), .ZN(n2334) );
  INV_X1 U2998 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2332) );
  INV_X1 U2999 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2331) );
  NAND2_X1 U3000 ( .A1(n2332), .A2(n2331), .ZN(n2333) );
  NAND2_X1 U3001 ( .A1(n2334), .A2(n2333), .ZN(n3084) );
  OR2_X1 U3002 ( .A1(n2763), .A2(n3084), .ZN(n2336) );
  INV_X1 U3003 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3012) );
  OR2_X1 U3004 ( .A1(n2319), .A2(n3012), .ZN(n2335) );
  INV_X1 U3005 ( .A(IR_REG_3__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3006 ( .A1(n2340), .A2(n2361), .ZN(n2341) );
  NAND2_X1 U3007 ( .A1(n2341), .A2(IR_REG_31__SCAN_IN), .ZN(n2342) );
  XNOR2_X1 U3008 ( .A(n2342), .B(IR_REG_4__SCAN_IN), .ZN(n4231) );
  MUX2_X1 U3009 ( .A(n4231), .B(DATAI_4_), .S(n3586), .Z(n2797) );
  OAI22_X1 U3010 ( .A1(n2796), .A2(n2339), .B1(n2713), .B2(n3083), .ZN(n2343)
         );
  XNOR2_X1 U3011 ( .A(n2343), .B(n2689), .ZN(n2350) );
  OR2_X1 U3012 ( .A1(n2796), .A2(n2703), .ZN(n2345) );
  NAND2_X1 U3013 ( .A1(n2797), .A2(n2611), .ZN(n2344) );
  NAND2_X1 U3014 ( .A1(n2345), .A2(n2344), .ZN(n2351) );
  XNOR2_X1 U3015 ( .A(n2350), .B(n2351), .ZN(n3052) );
  INV_X1 U3016 ( .A(n2346), .ZN(n2348) );
  NAND2_X1 U3017 ( .A1(n2348), .A2(n2347), .ZN(n3051) );
  AND2_X1 U3018 ( .A1(n3052), .A2(n3051), .ZN(n2349) );
  INV_X1 U3019 ( .A(n2350), .ZN(n2352) );
  NAND2_X1 U3020 ( .A1(n2352), .A2(n2351), .ZN(n2353) );
  NAND2_X1 U3021 ( .A1(n3053), .A2(n2353), .ZN(n3059) );
  NAND2_X1 U3022 ( .A1(n2915), .A2(REG0_REG_5__SCAN_IN), .ZN(n2360) );
  INV_X1 U3023 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2355) );
  OR2_X1 U3024 ( .A1(n2953), .A2(n2355), .ZN(n2359) );
  OAI21_X1 U3025 ( .B1(n2356), .B2(REG3_REG_5__SCAN_IN), .A(n2376), .ZN(n3128)
         );
  OR2_X1 U3026 ( .A1(n2763), .A2(n3128), .ZN(n2358) );
  INV_X1 U3027 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3129) );
  OR2_X1 U3028 ( .A1(n2319), .A2(n3129), .ZN(n2357) );
  NAND4_X1 U3029 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(n3688)
         );
  NAND2_X1 U3030 ( .A1(n3688), .A2(n2611), .ZN(n2366) );
  AND2_X1 U3031 ( .A1(n2362), .A2(n2361), .ZN(n2382) );
  NAND2_X1 U3032 ( .A1(n2363), .A2(IR_REG_31__SCAN_IN), .ZN(n2364) );
  XNOR2_X1 U3033 ( .A(n2364), .B(IR_REG_5__SCAN_IN), .ZN(n3007) );
  MUX2_X1 U3034 ( .A(n3007), .B(DATAI_5_), .S(n3586), .Z(n3127) );
  NAND2_X1 U3035 ( .A1(n3127), .A2(n2318), .ZN(n2365) );
  NAND2_X1 U3036 ( .A1(n2366), .A2(n2365), .ZN(n2367) );
  XNOR2_X1 U3037 ( .A(n2367), .B(n2716), .ZN(n2371) );
  AND2_X1 U3038 ( .A1(n3127), .A2(n2611), .ZN(n2368) );
  AOI21_X1 U3039 ( .B1(n3688), .B2(n2014), .A(n2368), .ZN(n2369) );
  XNOR2_X1 U3040 ( .A(n2371), .B(n2369), .ZN(n3060) );
  NAND2_X1 U3041 ( .A1(n3059), .A2(n3060), .ZN(n2373) );
  INV_X1 U3042 ( .A(n2369), .ZN(n2370) );
  NAND2_X1 U3043 ( .A1(n2371), .A2(n2370), .ZN(n2372) );
  NAND2_X1 U3044 ( .A1(n2915), .A2(REG0_REG_6__SCAN_IN), .ZN(n2381) );
  INV_X1 U3045 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2374) );
  OR2_X1 U3046 ( .A1(n2953), .A2(n2374), .ZN(n2380) );
  AND2_X1 U3047 ( .A1(n2376), .A2(n2375), .ZN(n2377) );
  OR2_X1 U3048 ( .A1(n2377), .A2(n2397), .ZN(n3158) );
  OR2_X1 U3049 ( .A1(n2763), .A2(n3158), .ZN(n2379) );
  INV_X1 U3050 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3159) );
  OR2_X1 U3051 ( .A1(n2319), .A2(n3159), .ZN(n2378) );
  NAND4_X1 U3052 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3687)
         );
  NAND2_X1 U3053 ( .A1(n3687), .A2(n2611), .ZN(n2389) );
  AND2_X1 U3054 ( .A1(n2383), .A2(n2382), .ZN(n2384) );
  NOR2_X1 U3055 ( .A1(n2384), .A2(n2759), .ZN(n2385) );
  MUX2_X1 U3056 ( .A(n2759), .B(n2385), .S(IR_REG_6__SCAN_IN), .Z(n2387) );
  OR2_X1 U3057 ( .A1(n2387), .A2(n2386), .ZN(n4264) );
  MUX2_X1 U3058 ( .A(n4486), .B(DATAI_6_), .S(n3586), .Z(n2883) );
  NAND2_X1 U3059 ( .A1(n2883), .A2(n2318), .ZN(n2388) );
  NAND2_X1 U3060 ( .A1(n2389), .A2(n2388), .ZN(n2390) );
  XNOR2_X1 U3061 ( .A(n2390), .B(n2716), .ZN(n2393) );
  NAND2_X1 U3062 ( .A1(n3687), .A2(n2014), .ZN(n2392) );
  NAND2_X1 U3063 ( .A1(n2883), .A2(n2611), .ZN(n2391) );
  NAND2_X1 U3064 ( .A1(n2392), .A2(n2391), .ZN(n2394) );
  AND2_X1 U3065 ( .A1(n2393), .A2(n2394), .ZN(n3090) );
  INV_X1 U3066 ( .A(n2393), .ZN(n2396) );
  INV_X1 U3067 ( .A(n2394), .ZN(n2395) );
  NAND2_X1 U3068 ( .A1(n2396), .A2(n2395), .ZN(n3091) );
  NAND2_X1 U3069 ( .A1(n2915), .A2(REG0_REG_7__SCAN_IN), .ZN(n2402) );
  INV_X1 U3070 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3004) );
  OR2_X1 U3071 ( .A1(n2953), .A2(n3004), .ZN(n2401) );
  OR2_X1 U3072 ( .A1(n2397), .A2(REG3_REG_7__SCAN_IN), .ZN(n2398) );
  NAND2_X1 U3073 ( .A1(n2415), .A2(n2398), .ZN(n3181) );
  OR2_X1 U3074 ( .A1(n2763), .A2(n3181), .ZN(n2400) );
  INV_X1 U3075 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3015) );
  OR2_X1 U3076 ( .A1(n2319), .A2(n3015), .ZN(n2399) );
  OR2_X1 U3077 ( .A1(n2386), .A2(n2759), .ZN(n2404) );
  INV_X1 U3078 ( .A(n2404), .ZN(n2403) );
  NAND2_X1 U3079 ( .A1(n2403), .A2(IR_REG_7__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3080 ( .A1(n2404), .A2(n2087), .ZN(n2423) );
  MUX2_X1 U3081 ( .A(n4230), .B(DATAI_7_), .S(n3586), .Z(n3180) );
  OAI22_X1 U3082 ( .A1(n3151), .A2(n2339), .B1(n2713), .B2(n3174), .ZN(n2406)
         );
  XNOR2_X1 U3083 ( .A(n2406), .B(n2716), .ZN(n2411) );
  OR2_X1 U3084 ( .A1(n3151), .A2(n2703), .ZN(n2408) );
  NAND2_X1 U3085 ( .A1(n3180), .A2(n2611), .ZN(n2407) );
  NAND2_X1 U3086 ( .A1(n2408), .A2(n2407), .ZN(n2410) );
  XNOR2_X1 U3087 ( .A(n2411), .B(n2410), .ZN(n3165) );
  NAND2_X1 U3088 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  NAND2_X1 U3089 ( .A1(n3166), .A2(n2412), .ZN(n3197) );
  NAND2_X1 U3090 ( .A1(n2915), .A2(REG0_REG_8__SCAN_IN), .ZN(n2422) );
  INV_X1 U3091 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2413) );
  OR2_X1 U3092 ( .A1(n2953), .A2(n2413), .ZN(n2421) );
  NAND2_X1 U3093 ( .A1(n2415), .A2(n2414), .ZN(n2416) );
  AND2_X1 U3094 ( .A1(n2431), .A2(n2416), .ZN(n4413) );
  INV_X1 U3095 ( .A(n4413), .ZN(n2417) );
  OR2_X1 U3096 ( .A1(n2763), .A2(n2417), .ZN(n2420) );
  INV_X1 U3097 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2418) );
  OR2_X1 U3098 ( .A1(n2319), .A2(n2418), .ZN(n2419) );
  NAND4_X1 U3099 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), .ZN(n3686)
         );
  NAND2_X1 U3100 ( .A1(n3686), .A2(n2014), .ZN(n2426) );
  NAND2_X1 U3101 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  XNOR2_X1 U3102 ( .A(n2424), .B(IR_REG_8__SCAN_IN), .ZN(n4265) );
  MUX2_X1 U3103 ( .A(n4265), .B(DATAI_8_), .S(n3586), .Z(n3198) );
  NAND2_X1 U3104 ( .A1(n3198), .A2(n2611), .ZN(n2425) );
  NAND2_X1 U3105 ( .A1(n2426), .A2(n2425), .ZN(n3195) );
  NAND2_X1 U3106 ( .A1(n3686), .A2(n2611), .ZN(n2428) );
  NAND2_X1 U3107 ( .A1(n3198), .A2(n2318), .ZN(n2427) );
  NAND2_X1 U3108 ( .A1(n2428), .A2(n2427), .ZN(n2429) );
  XNOR2_X1 U3109 ( .A(n2429), .B(n2716), .ZN(n3194) );
  NAND2_X1 U3110 ( .A1(n2915), .A2(REG0_REG_9__SCAN_IN), .ZN(n2437) );
  INV_X1 U3111 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2430) );
  OR2_X1 U3112 ( .A1(n2953), .A2(n2430), .ZN(n2436) );
  AND2_X1 U3113 ( .A1(n2431), .A2(n3219), .ZN(n2432) );
  OR2_X1 U3114 ( .A1(n2432), .A2(n2444), .ZN(n3211) );
  OR2_X1 U3115 ( .A1(n2763), .A2(n3211), .ZN(n2435) );
  INV_X1 U3116 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2433) );
  OR2_X1 U3117 ( .A1(n2319), .A2(n2433), .ZN(n2434) );
  NAND4_X1 U3118 ( .A1(n2437), .A2(n2436), .A3(n2435), .A4(n2434), .ZN(n3685)
         );
  NAND2_X1 U3119 ( .A1(n3685), .A2(n2611), .ZN(n2441) );
  NAND2_X1 U3120 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2439) );
  XNOR2_X1 U3121 ( .A(n2439), .B(IR_REG_9__SCAN_IN), .ZN(n4482) );
  MUX2_X1 U3122 ( .A(n4482), .B(DATAI_9_), .S(n3586), .Z(n3209) );
  NAND2_X1 U3123 ( .A1(n3209), .A2(n2318), .ZN(n2440) );
  NAND2_X1 U3124 ( .A1(n2441), .A2(n2440), .ZN(n2442) );
  XNOR2_X1 U3125 ( .A(n2442), .B(n2689), .ZN(n2458) );
  AND2_X1 U3126 ( .A1(n3209), .A2(n2611), .ZN(n2443) );
  AOI21_X1 U3127 ( .B1(n3685), .B2(n2014), .A(n2443), .ZN(n2457) );
  XNOR2_X1 U3128 ( .A(n2458), .B(n2457), .ZN(n3218) );
  NAND2_X1 U3129 ( .A1(n2915), .A2(REG0_REG_10__SCAN_IN), .ZN(n2451) );
  NOR2_X1 U3130 ( .A1(n2444), .A2(REG3_REG_10__SCAN_IN), .ZN(n2445) );
  OR2_X1 U3131 ( .A1(n2464), .A2(n2445), .ZN(n4405) );
  OR2_X1 U3132 ( .A1(n2763), .A2(n4405), .ZN(n2450) );
  INV_X1 U3133 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2446) );
  OR2_X1 U3134 ( .A1(n2953), .A2(n2446), .ZN(n2449) );
  INV_X1 U3135 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2447) );
  OR2_X1 U3136 ( .A1(n2319), .A2(n2447), .ZN(n2448) );
  NAND4_X1 U3137 ( .A1(n2451), .A2(n2450), .A3(n2449), .A4(n2448), .ZN(n4393)
         );
  NAND2_X1 U3138 ( .A1(n4393), .A2(n2611), .ZN(n2454) );
  NAND2_X1 U3139 ( .A1(n2506), .A2(IR_REG_31__SCAN_IN), .ZN(n2452) );
  XNOR2_X1 U3140 ( .A(n2452), .B(IR_REG_10__SCAN_IN), .ZN(n4287) );
  MUX2_X1 U3141 ( .A(n4287), .B(DATAI_10_), .S(n3586), .Z(n2884) );
  NAND2_X1 U3142 ( .A1(n2884), .A2(n2318), .ZN(n2453) );
  NAND2_X1 U3143 ( .A1(n2454), .A2(n2453), .ZN(n2455) );
  XNOR2_X1 U3144 ( .A(n2455), .B(n2716), .ZN(n2462) );
  AND2_X1 U3145 ( .A1(n2884), .A2(n2611), .ZN(n2456) );
  AOI21_X1 U3146 ( .B1(n4393), .B2(n2014), .A(n2456), .ZN(n2460) );
  XNOR2_X1 U3147 ( .A(n2462), .B(n2460), .ZN(n3229) );
  NAND2_X1 U31480 ( .A1(n2458), .A2(n2457), .ZN(n3227) );
  AND2_X1 U31490 ( .A1(n3229), .A2(n3227), .ZN(n2459) );
  INV_X1 U3150 ( .A(n2460), .ZN(n2461) );
  NAND2_X1 U3151 ( .A1(n2462), .A2(n2461), .ZN(n2463) );
  NAND2_X1 U3152 ( .A1(n3228), .A2(n2463), .ZN(n3252) );
  NAND2_X1 U3153 ( .A1(n2915), .A2(REG0_REG_11__SCAN_IN), .ZN(n2470) );
  OR2_X1 U3154 ( .A1(n2464), .A2(REG3_REG_11__SCAN_IN), .ZN(n2465) );
  AND2_X1 U3155 ( .A1(n2484), .A2(n2465), .ZN(n4399) );
  INV_X1 U3156 ( .A(n4399), .ZN(n3259) );
  OR2_X1 U3157 ( .A1(n2763), .A2(n3259), .ZN(n2469) );
  INV_X1 U3158 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2466) );
  OR2_X1 U3159 ( .A1(n2953), .A2(n2466), .ZN(n2468) );
  OR2_X1 U3160 ( .A1(n2319), .A2(n3719), .ZN(n2467) );
  NAND2_X1 U3161 ( .A1(n2471), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  INV_X1 U3162 ( .A(n2473), .ZN(n2472) );
  NAND2_X1 U3163 ( .A1(n2472), .A2(IR_REG_11__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3164 ( .A1(n2473), .A2(n2503), .ZN(n2491) );
  MUX2_X1 U3165 ( .A(n3710), .B(DATAI_11_), .S(n3586), .Z(n4402) );
  OAI22_X1 U3166 ( .A1(n3301), .A2(n2339), .B1(n2713), .B2(n4390), .ZN(n2475)
         );
  XNOR2_X1 U3167 ( .A(n2475), .B(n2689), .ZN(n2478) );
  OR2_X1 U3168 ( .A1(n3301), .A2(n2703), .ZN(n2477) );
  NAND2_X1 U3169 ( .A1(n4402), .A2(n2611), .ZN(n2476) );
  AND2_X1 U3170 ( .A1(n2477), .A2(n2476), .ZN(n2479) );
  NAND2_X1 U3171 ( .A1(n2478), .A2(n2479), .ZN(n3249) );
  INV_X1 U3172 ( .A(n2478), .ZN(n2481) );
  INV_X1 U3173 ( .A(n2479), .ZN(n2480) );
  NAND2_X1 U3174 ( .A1(n2481), .A2(n2480), .ZN(n3250) );
  NAND2_X1 U3175 ( .A1(n2915), .A2(REG0_REG_12__SCAN_IN), .ZN(n2490) );
  INV_X1 U3176 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2482) );
  OR2_X1 U3177 ( .A1(n2953), .A2(n2482), .ZN(n2489) );
  NAND2_X1 U3178 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  NAND2_X1 U3179 ( .A1(n2497), .A2(n2485), .ZN(n3262) );
  OR2_X1 U3180 ( .A1(n2763), .A2(n3262), .ZN(n2488) );
  INV_X1 U3181 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2486) );
  OR2_X1 U3182 ( .A1(n2955), .A2(n2486), .ZN(n2487) );
  NAND2_X1 U3183 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  XNOR2_X1 U3184 ( .A(n2492), .B(IR_REG_12__SCAN_IN), .ZN(n3722) );
  INV_X1 U3185 ( .A(DATAI_12_), .ZN(n2493) );
  MUX2_X1 U3186 ( .A(n4478), .B(n2493), .S(n3586), .Z(n3273) );
  OAI22_X1 U3187 ( .A1(n4391), .A2(n2339), .B1(n2713), .B2(n3273), .ZN(n2494)
         );
  XNOR2_X1 U3188 ( .A(n2494), .B(n2689), .ZN(n3327) );
  OR2_X1 U3189 ( .A1(n4391), .A2(n2703), .ZN(n2496) );
  INV_X1 U3190 ( .A(n3273), .ZN(n3267) );
  NAND2_X1 U3191 ( .A1(n3267), .A2(n2611), .ZN(n2495) );
  NAND2_X1 U3192 ( .A1(n2915), .A2(REG0_REG_13__SCAN_IN), .ZN(n2502) );
  INV_X1 U3193 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3700) );
  OR2_X1 U3194 ( .A1(n2953), .A2(n3700), .ZN(n2501) );
  NAND2_X1 U3195 ( .A1(n2497), .A2(n3336), .ZN(n2498) );
  NAND2_X1 U3196 ( .A1(n2522), .A2(n2498), .ZN(n3340) );
  OR2_X1 U3197 ( .A1(n2763), .A2(n3340), .ZN(n2500) );
  INV_X1 U3198 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3291) );
  OR2_X1 U3199 ( .A1(n2319), .A2(n3291), .ZN(n2499) );
  NAND4_X1 U3200 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(n3682)
         );
  NAND2_X1 U3201 ( .A1(n3682), .A2(n2611), .ZN(n2509) );
  NAND3_X1 U3202 ( .A1(n2504), .A2(n2503), .A3(n4107), .ZN(n2505) );
  NAND2_X1 U3203 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2507) );
  XNOR2_X1 U3204 ( .A(n2507), .B(IR_REG_13__SCAN_IN), .ZN(n3724) );
  MUX2_X1 U3205 ( .A(n3724), .B(DATAI_13_), .S(n3586), .Z(n3288) );
  NAND2_X1 U3206 ( .A1(n3288), .A2(n2318), .ZN(n2508) );
  NAND2_X1 U3207 ( .A1(n2509), .A2(n2508), .ZN(n2510) );
  XNOR2_X1 U3208 ( .A(n2510), .B(n2716), .ZN(n2513) );
  NAND2_X1 U3209 ( .A1(n3682), .A2(n2014), .ZN(n2512) );
  NAND2_X1 U32100 ( .A1(n3288), .A2(n2611), .ZN(n2511) );
  NAND2_X1 U32110 ( .A1(n2512), .A2(n2511), .ZN(n2514) );
  NAND2_X1 U32120 ( .A1(n2513), .A2(n2514), .ZN(n3332) );
  OAI21_X1 U32130 ( .B1(n3327), .B2(n3329), .A(n3332), .ZN(n2519) );
  NAND3_X1 U32140 ( .A1(n3327), .A2(n3329), .A3(n3332), .ZN(n2517) );
  INV_X1 U32150 ( .A(n2513), .ZN(n2516) );
  INV_X1 U32160 ( .A(n2514), .ZN(n2515) );
  NAND2_X1 U32170 ( .A1(n2516), .A2(n2515), .ZN(n3331) );
  AND2_X1 U32180 ( .A1(n2517), .A2(n3331), .ZN(n2518) );
  NAND2_X1 U32190 ( .A1(n2915), .A2(REG0_REG_14__SCAN_IN), .ZN(n2527) );
  INV_X1 U32200 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2520) );
  OR2_X1 U32210 ( .A1(n2953), .A2(n2520), .ZN(n2526) );
  AND2_X1 U32220 ( .A1(n2522), .A2(n2521), .ZN(n2523) );
  OR2_X1 U32230 ( .A1(n2523), .A2(n2537), .ZN(n3349) );
  OR2_X1 U32240 ( .A1(n2763), .A2(n3349), .ZN(n2525) );
  OR2_X1 U32250 ( .A1(n2319), .A2(n4331), .ZN(n2524) );
  OR2_X1 U32260 ( .A1(n2545), .A2(n2759), .ZN(n2529) );
  XNOR2_X1 U32270 ( .A(n2529), .B(IR_REG_14__SCAN_IN), .ZN(n3701) );
  MUX2_X1 U32280 ( .A(n3701), .B(DATAI_14_), .S(n3586), .Z(n3347) );
  INV_X1 U32290 ( .A(n3347), .ZN(n2814) );
  OAI22_X1 U32300 ( .A1(n2813), .A2(n2339), .B1(n2713), .B2(n2814), .ZN(n2530)
         );
  XNOR2_X1 U32310 ( .A(n2530), .B(n2689), .ZN(n3310) );
  OR2_X1 U32320 ( .A1(n2813), .A2(n2703), .ZN(n2532) );
  NAND2_X1 U32330 ( .A1(n3347), .A2(n2611), .ZN(n2531) );
  NAND2_X1 U32340 ( .A1(n2532), .A2(n2531), .ZN(n3311) );
  NAND2_X1 U32350 ( .A1(n2533), .A2(n3311), .ZN(n2536) );
  INV_X1 U32360 ( .A(n3313), .ZN(n2534) );
  NAND2_X1 U32370 ( .A1(n2534), .A2(n2179), .ZN(n2535) );
  NAND2_X1 U32380 ( .A1(n2915), .A2(REG0_REG_15__SCAN_IN), .ZN(n2543) );
  INV_X1 U32390 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3704) );
  OR2_X1 U32400 ( .A1(n2953), .A2(n3704), .ZN(n2542) );
  NOR2_X1 U32410 ( .A1(n2537), .A2(REG3_REG_15__SCAN_IN), .ZN(n2538) );
  OR2_X1 U32420 ( .A1(n2551), .A2(n2538), .ZN(n3361) );
  OR2_X1 U32430 ( .A1(n2763), .A2(n3361), .ZN(n2541) );
  INV_X1 U32440 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2539) );
  OR2_X1 U32450 ( .A1(n2955), .A2(n2539), .ZN(n2540) );
  NAND4_X1 U32460 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n3680)
         );
  NAND2_X1 U32470 ( .A1(n3680), .A2(n2611), .ZN(n2548) );
  NAND2_X1 U32480 ( .A1(n2545), .A2(n2544), .ZN(n2546) );
  NAND2_X1 U32490 ( .A1(n2546), .A2(IR_REG_31__SCAN_IN), .ZN(n2559) );
  XNOR2_X1 U32500 ( .A(n2559), .B(IR_REG_15__SCAN_IN), .ZN(n4472) );
  MUX2_X1 U32510 ( .A(n4472), .B(DATAI_15_), .S(n3586), .Z(n3400) );
  NAND2_X1 U32520 ( .A1(n3400), .A2(n2318), .ZN(n2547) );
  NAND2_X1 U32530 ( .A1(n2548), .A2(n2547), .ZN(n2549) );
  XNOR2_X1 U32540 ( .A(n2549), .B(n2716), .ZN(n2563) );
  AND2_X1 U32550 ( .A1(n3400), .A2(n2611), .ZN(n2550) );
  AOI21_X1 U32560 ( .B1(n3680), .B2(n2014), .A(n2550), .ZN(n3398) );
  NAND2_X1 U32570 ( .A1(n2915), .A2(REG0_REG_16__SCAN_IN), .ZN(n2557) );
  OR2_X1 U32580 ( .A1(n2551), .A2(REG3_REG_16__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32590 ( .A1(n2552), .A2(n2568), .ZN(n3375) );
  OR2_X1 U32600 ( .A1(n2763), .A2(n3375), .ZN(n2556) );
  INV_X1 U32610 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4166) );
  OR2_X1 U32620 ( .A1(n2953), .A2(n4166), .ZN(n2555) );
  INV_X1 U32630 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2553) );
  OR2_X1 U32640 ( .A1(n2955), .A2(n2553), .ZN(n2554) );
  NAND2_X1 U32650 ( .A1(n2559), .A2(n2558), .ZN(n2560) );
  NAND2_X1 U32660 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2561) );
  XNOR2_X1 U32670 ( .A(n2561), .B(IR_REG_16__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U32680 ( .A(n4470), .B(DATAI_16_), .S(n3586), .Z(n3390) );
  OAI22_X1 U32690 ( .A1(n3467), .A2(n2703), .B1(n2339), .B2(n3372), .ZN(n2565)
         );
  OAI22_X1 U32700 ( .A1(n3467), .A2(n2339), .B1(n2713), .B2(n3372), .ZN(n2562)
         );
  XNOR2_X1 U32710 ( .A(n2562), .B(n2716), .ZN(n2564) );
  XOR2_X1 U32720 ( .A(n2565), .B(n2564), .Z(n3388) );
  INV_X1 U32730 ( .A(n2564), .ZN(n2567) );
  INV_X1 U32740 ( .A(n3463), .ZN(n2579) );
  NAND2_X1 U32750 ( .A1(n2915), .A2(REG0_REG_17__SCAN_IN), .ZN(n2572) );
  INV_X1 U32760 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4162) );
  OR2_X1 U32770 ( .A1(n2953), .A2(n4162), .ZN(n2571) );
  XNOR2_X1 U32780 ( .A(REG3_REG_17__SCAN_IN), .B(n2580), .ZN(n3969) );
  OR2_X1 U32790 ( .A1(n2763), .A2(n3969), .ZN(n2570) );
  INV_X1 U32800 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3970) );
  OR2_X1 U32810 ( .A1(n2955), .A2(n3970), .ZN(n2569) );
  NAND2_X1 U32820 ( .A1(n2573), .A2(IR_REG_31__SCAN_IN), .ZN(n2574) );
  XNOR2_X1 U32830 ( .A(n2574), .B(IR_REG_17__SCAN_IN), .ZN(n3730) );
  MUX2_X1 U32840 ( .A(n3730), .B(DATAI_17_), .S(n3586), .Z(n2885) );
  INV_X1 U32850 ( .A(n2885), .ZN(n3966) );
  OAI22_X1 U32860 ( .A1(n3949), .A2(n2339), .B1(n2713), .B2(n3966), .ZN(n2575)
         );
  XOR2_X1 U32870 ( .A(n2716), .B(n2575), .Z(n3464) );
  OR2_X1 U32880 ( .A1(n3949), .A2(n2703), .ZN(n2577) );
  NAND2_X1 U32890 ( .A1(n2885), .A2(n2611), .ZN(n2576) );
  NAND2_X1 U32900 ( .A1(n2915), .A2(REG0_REG_18__SCAN_IN), .ZN(n2585) );
  INV_X1 U32910 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3707) );
  OR2_X1 U32920 ( .A1(n2953), .A2(n3707), .ZN(n2584) );
  OAI21_X1 U32930 ( .B1(n2581), .B2(REG3_REG_18__SCAN_IN), .A(n2593), .ZN(
        n3942) );
  OR2_X1 U32940 ( .A1(n2763), .A2(n3942), .ZN(n2583) );
  INV_X1 U32950 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3943) );
  OR2_X1 U32960 ( .A1(n2955), .A2(n3943), .ZN(n2582) );
  OR2_X1 U32970 ( .A1(n2586), .A2(n2759), .ZN(n2587) );
  XNOR2_X1 U32980 ( .A(n2587), .B(IR_REG_18__SCAN_IN), .ZN(n3731) );
  MUX2_X1 U32990 ( .A(n3731), .B(DATAI_18_), .S(n3586), .Z(n3946) );
  INV_X1 U33000 ( .A(n3946), .ZN(n3498) );
  OAI22_X1 U33010 ( .A1(n3959), .A2(n2339), .B1(n2713), .B2(n3498), .ZN(n2588)
         );
  XNOR2_X1 U33020 ( .A(n2588), .B(n2716), .ZN(n2592) );
  OR2_X1 U33030 ( .A1(n3959), .A2(n2703), .ZN(n2590) );
  NAND2_X1 U33040 ( .A1(n3946), .A2(n2611), .ZN(n2589) );
  NAND2_X1 U33050 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  NOR2_X1 U33060 ( .A1(n2592), .A2(n2591), .ZN(n3494) );
  NAND2_X1 U33070 ( .A1(n2915), .A2(REG0_REG_19__SCAN_IN), .ZN(n2598) );
  INV_X1 U33080 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4155) );
  OR2_X1 U33090 ( .A1(n2953), .A2(n4155), .ZN(n2597) );
  AND2_X1 U33100 ( .A1(n2593), .A2(n4083), .ZN(n2594) );
  OR2_X1 U33110 ( .A1(n2594), .A2(n2605), .ZN(n3932) );
  OR2_X1 U33120 ( .A1(n2763), .A2(n3932), .ZN(n2596) );
  INV_X1 U33130 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3933) );
  OR2_X1 U33140 ( .A1(n2955), .A2(n3933), .ZN(n2595) );
  NAND2_X1 U33150 ( .A1(n3947), .A2(n2611), .ZN(n2601) );
  INV_X1 U33160 ( .A(DATAI_19_), .ZN(n2599) );
  MUX2_X1 U33170 ( .A(n3736), .B(n2599), .S(n3586), .Z(n3929) );
  INV_X1 U33180 ( .A(n3929), .ZN(n2821) );
  NAND2_X1 U33190 ( .A1(n2821), .A2(n2318), .ZN(n2600) );
  NAND2_X1 U33200 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  XNOR2_X1 U33210 ( .A(n2602), .B(n2716), .ZN(n2604) );
  INV_X1 U33220 ( .A(n3947), .ZN(n2820) );
  OAI22_X1 U33230 ( .A1(n2820), .A2(n2703), .B1(n2339), .B2(n3929), .ZN(n2603)
         );
  XNOR2_X1 U33240 ( .A(n2604), .B(n2603), .ZN(n3435) );
  NAND2_X1 U33250 ( .A1(n2915), .A2(REG0_REG_20__SCAN_IN), .ZN(n2610) );
  INV_X1 U33260 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4151) );
  OR2_X1 U33270 ( .A1(n2953), .A2(n4151), .ZN(n2609) );
  OR2_X1 U33280 ( .A1(n2605), .A2(REG3_REG_20__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U33290 ( .A1(n2618), .A2(n2606), .ZN(n3908) );
  OR2_X1 U33300 ( .A1(n2763), .A2(n3908), .ZN(n2608) );
  INV_X1 U33310 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3909) );
  OR2_X1 U33320 ( .A1(n2955), .A2(n3909), .ZN(n2607) );
  NAND2_X1 U33330 ( .A1(n3884), .A2(n2611), .ZN(n2613) );
  OR2_X1 U33340 ( .A1(n3907), .A2(n2713), .ZN(n2612) );
  NAND2_X1 U33350 ( .A1(n2613), .A2(n2612), .ZN(n2614) );
  XNOR2_X1 U33360 ( .A(n2614), .B(n2689), .ZN(n2617) );
  NOR2_X1 U33370 ( .A1(n3907), .A2(n2339), .ZN(n2615) );
  AOI21_X1 U33380 ( .B1(n3884), .B2(n2014), .A(n2615), .ZN(n2616) );
  OR2_X1 U33390 ( .A1(n2617), .A2(n2616), .ZN(n3482) );
  NAND2_X1 U33400 ( .A1(n2617), .A2(n2616), .ZN(n3484) );
  NAND2_X1 U33410 ( .A1(n2915), .A2(REG0_REG_21__SCAN_IN), .ZN(n2623) );
  INV_X1 U33420 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4146) );
  OR2_X1 U33430 ( .A1(n2953), .A2(n4146), .ZN(n2622) );
  INV_X1 U33440 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3445) );
  NAND2_X1 U33450 ( .A1(n2618), .A2(n3445), .ZN(n2619) );
  NAND2_X1 U33460 ( .A1(n2632), .A2(n2619), .ZN(n3890) );
  OR2_X1 U33470 ( .A1(n2763), .A2(n3890), .ZN(n2621) );
  INV_X1 U33480 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3891) );
  OR2_X1 U33490 ( .A1(n2955), .A2(n3891), .ZN(n2620) );
  OAI22_X1 U33500 ( .A1(n3896), .A2(n2339), .B1(n2713), .B2(n3888), .ZN(n2624)
         );
  XNOR2_X1 U33510 ( .A(n2624), .B(n2716), .ZN(n3442) );
  OR2_X1 U33520 ( .A1(n3896), .A2(n2703), .ZN(n2626) );
  NAND2_X1 U3353 ( .A1(n2886), .A2(n2611), .ZN(n2625) );
  NAND2_X1 U33540 ( .A1(n2626), .A2(n2625), .ZN(n3441) );
  NOR2_X1 U3355 ( .A1(n3442), .A2(n3441), .ZN(n2629) );
  INV_X1 U3356 ( .A(n3442), .ZN(n2628) );
  INV_X1 U3357 ( .A(n3441), .ZN(n2627) );
  NAND2_X1 U3358 ( .A1(n2915), .A2(REG0_REG_22__SCAN_IN), .ZN(n2637) );
  INV_X1 U3359 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2630) );
  OR2_X1 U3360 ( .A1(n2953), .A2(n2630), .ZN(n2636) );
  INV_X1 U3361 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2631) );
  AND2_X1 U3362 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  OR2_X1 U3363 ( .A1(n2633), .A2(n2639), .ZN(n3864) );
  OR2_X1 U3364 ( .A1(n2763), .A2(n3864), .ZN(n2635) );
  INV_X1 U3365 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3865) );
  OR2_X1 U3366 ( .A1(n2955), .A2(n3865), .ZN(n2634) );
  INV_X1 U3367 ( .A(n3873), .ZN(n2825) );
  OAI22_X1 U3368 ( .A1(n3880), .A2(n2339), .B1(n2713), .B2(n2825), .ZN(n2638)
         );
  XNOR2_X1 U3369 ( .A(n2638), .B(n2716), .ZN(n2649) );
  OAI22_X1 U3370 ( .A1(n3880), .A2(n2703), .B1(n2339), .B2(n2825), .ZN(n2648)
         );
  XNOR2_X1 U3371 ( .A(n2649), .B(n2648), .ZN(n3408) );
  NAND2_X1 U3372 ( .A1(n2915), .A2(REG0_REG_23__SCAN_IN), .ZN(n2644) );
  INV_X1 U3373 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4137) );
  OR2_X1 U3374 ( .A1(n2953), .A2(n4137), .ZN(n2643) );
  NOR2_X1 U3375 ( .A1(n2639), .A2(REG3_REG_23__SCAN_IN), .ZN(n2640) );
  OR2_X1 U3376 ( .A1(n2654), .A2(n2640), .ZN(n3854) );
  OR2_X1 U3377 ( .A1(n2763), .A2(n3854), .ZN(n2642) );
  INV_X1 U3378 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3855) );
  OR2_X1 U3379 ( .A1(n2955), .A2(n3855), .ZN(n2641) );
  OAI22_X1 U3380 ( .A1(n3872), .A2(n2339), .B1(n2713), .B2(n3853), .ZN(n2645)
         );
  XNOR2_X1 U3381 ( .A(n2645), .B(n2716), .ZN(n2650) );
  OR2_X1 U3382 ( .A1(n3872), .A2(n2703), .ZN(n2647) );
  NAND2_X1 U3383 ( .A1(n3847), .A2(n2611), .ZN(n2646) );
  NAND2_X1 U3384 ( .A1(n2647), .A2(n2646), .ZN(n2651) );
  XNOR2_X1 U3385 ( .A(n2650), .B(n2651), .ZN(n3427) );
  NOR2_X1 U3386 ( .A1(n2649), .A2(n2648), .ZN(n3428) );
  INV_X1 U3387 ( .A(n2650), .ZN(n2653) );
  INV_X1 U3388 ( .A(n2651), .ZN(n2652) );
  NOR2_X1 U3389 ( .A1(n2653), .A2(n2652), .ZN(n2667) );
  INV_X1 U3390 ( .A(n2667), .ZN(n2663) );
  NAND2_X1 U3391 ( .A1(n2915), .A2(REG0_REG_24__SCAN_IN), .ZN(n2659) );
  INV_X1 U3392 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4133) );
  OR2_X1 U3393 ( .A1(n2953), .A2(n4133), .ZN(n2658) );
  OR2_X1 U3394 ( .A1(n2654), .A2(REG3_REG_24__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3395 ( .A1(n2669), .A2(n2655), .ZN(n3833) );
  INV_X1 U3396 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3834) );
  OR2_X1 U3397 ( .A1(n2955), .A2(n3834), .ZN(n2656) );
  NAND2_X1 U3398 ( .A1(n3848), .A2(n2014), .ZN(n2661) );
  NAND2_X1 U3399 ( .A1(n3586), .A2(DATAI_24_), .ZN(n3832) );
  OR2_X1 U3400 ( .A1(n3832), .A2(n2339), .ZN(n2660) );
  NAND2_X1 U3401 ( .A1(n2661), .A2(n2660), .ZN(n2666) );
  INV_X1 U3402 ( .A(n2666), .ZN(n2662) );
  OAI22_X1 U3403 ( .A1(n3807), .A2(n2339), .B1(n2713), .B2(n3832), .ZN(n2665)
         );
  XOR2_X1 U3404 ( .A(n2716), .B(n2665), .Z(n3473) );
  NAND2_X1 U3405 ( .A1(n2915), .A2(REG0_REG_25__SCAN_IN), .ZN(n2674) );
  INV_X1 U3406 ( .A(REG1_REG_25__SCAN_IN), .ZN(n2668) );
  OR2_X1 U3407 ( .A1(n2953), .A2(n2668), .ZN(n2673) );
  INV_X1 U3408 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U3409 ( .A1(n2669), .A2(n3456), .ZN(n2670) );
  NAND2_X1 U3410 ( .A1(n2680), .A2(n2670), .ZN(n3815) );
  INV_X1 U3411 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3816) );
  OR2_X1 U3412 ( .A1(n2319), .A2(n3816), .ZN(n2671) );
  INV_X1 U3413 ( .A(n3812), .ZN(n3457) );
  OAI22_X1 U3414 ( .A1(n3824), .A2(n2339), .B1(n2713), .B2(n3457), .ZN(n2675)
         );
  XNOR2_X1 U3415 ( .A(n2675), .B(n2689), .ZN(n2679) );
  OR2_X1 U3416 ( .A1(n3824), .A2(n2703), .ZN(n2677) );
  NAND2_X1 U3417 ( .A1(n3812), .A2(n2611), .ZN(n2676) );
  AND2_X1 U3418 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  NAND2_X1 U3419 ( .A1(n2679), .A2(n2678), .ZN(n3452) );
  NOR2_X1 U3420 ( .A1(n2679), .A2(n2678), .ZN(n3454) );
  NAND2_X1 U3421 ( .A1(n2915), .A2(REG0_REG_26__SCAN_IN), .ZN(n2686) );
  INV_X1 U3422 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4050) );
  OR2_X1 U3423 ( .A1(n2953), .A2(n4050), .ZN(n2685) );
  INV_X1 U3424 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3510) );
  NAND2_X1 U3425 ( .A1(n2680), .A2(n3510), .ZN(n2681) );
  NAND2_X1 U3426 ( .A1(n2697), .A2(n2681), .ZN(n3509) );
  INV_X1 U3427 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2682) );
  OR2_X1 U3428 ( .A1(n2955), .A2(n2682), .ZN(n2683) );
  NAND2_X1 U3429 ( .A1(n3805), .A2(n2611), .ZN(n2688) );
  NAND2_X1 U3430 ( .A1(n3586), .A2(DATAI_26_), .ZN(n3513) );
  OR2_X1 U3431 ( .A1(n3513), .A2(n2713), .ZN(n2687) );
  NAND2_X1 U3432 ( .A1(n2688), .A2(n2687), .ZN(n2690) );
  XNOR2_X1 U3433 ( .A(n2690), .B(n2689), .ZN(n2695) );
  INV_X1 U3434 ( .A(n2695), .ZN(n2693) );
  NOR2_X1 U3435 ( .A1(n3513), .A2(n2339), .ZN(n2691) );
  AOI21_X1 U3436 ( .B1(n3805), .B2(n2014), .A(n2691), .ZN(n2694) );
  INV_X1 U3437 ( .A(n2694), .ZN(n2692) );
  NAND2_X1 U3438 ( .A1(n2693), .A2(n2692), .ZN(n3506) );
  AND2_X1 U3439 ( .A1(n2695), .A2(n2694), .ZN(n3505) );
  AOI21_X1 U3440 ( .B1(n3504), .B2(n3506), .A(n3505), .ZN(n2784) );
  NAND2_X1 U3441 ( .A1(n2915), .A2(REG0_REG_27__SCAN_IN), .ZN(n2702) );
  INV_X1 U3442 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2696) );
  OR2_X1 U3443 ( .A1(n2953), .A2(n2696), .ZN(n2701) );
  INV_X1 U3444 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4076) );
  AND2_X1 U3445 ( .A1(n2697), .A2(n4076), .ZN(n2698) );
  INV_X1 U3446 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3769) );
  OR2_X1 U3447 ( .A1(n2955), .A2(n3769), .ZN(n2699) );
  NAND2_X1 U3448 ( .A1(n3586), .A2(DATAI_27_), .ZN(n2867) );
  OAI22_X1 U3449 ( .A1(n3511), .A2(n2703), .B1(n2339), .B2(n2867), .ZN(n2747)
         );
  OAI22_X1 U3450 ( .A1(n3511), .A2(n2339), .B1(n2713), .B2(n2867), .ZN(n2704)
         );
  XNOR2_X1 U3451 ( .A(n2704), .B(n2716), .ZN(n2748) );
  XOR2_X1 U3452 ( .A(n2747), .B(n2748), .Z(n2783) );
  NAND2_X1 U3453 ( .A1(n2784), .A2(n2783), .ZN(n2782) );
  NAND2_X1 U3454 ( .A1(n2915), .A2(REG0_REG_28__SCAN_IN), .ZN(n2712) );
  INV_X1 U3455 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2881) );
  OR2_X1 U3456 ( .A1(n2953), .A2(n2881), .ZN(n2711) );
  NAND2_X1 U3457 ( .A1(n2705), .A2(REG3_REG_28__SCAN_IN), .ZN(n3741) );
  INV_X1 U34580 ( .A(n2705), .ZN(n2707) );
  INV_X1 U34590 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U3460 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  NAND2_X1 U3461 ( .A1(n3741), .A2(n2708), .ZN(n3416) );
  INV_X1 U3462 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3417) );
  OR2_X1 U3463 ( .A1(n2319), .A2(n3417), .ZN(n2709) );
  NAND2_X1 U3464 ( .A1(n3776), .A2(n2611), .ZN(n2715) );
  NAND2_X1 U3465 ( .A1(n3586), .A2(DATAI_28_), .ZN(n2887) );
  OR2_X1 U3466 ( .A1(n2887), .A2(n2713), .ZN(n2714) );
  NAND2_X1 U34670 ( .A1(n2715), .A2(n2714), .ZN(n2717) );
  XNOR2_X1 U3468 ( .A(n2717), .B(n2716), .ZN(n2720) );
  NOR2_X1 U34690 ( .A1(n2887), .A2(n2339), .ZN(n2718) );
  AOI21_X1 U3470 ( .B1(n3776), .B2(n2014), .A(n2718), .ZN(n2719) );
  XNOR2_X1 U34710 ( .A(n2720), .B(n2719), .ZN(n2749) );
  INV_X1 U3472 ( .A(n2749), .ZN(n2746) );
  NAND2_X1 U34730 ( .A1(n2721), .A2(n2913), .ZN(n2722) );
  MUX2_X1 U3474 ( .A(n2721), .B(n2722), .S(B_REG_SCAN_IN), .Z(n2723) );
  INV_X1 U34750 ( .A(n2910), .ZN(n2726) );
  INV_X1 U3476 ( .A(D_REG_0__SCAN_IN), .ZN(n3415) );
  INV_X1 U34770 ( .A(n2912), .ZN(n2724) );
  NOR2_X1 U3478 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_9__SCAN_IN), .ZN(n4114) );
  NOR4_X1 U34790 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2729) );
  NOR4_X1 U3480 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2728) );
  NOR4_X1 U34810 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2727) );
  AND4_X1 U3482 ( .A1(n4114), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(n2735)
         );
  NOR4_X1 U34830 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2733) );
  NOR4_X1 U3484 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2732) );
  NOR4_X1 U34850 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2731) );
  NOR4_X1 U3486 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2730) );
  AND4_X1 U34870 ( .A1(n2733), .A2(n2732), .A3(n2731), .A4(n2730), .ZN(n2734)
         );
  AND2_X1 U3488 ( .A1(n2735), .A2(n2734), .ZN(n2736) );
  NOR2_X1 U34890 ( .A1(n2910), .A2(n2736), .ZN(n2879) );
  INV_X1 U3490 ( .A(n2913), .ZN(n4227) );
  OAI22_X1 U34910 ( .A1(n2910), .A2(D_REG_1__SCAN_IN), .B1(n2912), .B2(n4227), 
        .ZN(n3068) );
  NOR2_X1 U3492 ( .A1(n2879), .A2(n3068), .ZN(n2737) );
  NAND2_X1 U34930 ( .A1(n2919), .A2(STATE_REG_SCAN_IN), .ZN(n4464) );
  AND2_X1 U3494 ( .A1(n2769), .A2(n3736), .ZN(n2752) );
  INV_X1 U34950 ( .A(n2752), .ZN(n2741) );
  NAND2_X1 U3496 ( .A1(n4448), .A2(n2741), .ZN(n2743) );
  NAND2_X1 U34970 ( .A1(n3670), .A2(n2742), .ZN(n2871) );
  NAND2_X1 U3498 ( .A1(n2743), .A2(n2871), .ZN(n2744) );
  NOR2_X1 U34990 ( .A1(n2918), .A2(n2744), .ZN(n2745) );
  NAND2_X1 U3500 ( .A1(n2746), .A2(n3496), .ZN(n2781) );
  NAND2_X1 U35010 ( .A1(n2748), .A2(n2747), .ZN(n2750) );
  NAND2_X1 U3502 ( .A1(n2782), .A2(n2040), .ZN(n2780) );
  NOR3_X1 U35030 ( .A1(n2750), .A2(n2749), .A3(n3520), .ZN(n2778) );
  INV_X1 U3504 ( .A(n2774), .ZN(n2771) );
  AND2_X1 U35050 ( .A1(n2769), .A2(n4229), .ZN(n4451) );
  NAND2_X1 U35060 ( .A1(n4538), .A2(n2751), .ZN(n2877) );
  NAND2_X1 U35070 ( .A1(n2771), .A2(n2877), .ZN(n2988) );
  NOR2_X1 U35080 ( .A1(n2871), .A2(n2752), .ZN(n2878) );
  INV_X1 U35090 ( .A(n2919), .ZN(n2753) );
  NOR2_X1 U35100 ( .A1(n2878), .A2(n2753), .ZN(n2754) );
  AND2_X1 U35110 ( .A1(n2256), .A2(n2754), .ZN(n2755) );
  NAND2_X1 U35120 ( .A1(n2988), .A2(n2755), .ZN(n2756) );
  NAND3_X1 U35130 ( .A1(n2757), .A2(n3670), .A3(n3736), .ZN(n2758) );
  OR2_X1 U35140 ( .A1(n2339), .A2(n2758), .ZN(n3669) );
  OR2_X1 U35150 ( .A1(n2055), .A2(n2759), .ZN(n2761) );
  XNOR2_X1 U35160 ( .A(n2761), .B(n2760), .ZN(n4234) );
  INV_X1 U35170 ( .A(n4234), .ZN(n2963) );
  NOR2_X1 U35180 ( .A1(n3669), .A2(n2963), .ZN(n2762) );
  NAND2_X1 U35190 ( .A1(n2295), .A2(REG1_REG_29__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U35200 ( .A1(n2915), .A2(REG0_REG_29__SCAN_IN), .ZN(n2767) );
  OR2_X1 U35210 ( .A1(n2763), .A2(n3741), .ZN(n2766) );
  INV_X1 U35220 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2764) );
  OR2_X1 U35230 ( .A1(n2955), .A2(n2764), .ZN(n2765) );
  NAND4_X1 U35240 ( .A1(n2768), .A2(n2767), .A3(n2766), .A4(n2765), .ZN(n3675)
         );
  INV_X1 U35250 ( .A(n2769), .ZN(n3664) );
  NAND2_X1 U35260 ( .A1(n4448), .A2(n3664), .ZN(n4389) );
  OR2_X1 U35270 ( .A1(n2918), .A2(n4389), .ZN(n2770) );
  OR2_X1 U35280 ( .A1(n2771), .A2(n2770), .ZN(n2772) );
  NAND2_X1 U35290 ( .A1(n2772), .A2(n4457), .ZN(n3487) );
  INV_X1 U35300 ( .A(n2887), .ZN(n3754) );
  AOI22_X1 U35310 ( .A1(n3500), .A2(n3675), .B1(n3487), .B2(n3754), .ZN(n2776)
         );
  NOR2_X1 U35320 ( .A1(n3669), .A2(n4234), .ZN(n2773) );
  AOI22_X1 U35330 ( .A1(n3488), .A2(n3788), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2775) );
  OAI211_X1 U35340 ( .C1(n3503), .C2(n3416), .A(n2776), .B(n2775), .ZN(n2777)
         );
  NOR2_X1 U35350 ( .A1(n2778), .A2(n2777), .ZN(n2779) );
  OAI211_X1 U35360 ( .C1(n2782), .C2(n2781), .A(n2780), .B(n2779), .ZN(U3217)
         );
  XNOR2_X1 U35370 ( .A(n2784), .B(n2783), .ZN(n2789) );
  AOI22_X1 U35380 ( .A1(n3488), .A2(n3805), .B1(n3487), .B2(n3775), .ZN(n2786)
         );
  AOI22_X1 U35390 ( .A1(n3500), .A2(n3776), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n2785) );
  OAI211_X1 U35400 ( .C1(n3768), .C2(n3503), .A(n2786), .B(n2785), .ZN(n2787)
         );
  INV_X1 U35410 ( .A(n2787), .ZN(n2788) );
  OAI21_X1 U35420 ( .B1(n2789), .B2(n3520), .A(n2788), .ZN(U3211) );
  NAND2_X1 U35430 ( .A1(n4436), .A2(n2790), .ZN(n3538) );
  AND2_X1 U35440 ( .A1(n2840), .A2(n2882), .ZN(n4429) );
  NAND2_X1 U35450 ( .A1(n2790), .A2(n4421), .ZN(n2791) );
  NAND2_X1 U35460 ( .A1(n4428), .A2(n2791), .ZN(n3100) );
  INV_X1 U35470 ( .A(n3100), .ZN(n2792) );
  NAND2_X1 U35480 ( .A1(n4424), .A2(n3027), .ZN(n3541) );
  NAND2_X1 U35490 ( .A1(n3137), .A2(n3027), .ZN(n2793) );
  NOR2_X1 U35500 ( .A1(n3690), .A2(n3544), .ZN(n2795) );
  NAND2_X1 U35510 ( .A1(n3690), .A2(n3544), .ZN(n2794) );
  NAND2_X1 U35520 ( .A1(n2796), .A2(n2797), .ZN(n3546) );
  NAND2_X1 U35530 ( .A1(n3123), .A2(n3083), .ZN(n3549) );
  NAND2_X1 U35540 ( .A1(n3546), .A2(n3549), .ZN(n3620) );
  NAND2_X1 U35550 ( .A1(n3066), .A2(n3620), .ZN(n2799) );
  NAND2_X1 U35560 ( .A1(n3123), .A2(n2797), .ZN(n2798) );
  AND2_X1 U35570 ( .A1(n3688), .A2(n3127), .ZN(n2800) );
  NOR2_X1 U35580 ( .A1(n3687), .A2(n2883), .ZN(n2802) );
  NAND2_X1 U35590 ( .A1(n3687), .A2(n2883), .ZN(n2801) );
  NAND2_X1 U35600 ( .A1(n3151), .A2(n3180), .ZN(n2849) );
  NAND2_X1 U35610 ( .A1(n3240), .A2(n3174), .ZN(n3559) );
  NAND2_X1 U35620 ( .A1(n2849), .A2(n3559), .ZN(n3621) );
  NAND2_X1 U35630 ( .A1(n3183), .A2(n3621), .ZN(n2804) );
  NAND2_X1 U35640 ( .A1(n3240), .A2(n3180), .ZN(n2803) );
  AND2_X1 U35650 ( .A1(n3686), .A2(n3198), .ZN(n2806) );
  NAND2_X1 U35660 ( .A1(n3221), .A2(n3237), .ZN(n2805) );
  NOR2_X1 U35670 ( .A1(n3685), .A2(n3209), .ZN(n2807) );
  INV_X1 U35680 ( .A(n3209), .ZN(n3220) );
  AND2_X1 U35690 ( .A1(n4393), .A2(n2884), .ZN(n2809) );
  INV_X1 U35700 ( .A(n4393), .ZN(n3255) );
  INV_X1 U35710 ( .A(n2884), .ZN(n3300) );
  NAND2_X1 U35720 ( .A1(n3255), .A2(n3300), .ZN(n2808) );
  OAI21_X2 U35730 ( .B1(n3298), .B2(n2809), .A(n2808), .ZN(n4386) );
  NAND2_X1 U35740 ( .A1(n3301), .A2(n4402), .ZN(n3528) );
  NAND2_X1 U35750 ( .A1(n3684), .A2(n4390), .ZN(n3526) );
  NAND2_X1 U35760 ( .A1(n3528), .A2(n3526), .ZN(n4387) );
  NOR2_X1 U35770 ( .A1(n3684), .A2(n4402), .ZN(n2810) );
  NAND2_X1 U35780 ( .A1(n3682), .A2(n3288), .ZN(n2812) );
  NOR2_X1 U35790 ( .A1(n3682), .A2(n3288), .ZN(n2811) );
  NAND2_X1 U35800 ( .A1(n2813), .A2(n3347), .ZN(n3534) );
  NAND2_X1 U35810 ( .A1(n3681), .A2(n2814), .ZN(n3522) );
  NOR2_X1 U3582 ( .A1(n3680), .A2(n3400), .ZN(n2817) );
  INV_X1 U3583 ( .A(n3680), .ZN(n3315) );
  INV_X1 U3584 ( .A(n3400), .ZN(n3356) );
  NAND2_X1 U3585 ( .A1(n3467), .A2(n3390), .ZN(n3641) );
  NAND2_X1 U3586 ( .A1(n3645), .A2(n3641), .ZN(n3604) );
  INV_X1 U3587 ( .A(n3467), .ZN(n3961) );
  INV_X1 U3588 ( .A(n3949), .ZN(n3679) );
  NAND2_X1 U3589 ( .A1(n3959), .A2(n3946), .ZN(n3919) );
  INV_X1 U3590 ( .A(n3959), .ZN(n3926) );
  NAND2_X1 U3591 ( .A1(n3926), .A2(n3498), .ZN(n3920) );
  NAND2_X1 U3592 ( .A1(n3919), .A2(n3920), .ZN(n3945) );
  NAND2_X1 U3593 ( .A1(n2820), .A2(n3929), .ZN(n2823) );
  AOI21_X2 U3594 ( .B1(n3914), .B2(n2823), .A(n2822), .ZN(n3904) );
  INV_X1 U3595 ( .A(n3907), .ZN(n3486) );
  NAND2_X1 U3596 ( .A1(n3884), .A2(n3486), .ZN(n3593) );
  NOR2_X1 U3597 ( .A1(n3884), .A2(n3486), .ZN(n3594) );
  NOR2_X1 U3598 ( .A1(n3896), .A2(n3888), .ZN(n2824) );
  NAND2_X1 U3599 ( .A1(n3880), .A2(n3873), .ZN(n3843) );
  INV_X1 U3600 ( .A(n3880), .ZN(n3677) );
  INV_X1 U3601 ( .A(n2863), .ZN(n2826) );
  INV_X1 U3602 ( .A(n3872), .ZN(n3676) );
  NOR2_X1 U3603 ( .A1(n3676), .A2(n3847), .ZN(n2829) );
  NAND2_X1 U3604 ( .A1(n3677), .A2(n3873), .ZN(n3839) );
  OAI22_X1 U3605 ( .A1(n2829), .A2(n3839), .B1(n3872), .B2(n3853), .ZN(n2830)
         );
  INV_X1 U3606 ( .A(n3832), .ZN(n3474) );
  INV_X1 U3607 ( .A(n3824), .ZN(n3789) );
  NOR2_X1 U3608 ( .A1(n3789), .A2(n3812), .ZN(n2835) );
  NOR2_X1 U3609 ( .A1(n3779), .A2(n3513), .ZN(n2836) );
  NOR2_X1 U3610 ( .A1(n3788), .A2(n3775), .ZN(n2837) );
  NOR2_X1 U3611 ( .A1(n3776), .A2(n2887), .ZN(n3743) );
  OR2_X1 U3612 ( .A1(n3742), .A2(n3743), .ZN(n3752) );
  XNOR2_X1 U3613 ( .A(n3753), .B(n3752), .ZN(n3422) );
  INV_X1 U3614 ( .A(n3422), .ZN(n2876) );
  XNOR2_X1 U3615 ( .A(n3073), .B(n2838), .ZN(n2839) );
  NAND2_X1 U3616 ( .A1(n2839), .A2(n3736), .ZN(n4430) );
  INV_X1 U3617 ( .A(n4538), .ZN(n4498) );
  INV_X1 U3618 ( .A(n2840), .ZN(n4427) );
  NAND2_X1 U3619 ( .A1(n4427), .A2(n2882), .ZN(n3623) );
  INV_X1 U3620 ( .A(n3623), .ZN(n2842) );
  NAND2_X1 U3621 ( .A1(n2845), .A2(n3105), .ZN(n3104) );
  NAND2_X1 U3622 ( .A1(n3104), .A2(n3539), .ZN(n2846) );
  XNOR2_X1 U3623 ( .A(n3690), .B(n3544), .ZN(n3133) );
  INV_X1 U3624 ( .A(n3690), .ZN(n3543) );
  NAND2_X1 U3625 ( .A1(n3543), .A2(n3544), .ZN(n3545) );
  INV_X1 U3626 ( .A(n3546), .ZN(n2847) );
  INV_X1 U3627 ( .A(n3127), .ZN(n3121) );
  AND2_X1 U3628 ( .A1(n3688), .A2(n3121), .ZN(n3119) );
  INV_X1 U3629 ( .A(n3688), .ZN(n3095) );
  NAND2_X1 U3630 ( .A1(n3095), .A2(n3127), .ZN(n3555) );
  INV_X1 U3631 ( .A(n2883), .ZN(n3157) );
  NAND2_X1 U3632 ( .A1(n3687), .A2(n3157), .ZN(n3554) );
  NAND2_X1 U3633 ( .A1(n3150), .A2(n3554), .ZN(n2848) );
  INV_X1 U3634 ( .A(n3687), .ZN(n3168) );
  NAND2_X1 U3635 ( .A1(n3168), .A2(n2883), .ZN(n3551) );
  NAND2_X1 U3636 ( .A1(n3221), .A2(n3198), .ZN(n3566) );
  NAND2_X1 U3637 ( .A1(n3236), .A2(n3566), .ZN(n2850) );
  NAND2_X1 U3638 ( .A1(n3686), .A2(n3237), .ZN(n3560) );
  AND2_X1 U3639 ( .A1(n3685), .A2(n3220), .ZN(n3203) );
  NAND2_X1 U3640 ( .A1(n3238), .A2(n3209), .ZN(n3567) );
  NAND2_X1 U3641 ( .A1(n4393), .A2(n3300), .ZN(n3525) );
  NAND2_X1 U3642 ( .A1(n3255), .A2(n2884), .ZN(n3524) );
  NAND2_X1 U3643 ( .A1(n2851), .A2(n3524), .ZN(n4388) );
  NAND2_X1 U3644 ( .A1(n4388), .A2(n3526), .ZN(n2852) );
  NAND2_X1 U3645 ( .A1(n2852), .A2(n3528), .ZN(n3268) );
  NOR2_X1 U3646 ( .A1(n3683), .A2(n3273), .ZN(n3530) );
  NAND2_X1 U3647 ( .A1(n3682), .A2(n2136), .ZN(n3282) );
  NAND2_X1 U3648 ( .A1(n3683), .A2(n3273), .ZN(n3280) );
  NAND2_X1 U3649 ( .A1(n3281), .A2(n3529), .ZN(n2853) );
  INV_X1 U3650 ( .A(n3682), .ZN(n3345) );
  NAND2_X1 U3651 ( .A1(n3345), .A2(n3288), .ZN(n3533) );
  NAND2_X1 U3652 ( .A1(n2853), .A2(n3533), .ZN(n3640) );
  NAND2_X1 U3653 ( .A1(n3640), .A2(n3617), .ZN(n3354) );
  NAND2_X1 U3654 ( .A1(n3315), .A2(n3400), .ZN(n3532) );
  NAND2_X1 U3655 ( .A1(n3680), .A2(n3356), .ZN(n3523) );
  NAND2_X1 U3656 ( .A1(n3532), .A2(n3523), .ZN(n3625) );
  INV_X1 U3657 ( .A(n3534), .ZN(n3639) );
  NOR2_X1 U3658 ( .A1(n3625), .A2(n3639), .ZN(n2854) );
  INV_X1 U3659 ( .A(n3915), .ZN(n2857) );
  NAND2_X1 U3660 ( .A1(n3947), .A2(n3929), .ZN(n2855) );
  AND2_X1 U3661 ( .A1(n3920), .A2(n2855), .ZN(n2859) );
  OR2_X1 U3662 ( .A1(n3949), .A2(n2885), .ZN(n3916) );
  NAND2_X1 U3663 ( .A1(n2859), .A2(n3916), .ZN(n3644) );
  NAND2_X1 U3664 ( .A1(n3949), .A2(n2885), .ZN(n3917) );
  NAND2_X1 U3665 ( .A1(n3919), .A2(n3917), .ZN(n2860) );
  NOR2_X1 U3666 ( .A1(n3947), .A2(n3929), .ZN(n2858) );
  AOI21_X1 U3667 ( .B1(n2860), .B2(n2859), .A(n2858), .ZN(n3897) );
  INV_X1 U3668 ( .A(n3884), .ZN(n3924) );
  NAND2_X1 U3669 ( .A1(n3924), .A2(n3486), .ZN(n2861) );
  AND2_X1 U3670 ( .A1(n3897), .A2(n2861), .ZN(n3649) );
  NOR2_X1 U3671 ( .A1(n3649), .A2(n3650), .ZN(n3576) );
  NAND2_X1 U3672 ( .A1(n3896), .A2(n2886), .ZN(n3841) );
  AND2_X1 U3673 ( .A1(n3843), .A2(n3841), .ZN(n3647) );
  NOR2_X1 U3674 ( .A1(n3896), .A2(n2886), .ZN(n3842) );
  NOR2_X1 U3675 ( .A1(n3872), .A2(n3847), .ZN(n3607) );
  NOR2_X1 U3676 ( .A1(n3607), .A2(n2863), .ZN(n3580) );
  INV_X1 U3677 ( .A(n3580), .ZN(n2864) );
  AOI21_X1 U3678 ( .B1(n3842), .B2(n3843), .A(n2864), .ZN(n3652) );
  INV_X1 U3679 ( .A(n3652), .ZN(n2865) );
  NAND2_X1 U3680 ( .A1(n3872), .A2(n3847), .ZN(n3606) );
  NAND2_X1 U3681 ( .A1(n3807), .A2(n3474), .ZN(n3608) );
  NAND2_X1 U3682 ( .A1(n3606), .A2(n3608), .ZN(n3653) );
  NAND2_X1 U3683 ( .A1(n3824), .A2(n3812), .ZN(n3784) );
  NAND2_X1 U3684 ( .A1(n3779), .A2(n3793), .ZN(n3624) );
  NAND2_X1 U3685 ( .A1(n3784), .A2(n3624), .ZN(n3636) );
  INV_X1 U3686 ( .A(n3636), .ZN(n2866) );
  OR2_X1 U3687 ( .A1(n3824), .A2(n3812), .ZN(n3597) );
  NAND2_X1 U3688 ( .A1(n3848), .A2(n3832), .ZN(n3802) );
  AND2_X1 U3689 ( .A1(n3597), .A2(n3802), .ZN(n3783) );
  NAND2_X1 U3690 ( .A1(n3805), .A2(n3513), .ZN(n3633) );
  OAI21_X1 U3691 ( .B1(n3783), .B2(n3636), .A(n3633), .ZN(n3583) );
  AOI21_X1 U3692 ( .B1(n3801), .B2(n2866), .A(n3583), .ZN(n3773) );
  AND2_X1 U3693 ( .A1(n3788), .A2(n2867), .ZN(n3585) );
  NOR2_X1 U3694 ( .A1(n3788), .A2(n2867), .ZN(n3637) );
  NAND2_X1 U3695 ( .A1(n3773), .A2(n3772), .ZN(n3771) );
  INV_X1 U3696 ( .A(n3637), .ZN(n2868) );
  XOR2_X1 U3697 ( .A(n3752), .B(n3745), .Z(n2874) );
  NAND2_X1 U3698 ( .A1(n3670), .A2(n4229), .ZN(n2870) );
  NAND2_X1 U3699 ( .A1(n3664), .A2(n2742), .ZN(n2869) );
  INV_X1 U3700 ( .A(n2871), .ZN(n2920) );
  AOI22_X1 U3701 ( .A1(n3675), .A2(n4423), .B1(n4422), .B2(n3754), .ZN(n2872)
         );
  OAI21_X1 U3702 ( .B1(n3511), .B2(n4426), .A(n2872), .ZN(n2873) );
  INV_X1 U3703 ( .A(n3418), .ZN(n2875) );
  NAND2_X1 U3704 ( .A1(n3068), .A2(n2877), .ZN(n2880) );
  MUX2_X1 U3705 ( .A(n2881), .B(n2894), .S(n4558), .Z(n2891) );
  NAND2_X1 U3706 ( .A1(n4450), .A2(n4436), .ZN(n4435) );
  NAND2_X1 U3707 ( .A1(n3178), .A2(n3237), .ZN(n3234) );
  NAND2_X1 U3708 ( .A1(n3373), .A2(n3372), .ZN(n3964) );
  NAND2_X1 U3709 ( .A1(n3851), .A2(n3832), .ZN(n3831) );
  OR2_X1 U3710 ( .A1(n3767), .A2(n2887), .ZN(n2888) );
  NAND2_X1 U3711 ( .A1(n2891), .A2(n2890), .ZN(U3546) );
  INV_X1 U3712 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2895) );
  INV_X1 U3713 ( .A(n2892), .ZN(n3069) );
  MUX2_X1 U3714 ( .A(n2895), .B(n2894), .S(n4544), .Z(n2898) );
  NAND2_X1 U3715 ( .A1(n2898), .A2(n2897), .ZN(U3514) );
  INV_X1 U3716 ( .A(DATAI_1_), .ZN(n2899) );
  MUX2_X1 U3717 ( .A(n2938), .B(n2899), .S(U3149), .Z(n2900) );
  INV_X1 U3718 ( .A(n2900), .ZN(U3351) );
  INV_X1 U3719 ( .A(DATAI_3_), .ZN(n2901) );
  MUX2_X1 U3720 ( .A(n2901), .B(n2147), .S(STATE_REG_SCAN_IN), .Z(n2902) );
  INV_X1 U3721 ( .A(n2902), .ZN(U3349) );
  INV_X1 U3722 ( .A(DATAI_26_), .ZN(n2904) );
  NAND2_X1 U3723 ( .A1(n2912), .A2(STATE_REG_SCAN_IN), .ZN(n2903) );
  OAI21_X1 U3724 ( .B1(STATE_REG_SCAN_IN), .B2(n2904), .A(n2903), .ZN(U3326)
         );
  INV_X1 U3725 ( .A(DATAI_22_), .ZN(n2906) );
  NAND2_X1 U3726 ( .A1(n3670), .A2(STATE_REG_SCAN_IN), .ZN(n2905) );
  OAI21_X1 U3727 ( .B1(STATE_REG_SCAN_IN), .B2(n2906), .A(n2905), .ZN(U3330)
         );
  INV_X1 U3728 ( .A(DATAI_21_), .ZN(n2908) );
  NAND2_X1 U3729 ( .A1(n2742), .A2(STATE_REG_SCAN_IN), .ZN(n2907) );
  OAI21_X1 U3730 ( .B1(STATE_REG_SCAN_IN), .B2(n2908), .A(n2907), .ZN(U3331)
         );
  INV_X1 U3731 ( .A(DATAI_20_), .ZN(n4072) );
  NAND2_X1 U3732 ( .A1(n3664), .A2(STATE_REG_SCAN_IN), .ZN(n2909) );
  OAI21_X1 U3733 ( .B1(STATE_REG_SCAN_IN), .B2(n4072), .A(n2909), .ZN(U3332)
         );
  INV_X1 U3734 ( .A(n2918), .ZN(n2911) );
  INV_X1 U3735 ( .A(D_REG_1__SCAN_IN), .ZN(n2914) );
  NOR2_X1 U3736 ( .A1(n2912), .A2(n4464), .ZN(n3414) );
  AOI22_X1 U3737 ( .A1(n4460), .A2(n2914), .B1(n3414), .B2(n2913), .ZN(U3459)
         );
  AOI222_X1 U3738 ( .A1(n2295), .A2(REG1_REG_30__SCAN_IN), .B1(n2916), .B2(
        REG2_REG_30__SCAN_IN), .C1(n2915), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n3748) );
  NAND2_X1 U3739 ( .A1(n3689), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2917) );
  OAI21_X1 U3740 ( .B1(n3748), .B2(n3689), .A(n2917), .ZN(U3580) );
  OR2_X1 U3741 ( .A1(n2919), .A2(U3149), .ZN(n3673) );
  NAND2_X1 U3742 ( .A1(n2918), .A2(n3673), .ZN(n2934) );
  NAND2_X1 U3743 ( .A1(n2920), .A2(n2919), .ZN(n2921) );
  AND2_X1 U3744 ( .A1(n3586), .A2(n2921), .ZN(n2933) );
  NAND2_X1 U3745 ( .A1(n2934), .A2(n2933), .ZN(n4245) );
  NOR2_X1 U3746 ( .A1(n2015), .A2(n2277), .ZN(n2964) );
  INV_X1 U3747 ( .A(n2964), .ZN(n2923) );
  AOI21_X1 U3748 ( .B1(n2923), .B2(n2922), .A(n2974), .ZN(n2932) );
  XNOR2_X1 U3749 ( .A(n2925), .B(n2924), .ZN(n3747) );
  OR2_X1 U3750 ( .A1(n4234), .A2(n3747), .ZN(n3668) );
  NOR2_X2 U3751 ( .A1(n4245), .A2(n3668), .ZN(n4358) );
  NAND2_X1 U3752 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2930) );
  INV_X1 U3753 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4546) );
  MUX2_X1 U3754 ( .A(n4546), .B(REG1_REG_1__SCAN_IN), .S(n2938), .Z(n2927) );
  INV_X1 U3755 ( .A(n2927), .ZN(n2929) );
  INV_X1 U3756 ( .A(n2930), .ZN(n2926) );
  NAND2_X1 U3757 ( .A1(n2927), .A2(n2926), .ZN(n2943) );
  INV_X1 U3758 ( .A(n2943), .ZN(n2928) );
  INV_X1 U3759 ( .A(n3747), .ZN(n4242) );
  AOI211_X1 U3760 ( .C1(n2930), .C2(n2929), .A(n2928), .B(n4354), .ZN(n2931)
         );
  AOI21_X1 U3761 ( .B1(n2932), .B2(n4358), .A(n2931), .ZN(n2937) );
  INV_X1 U3762 ( .A(n2933), .ZN(n2935) );
  AOI22_X1 U3763 ( .A1(n4378), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n2936) );
  OAI211_X1 U3764 ( .C1(n2938), .C2(n4385), .A(n2937), .B(n2936), .ZN(U3241)
         );
  INV_X1 U3765 ( .A(n4232), .ZN(n2940) );
  NOR2_X1 U3766 ( .A1(n2938), .A2(n2235), .ZN(n2969) );
  MUX2_X1 U3767 ( .A(n2296), .B(REG2_REG_2__SCAN_IN), .S(n4232), .Z(n2971) );
  INV_X1 U3768 ( .A(n2971), .ZN(n2939) );
  OAI21_X1 U3769 ( .B1(n2974), .B2(n2969), .A(n2939), .ZN(n2972) );
  XNOR2_X1 U3770 ( .A(n3009), .B(REG2_REG_3__SCAN_IN), .ZN(n2947) );
  INV_X1 U3771 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U3772 ( .A1(n2941), .A2(REG1_REG_1__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3773 ( .A1(n2943), .A2(n2942), .ZN(n2976) );
  INV_X1 U3774 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4548) );
  MUX2_X1 U3775 ( .A(REG1_REG_2__SCAN_IN), .B(n4548), .S(n4232), .Z(n2977) );
  NAND2_X1 U3776 ( .A1(n2976), .A2(n2977), .ZN(n2975) );
  NAND2_X1 U3777 ( .A1(n4232), .A2(REG1_REG_2__SCAN_IN), .ZN(n2944) );
  AOI211_X1 U3778 ( .C1(n4550), .C2(n2945), .A(n2997), .B(n4354), .ZN(n2946)
         );
  AOI21_X1 U3779 ( .B1(n4358), .B2(n2947), .A(n2946), .ZN(n2949) );
  NOR2_X1 U3780 ( .A1(STATE_REG_SCAN_IN), .A2(n2332), .ZN(n3048) );
  AOI21_X1 U3781 ( .B1(n4378), .B2(ADDR_REG_3__SCAN_IN), .A(n3048), .ZN(n2948)
         );
  OAI211_X1 U3782 ( .C1(n2147), .C2(n4385), .A(n2949), .B(n2948), .ZN(U3243)
         );
  NOR2_X1 U3783 ( .A1(n4378), .A2(U4043), .ZN(U3148) );
  INV_X1 U3784 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4119) );
  NAND2_X1 U3785 ( .A1(n3123), .A2(U4043), .ZN(n2950) );
  OAI21_X1 U3786 ( .B1(U4043), .B2(n4119), .A(n2950), .ZN(U3554) );
  INV_X1 U3787 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4120) );
  NAND2_X1 U3788 ( .A1(n3240), .A2(U4043), .ZN(n2951) );
  OAI21_X1 U3789 ( .B1(U4043), .B2(n4120), .A(n2951), .ZN(U3557) );
  INV_X1 U3790 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4015) );
  NAND2_X1 U3791 ( .A1(n2915), .A2(REG0_REG_31__SCAN_IN), .ZN(n2958) );
  INV_X1 U3792 ( .A(REG1_REG_31__SCAN_IN), .ZN(n2952) );
  OR2_X1 U3793 ( .A1(n2953), .A2(n2952), .ZN(n2957) );
  INV_X1 U3794 ( .A(REG2_REG_31__SCAN_IN), .ZN(n2954) );
  OR2_X1 U3795 ( .A1(n2955), .A2(n2954), .ZN(n2956) );
  AND3_X1 U3796 ( .A1(n2958), .A2(n2957), .A3(n2956), .ZN(n3979) );
  INV_X1 U3797 ( .A(n3979), .ZN(n3588) );
  NAND2_X1 U3798 ( .A1(n3588), .A2(U4043), .ZN(n2959) );
  OAI21_X1 U3799 ( .B1(U4043), .B2(n4015), .A(n2959), .ZN(U3581) );
  INV_X1 U3800 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U3801 ( .A1(n2840), .A2(U4043), .ZN(n2960) );
  OAI21_X1 U3802 ( .B1(U4043), .B2(n4118), .A(n2960), .ZN(U3550) );
  AOI21_X1 U3803 ( .B1(n4242), .B2(n2277), .A(n4234), .ZN(n4241) );
  XNOR2_X1 U3804 ( .A(n2961), .B(n2962), .ZN(n2996) );
  NAND3_X1 U3805 ( .A1(n2996), .A2(n2963), .A3(n3747), .ZN(n2967) );
  INV_X1 U3806 ( .A(n3668), .ZN(n2965) );
  AOI21_X1 U3807 ( .B1(n2965), .B2(n2964), .A(n3689), .ZN(n2966) );
  OAI211_X1 U3808 ( .C1(IR_REG_0__SCAN_IN), .C2(n4241), .A(n2967), .B(n2966), 
        .ZN(n3035) );
  INV_X1 U3809 ( .A(n4385), .ZN(n2982) );
  NAND2_X1 U3810 ( .A1(n4378), .A2(ADDR_REG_2__SCAN_IN), .ZN(n2968) );
  OAI21_X1 U3811 ( .B1(STATE_REG_SCAN_IN), .B2(n3103), .A(n2968), .ZN(n2981)
         );
  INV_X1 U3812 ( .A(n2969), .ZN(n2970) );
  NAND2_X1 U3813 ( .A1(n2971), .A2(n2970), .ZN(n2973) );
  OAI211_X1 U3814 ( .C1(n2974), .C2(n2973), .A(n4358), .B(n2972), .ZN(n2979)
         );
  OAI211_X1 U3815 ( .C1(n2977), .C2(n2976), .A(n4380), .B(n2975), .ZN(n2978)
         );
  NAND2_X1 U3816 ( .A1(n2979), .A2(n2978), .ZN(n2980) );
  AOI211_X1 U3817 ( .C1(n4232), .C2(n2982), .A(n2981), .B(n2980), .ZN(n2983)
         );
  NAND2_X1 U3818 ( .A1(n3035), .A2(n2983), .ZN(U3242) );
  XNOR2_X1 U3819 ( .A(n2985), .B(n2984), .ZN(n2992) );
  INV_X1 U3820 ( .A(n2986), .ZN(n2987) );
  NAND2_X1 U3821 ( .A1(n2988), .A2(n2987), .ZN(n3029) );
  AOI22_X1 U3822 ( .A1(n4424), .A2(n3500), .B1(n3488), .B2(n2840), .ZN(n2989)
         );
  OAI21_X1 U3823 ( .B1(n3514), .B2(n4436), .A(n2989), .ZN(n2990) );
  AOI21_X1 U3824 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3029), .A(n2990), .ZN(n2991)
         );
  OAI21_X1 U3825 ( .B1(n2992), .B2(n3520), .A(n2991), .ZN(U3219) );
  OAI22_X1 U3826 ( .A1(n2993), .A2(n3512), .B1(n3514), .B2(n4450), .ZN(n2994)
         );
  AOI21_X1 U3827 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3029), .A(n2994), .ZN(n2995)
         );
  OAI21_X1 U3828 ( .B1(n3520), .B2(n2996), .A(n2995), .ZN(U3229) );
  XNOR2_X1 U3829 ( .A(n2999), .B(n4231), .ZN(n3032) );
  INV_X1 U3830 ( .A(n2999), .ZN(n3000) );
  INV_X1 U3831 ( .A(n3007), .ZN(n4489) );
  AOI22_X1 U3832 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4489), .B1(n3007), .B2(n2355), .ZN(n4248) );
  NOR2_X1 U3833 ( .A1(n3002), .A2(n4264), .ZN(n3003) );
  MUX2_X1 U3834 ( .A(n3004), .B(REG1_REG_7__SCAN_IN), .S(n4230), .Z(n3006) );
  OAI21_X1 U3835 ( .B1(n3691), .B2(n3006), .A(n4380), .ZN(n3005) );
  AOI21_X1 U3836 ( .B1(n3691), .B2(n3006), .A(n3005), .ZN(n3021) );
  INV_X1 U3837 ( .A(n4230), .ZN(n3712) );
  AOI22_X1 U3838 ( .A1(REG2_REG_5__SCAN_IN), .A2(n3007), .B1(n4489), .B2(n3129), .ZN(n4253) );
  INV_X1 U3839 ( .A(n3010), .ZN(n3011) );
  INV_X1 U3840 ( .A(n4231), .ZN(n3041) );
  NAND2_X1 U3841 ( .A1(n4253), .A2(n4252), .ZN(n4251) );
  NAND2_X1 U3842 ( .A1(n4486), .A2(n3013), .ZN(n3014) );
  NAND2_X1 U3843 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4261), .ZN(n4260) );
  NAND2_X1 U3844 ( .A1(n3014), .A2(n4260), .ZN(n3017) );
  MUX2_X1 U3845 ( .A(REG2_REG_7__SCAN_IN), .B(n3015), .S(n4230), .Z(n3016) );
  NAND2_X1 U3846 ( .A1(n3017), .A2(n3016), .ZN(n3711) );
  OAI211_X1 U3847 ( .C1(n3017), .C2(n3016), .A(n4358), .B(n3711), .ZN(n3019)
         );
  AND2_X1 U3848 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3170) );
  AOI21_X1 U3849 ( .B1(n4378), .B2(ADDR_REG_7__SCAN_IN), .A(n3170), .ZN(n3018)
         );
  OAI211_X1 U3850 ( .C1(n4385), .C2(n3712), .A(n3019), .B(n3018), .ZN(n3020)
         );
  OR2_X1 U3851 ( .A1(n3021), .A2(n3020), .ZN(U3247) );
  INV_X1 U3852 ( .A(n3023), .ZN(n3024) );
  AOI21_X1 U3853 ( .B1(n3022), .B2(n3025), .A(n3024), .ZN(n3031) );
  AOI22_X1 U3854 ( .A1(n2790), .A2(n3488), .B1(n3500), .B2(n3690), .ZN(n3026)
         );
  OAI21_X1 U3855 ( .B1(n3514), .B2(n3027), .A(n3026), .ZN(n3028) );
  AOI21_X1 U3856 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3029), .A(n3028), .ZN(n3030)
         );
  OAI21_X1 U3857 ( .B1(n3031), .B2(n3520), .A(n3030), .ZN(U3234) );
  AND2_X1 U3858 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3056) );
  OAI21_X1 U3859 ( .B1(REG1_REG_4__SCAN_IN), .B2(n3032), .A(n4380), .ZN(n3037)
         );
  XNOR2_X1 U3860 ( .A(REG2_REG_4__SCAN_IN), .B(n3033), .ZN(n3034) );
  NAND2_X1 U3861 ( .A1(n4358), .A2(n3034), .ZN(n3036) );
  OAI211_X1 U3862 ( .C1(n3038), .C2(n3037), .A(n3036), .B(n3035), .ZN(n3039)
         );
  AOI211_X1 U3863 ( .C1(n4378), .C2(ADDR_REG_4__SCAN_IN), .A(n3056), .B(n3039), 
        .ZN(n3040) );
  OAI21_X1 U3864 ( .B1(n3041), .B2(n4385), .A(n3040), .ZN(U3244) );
  OAI21_X1 U3865 ( .B1(n3044), .B2(n3043), .A(n3042), .ZN(n3045) );
  NAND2_X1 U3866 ( .A1(n3045), .A2(n3496), .ZN(n3050) );
  INV_X1 U3867 ( .A(n3544), .ZN(n3046) );
  OAI22_X1 U3868 ( .A1(n3137), .A2(n3515), .B1(n3514), .B2(n3046), .ZN(n3047)
         );
  AOI211_X1 U3869 ( .C1(n3500), .C2(n3123), .A(n3048), .B(n3047), .ZN(n3049)
         );
  OAI211_X1 U3870 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3503), .A(n3050), .B(n3049), 
        .ZN(U3215) );
  AND2_X1 U3871 ( .A1(n3042), .A2(n3051), .ZN(n3054) );
  OAI211_X1 U3872 ( .C1(n3054), .C2(n3052), .A(n3496), .B(n3053), .ZN(n3058)
         );
  OAI22_X1 U3873 ( .A1(n3543), .A2(n3515), .B1(n3514), .B2(n3083), .ZN(n3055)
         );
  AOI211_X1 U3874 ( .C1(n3500), .C2(n3688), .A(n3056), .B(n3055), .ZN(n3057)
         );
  OAI211_X1 U3875 ( .C1(n3503), .C2(n3084), .A(n3058), .B(n3057), .ZN(U3227)
         );
  XOR2_X1 U3876 ( .A(n3059), .B(n3060), .Z(n3061) );
  NAND2_X1 U3877 ( .A1(n3061), .A2(n3496), .ZN(n3065) );
  INV_X1 U3878 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3062) );
  NOR2_X1 U3879 ( .A1(STATE_REG_SCAN_IN), .A2(n3062), .ZN(n4249) );
  OAI22_X1 U3880 ( .A1(n2796), .A2(n3515), .B1(n3514), .B2(n3121), .ZN(n3063)
         );
  AOI211_X1 U3881 ( .C1(n3500), .C2(n3687), .A(n4249), .B(n3063), .ZN(n3064)
         );
  OAI211_X1 U3882 ( .C1(n3503), .C2(n3128), .A(n3065), .B(n3064), .ZN(U3224)
         );
  INV_X1 U3883 ( .A(n3620), .ZN(n3075) );
  XNOR2_X1 U3884 ( .A(n3066), .B(n3075), .ZN(n4514) );
  INV_X1 U3885 ( .A(n4514), .ZN(n3088) );
  INV_X1 U3886 ( .A(n3067), .ZN(n3071) );
  INV_X1 U3887 ( .A(n3068), .ZN(n3070) );
  NAND3_X1 U3888 ( .A1(n3071), .A2(n3070), .A3(n3069), .ZN(n3072) );
  NAND2_X2 U3889 ( .A1(n3072), .A2(n4457), .ZN(n4453) );
  AND2_X1 U3890 ( .A1(n3073), .A2(n4229), .ZN(n3074) );
  NAND2_X1 U3891 ( .A1(n4453), .A2(n3074), .ZN(n3117) );
  NAND2_X1 U3892 ( .A1(n4514), .A2(n4445), .ZN(n3082) );
  XNOR2_X1 U3893 ( .A(n3076), .B(n3075), .ZN(n3080) );
  NAND2_X1 U3894 ( .A1(n3690), .A2(n4394), .ZN(n3078) );
  NAND2_X1 U3895 ( .A1(n3688), .A2(n4423), .ZN(n3077) );
  OAI211_X1 U3896 ( .C1(n4389), .C2(n3083), .A(n3078), .B(n3077), .ZN(n3079)
         );
  AOI21_X1 U3897 ( .B1(n3080), .B2(n4444), .A(n3079), .ZN(n3081) );
  NAND2_X1 U3898 ( .A1(n3082), .A2(n3081), .ZN(n4518) );
  OAI211_X1 U3899 ( .C1(n3145), .C2(n3083), .A(n4537), .B(n3126), .ZN(n4515)
         );
  OAI22_X1 U3900 ( .A1(n4515), .A2(n4229), .B1(n4457), .B2(n3084), .ZN(n3085)
         );
  OAI21_X1 U3901 ( .B1(n4518), .B2(n3085), .A(n4453), .ZN(n3087) );
  NAND2_X1 U3902 ( .A1(n4442), .A2(REG2_REG_4__SCAN_IN), .ZN(n3086) );
  OAI211_X1 U3903 ( .C1(n3088), .C2(n3117), .A(n3087), .B(n3086), .ZN(U3286)
         );
  INV_X1 U3904 ( .A(n3090), .ZN(n3092) );
  NAND2_X1 U3905 ( .A1(n3092), .A2(n3091), .ZN(n3093) );
  XNOR2_X1 U3906 ( .A(n3089), .B(n3093), .ZN(n3094) );
  NAND2_X1 U3907 ( .A1(n3094), .A2(n3496), .ZN(n3098) );
  AND2_X1 U3908 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n4259) );
  OAI22_X1 U3909 ( .A1(n3095), .A2(n3515), .B1(n3514), .B2(n3157), .ZN(n3096)
         );
  AOI211_X1 U3910 ( .C1(n3500), .C2(n3240), .A(n4259), .B(n3096), .ZN(n3097)
         );
  OAI211_X1 U3911 ( .C1(n3503), .C2(n3158), .A(n3098), .B(n3097), .ZN(U3236)
         );
  INV_X1 U3912 ( .A(n3117), .ZN(n4443) );
  NAND2_X1 U3913 ( .A1(n3100), .A2(n3105), .ZN(n3101) );
  NAND2_X1 U3914 ( .A1(n3099), .A2(n3101), .ZN(n4507) );
  NAND2_X1 U3915 ( .A1(n4435), .A2(n3107), .ZN(n4503) );
  NAND3_X1 U3916 ( .A1(n4438), .A2(n4504), .A3(n4503), .ZN(n3102) );
  OAI21_X1 U3917 ( .B1(n4457), .B2(n3103), .A(n3102), .ZN(n3114) );
  NAND2_X1 U3918 ( .A1(n3104), .A2(n3106), .ZN(n3110) );
  AOI22_X1 U3919 ( .A1(n3690), .A2(n4423), .B1(n3107), .B2(n4422), .ZN(n3108)
         );
  OAI21_X1 U3920 ( .B1(n2993), .B2(n4426), .A(n3108), .ZN(n3109) );
  AOI21_X1 U3921 ( .B1(n3110), .B2(n4444), .A(n3109), .ZN(n3112) );
  NAND2_X1 U3922 ( .A1(n4507), .A2(n4445), .ZN(n3111) );
  NAND2_X1 U3923 ( .A1(n3112), .A2(n3111), .ZN(n4505) );
  MUX2_X1 U3924 ( .A(REG2_REG_2__SCAN_IN), .B(n4505), .S(n4453), .Z(n3113) );
  AOI211_X1 U3925 ( .C1(n4443), .C2(n4507), .A(n3114), .B(n3113), .ZN(n3115)
         );
  INV_X1 U3926 ( .A(n3115), .ZN(U3288) );
  NAND2_X1 U3927 ( .A1(n4453), .A2(n4445), .ZN(n3116) );
  INV_X1 U3928 ( .A(n3119), .ZN(n3548) );
  NAND2_X1 U3929 ( .A1(n3548), .A2(n3555), .ZN(n3612) );
  XNOR2_X1 U3930 ( .A(n3118), .B(n3612), .ZN(n4521) );
  XOR2_X1 U3931 ( .A(n3612), .B(n3120), .Z(n3125) );
  OAI22_X1 U3932 ( .A1(n3168), .A2(n4447), .B1(n4389), .B2(n3121), .ZN(n3122)
         );
  AOI21_X1 U3933 ( .B1(n4394), .B2(n3123), .A(n3122), .ZN(n3124) );
  OAI21_X1 U3934 ( .B1(n3125), .B2(n4396), .A(n3124), .ZN(n4522) );
  NAND2_X1 U3935 ( .A1(n4522), .A2(n4453), .ZN(n3132) );
  AOI21_X1 U3936 ( .B1(n3127), .B2(n3126), .A(n2050), .ZN(n4524) );
  OAI22_X1 U3937 ( .A1(n4453), .A2(n3129), .B1(n3128), .B2(n4457), .ZN(n3130)
         );
  AOI21_X1 U3938 ( .B1(n4524), .B2(n4438), .A(n3130), .ZN(n3131) );
  OAI211_X1 U3939 ( .C1(n3974), .C2(n4521), .A(n3132), .B(n3131), .ZN(U3285)
         );
  INV_X1 U3940 ( .A(n3133), .ZN(n3630) );
  XNOR2_X1 U3941 ( .A(n3134), .B(n3630), .ZN(n4510) );
  NAND2_X1 U3942 ( .A1(n4510), .A2(n4445), .ZN(n3143) );
  NAND3_X1 U3943 ( .A1(n3104), .A2(n3539), .A3(n3630), .ZN(n3135) );
  NAND2_X1 U3944 ( .A1(n3136), .A2(n3135), .ZN(n3141) );
  OR2_X1 U3945 ( .A1(n3137), .A2(n4426), .ZN(n3139) );
  NAND2_X1 U3946 ( .A1(n3544), .A2(n4422), .ZN(n3138) );
  OAI211_X1 U3947 ( .C1(n2796), .C2(n4447), .A(n3139), .B(n3138), .ZN(n3140)
         );
  AOI21_X1 U3948 ( .B1(n3141), .B2(n4444), .A(n3140), .ZN(n3142) );
  AND2_X1 U3949 ( .A1(n3143), .A2(n3142), .ZN(n4512) );
  AND2_X1 U3950 ( .A1(n4504), .A2(n3544), .ZN(n3144) );
  NOR2_X1 U3951 ( .A1(n3145), .A2(n3144), .ZN(n4509) );
  INV_X1 U3952 ( .A(n4509), .ZN(n3147) );
  INV_X1 U3953 ( .A(n4457), .ZN(n4434) );
  AOI22_X1 U3954 ( .A1(n4442), .A2(REG2_REG_3__SCAN_IN), .B1(n4434), .B2(n2332), .ZN(n3146) );
  OAI21_X1 U3955 ( .B1(n3968), .B2(n3147), .A(n3146), .ZN(n3148) );
  AOI21_X1 U3956 ( .B1(n4510), .B2(n4443), .A(n3148), .ZN(n3149) );
  OAI21_X1 U3957 ( .B1(n4512), .B2(n4442), .A(n3149), .ZN(U3287) );
  NAND2_X1 U3958 ( .A1(n3551), .A2(n3554), .ZN(n3619) );
  XNOR2_X1 U3959 ( .A(n3150), .B(n3619), .ZN(n3154) );
  OAI22_X1 U3960 ( .A1(n3151), .A2(n4447), .B1(n4389), .B2(n3157), .ZN(n3152)
         );
  AOI21_X1 U3961 ( .B1(n4394), .B2(n3688), .A(n3152), .ZN(n3153) );
  OAI21_X1 U3962 ( .B1(n3154), .B2(n4396), .A(n3153), .ZN(n3187) );
  INV_X1 U3963 ( .A(n3187), .ZN(n3163) );
  XNOR2_X1 U3964 ( .A(n3155), .B(n3619), .ZN(n3188) );
  INV_X1 U3965 ( .A(n3156), .ZN(n3179) );
  OAI21_X1 U3966 ( .B1(n2050), .B2(n3157), .A(n3179), .ZN(n3193) );
  NOR2_X1 U3967 ( .A1(n3193), .A2(n3968), .ZN(n3161) );
  OAI22_X1 U3968 ( .A1(n4453), .A2(n3159), .B1(n3158), .B2(n4457), .ZN(n3160)
         );
  AOI211_X1 U3969 ( .C1(n3188), .C2(n3905), .A(n3161), .B(n3160), .ZN(n3162)
         );
  OAI21_X1 U3970 ( .B1(n3163), .B2(n4442), .A(n3162), .ZN(U3284) );
  AOI21_X1 U3971 ( .B1(n3164), .B2(n3165), .A(n3520), .ZN(n3167) );
  NAND2_X1 U3972 ( .A1(n3167), .A2(n3166), .ZN(n3172) );
  OAI22_X1 U3973 ( .A1(n3168), .A2(n3515), .B1(n3514), .B2(n3174), .ZN(n3169)
         );
  AOI211_X1 U3974 ( .C1(n3500), .C2(n3686), .A(n3170), .B(n3169), .ZN(n3171)
         );
  OAI211_X1 U3975 ( .C1(n3503), .C2(n3181), .A(n3172), .B(n3171), .ZN(U3210)
         );
  XNOR2_X1 U3976 ( .A(n3173), .B(n3621), .ZN(n3177) );
  OAI22_X1 U3977 ( .A1(n3221), .A2(n4447), .B1(n4389), .B2(n3174), .ZN(n3175)
         );
  AOI21_X1 U3978 ( .B1(n4394), .B2(n3687), .A(n3175), .ZN(n3176) );
  OAI21_X1 U3979 ( .B1(n3177), .B2(n4396), .A(n3176), .ZN(n4526) );
  INV_X1 U3980 ( .A(n4526), .ZN(n3186) );
  AOI211_X1 U3981 ( .C1(n3180), .C2(n3179), .A(n3992), .B(n3178), .ZN(n4527)
         );
  OAI22_X1 U3982 ( .A1(n4453), .A2(n3015), .B1(n3181), .B2(n4457), .ZN(n3182)
         );
  AOI21_X1 U3983 ( .B1(n4527), .B2(n3954), .A(n3182), .ZN(n3185) );
  XOR2_X1 U3984 ( .A(n3183), .B(n3621), .Z(n4528) );
  NAND2_X1 U3985 ( .A1(n4528), .A2(n3905), .ZN(n3184) );
  OAI211_X1 U3986 ( .C1(n3186), .C2(n4442), .A(n3185), .B(n3184), .ZN(U3283)
         );
  AOI21_X1 U3987 ( .B1(n4534), .B2(n3188), .A(n3187), .ZN(n3190) );
  MUX2_X1 U3988 ( .A(n2374), .B(n3190), .S(n4558), .Z(n3189) );
  OAI21_X1 U3989 ( .B1(n3193), .B2(n4168), .A(n3189), .ZN(U3524) );
  INV_X1 U3990 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3191) );
  MUX2_X1 U3991 ( .A(n3191), .B(n3190), .S(n4544), .Z(n3192) );
  OAI21_X1 U3992 ( .B1(n3193), .B2(n4221), .A(n3192), .ZN(U3479) );
  XOR2_X1 U3993 ( .A(n3195), .B(n3194), .Z(n3196) );
  XNOR2_X1 U3994 ( .A(n3197), .B(n3196), .ZN(n3202) );
  AOI22_X1 U3995 ( .A1(n3240), .A2(n3488), .B1(n3487), .B2(n3198), .ZN(n3199)
         );
  NAND2_X1 U3996 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4268) );
  OAI211_X1 U3997 ( .C1(n3238), .C2(n3512), .A(n3199), .B(n4268), .ZN(n3200)
         );
  AOI21_X1 U3998 ( .B1(n4413), .B2(n3518), .A(n3200), .ZN(n3201) );
  OAI21_X1 U3999 ( .B1(n3202), .B2(n3520), .A(n3201), .ZN(U3218) );
  INV_X1 U4000 ( .A(n3203), .ZN(n3568) );
  NAND2_X1 U4001 ( .A1(n3568), .A2(n3567), .ZN(n3613) );
  XNOR2_X1 U4002 ( .A(n3204), .B(n3613), .ZN(n3207) );
  AOI22_X1 U4003 ( .A1(n4393), .A2(n4423), .B1(n4422), .B2(n3209), .ZN(n3205)
         );
  OAI21_X1 U4004 ( .B1(n3221), .B2(n4426), .A(n3205), .ZN(n3206) );
  AOI21_X1 U4005 ( .B1(n3207), .B2(n4444), .A(n3206), .ZN(n4530) );
  XNOR2_X1 U4006 ( .A(n3208), .B(n3613), .ZN(n4533) );
  NAND2_X1 U4007 ( .A1(n3234), .A2(n3209), .ZN(n3210) );
  NAND2_X1 U4008 ( .A1(n3295), .A2(n3210), .ZN(n4531) );
  INV_X1 U4009 ( .A(n3211), .ZN(n3223) );
  AOI22_X1 U4010 ( .A1(n4442), .A2(REG2_REG_9__SCAN_IN), .B1(n3223), .B2(n4434), .ZN(n3212) );
  OAI21_X1 U4011 ( .B1(n4531), .B2(n3968), .A(n3212), .ZN(n3213) );
  AOI21_X1 U4012 ( .B1(n4533), .B2(n3905), .A(n3213), .ZN(n3214) );
  OAI21_X1 U4013 ( .B1(n4530), .B2(n4442), .A(n3214), .ZN(U3281) );
  INV_X1 U4014 ( .A(n3215), .ZN(n3216) );
  AOI21_X1 U4015 ( .B1(n3218), .B2(n3217), .A(n3216), .ZN(n3226) );
  NOR2_X1 U4016 ( .A1(STATE_REG_SCAN_IN), .A2(n3219), .ZN(n4285) );
  OAI22_X1 U4017 ( .A1(n3221), .A2(n3515), .B1(n3514), .B2(n3220), .ZN(n3222)
         );
  AOI211_X1 U4018 ( .C1(n3500), .C2(n4393), .A(n4285), .B(n3222), .ZN(n3225)
         );
  NAND2_X1 U4019 ( .A1(n3518), .A2(n3223), .ZN(n3224) );
  OAI211_X1 U4020 ( .C1(n3226), .C2(n3520), .A(n3225), .B(n3224), .ZN(U3228)
         );
  AND2_X1 U4021 ( .A1(n3215), .A2(n3227), .ZN(n3230) );
  OAI211_X1 U4022 ( .C1(n3230), .C2(n3229), .A(n3496), .B(n3228), .ZN(n3233)
         );
  INV_X1 U4023 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4096) );
  NOR2_X1 U4024 ( .A1(STATE_REG_SCAN_IN), .A2(n4096), .ZN(n4295) );
  OAI22_X1 U4025 ( .A1(n3238), .A2(n3515), .B1(n3514), .B2(n3300), .ZN(n3231)
         );
  AOI211_X1 U4026 ( .C1(n3500), .C2(n3684), .A(n4295), .B(n3231), .ZN(n3232)
         );
  OAI211_X1 U4027 ( .C1(n3503), .C2(n4405), .A(n3233), .B(n3232), .ZN(U3214)
         );
  OAI21_X1 U4028 ( .B1(n3178), .B2(n3237), .A(n3234), .ZN(n4414) );
  NAND2_X1 U4029 ( .A1(n3566), .A2(n3560), .ZN(n3611) );
  XOR2_X1 U4030 ( .A(n3611), .B(n3235), .Z(n4416) );
  XOR2_X1 U4031 ( .A(n3611), .B(n3236), .Z(n3242) );
  OAI22_X1 U4032 ( .A1(n3238), .A2(n4447), .B1(n4389), .B2(n3237), .ZN(n3239)
         );
  AOI21_X1 U4033 ( .B1(n4394), .B2(n3240), .A(n3239), .ZN(n3241) );
  OAI21_X1 U4034 ( .B1(n3242), .B2(n4396), .A(n3241), .ZN(n3243) );
  AOI21_X1 U4035 ( .B1(n4445), .B2(n4416), .A(n3243), .ZN(n4419) );
  INV_X1 U4036 ( .A(n4419), .ZN(n3244) );
  AOI21_X1 U4037 ( .B1(n4538), .B2(n4416), .A(n3244), .ZN(n3246) );
  MUX2_X1 U4038 ( .A(n2413), .B(n3246), .S(n4558), .Z(n3245) );
  OAI21_X1 U4039 ( .B1(n4414), .B2(n4168), .A(n3245), .ZN(U3526) );
  INV_X1 U4040 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3247) );
  MUX2_X1 U4041 ( .A(n3247), .B(n3246), .S(n4544), .Z(n3248) );
  OAI21_X1 U4042 ( .B1(n4414), .B2(n4221), .A(n3248), .ZN(U3483) );
  NAND2_X1 U40430 ( .A1(n3250), .A2(n3249), .ZN(n3251) );
  XNOR2_X1 U4044 ( .A(n3252), .B(n3251), .ZN(n3253) );
  NAND2_X1 U4045 ( .A1(n3253), .A2(n3496), .ZN(n3258) );
  INV_X1 U4046 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3254) );
  NOR2_X1 U4047 ( .A1(STATE_REG_SCAN_IN), .A2(n3254), .ZN(n4306) );
  OAI22_X1 U4048 ( .A1(n3255), .A2(n3515), .B1(n3514), .B2(n4390), .ZN(n3256)
         );
  AOI211_X1 U4049 ( .C1(n3500), .C2(n3683), .A(n4306), .B(n3256), .ZN(n3257)
         );
  OAI211_X1 U4050 ( .C1(n3503), .C2(n3259), .A(n3258), .B(n3257), .ZN(U3233)
         );
  INV_X1 U4051 ( .A(n3327), .ZN(n3326) );
  XNOR2_X1 U4052 ( .A(n3326), .B(n3329), .ZN(n3261) );
  XNOR2_X1 U4053 ( .A(n3260), .B(n3261), .ZN(n3266) );
  INV_X1 U4054 ( .A(n3262), .ZN(n3275) );
  AOI22_X1 U4055 ( .A1(n3684), .A2(n3488), .B1(n3487), .B2(n3267), .ZN(n3263)
         );
  NAND2_X1 U4056 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4310) );
  OAI211_X1 U4057 ( .C1(n3345), .C2(n3512), .A(n3263), .B(n4310), .ZN(n3264)
         );
  AOI21_X1 U4058 ( .B1(n3275), .B2(n3518), .A(n3264), .ZN(n3265) );
  OAI21_X1 U4059 ( .B1(n3266), .B2(n3520), .A(n3265), .ZN(U3221) );
  XNOR2_X1 U4060 ( .A(n4391), .B(n3267), .ZN(n3629) );
  XNOR2_X1 U4061 ( .A(n3268), .B(n3629), .ZN(n3271) );
  OAI22_X1 U4062 ( .A1(n3345), .A2(n4447), .B1(n4389), .B2(n3273), .ZN(n3269)
         );
  AOI21_X1 U4063 ( .B1(n4394), .B2(n3684), .A(n3269), .ZN(n3270) );
  OAI21_X1 U4064 ( .B1(n3271), .B2(n4396), .A(n3270), .ZN(n3320) );
  INV_X1 U4065 ( .A(n3320), .ZN(n3279) );
  XOR2_X1 U4066 ( .A(n3629), .B(n3272), .Z(n3321) );
  OR2_X1 U4067 ( .A1(n4400), .A2(n3273), .ZN(n3274) );
  NAND2_X1 U4068 ( .A1(n3289), .A2(n3274), .ZN(n3325) );
  AOI22_X1 U4069 ( .A1(n4442), .A2(REG2_REG_12__SCAN_IN), .B1(n3275), .B2(
        n4434), .ZN(n3276) );
  OAI21_X1 U4070 ( .B1(n3325), .B2(n3968), .A(n3276), .ZN(n3277) );
  AOI21_X1 U4071 ( .B1(n3321), .B2(n3905), .A(n3277), .ZN(n3278) );
  OAI21_X1 U4072 ( .B1(n4442), .B2(n3279), .A(n3278), .ZN(U3278) );
  NAND2_X1 U4073 ( .A1(n3281), .A2(n3280), .ZN(n3283) );
  NAND2_X1 U4074 ( .A1(n3533), .A2(n3282), .ZN(n3610) );
  XNOR2_X1 U4075 ( .A(n3283), .B(n3610), .ZN(n3286) );
  AOI22_X1 U4076 ( .A1(n3681), .A2(n4423), .B1(n4422), .B2(n3288), .ZN(n3284)
         );
  OAI21_X1 U4077 ( .B1(n4391), .B2(n4426), .A(n3284), .ZN(n3285) );
  AOI21_X1 U4078 ( .B1(n3286), .B2(n4444), .A(n3285), .ZN(n4176) );
  XNOR2_X1 U4079 ( .A(n3287), .B(n3610), .ZN(n4175) );
  NAND2_X1 U4080 ( .A1(n3289), .A2(n3288), .ZN(n3290) );
  NAND2_X1 U4081 ( .A1(n3348), .A2(n3290), .ZN(n4178) );
  NOR2_X1 U4082 ( .A1(n4178), .A2(n3968), .ZN(n3293) );
  OAI22_X1 U4083 ( .A1(n4453), .A2(n3291), .B1(n3340), .B2(n4457), .ZN(n3292)
         );
  AOI211_X1 U4084 ( .C1(n4175), .C2(n3905), .A(n3293), .B(n3292), .ZN(n3294)
         );
  OAI21_X1 U4085 ( .B1(n4442), .B2(n4176), .A(n3294), .ZN(U3277) );
  INV_X1 U4086 ( .A(n3295), .ZN(n3297) );
  INV_X1 U4087 ( .A(n3296), .ZN(n4401) );
  OAI21_X1 U4088 ( .B1(n3297), .B2(n3300), .A(n4401), .ZN(n4407) );
  NAND2_X1 U4089 ( .A1(n3524), .A2(n3525), .ZN(n3609) );
  XOR2_X1 U4090 ( .A(n3609), .B(n3298), .Z(n4409) );
  XNOR2_X1 U4091 ( .A(n3299), .B(n3609), .ZN(n3304) );
  OAI22_X1 U4092 ( .A1(n3301), .A2(n4447), .B1(n4389), .B2(n3300), .ZN(n3302)
         );
  AOI21_X1 U4093 ( .B1(n4394), .B2(n3685), .A(n3302), .ZN(n3303) );
  OAI21_X1 U4094 ( .B1(n3304), .B2(n4396), .A(n3303), .ZN(n3305) );
  AOI21_X1 U4095 ( .B1(n4409), .B2(n4445), .A(n3305), .ZN(n4412) );
  INV_X1 U4096 ( .A(n4412), .ZN(n3306) );
  AOI21_X1 U4097 ( .B1(n4538), .B2(n4409), .A(n3306), .ZN(n3308) );
  MUX2_X1 U4098 ( .A(n2446), .B(n3308), .S(n4558), .Z(n3307) );
  OAI21_X1 U4099 ( .B1(n4407), .B2(n4168), .A(n3307), .ZN(U3528) );
  INV_X1 U4100 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4039) );
  MUX2_X1 U4101 ( .A(n4039), .B(n3308), .S(n4544), .Z(n3309) );
  OAI21_X1 U4102 ( .B1(n4407), .B2(n4221), .A(n3309), .ZN(U3487) );
  XOR2_X1 U4103 ( .A(n3311), .B(n3310), .Z(n3312) );
  XNOR2_X1 U4104 ( .A(n3313), .B(n3312), .ZN(n3319) );
  INV_X1 U4105 ( .A(n3349), .ZN(n3317) );
  AOI22_X1 U4106 ( .A1(n3488), .A2(n3682), .B1(n3487), .B2(n3347), .ZN(n3314)
         );
  NAND2_X1 U4107 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4328) );
  OAI211_X1 U4108 ( .C1(n3315), .C2(n3512), .A(n3314), .B(n4328), .ZN(n3316)
         );
  AOI21_X1 U4109 ( .B1(n3317), .B2(n3518), .A(n3316), .ZN(n3318) );
  OAI21_X1 U4110 ( .B1(n3319), .B2(n3520), .A(n3318), .ZN(U3212) );
  INV_X1 U4111 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4046) );
  AOI21_X1 U4112 ( .B1(n3321), .B2(n4534), .A(n3320), .ZN(n3323) );
  MUX2_X1 U4113 ( .A(n4046), .B(n3323), .S(n4544), .Z(n3322) );
  OAI21_X1 U4114 ( .B1(n3325), .B2(n4221), .A(n3322), .ZN(U3491) );
  MUX2_X1 U4115 ( .A(n2482), .B(n3323), .S(n4558), .Z(n3324) );
  OAI21_X1 U4116 ( .B1(n3325), .B2(n4168), .A(n3324), .ZN(U3530) );
  NOR2_X1 U4117 ( .A1(n3260), .A2(n3326), .ZN(n3330) );
  INV_X1 U4118 ( .A(n3260), .ZN(n3328) );
  OAI22_X1 U4119 ( .A1(n3330), .A2(n3329), .B1(n3328), .B2(n3327), .ZN(n3334)
         );
  NAND2_X1 U4120 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  XNOR2_X1 U4121 ( .A(n3334), .B(n3333), .ZN(n3335) );
  NAND2_X1 U4122 ( .A1(n3335), .A2(n3496), .ZN(n3339) );
  NOR2_X1 U4123 ( .A1(STATE_REG_SCAN_IN), .A2(n3336), .ZN(n4322) );
  OAI22_X1 U4124 ( .A1(n4391), .A2(n3515), .B1(n3514), .B2(n2136), .ZN(n3337)
         );
  AOI211_X1 U4125 ( .C1(n3500), .C2(n3681), .A(n4322), .B(n3337), .ZN(n3338)
         );
  OAI211_X1 U4126 ( .C1(n3503), .C2(n3340), .A(n3339), .B(n3338), .ZN(U3231)
         );
  XNOR2_X1 U4127 ( .A(n3341), .B(n3617), .ZN(n4169) );
  OAI21_X1 U4128 ( .B1(n3617), .B2(n3640), .A(n3354), .ZN(n3342) );
  NAND2_X1 U4129 ( .A1(n3342), .A2(n4444), .ZN(n3344) );
  AOI22_X1 U4130 ( .A1(n3680), .A2(n4423), .B1(n4422), .B2(n3347), .ZN(n3343)
         );
  OAI211_X1 U4131 ( .C1(n3345), .C2(n4426), .A(n3344), .B(n3343), .ZN(n3346)
         );
  AOI21_X1 U4132 ( .B1(n4169), .B2(n4445), .A(n3346), .ZN(n4173) );
  NAND2_X1 U4133 ( .A1(n3348), .A2(n3347), .ZN(n4170) );
  AND3_X1 U4134 ( .A1(n4171), .A2(n4438), .A3(n4170), .ZN(n3351) );
  OAI22_X1 U4135 ( .A1(n4453), .A2(n4331), .B1(n3349), .B2(n4457), .ZN(n3350)
         );
  AOI211_X1 U4136 ( .C1(n4169), .C2(n4443), .A(n3351), .B(n3350), .ZN(n3352)
         );
  OAI21_X1 U4137 ( .B1(n4173), .B2(n4442), .A(n3352), .ZN(U3276) );
  XNOR2_X1 U4138 ( .A(n3353), .B(n3625), .ZN(n3381) );
  INV_X1 U4139 ( .A(n3381), .ZN(n3365) );
  NAND2_X1 U4140 ( .A1(n3354), .A2(n3534), .ZN(n3355) );
  XNOR2_X1 U4141 ( .A(n3355), .B(n3625), .ZN(n3359) );
  OAI22_X1 U4142 ( .A1(n3467), .A2(n4447), .B1(n4389), .B2(n3356), .ZN(n3357)
         );
  AOI21_X1 U4143 ( .B1(n4394), .B2(n3681), .A(n3357), .ZN(n3358) );
  OAI21_X1 U4144 ( .B1(n3359), .B2(n4396), .A(n3358), .ZN(n3380) );
  AND2_X1 U4145 ( .A1(n4171), .A2(n3400), .ZN(n3360) );
  OR2_X1 U4146 ( .A1(n3360), .A2(n3373), .ZN(n3386) );
  INV_X1 U4147 ( .A(n3361), .ZN(n3403) );
  AOI22_X1 U4148 ( .A1(n4442), .A2(REG2_REG_15__SCAN_IN), .B1(n3403), .B2(
        n4434), .ZN(n3362) );
  OAI21_X1 U4149 ( .B1(n3386), .B2(n3968), .A(n3362), .ZN(n3363) );
  AOI21_X1 U4150 ( .B1(n3380), .B2(n4453), .A(n3363), .ZN(n3364) );
  OAI21_X1 U4151 ( .B1(n3365), .B2(n3974), .A(n3364), .ZN(U3275) );
  XNOR2_X1 U4152 ( .A(n3366), .B(n3368), .ZN(n4165) );
  INV_X1 U4153 ( .A(n4165), .ZN(n3379) );
  XNOR2_X1 U4154 ( .A(n3367), .B(n3368), .ZN(n3371) );
  OAI22_X1 U4155 ( .A1(n3949), .A2(n4447), .B1(n4389), .B2(n3372), .ZN(n3369)
         );
  AOI21_X1 U4156 ( .B1(n4394), .B2(n3680), .A(n3369), .ZN(n3370) );
  OAI21_X1 U4157 ( .B1(n3371), .B2(n4396), .A(n3370), .ZN(n4164) );
  OR2_X1 U4158 ( .A1(n3373), .A2(n3372), .ZN(n3374) );
  NAND2_X1 U4159 ( .A1(n3964), .A2(n3374), .ZN(n4222) );
  INV_X1 U4160 ( .A(n3375), .ZN(n3393) );
  AOI22_X1 U4161 ( .A1(n4442), .A2(REG2_REG_16__SCAN_IN), .B1(n3393), .B2(
        n4434), .ZN(n3376) );
  OAI21_X1 U4162 ( .B1(n4222), .B2(n3968), .A(n3376), .ZN(n3377) );
  AOI21_X1 U4163 ( .B1(n4164), .B2(n4453), .A(n3377), .ZN(n3378) );
  OAI21_X1 U4164 ( .B1(n3379), .B2(n3974), .A(n3378), .ZN(U3274) );
  INV_X1 U4165 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3382) );
  AOI21_X1 U4166 ( .B1(n3381), .B2(n4534), .A(n3380), .ZN(n3384) );
  MUX2_X1 U4167 ( .A(n3382), .B(n3384), .S(n4544), .Z(n3383) );
  OAI21_X1 U4168 ( .B1(n3386), .B2(n4221), .A(n3383), .ZN(U3497) );
  MUX2_X1 U4169 ( .A(n3704), .B(n3384), .S(n4558), .Z(n3385) );
  OAI21_X1 U4170 ( .B1(n4168), .B2(n3386), .A(n3385), .ZN(U3533) );
  AOI21_X1 U4171 ( .B1(n3398), .B2(n3396), .A(n3387), .ZN(n3389) );
  XNOR2_X1 U4172 ( .A(n3389), .B(n3388), .ZN(n3395) );
  AOI22_X1 U4173 ( .A1(n3488), .A2(n3680), .B1(n3487), .B2(n3390), .ZN(n3391)
         );
  NAND2_X1 U4174 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4359) );
  OAI211_X1 U4175 ( .C1(n3949), .C2(n3512), .A(n3391), .B(n4359), .ZN(n3392)
         );
  AOI21_X1 U4176 ( .B1(n3393), .B2(n3518), .A(n3392), .ZN(n3394) );
  OAI21_X1 U4177 ( .B1(n3395), .B2(n3520), .A(n3394), .ZN(U3223) );
  INV_X1 U4178 ( .A(n3387), .ZN(n3397) );
  NAND2_X1 U4179 ( .A1(n3397), .A2(n3396), .ZN(n3399) );
  XNOR2_X1 U4180 ( .A(n3399), .B(n3398), .ZN(n3405) );
  AOI22_X1 U4181 ( .A1(n3681), .A2(n3488), .B1(n3487), .B2(n3400), .ZN(n3401)
         );
  NAND2_X1 U4182 ( .A1(REG3_REG_15__SCAN_IN), .A2(U3149), .ZN(n4338) );
  OAI211_X1 U4183 ( .C1(n3467), .C2(n3512), .A(n3401), .B(n4338), .ZN(n3402)
         );
  AOI21_X1 U4184 ( .B1(n3403), .B2(n3518), .A(n3402), .ZN(n3404) );
  OAI21_X1 U4185 ( .B1(n3405), .B2(n3520), .A(n3404), .ZN(U3238) );
  AOI21_X1 U4186 ( .B1(n3408), .B2(n3407), .A(n3406), .ZN(n3413) );
  AOI22_X1 U4187 ( .A1(n3676), .A2(n3500), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3410) );
  INV_X1 U4188 ( .A(n3896), .ZN(n3678) );
  AOI22_X1 U4189 ( .A1(n3678), .A2(n3488), .B1(n3487), .B2(n3873), .ZN(n3409)
         );
  OAI211_X1 U4190 ( .C1(n3864), .C2(n3503), .A(n3410), .B(n3409), .ZN(n3411)
         );
  INV_X1 U4191 ( .A(n3411), .ZN(n3412) );
  OAI21_X1 U4192 ( .B1(n3413), .B2(n3520), .A(n3412), .ZN(U3232) );
  AOI22_X1 U4193 ( .A1(n4460), .A2(n3415), .B1(n3414), .B2(n2721), .ZN(U3458)
         );
  OAI22_X1 U4194 ( .A1(n4453), .A2(n3417), .B1(n3416), .B2(n4457), .ZN(n3420)
         );
  NOR2_X1 U4195 ( .A1(n3418), .A2(n4442), .ZN(n3419) );
  OAI21_X1 U4196 ( .B1(n3422), .B2(n3974), .A(n3421), .ZN(U3262) );
  NAND3_X1 U4197 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n2230), 
        .ZN(n3425) );
  INV_X1 U4198 ( .A(DATAI_31_), .ZN(n3424) );
  OAI22_X1 U4199 ( .A1(n3423), .A2(n3425), .B1(STATE_REG_SCAN_IN), .B2(n3424), 
        .ZN(U3321) );
  OAI21_X1 U4200 ( .B1(n3406), .B2(n3428), .A(n3427), .ZN(n3429) );
  NAND3_X1 U4201 ( .A1(n3430), .A2(n3496), .A3(n3429), .ZN(n3434) );
  NOR2_X1 U4202 ( .A1(n3512), .A2(n3807), .ZN(n3432) );
  OAI22_X1 U4203 ( .A1(n3880), .A2(n3515), .B1(n3514), .B2(n3853), .ZN(n3431)
         );
  AOI211_X1 U4204 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3432), .B(n3431), .ZN(n3433) );
  OAI211_X1 U4205 ( .C1(n3503), .C2(n3854), .A(n3434), .B(n3433), .ZN(U3213)
         );
  XNOR2_X1 U4206 ( .A(n3436), .B(n3435), .ZN(n3437) );
  NAND2_X1 U4207 ( .A1(n3437), .A2(n3496), .ZN(n3440) );
  NOR2_X1 U4208 ( .A1(n4083), .A2(STATE_REG_SCAN_IN), .ZN(n3734) );
  OAI22_X1 U4209 ( .A1(n3959), .A2(n3515), .B1(n3514), .B2(n3929), .ZN(n3438)
         );
  AOI211_X1 U4210 ( .C1(n3500), .C2(n3884), .A(n3734), .B(n3438), .ZN(n3439)
         );
  OAI211_X1 U4211 ( .C1(n3503), .C2(n3932), .A(n3440), .B(n3439), .ZN(U3216)
         );
  XNOR2_X1 U4212 ( .A(n3442), .B(n3441), .ZN(n3443) );
  XNOR2_X1 U4213 ( .A(n3444), .B(n3443), .ZN(n3450) );
  INV_X1 U4214 ( .A(n3890), .ZN(n3448) );
  OAI22_X1 U4215 ( .A1(n3512), .A2(n3880), .B1(STATE_REG_SCAN_IN), .B2(n3445), 
        .ZN(n3447) );
  OAI22_X1 U4216 ( .A1(n3924), .A2(n3515), .B1(n3514), .B2(n3888), .ZN(n3446)
         );
  AOI211_X1 U4217 ( .C1(n3448), .C2(n3518), .A(n3447), .B(n3446), .ZN(n3449)
         );
  OAI21_X1 U4218 ( .B1(n3450), .B2(n3520), .A(n3449), .ZN(U3220) );
  INV_X1 U4219 ( .A(n3452), .ZN(n3453) );
  NOR2_X1 U4220 ( .A1(n3454), .A2(n3453), .ZN(n3455) );
  XNOR2_X1 U4221 ( .A(n3451), .B(n3455), .ZN(n3462) );
  INV_X1 U4222 ( .A(n3815), .ZN(n3460) );
  OAI22_X1 U4223 ( .A1(n3512), .A2(n3779), .B1(STATE_REG_SCAN_IN), .B2(n3456), 
        .ZN(n3459) );
  OAI22_X1 U4224 ( .A1(n3807), .A2(n3515), .B1(n3514), .B2(n3457), .ZN(n3458)
         );
  AOI211_X1 U4225 ( .C1(n3460), .C2(n3518), .A(n3459), .B(n3458), .ZN(n3461)
         );
  OAI21_X1 U4226 ( .B1(n3462), .B2(n3520), .A(n3461), .ZN(U3222) );
  XNOR2_X1 U4227 ( .A(n3464), .B(n2214), .ZN(n3465) );
  XNOR2_X1 U4228 ( .A(n3463), .B(n3465), .ZN(n3466) );
  NAND2_X1 U4229 ( .A1(n3466), .A2(n3496), .ZN(n3470) );
  AND2_X1 U4230 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4367) );
  OAI22_X1 U4231 ( .A1(n3467), .A2(n3515), .B1(n3514), .B2(n3966), .ZN(n3468)
         );
  AOI211_X1 U4232 ( .C1(n3500), .C2(n3926), .A(n4367), .B(n3468), .ZN(n3469)
         );
  OAI211_X1 U4233 ( .C1(n3969), .C2(n3503), .A(n3470), .B(n3469), .ZN(U3225)
         );
  NAND2_X1 U4234 ( .A1(n2017), .A2(n3471), .ZN(n3472) );
  XOR2_X1 U4235 ( .A(n3473), .B(n3472), .Z(n3478) );
  AOI22_X1 U4236 ( .A1(n3789), .A2(n3500), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3476) );
  AOI22_X1 U4237 ( .A1(n3676), .A2(n3488), .B1(n3487), .B2(n3474), .ZN(n3475)
         );
  OAI211_X1 U4238 ( .C1(n3833), .C2(n3503), .A(n3476), .B(n3475), .ZN(n3477)
         );
  AOI21_X1 U4239 ( .B1(n3478), .B2(n3496), .A(n3477), .ZN(n3479) );
  INV_X1 U4240 ( .A(n3479), .ZN(U3226) );
  INV_X1 U4241 ( .A(n3480), .ZN(n3485) );
  AOI21_X1 U4242 ( .B1(n3484), .B2(n3482), .A(n3481), .ZN(n3483) );
  AOI21_X1 U4243 ( .B1(n3485), .B2(n3484), .A(n3483), .ZN(n3493) );
  AOI22_X1 U4244 ( .A1(n3678), .A2(n3500), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3490) );
  AOI22_X1 U4245 ( .A1(n3488), .A2(n3947), .B1(n3487), .B2(n3486), .ZN(n3489)
         );
  OAI211_X1 U4246 ( .C1(n3908), .C2(n3503), .A(n3490), .B(n3489), .ZN(n3491)
         );
  INV_X1 U4247 ( .A(n3491), .ZN(n3492) );
  OAI21_X1 U4248 ( .B1(n3493), .B2(n3520), .A(n3492), .ZN(U3230) );
  NOR2_X1 U4249 ( .A1(n3494), .A2(n2048), .ZN(n3495) );
  XNOR2_X1 U4250 ( .A(n2039), .B(n3495), .ZN(n3497) );
  NAND2_X1 U4251 ( .A1(n3497), .A2(n3496), .ZN(n3502) );
  AND2_X1 U4252 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4377) );
  OAI22_X1 U4253 ( .A1(n3949), .A2(n3515), .B1(n3514), .B2(n3498), .ZN(n3499)
         );
  AOI211_X1 U4254 ( .C1(n3500), .C2(n3947), .A(n4377), .B(n3499), .ZN(n3501)
         );
  OAI211_X1 U4255 ( .C1(n3503), .C2(n3942), .A(n3502), .B(n3501), .ZN(U3235)
         );
  INV_X1 U4256 ( .A(n3505), .ZN(n3507) );
  NAND2_X1 U4257 ( .A1(n3507), .A2(n3506), .ZN(n3508) );
  XNOR2_X1 U4258 ( .A(n3504), .B(n3508), .ZN(n3521) );
  INV_X1 U4259 ( .A(n3509), .ZN(n3796) );
  OAI22_X1 U4260 ( .A1(n3512), .A2(n3511), .B1(STATE_REG_SCAN_IN), .B2(n3510), 
        .ZN(n3517) );
  OAI22_X1 U4261 ( .A1(n3824), .A2(n3515), .B1(n3514), .B2(n3513), .ZN(n3516)
         );
  AOI211_X1 U4262 ( .C1(n3796), .C2(n3518), .A(n3517), .B(n3516), .ZN(n3519)
         );
  OAI21_X1 U4263 ( .B1(n3521), .B2(n3520), .A(n3519), .ZN(U3237) );
  INV_X1 U4264 ( .A(n3532), .ZN(n3638) );
  AND2_X1 U4265 ( .A1(n3523), .A2(n3522), .ZN(n3564) );
  NOR2_X1 U4266 ( .A1(n3638), .A2(n3564), .ZN(n3642) );
  INV_X1 U4267 ( .A(n3524), .ZN(n3537) );
  AND2_X1 U4268 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  AND2_X1 U4269 ( .A1(n3529), .A2(n3527), .ZN(n3569) );
  INV_X1 U4270 ( .A(n3528), .ZN(n3531) );
  OAI21_X1 U4271 ( .B1(n3531), .B2(n3530), .A(n3529), .ZN(n3535) );
  NAND4_X1 U4272 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3536)
         );
  AOI21_X1 U4273 ( .B1(n3537), .B2(n3569), .A(n3536), .ZN(n3573) );
  NAND2_X1 U4274 ( .A1(n2840), .A2(n4450), .ZN(n3622) );
  OAI211_X1 U4275 ( .C1(n2842), .C2(n2742), .A(n3622), .B(n3538), .ZN(n3540)
         );
  NAND3_X1 U4276 ( .A1(n3540), .A2(n3539), .A3(n2843), .ZN(n3542) );
  OAI211_X1 U4277 ( .C1(n3544), .C2(n3543), .A(n3542), .B(n3541), .ZN(n3547)
         );
  NAND3_X1 U4278 ( .A1(n3547), .A2(n3546), .A3(n3545), .ZN(n3550) );
  NAND4_X1 U4279 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3554), .ZN(n3553)
         );
  INV_X1 U4280 ( .A(n3621), .ZN(n3552) );
  NAND3_X1 U4281 ( .A1(n3553), .A2(n3552), .A3(n3551), .ZN(n3558) );
  INV_X1 U4282 ( .A(n3554), .ZN(n3556) );
  NOR3_X1 U4283 ( .A1(n3642), .A2(n3556), .A3(n3555), .ZN(n3557) );
  AOI21_X1 U4284 ( .B1(n3558), .B2(n3564), .A(n3557), .ZN(n3563) );
  INV_X1 U4285 ( .A(n3559), .ZN(n3562) );
  INV_X1 U4286 ( .A(n3560), .ZN(n3561) );
  NOR3_X1 U4287 ( .A1(n3563), .A2(n3562), .A3(n3561), .ZN(n3571) );
  INV_X1 U4288 ( .A(n3564), .ZN(n3565) );
  AOI21_X1 U4289 ( .B1(n3567), .B2(n3566), .A(n3565), .ZN(n3570) );
  OAI211_X1 U4290 ( .C1(n3571), .C2(n3570), .A(n3569), .B(n3568), .ZN(n3572)
         );
  OAI21_X1 U4291 ( .B1(n3642), .B2(n3573), .A(n3572), .ZN(n3574) );
  NAND2_X1 U4292 ( .A1(n3645), .A2(n3574), .ZN(n3575) );
  AOI211_X1 U4293 ( .C1(n3641), .C2(n3575), .A(n3650), .B(n3644), .ZN(n3577)
         );
  NOR2_X1 U4294 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  OAI21_X1 U4295 ( .B1(n3842), .B2(n3578), .A(n3647), .ZN(n3579) );
  AOI211_X1 U4296 ( .C1(n3580), .C2(n3579), .A(n3653), .B(n3636), .ZN(n3584)
         );
  NAND2_X1 U4297 ( .A1(n3586), .A2(DATAI_29_), .ZN(n3759) );
  AND2_X1 U4298 ( .A1(n3675), .A2(n3759), .ZN(n3581) );
  NOR2_X1 U4299 ( .A1(n3742), .A2(n3581), .ZN(n3634) );
  INV_X1 U4300 ( .A(n3634), .ZN(n3582) );
  OR4_X1 U4301 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3592) );
  OR2_X1 U4302 ( .A1(n3743), .A2(n3637), .ZN(n3587) );
  AND2_X1 U4303 ( .A1(n3586), .A2(DATAI_30_), .ZN(n3987) );
  NAND2_X1 U4304 ( .A1(n3748), .A2(n3987), .ZN(n3599) );
  NAND2_X1 U4305 ( .A1(n3586), .A2(DATAI_31_), .ZN(n3977) );
  AND2_X1 U4306 ( .A1(n3588), .A2(n3977), .ZN(n3598) );
  INV_X1 U4307 ( .A(n3598), .ZN(n3591) );
  OAI211_X1 U4308 ( .C1(n3675), .C2(n3759), .A(n3599), .B(n3591), .ZN(n3635)
         );
  AOI21_X1 U4309 ( .B1(n3587), .B2(n3634), .A(n3635), .ZN(n3657) );
  NOR2_X1 U4310 ( .A1(n3748), .A2(n3987), .ZN(n3661) );
  INV_X1 U4311 ( .A(n3661), .ZN(n3602) );
  NOR2_X1 U4312 ( .A1(n3588), .A2(n3977), .ZN(n3660) );
  INV_X1 U4313 ( .A(n3660), .ZN(n3589) );
  NAND2_X1 U4314 ( .A1(n3602), .A2(n3589), .ZN(n3590) );
  AOI22_X1 U4315 ( .A1(n3592), .A2(n3657), .B1(n3591), .B2(n3590), .ZN(n3666)
         );
  INV_X1 U4316 ( .A(n3593), .ZN(n3595) );
  NOR2_X1 U4317 ( .A1(n3595), .A2(n3594), .ZN(n3903) );
  INV_X1 U4318 ( .A(n3841), .ZN(n3596) );
  OR2_X1 U4319 ( .A1(n3842), .A2(n3596), .ZN(n3886) );
  XNOR2_X1 U4320 ( .A(n3947), .B(n3929), .ZN(n3923) );
  NAND2_X1 U4321 ( .A1(n3916), .A2(n3917), .ZN(n3958) );
  NOR4_X1 U4322 ( .A1(n3903), .A2(n3886), .A3(n3923), .A4(n3958), .ZN(n3601)
         );
  NAND2_X1 U4323 ( .A1(n3597), .A2(n3784), .ZN(n3810) );
  NOR3_X1 U4324 ( .A1(n3810), .A2(n3598), .A3(n3660), .ZN(n3600) );
  NAND4_X1 U4325 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3605)
         );
  NOR3_X1 U4326 ( .A1(n3605), .A2(n3604), .A3(n3603), .ZN(n3616) );
  INV_X1 U4327 ( .A(n3606), .ZN(n3821) );
  OR2_X1 U4328 ( .A1(n3821), .A2(n3607), .ZN(n3845) );
  NAND2_X1 U4329 ( .A1(n3608), .A2(n3802), .ZN(n3829) );
  NOR4_X1 U4330 ( .A1(n3845), .A2(n3610), .A3(n3609), .A4(n3829), .ZN(n3615)
         );
  NOR4_X1 U4331 ( .A1(n3613), .A2(n3612), .A3(n3945), .A4(n3611), .ZN(n3614)
         );
  NAND3_X1 U4332 ( .A1(n3616), .A2(n3615), .A3(n3614), .ZN(n3632) );
  INV_X1 U4333 ( .A(n3617), .ZN(n3618) );
  NOR4_X1 U4334 ( .A1(n3618), .A2(n2844), .A3(n2828), .A4(n2841), .ZN(n3628)
         );
  XNOR2_X1 U4335 ( .A(n3675), .B(n3759), .ZN(n3756) );
  NOR4_X1 U4336 ( .A1(n4387), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3627)
         );
  NAND2_X1 U4337 ( .A1(n3623), .A2(n3622), .ZN(n4494) );
  NAND2_X1 U4338 ( .A1(n3624), .A2(n3633), .ZN(n3786) );
  NOR4_X1 U4339 ( .A1(n3752), .A2(n3625), .A3(n4494), .A4(n3786), .ZN(n3626)
         );
  NAND4_X1 U4340 ( .A1(n3628), .A2(n3757), .A3(n3627), .A4(n3626), .ZN(n3631)
         );
  NOR4_X1 U4341 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3663)
         );
  INV_X1 U4342 ( .A(n3977), .ZN(n3980) );
  NAND3_X1 U4343 ( .A1(n3772), .A2(n3634), .A3(n3633), .ZN(n3656) );
  NOR4_X1 U4344 ( .A1(n3743), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3655)
         );
  NOR3_X1 U4345 ( .A1(n3640), .A2(n3639), .A3(n3638), .ZN(n3643) );
  OAI21_X1 U4346 ( .B1(n3643), .B2(n3642), .A(n3641), .ZN(n3646) );
  NAND3_X1 U4347 ( .A1(n3646), .A2(n2856), .A3(n3645), .ZN(n3648) );
  OAI221_X1 U4348 ( .B1(n3650), .B2(n3649), .C1(n3650), .C2(n3648), .A(n3647), 
        .ZN(n3651) );
  OAI221_X1 U4349 ( .B1(n3653), .B2(n3652), .C1(n3653), .C2(n3651), .A(n3783), 
        .ZN(n3654) );
  AOI22_X1 U4350 ( .A1(n3657), .A2(n3656), .B1(n3655), .B2(n3654), .ZN(n3658)
         );
  AOI21_X1 U4351 ( .B1(n3987), .B2(n3979), .A(n3658), .ZN(n3659) );
  AOI211_X1 U4352 ( .C1(n3980), .C2(n3661), .A(n3660), .B(n3659), .ZN(n3662)
         );
  MUX2_X1 U4353 ( .A(n3663), .B(n3662), .S(n2742), .Z(n3665) );
  MUX2_X1 U4354 ( .A(n3666), .B(n3665), .S(n3664), .Z(n3667) );
  XNOR2_X1 U4355 ( .A(n3667), .B(n4229), .ZN(n3674) );
  NOR2_X1 U4356 ( .A1(n3669), .A2(n3668), .ZN(n3672) );
  OAI21_X1 U4357 ( .B1(n3673), .B2(n3670), .A(B_REG_SCAN_IN), .ZN(n3671) );
  OAI22_X1 U4358 ( .A1(n3674), .A2(n3673), .B1(n3672), .B2(n3671), .ZN(U3239)
         );
  MUX2_X1 U4359 ( .A(n3675), .B(DATAO_REG_29__SCAN_IN), .S(n3689), .Z(U3579)
         );
  MUX2_X1 U4360 ( .A(n3776), .B(DATAO_REG_28__SCAN_IN), .S(n3689), .Z(U3578)
         );
  MUX2_X1 U4361 ( .A(n3788), .B(DATAO_REG_27__SCAN_IN), .S(n3689), .Z(U3577)
         );
  MUX2_X1 U4362 ( .A(n3805), .B(DATAO_REG_26__SCAN_IN), .S(n3689), .Z(U3576)
         );
  MUX2_X1 U4363 ( .A(DATAO_REG_25__SCAN_IN), .B(n3789), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4364 ( .A(n3848), .B(DATAO_REG_24__SCAN_IN), .S(n3689), .Z(U3574)
         );
  MUX2_X1 U4365 ( .A(DATAO_REG_23__SCAN_IN), .B(n3676), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4366 ( .A(DATAO_REG_22__SCAN_IN), .B(n3677), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4367 ( .A(DATAO_REG_21__SCAN_IN), .B(n3678), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4368 ( .A(n3884), .B(DATAO_REG_20__SCAN_IN), .S(n3689), .Z(U3570)
         );
  MUX2_X1 U4369 ( .A(n3947), .B(DATAO_REG_19__SCAN_IN), .S(n3689), .Z(U3569)
         );
  MUX2_X1 U4370 ( .A(DATAO_REG_18__SCAN_IN), .B(n3926), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4371 ( .A(DATAO_REG_17__SCAN_IN), .B(n3679), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4372 ( .A(DATAO_REG_16__SCAN_IN), .B(n3961), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4373 ( .A(n3680), .B(DATAO_REG_15__SCAN_IN), .S(n3689), .Z(U3565)
         );
  MUX2_X1 U4374 ( .A(DATAO_REG_14__SCAN_IN), .B(n3681), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4375 ( .A(n3682), .B(DATAO_REG_13__SCAN_IN), .S(n3689), .Z(U3563)
         );
  MUX2_X1 U4376 ( .A(DATAO_REG_12__SCAN_IN), .B(n3683), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4377 ( .A(DATAO_REG_11__SCAN_IN), .B(n3684), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4378 ( .A(n4393), .B(DATAO_REG_10__SCAN_IN), .S(n3689), .Z(U3560)
         );
  MUX2_X1 U4379 ( .A(n3685), .B(DATAO_REG_9__SCAN_IN), .S(n3689), .Z(U3559) );
  MUX2_X1 U4380 ( .A(n3686), .B(DATAO_REG_8__SCAN_IN), .S(n3689), .Z(U3558) );
  MUX2_X1 U4381 ( .A(n3687), .B(DATAO_REG_6__SCAN_IN), .S(n3689), .Z(U3556) );
  MUX2_X1 U4382 ( .A(n3688), .B(DATAO_REG_5__SCAN_IN), .S(n3689), .Z(U3555) );
  MUX2_X1 U4383 ( .A(n3690), .B(DATAO_REG_3__SCAN_IN), .S(n3689), .Z(U3553) );
  MUX2_X1 U4384 ( .A(DATAO_REG_2__SCAN_IN), .B(n4424), .S(U4043), .Z(U3552) );
  MUX2_X1 U4385 ( .A(DATAO_REG_1__SCAN_IN), .B(n2790), .S(U4043), .Z(U3551) );
  INV_X1 U4386 ( .A(n3731), .ZN(n4467) );
  INV_X1 U4387 ( .A(n4472), .ZN(n4348) );
  AOI22_X1 U4388 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4472), .B1(n4348), .B2(
        n3704), .ZN(n4345) );
  INV_X1 U4389 ( .A(n3724), .ZN(n4477) );
  AOI22_X1 U4390 ( .A1(n3724), .A2(REG1_REG_13__SCAN_IN), .B1(n3700), .B2(
        n4477), .ZN(n4325) );
  AOI22_X1 U4391 ( .A1(n3710), .A2(REG1_REG_11__SCAN_IN), .B1(n2466), .B2(
        n4480), .ZN(n4299) );
  NAND2_X1 U4392 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4482), .ZN(n3694) );
  INV_X1 U4393 ( .A(n4482), .ZN(n4283) );
  AOI22_X1 U4394 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4482), .B1(n4283), .B2(n2430), .ZN(n4277) );
  NAND2_X1 U4395 ( .A1(n4272), .A2(REG1_REG_8__SCAN_IN), .ZN(n4271) );
  NAND2_X1 U4396 ( .A1(n4265), .A2(n3692), .ZN(n3693) );
  NAND2_X1 U4397 ( .A1(n4287), .A2(n3695), .ZN(n3696) );
  NAND2_X1 U4398 ( .A1(n3696), .A2(n4288), .ZN(n4298) );
  NAND2_X1 U4399 ( .A1(n4299), .A2(n4298), .ZN(n4297) );
  NAND2_X1 U4400 ( .A1(n3710), .A2(REG1_REG_11__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U4401 ( .A1(n3722), .A2(n3698), .ZN(n3699) );
  NAND2_X1 U4402 ( .A1(n3699), .A2(n4313), .ZN(n4324) );
  NAND2_X1 U4403 ( .A1(n4325), .A2(n4324), .ZN(n4323) );
  NAND2_X1 U4404 ( .A1(n3701), .A2(n3702), .ZN(n3703) );
  INV_X1 U4405 ( .A(n3701), .ZN(n4475) );
  NOR2_X1 U4406 ( .A1(n4470), .A2(n3705), .ZN(n3706) );
  INV_X1 U4407 ( .A(n4470), .ZN(n4353) );
  INV_X1 U4408 ( .A(n3730), .ZN(n4469) );
  AOI22_X1 U4409 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4469), .B1(n3730), .B2(
        n4162), .ZN(n4368) );
  AOI22_X1 U4410 ( .A1(n3731), .A2(REG1_REG_18__SCAN_IN), .B1(n3707), .B2(
        n4467), .ZN(n4382) );
  OAI21_X1 U4411 ( .B1(n3707), .B2(n4467), .A(n4379), .ZN(n3709) );
  XNOR2_X1 U4412 ( .A(n3736), .B(REG1_REG_19__SCAN_IN), .ZN(n3708) );
  XNOR2_X1 U4413 ( .A(n3709), .B(n3708), .ZN(n3740) );
  AOI22_X1 U4414 ( .A1(n3731), .A2(n3943), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4467), .ZN(n4375) );
  AOI22_X1 U4415 ( .A1(REG2_REG_17__SCAN_IN), .A2(n3730), .B1(n4469), .B2(
        n3970), .ZN(n4365) );
  INV_X1 U4416 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4417 ( .A1(n3710), .A2(REG2_REG_11__SCAN_IN), .B1(n3719), .B2(
        n4480), .ZN(n4302) );
  AOI22_X1 U4418 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4482), .B1(n4283), .B2(n2433), .ZN(n4280) );
  NAND2_X1 U4419 ( .A1(n4265), .A2(n3713), .ZN(n3714) );
  NAND2_X1 U4420 ( .A1(n4280), .A2(n4279), .ZN(n4278) );
  NAND2_X1 U4421 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4482), .ZN(n3715) );
  NAND2_X1 U4422 ( .A1(n4287), .A2(n3717), .ZN(n3718) );
  NAND2_X1 U4423 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4291), .ZN(n4290) );
  NAND2_X1 U4424 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4309), .ZN(n4308) );
  NAND2_X1 U4425 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  NOR2_X1 U4426 ( .A1(n4477), .A2(n3291), .ZN(n4317) );
  NOR2_X1 U4427 ( .A1(n4475), .A2(n3725), .ZN(n3726) );
  INV_X1 U4428 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4331) );
  NAND2_X1 U4429 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4472), .ZN(n3727) );
  OAI21_X1 U4430 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4472), .A(n3727), .ZN(n4340) );
  AOI21_X1 U4431 ( .B1(n4472), .B2(REG2_REG_15__SCAN_IN), .A(n4339), .ZN(n3728) );
  NAND2_X1 U4432 ( .A1(n3728), .A2(n4353), .ZN(n3729) );
  XNOR2_X1 U4433 ( .A(n4470), .B(n3728), .ZN(n4350) );
  NOR2_X1 U4434 ( .A1(n4373), .A2(n2213), .ZN(n3733) );
  MUX2_X1 U4435 ( .A(n3933), .B(REG2_REG_19__SCAN_IN), .S(n3736), .Z(n3732) );
  XNOR2_X1 U4436 ( .A(n3733), .B(n3732), .ZN(n3738) );
  AOI21_X1 U4437 ( .B1(n4378), .B2(ADDR_REG_19__SCAN_IN), .A(n3734), .ZN(n3735) );
  OAI21_X1 U4438 ( .B1(n3736), .B2(n4385), .A(n3735), .ZN(n3737) );
  AOI21_X1 U4439 ( .B1(n3738), .B2(n4358), .A(n3737), .ZN(n3739) );
  OAI21_X1 U4440 ( .B1(n3740), .B2(n4354), .A(n3739), .ZN(U3259) );
  INV_X1 U4441 ( .A(n3741), .ZN(n3751) );
  INV_X1 U4442 ( .A(n3742), .ZN(n3744) );
  INV_X1 U4443 ( .A(B_REG_SCAN_IN), .ZN(n3746) );
  OAI21_X1 U4444 ( .B1(n3747), .B2(n3746), .A(n4423), .ZN(n3978) );
  OAI22_X1 U4445 ( .A1(n3748), .A2(n3978), .B1(n4389), .B2(n3759), .ZN(n3749)
         );
  AOI21_X1 U4446 ( .B1(n4394), .B2(n3776), .A(n3749), .ZN(n3750) );
  AOI21_X1 U4447 ( .B1(n3751), .B2(n4434), .A(n3993), .ZN(n3764) );
  XNOR2_X1 U4448 ( .A(n3758), .B(n3757), .ZN(n3990) );
  NAND2_X1 U4449 ( .A1(n3990), .A2(n3905), .ZN(n3763) );
  INV_X1 U4450 ( .A(n3759), .ZN(n3761) );
  AOI21_X1 U4451 ( .B1(n3761), .B2(n3760), .A(n3982), .ZN(n3991) );
  AOI22_X1 U4452 ( .A1(n3991), .A2(n4438), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4442), .ZN(n3762) );
  OAI211_X1 U4453 ( .C1(n4442), .C2(n3764), .A(n3763), .B(n3762), .ZN(U3354)
         );
  XNOR2_X1 U4454 ( .A(n3765), .B(n3772), .ZN(n3998) );
  AND2_X1 U4455 ( .A1(n3795), .A2(n3775), .ZN(n3766) );
  NOR2_X1 U4456 ( .A1(n3767), .A2(n3766), .ZN(n3996) );
  OAI22_X1 U4457 ( .A1(n4453), .A2(n3769), .B1(n3768), .B2(n4457), .ZN(n3770)
         );
  AOI21_X1 U4458 ( .B1(n3996), .B2(n4438), .A(n3770), .ZN(n3781) );
  OAI21_X1 U4459 ( .B1(n3773), .B2(n3772), .A(n3771), .ZN(n3774) );
  NAND2_X1 U4460 ( .A1(n3774), .A2(n4444), .ZN(n3778) );
  AOI22_X1 U4461 ( .A1(n3776), .A2(n4423), .B1(n3775), .B2(n4422), .ZN(n3777)
         );
  OAI211_X1 U4462 ( .C1(n3779), .C2(n4426), .A(n3778), .B(n3777), .ZN(n3995)
         );
  NAND2_X1 U4463 ( .A1(n3995), .A2(n4453), .ZN(n3780) );
  OAI211_X1 U4464 ( .C1(n3998), .C2(n3974), .A(n3781), .B(n3780), .ZN(U3263)
         );
  XOR2_X1 U4465 ( .A(n3786), .B(n3782), .Z(n4000) );
  INV_X1 U4466 ( .A(n4000), .ZN(n3800) );
  INV_X1 U4467 ( .A(n3783), .ZN(n3785) );
  OAI21_X1 U4468 ( .B1(n3801), .B2(n3785), .A(n3784), .ZN(n3787) );
  XNOR2_X1 U4469 ( .A(n3787), .B(n3786), .ZN(n3792) );
  AOI22_X1 U4470 ( .A1(n3788), .A2(n4423), .B1(n3793), .B2(n4422), .ZN(n3791)
         );
  NAND2_X1 U4471 ( .A1(n3789), .A2(n4394), .ZN(n3790) );
  OAI211_X1 U4472 ( .C1(n3792), .C2(n4396), .A(n3791), .B(n3790), .ZN(n3999)
         );
  NAND2_X1 U4473 ( .A1(n3814), .A2(n3793), .ZN(n3794) );
  NAND2_X1 U4474 ( .A1(n3795), .A2(n3794), .ZN(n4190) );
  AOI22_X1 U4475 ( .A1(n4442), .A2(REG2_REG_26__SCAN_IN), .B1(n3796), .B2(
        n4434), .ZN(n3797) );
  OAI21_X1 U4476 ( .B1(n4190), .B2(n3968), .A(n3797), .ZN(n3798) );
  AOI21_X1 U4477 ( .B1(n3999), .B2(n4453), .A(n3798), .ZN(n3799) );
  OAI21_X1 U4478 ( .B1(n3800), .B2(n3974), .A(n3799), .ZN(U3264) );
  INV_X1 U4479 ( .A(n3801), .ZN(n3803) );
  NAND2_X1 U4480 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  XNOR2_X1 U4481 ( .A(n3804), .B(n3810), .ZN(n3809) );
  AOI22_X1 U4482 ( .A1(n3805), .A2(n4423), .B1(n4422), .B2(n3812), .ZN(n3806)
         );
  OAI21_X1 U4483 ( .B1(n3807), .B2(n4426), .A(n3806), .ZN(n3808) );
  AOI21_X1 U4484 ( .B1(n3809), .B2(n4444), .A(n3808), .ZN(n4003) );
  XNOR2_X1 U4485 ( .A(n3811), .B(n3810), .ZN(n4002) );
  NAND2_X1 U4486 ( .A1(n4002), .A2(n3905), .ZN(n3820) );
  NAND2_X1 U4487 ( .A1(n3831), .A2(n3812), .ZN(n3813) );
  NAND2_X1 U4488 ( .A1(n3814), .A2(n3813), .ZN(n4005) );
  INV_X1 U4489 ( .A(n4005), .ZN(n3818) );
  OAI22_X1 U4490 ( .A1(n4453), .A2(n3816), .B1(n3815), .B2(n4457), .ZN(n3817)
         );
  AOI21_X1 U4491 ( .B1(n3818), .B2(n4438), .A(n3817), .ZN(n3819) );
  OAI211_X1 U4492 ( .C1(n4442), .C2(n4003), .A(n3820), .B(n3819), .ZN(U3265)
         );
  NOR2_X1 U4493 ( .A1(n3822), .A2(n3821), .ZN(n3823) );
  XNOR2_X1 U4494 ( .A(n3823), .B(n3829), .ZN(n3827) );
  NOR2_X1 U4495 ( .A1(n3872), .A2(n4426), .ZN(n3826) );
  OAI22_X1 U4496 ( .A1(n3824), .A2(n4447), .B1(n4389), .B2(n3832), .ZN(n3825)
         );
  AOI211_X1 U4497 ( .C1(n3827), .C2(n4444), .A(n3826), .B(n3825), .ZN(n4130)
         );
  XNOR2_X1 U4498 ( .A(n3830), .B(n3829), .ZN(n4132) );
  NAND2_X1 U4499 ( .A1(n4132), .A2(n3905), .ZN(n3838) );
  OAI21_X1 U4500 ( .B1(n3851), .B2(n3832), .A(n3831), .ZN(n4195) );
  INV_X1 U4501 ( .A(n4195), .ZN(n3836) );
  OAI22_X1 U4502 ( .A1(n4453), .A2(n3834), .B1(n3833), .B2(n4457), .ZN(n3835)
         );
  AOI21_X1 U4503 ( .B1(n3836), .B2(n4438), .A(n3835), .ZN(n3837) );
  OAI211_X1 U4504 ( .C1(n4442), .C2(n4130), .A(n3838), .B(n3837), .ZN(U3266)
         );
  OR2_X1 U4505 ( .A1(n3860), .A2(n3868), .ZN(n3861) );
  NAND2_X1 U4506 ( .A1(n3861), .A2(n3839), .ZN(n3840) );
  XOR2_X1 U4507 ( .A(n3845), .B(n3840), .Z(n4136) );
  INV_X1 U4508 ( .A(n4136), .ZN(n3859) );
  OAI21_X1 U4509 ( .B1(n2025), .B2(n3842), .A(n3841), .ZN(n3869) );
  NAND2_X1 U4510 ( .A1(n3869), .A2(n3868), .ZN(n3871) );
  NAND2_X1 U4511 ( .A1(n3871), .A2(n3843), .ZN(n3844) );
  XOR2_X1 U4512 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND2_X1 U4513 ( .A1(n3846), .A2(n4444), .ZN(n3850) );
  AOI22_X1 U4514 ( .A1(n3848), .A2(n4423), .B1(n3847), .B2(n4422), .ZN(n3849)
         );
  OAI211_X1 U4515 ( .C1(n3880), .C2(n4426), .A(n3850), .B(n3849), .ZN(n4135)
         );
  INV_X1 U4516 ( .A(n3851), .ZN(n3852) );
  OAI21_X1 U4517 ( .B1(n3863), .B2(n3853), .A(n3852), .ZN(n4199) );
  NOR2_X1 U4518 ( .A1(n4199), .A2(n3968), .ZN(n3857) );
  OAI22_X1 U4519 ( .A1(n4453), .A2(n3855), .B1(n3854), .B2(n4457), .ZN(n3856)
         );
  AOI211_X1 U4520 ( .C1(n4135), .C2(n4453), .A(n3857), .B(n3856), .ZN(n3858)
         );
  OAI21_X1 U4521 ( .B1(n3859), .B2(n3974), .A(n3858), .ZN(U3267) );
  INV_X1 U4522 ( .A(n3860), .ZN(n3862) );
  OAI21_X1 U4523 ( .B1(n3862), .B2(n2828), .A(n3861), .ZN(n4142) );
  NAND2_X1 U4524 ( .A1(n3887), .A2(n3873), .ZN(n4139) );
  AND2_X1 U4525 ( .A1(n4139), .A2(n4438), .ZN(n3867) );
  OAI22_X1 U4526 ( .A1(n4453), .A2(n3865), .B1(n3864), .B2(n4457), .ZN(n3866)
         );
  AOI21_X1 U4527 ( .B1(n2132), .B2(n3867), .A(n3866), .ZN(n3879) );
  OR2_X1 U4528 ( .A1(n3869), .A2(n3868), .ZN(n3870) );
  NAND2_X1 U4529 ( .A1(n3871), .A2(n3870), .ZN(n3877) );
  OR2_X1 U4530 ( .A1(n3872), .A2(n4447), .ZN(n3875) );
  NAND2_X1 U4531 ( .A1(n3873), .A2(n4422), .ZN(n3874) );
  OAI211_X1 U4532 ( .C1(n3896), .C2(n4426), .A(n3875), .B(n3874), .ZN(n3876)
         );
  AOI21_X1 U4533 ( .B1(n3877), .B2(n4444), .A(n3876), .ZN(n4141) );
  OR2_X1 U4534 ( .A1(n4141), .A2(n4442), .ZN(n3878) );
  OAI211_X1 U4535 ( .C1(n4142), .C2(n3974), .A(n3879), .B(n3878), .ZN(U3268)
         );
  OAI22_X1 U4536 ( .A1(n3880), .A2(n4447), .B1(n4389), .B2(n3888), .ZN(n3883)
         );
  XOR2_X1 U4537 ( .A(n3886), .B(n2025), .Z(n3881) );
  NOR2_X1 U4538 ( .A1(n3881), .A2(n4396), .ZN(n3882) );
  AOI211_X1 U4539 ( .C1(n4394), .C2(n3884), .A(n3883), .B(n3882), .ZN(n4143)
         );
  XOR2_X1 U4540 ( .A(n3886), .B(n3885), .Z(n4145) );
  NAND2_X1 U4541 ( .A1(n4145), .A2(n3905), .ZN(n3895) );
  INV_X1 U4542 ( .A(n3906), .ZN(n3889) );
  OAI21_X1 U4543 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(n4204) );
  INV_X1 U4544 ( .A(n4204), .ZN(n3893) );
  OAI22_X1 U4545 ( .A1(n4453), .A2(n3891), .B1(n3890), .B2(n4457), .ZN(n3892)
         );
  AOI21_X1 U4546 ( .B1(n3893), .B2(n4438), .A(n3892), .ZN(n3894) );
  OAI211_X1 U4547 ( .C1(n4442), .C2(n4143), .A(n3895), .B(n3894), .ZN(U3269)
         );
  OAI22_X1 U4548 ( .A1(n3896), .A2(n4447), .B1(n4389), .B2(n3907), .ZN(n3902)
         );
  NAND2_X1 U4549 ( .A1(n3898), .A2(n3897), .ZN(n3899) );
  XNOR2_X1 U4550 ( .A(n3899), .B(n3903), .ZN(n3900) );
  NOR2_X1 U4551 ( .A1(n3900), .A2(n4396), .ZN(n3901) );
  AOI211_X1 U4552 ( .C1(n4394), .C2(n3947), .A(n3902), .B(n3901), .ZN(n4148)
         );
  XNOR2_X1 U4553 ( .A(n3904), .B(n3903), .ZN(n4150) );
  NAND2_X1 U4554 ( .A1(n4150), .A2(n3905), .ZN(n3913) );
  OAI21_X1 U4555 ( .B1(n3931), .B2(n3907), .A(n3906), .ZN(n4208) );
  INV_X1 U4556 ( .A(n4208), .ZN(n3911) );
  OAI22_X1 U4557 ( .A1(n4453), .A2(n3909), .B1(n3908), .B2(n4457), .ZN(n3910)
         );
  AOI21_X1 U4558 ( .B1(n3911), .B2(n4438), .A(n3910), .ZN(n3912) );
  OAI211_X1 U4559 ( .C1(n4442), .C2(n4148), .A(n3913), .B(n3912), .ZN(U3270)
         );
  XOR2_X1 U4560 ( .A(n3923), .B(n3914), .Z(n4154) );
  INV_X1 U4561 ( .A(n4154), .ZN(n3937) );
  INV_X1 U4562 ( .A(n3916), .ZN(n3918) );
  OAI21_X1 U4563 ( .B1(n3915), .B2(n3918), .A(n3917), .ZN(n3944) );
  INV_X1 U4564 ( .A(n3919), .ZN(n3921) );
  OAI21_X1 U4565 ( .B1(n3944), .B2(n3921), .A(n3920), .ZN(n3922) );
  XOR2_X1 U4566 ( .A(n3923), .B(n3922), .Z(n3928) );
  OAI22_X1 U4567 ( .A1(n3924), .A2(n4447), .B1(n4389), .B2(n3929), .ZN(n3925)
         );
  AOI21_X1 U4568 ( .B1(n4394), .B2(n3926), .A(n3925), .ZN(n3927) );
  OAI21_X1 U4569 ( .B1(n3928), .B2(n4396), .A(n3927), .ZN(n4153) );
  NOR2_X1 U4570 ( .A1(n3940), .A2(n3929), .ZN(n3930) );
  OR2_X1 U4571 ( .A1(n3931), .A2(n3930), .ZN(n4212) );
  NOR2_X1 U4572 ( .A1(n4212), .A2(n3968), .ZN(n3935) );
  OAI22_X1 U4573 ( .A1(n4453), .A2(n3933), .B1(n3932), .B2(n4457), .ZN(n3934)
         );
  AOI211_X1 U4574 ( .C1(n4153), .C2(n4453), .A(n3935), .B(n3934), .ZN(n3936)
         );
  OAI21_X1 U4575 ( .B1(n3937), .B2(n3974), .A(n3936), .ZN(U3271) );
  XOR2_X1 U4576 ( .A(n3945), .B(n3938), .Z(n4159) );
  NAND2_X1 U4577 ( .A1(n3965), .A2(n3946), .ZN(n3939) );
  NAND2_X1 U4578 ( .A1(n3939), .A2(n4537), .ZN(n3941) );
  OR2_X1 U4579 ( .A1(n3941), .A2(n3940), .ZN(n4157) );
  INV_X1 U4580 ( .A(n4157), .ZN(n3955) );
  OAI22_X1 U4581 ( .A1(n4453), .A2(n3943), .B1(n3942), .B2(n4457), .ZN(n3953)
         );
  XOR2_X1 U4582 ( .A(n3945), .B(n3944), .Z(n3951) );
  AOI22_X1 U4583 ( .A1(n3947), .A2(n4423), .B1(n3946), .B2(n4422), .ZN(n3948)
         );
  OAI21_X1 U4584 ( .B1(n3949), .B2(n4426), .A(n3948), .ZN(n3950) );
  AOI21_X1 U4585 ( .B1(n3951), .B2(n4444), .A(n3950), .ZN(n4158) );
  NOR2_X1 U4586 ( .A1(n4158), .A2(n4442), .ZN(n3952) );
  AOI211_X1 U4587 ( .C1(n3955), .C2(n3954), .A(n3953), .B(n3952), .ZN(n3956)
         );
  OAI21_X1 U4588 ( .B1(n4159), .B2(n3974), .A(n3956), .ZN(U3272) );
  XNOR2_X1 U4589 ( .A(n3957), .B(n3958), .ZN(n4161) );
  INV_X1 U4590 ( .A(n4161), .ZN(n3975) );
  XOR2_X1 U4591 ( .A(n3958), .B(n3915), .Z(n3963) );
  OAI22_X1 U4592 ( .A1(n3959), .A2(n4447), .B1(n4389), .B2(n3966), .ZN(n3960)
         );
  AOI21_X1 U4593 ( .B1(n4394), .B2(n3961), .A(n3960), .ZN(n3962) );
  OAI21_X1 U4594 ( .B1(n3963), .B2(n4396), .A(n3962), .ZN(n4160) );
  INV_X1 U4595 ( .A(n3964), .ZN(n3967) );
  OAI21_X1 U4596 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n4217) );
  NOR2_X1 U4597 ( .A1(n4217), .A2(n3968), .ZN(n3972) );
  OAI22_X1 U4598 ( .A1(n4453), .A2(n3970), .B1(n3969), .B2(n4457), .ZN(n3971)
         );
  AOI211_X1 U4599 ( .C1(n4160), .C2(n4453), .A(n3972), .B(n3971), .ZN(n3973)
         );
  OAI21_X1 U4600 ( .B1(n3975), .B2(n3974), .A(n3973), .ZN(U3273) );
  INV_X1 U4601 ( .A(n3987), .ZN(n3976) );
  NAND2_X1 U4602 ( .A1(n3982), .A2(n3976), .ZN(n3983) );
  XNOR2_X1 U4603 ( .A(n3983), .B(n3977), .ZN(n4235) );
  INV_X1 U4604 ( .A(n4235), .ZN(n4181) );
  NOR2_X1 U4605 ( .A1(n3979), .A2(n3978), .ZN(n3986) );
  AOI21_X1 U4606 ( .B1(n3980), .B2(n4422), .A(n3986), .ZN(n4237) );
  MUX2_X1 U4607 ( .A(n2952), .B(n4237), .S(n4558), .Z(n3981) );
  OAI21_X1 U4608 ( .B1(n4181), .B2(n4168), .A(n3981), .ZN(U3549) );
  INV_X1 U4609 ( .A(n3982), .ZN(n3985) );
  INV_X1 U4610 ( .A(n3983), .ZN(n3984) );
  AOI21_X1 U4611 ( .B1(n3987), .B2(n3985), .A(n3984), .ZN(n4238) );
  INV_X1 U4612 ( .A(n4238), .ZN(n4184) );
  INV_X1 U4613 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3988) );
  AOI21_X1 U4614 ( .B1(n3987), .B2(n4422), .A(n3986), .ZN(n4240) );
  MUX2_X1 U4615 ( .A(n3988), .B(n4240), .S(n4558), .Z(n3989) );
  OAI21_X1 U4616 ( .B1(n4184), .B2(n4168), .A(n3989), .ZN(U3548) );
  NAND2_X1 U4617 ( .A1(n3990), .A2(n4534), .ZN(n3994) );
  MUX2_X1 U4618 ( .A(REG1_REG_29__SCAN_IN), .B(n4185), .S(n4558), .Z(U3547) );
  INV_X1 U4619 ( .A(n4534), .ZN(n4520) );
  AOI21_X1 U4620 ( .B1(n4537), .B2(n3996), .A(n3995), .ZN(n3997) );
  OAI21_X1 U4621 ( .B1(n3998), .B2(n4520), .A(n3997), .ZN(n4186) );
  MUX2_X1 U4622 ( .A(REG1_REG_27__SCAN_IN), .B(n4186), .S(n4558), .Z(U3545) );
  AOI21_X1 U4623 ( .B1(n4000), .B2(n4534), .A(n3999), .ZN(n4187) );
  MUX2_X1 U4624 ( .A(n4050), .B(n4187), .S(n4558), .Z(n4001) );
  OAI21_X1 U4625 ( .B1(n4168), .B2(n4190), .A(n4001), .ZN(U3544) );
  NAND2_X1 U4626 ( .A1(n4002), .A2(n4534), .ZN(n4004) );
  OAI211_X1 U4627 ( .C1(n3992), .C2(n4005), .A(n4004), .B(n4003), .ZN(n4191)
         );
  MUX2_X1 U4628 ( .A(REG1_REG_25__SCAN_IN), .B(n4191), .S(n4558), .Z(n4129) );
  XNOR2_X1 U4629 ( .A(keyinput21), .B(DATAO_REG_22__SCAN_IN), .ZN(n4009) );
  XNOR2_X1 U4630 ( .A(keyinput2), .B(DATAO_REG_25__SCAN_IN), .ZN(n4008) );
  XNOR2_X1 U4631 ( .A(keyinput58), .B(DATAO_REG_14__SCAN_IN), .ZN(n4007) );
  XNOR2_X1 U4632 ( .A(keyinput17), .B(DATAO_REG_10__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4633 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4070)
         );
  XNOR2_X1 U4634 ( .A(keyinput61), .B(ADDR_REG_1__SCAN_IN), .ZN(n4013) );
  XNOR2_X1 U4635 ( .A(keyinput24), .B(DATAO_REG_0__SCAN_IN), .ZN(n4012) );
  XNOR2_X1 U4636 ( .A(keyinput35), .B(ADDR_REG_6__SCAN_IN), .ZN(n4011) );
  XNOR2_X1 U4637 ( .A(keyinput33), .B(ADDR_REG_16__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4638 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4069)
         );
  OAI22_X1 U4639 ( .A1(n3103), .A2(keyinput28), .B1(n4015), .B2(keyinput11), 
        .ZN(n4014) );
  AOI221_X1 U4640 ( .B1(n3103), .B2(keyinput28), .C1(keyinput11), .C2(n4015), 
        .A(n4014), .ZN(n4023) );
  XOR2_X1 U4641 ( .A(keyinput59), .B(DATAO_REG_9__SCAN_IN), .Z(n4019) );
  XOR2_X1 U4642 ( .A(keyinput55), .B(DATAO_REG_8__SCAN_IN), .Z(n4018) );
  XOR2_X1 U4643 ( .A(keyinput39), .B(DATAO_REG_7__SCAN_IN), .Z(n4017) );
  XOR2_X1 U4644 ( .A(keyinput16), .B(DATAO_REG_4__SCAN_IN), .Z(n4016) );
  NOR4_X1 U4645 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4022)
         );
  XNOR2_X1 U4646 ( .A(D_REG_9__SCAN_IN), .B(keyinput60), .ZN(n4021) );
  XNOR2_X1 U4647 ( .A(keyinput49), .B(DATAO_REG_26__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4648 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4068)
         );
  XOR2_X1 U4649 ( .A(n2504), .B(keyinput34), .Z(n4028) );
  INV_X1 U4650 ( .A(IR_REG_22__SCAN_IN), .ZN(n4024) );
  XOR2_X1 U4651 ( .A(n4024), .B(keyinput20), .Z(n4027) );
  XNOR2_X1 U4652 ( .A(IR_REG_23__SCAN_IN), .B(keyinput40), .ZN(n4026) );
  XNOR2_X1 U4653 ( .A(IR_REG_21__SCAN_IN), .B(keyinput0), .ZN(n4025) );
  NAND4_X1 U4654 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4034)
         );
  XNOR2_X1 U4655 ( .A(IR_REG_10__SCAN_IN), .B(keyinput43), .ZN(n4032) );
  XNOR2_X1 U4656 ( .A(IR_REG_8__SCAN_IN), .B(keyinput63), .ZN(n4031) );
  XNOR2_X1 U4657 ( .A(IR_REG_17__SCAN_IN), .B(keyinput45), .ZN(n4030) );
  XNOR2_X1 U4658 ( .A(IR_REG_13__SCAN_IN), .B(keyinput18), .ZN(n4029) );
  NAND4_X1 U4659 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4033)
         );
  NOR2_X1 U4660 ( .A1(n4034), .A2(n4033), .ZN(n4066) );
  INV_X1 U4661 ( .A(D_REG_2__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U4662 ( .A1(n4462), .A2(keyinput3), .B1(keyinput30), .B2(n2230), 
        .ZN(n4035) );
  OAI221_X1 U4663 ( .B1(n4462), .B2(keyinput3), .C1(n2230), .C2(keyinput30), 
        .A(n4035), .ZN(n4043) );
  INV_X1 U4664 ( .A(D_REG_12__SCAN_IN), .ZN(n4459) );
  INV_X1 U4665 ( .A(D_REG_3__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U4666 ( .A1(n4459), .A2(keyinput1), .B1(n4461), .B2(keyinput5), 
        .ZN(n4036) );
  OAI221_X1 U4667 ( .B1(n4459), .B2(keyinput1), .C1(n4461), .C2(keyinput5), 
        .A(n4036), .ZN(n4042) );
  INV_X1 U4668 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4495) );
  INV_X1 U4669 ( .A(D_REG_31__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U4670 ( .A1(n4495), .A2(keyinput27), .B1(n4458), .B2(keyinput15), 
        .ZN(n4037) );
  OAI221_X1 U4671 ( .B1(n4495), .B2(keyinput27), .C1(n4458), .C2(keyinput15), 
        .A(n4037), .ZN(n4041) );
  INV_X1 U4672 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4508) );
  AOI22_X1 U4673 ( .A1(n4508), .A2(keyinput62), .B1(n4039), .B2(keyinput44), 
        .ZN(n4038) );
  OAI221_X1 U4674 ( .B1(n4508), .B2(keyinput62), .C1(n4039), .C2(keyinput44), 
        .A(n4038), .ZN(n4040) );
  NOR4_X1 U4675 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4065)
         );
  INV_X1 U4676 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4677 ( .A1(n4046), .A2(keyinput36), .B1(keyinput47), .B2(n4045), 
        .ZN(n4044) );
  OAI221_X1 U4678 ( .B1(n4046), .B2(keyinput36), .C1(n4045), .C2(keyinput47), 
        .A(n4044), .ZN(n4054) );
  INV_X1 U4679 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4210) );
  INV_X1 U4680 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U4681 ( .A1(n4210), .A2(keyinput50), .B1(n4193), .B2(keyinput26), 
        .ZN(n4047) );
  OAI221_X1 U4682 ( .B1(n4210), .B2(keyinput50), .C1(n4193), .C2(keyinput26), 
        .A(n4047), .ZN(n4053) );
  AOI22_X1 U4683 ( .A1(n2466), .A2(keyinput4), .B1(n4151), .B2(keyinput12), 
        .ZN(n4048) );
  OAI221_X1 U4684 ( .B1(n2466), .B2(keyinput4), .C1(n4151), .C2(keyinput12), 
        .A(n4048), .ZN(n4052) );
  AOI22_X1 U4685 ( .A1(n4050), .A2(keyinput22), .B1(keyinput53), .B2(n4146), 
        .ZN(n4049) );
  OAI221_X1 U4686 ( .B1(n4050), .B2(keyinput22), .C1(n4146), .C2(keyinput53), 
        .A(n4049), .ZN(n4051) );
  NOR4_X1 U4687 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4064)
         );
  AOI22_X1 U4688 ( .A1(n2277), .A2(keyinput38), .B1(keyinput7), .B2(n2952), 
        .ZN(n4055) );
  OAI221_X1 U4689 ( .B1(n2277), .B2(keyinput38), .C1(n2952), .C2(keyinput7), 
        .A(n4055), .ZN(n4062) );
  AOI22_X1 U4690 ( .A1(n3008), .A2(keyinput52), .B1(n3015), .B2(keyinput29), 
        .ZN(n4056) );
  OAI221_X1 U4691 ( .B1(n3008), .B2(keyinput52), .C1(n3015), .C2(keyinput29), 
        .A(n4056), .ZN(n4061) );
  AOI22_X1 U4692 ( .A1(n2418), .A2(keyinput14), .B1(n2447), .B2(keyinput42), 
        .ZN(n4057) );
  OAI221_X1 U4693 ( .B1(n2418), .B2(keyinput14), .C1(n2447), .C2(keyinput42), 
        .A(n4057), .ZN(n4060) );
  AOI22_X1 U4694 ( .A1(n3816), .A2(keyinput6), .B1(keyinput31), .B2(n3891), 
        .ZN(n4058) );
  OAI221_X1 U4695 ( .B1(n3816), .B2(keyinput6), .C1(n3891), .C2(keyinput31), 
        .A(n4058), .ZN(n4059) );
  NOR4_X1 U4696 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  NAND4_X1 U4697 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NOR4_X1 U4698 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4094)
         );
  INV_X1 U4699 ( .A(DATAI_28_), .ZN(n4233) );
  AOI22_X1 U4700 ( .A1(n4233), .A2(keyinput46), .B1(keyinput13), .B2(n4072), 
        .ZN(n4071) );
  OAI221_X1 U4701 ( .B1(n4233), .B2(keyinput46), .C1(n4072), .C2(keyinput13), 
        .A(n4071), .ZN(n4080) );
  INV_X1 U4702 ( .A(DATAI_13_), .ZN(n4476) );
  AOI22_X1 U4703 ( .A1(n4476), .A2(keyinput32), .B1(n2599), .B2(keyinput10), 
        .ZN(n4073) );
  OAI221_X1 U4704 ( .B1(n4476), .B2(keyinput32), .C1(n2599), .C2(keyinput10), 
        .A(n4073), .ZN(n4079) );
  INV_X1 U4705 ( .A(DATAI_5_), .ZN(n4488) );
  AOI22_X1 U4706 ( .A1(n4488), .A2(keyinput57), .B1(n2493), .B2(keyinput19), 
        .ZN(n4074) );
  OAI221_X1 U4707 ( .B1(n4488), .B2(keyinput57), .C1(n2493), .C2(keyinput19), 
        .A(n4074), .ZN(n4078) );
  INV_X1 U4708 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4709 ( .A1(n4076), .A2(keyinput23), .B1(n4095), .B2(keyinput25), 
        .ZN(n4075) );
  OAI221_X1 U4710 ( .B1(n4076), .B2(keyinput23), .C1(n4095), .C2(keyinput25), 
        .A(n4075), .ZN(n4077) );
  NOR4_X1 U4711 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4093)
         );
  AOI22_X1 U4712 ( .A1(n2276), .A2(keyinput54), .B1(n2237), .B2(keyinput51), 
        .ZN(n4081) );
  OAI221_X1 U4713 ( .B1(n2276), .B2(keyinput54), .C1(n2237), .C2(keyinput51), 
        .A(n4081), .ZN(n4091) );
  AOI22_X1 U4714 ( .A1(n4083), .A2(keyinput48), .B1(keyinput37), .B2(n4096), 
        .ZN(n4082) );
  OAI221_X1 U4715 ( .B1(n4083), .B2(keyinput48), .C1(n4096), .C2(keyinput37), 
        .A(n4082), .ZN(n4090) );
  AOI22_X1 U4716 ( .A1(n2015), .A2(keyinput8), .B1(n4108), .B2(keyinput56), 
        .ZN(n4084) );
  OAI221_X1 U4717 ( .B1(n2015), .B2(keyinput8), .C1(n4108), .C2(keyinput56), 
        .A(n4084), .ZN(n4089) );
  INV_X1 U4718 ( .A(IR_REG_6__SCAN_IN), .ZN(n4085) );
  XOR2_X1 U4719 ( .A(n4085), .B(keyinput41), .Z(n4087) );
  XNOR2_X1 U4720 ( .A(IR_REG_5__SCAN_IN), .B(keyinput9), .ZN(n4086) );
  NAND2_X1 U4721 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  NOR4_X1 U4722 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  NAND3_X1 U4723 ( .A1(n4094), .A2(n4093), .A3(n4092), .ZN(n4127) );
  NOR4_X1 U4724 ( .A1(REG0_REG_24__SCAN_IN), .A2(REG2_REG_25__SCAN_IN), .A3(
        n4095), .A4(n4151), .ZN(n4106) );
  NAND4_X1 U4725 ( .A1(IR_REG_30__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        REG3_REG_19__SCAN_IN), .A4(n4096), .ZN(n4099) );
  NAND4_X1 U4726 ( .A1(DATAI_20_), .A2(REG0_REG_19__SCAN_IN), .A3(DATAI_19_), 
        .A4(DATAI_13_), .ZN(n4098) );
  NAND3_X1 U4727 ( .A1(DATAI_12_), .A2(REG1_REG_11__SCAN_IN), .A3(
        REG2_REG_10__SCAN_IN), .ZN(n4097) );
  NOR4_X1 U4728 ( .A1(REG0_REG_10__SCAN_IN), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4105) );
  NOR4_X1 U4729 ( .A1(REG2_REG_8__SCAN_IN), .A2(DATAI_5_), .A3(
        REG0_REG_2__SCAN_IN), .A4(n3015), .ZN(n4104) );
  NAND4_X1 U4730 ( .A1(REG0_REG_0__SCAN_IN), .A2(REG3_REG_0__SCAN_IN), .A3(
        n3103), .A4(n2237), .ZN(n4102) );
  NAND4_X1 U4731 ( .A1(REG2_REG_3__SCAN_IN), .A2(REG0_REG_12__SCAN_IN), .A3(
        REG0_REG_13__SCAN_IN), .A4(n2277), .ZN(n4101) );
  NAND3_X1 U4732 ( .A1(DATAI_28_), .A2(REG1_REG_26__SCAN_IN), .A3(
        REG2_REG_21__SCAN_IN), .ZN(n4100) );
  NOR4_X1 U4733 ( .A1(REG1_REG_21__SCAN_IN), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4103) );
  NAND4_X1 U4734 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4117)
         );
  NAND4_X1 U4735 ( .A1(n2086), .A2(n2217), .A3(n4107), .A4(IR_REG_6__SCAN_IN), 
        .ZN(n4110) );
  NAND3_X1 U4736 ( .A1(n2223), .A2(IR_REG_13__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .ZN(n4109) );
  NOR4_X1 U4737 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n2015), .ZN(n4112)
         );
  NOR3_X1 U4738 ( .A1(DATAO_REG_14__SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        DATAO_REG_31__SCAN_IN), .ZN(n4111) );
  NAND2_X1 U4739 ( .A1(n4112), .A2(n4111), .ZN(n4116) );
  NOR4_X1 U4740 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(n4462), .ZN(n4113) );
  NAND4_X1 U4741 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .A3(n4114), .A4(n4113), .ZN(n4115) );
  NOR3_X1 U4742 ( .A1(n4117), .A2(n4116), .A3(n4115), .ZN(n4125) );
  NAND3_X1 U4743 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG1_REG_31__SCAN_IN), .A3(
        DATAO_REG_25__SCAN_IN), .ZN(n4123) );
  INV_X1 U4744 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4362) );
  NAND4_X1 U4745 ( .A1(ADDR_REG_1__SCAN_IN), .A2(ADDR_REG_6__SCAN_IN), .A3(
        n4118), .A4(n4362), .ZN(n4122) );
  NAND4_X1 U4746 ( .A1(DATAO_REG_8__SCAN_IN), .A2(DATAO_REG_9__SCAN_IN), .A3(
        n4120), .A4(n4119), .ZN(n4121) );
  NOR4_X1 U4747 ( .A1(DATAO_REG_22__SCAN_IN), .A2(n4123), .A3(n4122), .A4(
        n4121), .ZN(n4124) );
  NAND2_X1 U4748 ( .A1(n4125), .A2(n4124), .ZN(n4126) );
  XNOR2_X1 U4749 ( .A(n4127), .B(n4126), .ZN(n4128) );
  XNOR2_X1 U4750 ( .A(n4129), .B(n4128), .ZN(U3543) );
  INV_X1 U4751 ( .A(n4130), .ZN(n4131) );
  AOI21_X1 U4752 ( .B1(n4132), .B2(n4534), .A(n4131), .ZN(n4192) );
  MUX2_X1 U4753 ( .A(n4133), .B(n4192), .S(n4558), .Z(n4134) );
  OAI21_X1 U4754 ( .B1(n4168), .B2(n4195), .A(n4134), .ZN(U3542) );
  AOI21_X1 U4755 ( .B1(n4136), .B2(n4534), .A(n4135), .ZN(n4196) );
  MUX2_X1 U4756 ( .A(n4137), .B(n4196), .S(n4558), .Z(n4138) );
  OAI21_X1 U4757 ( .B1(n4168), .B2(n4199), .A(n4138), .ZN(U3541) );
  NAND3_X1 U4758 ( .A1(n2132), .A2(n4537), .A3(n4139), .ZN(n4140) );
  OAI211_X1 U4759 ( .C1(n4142), .C2(n4520), .A(n4141), .B(n4140), .ZN(n4200)
         );
  MUX2_X1 U4760 ( .A(REG1_REG_22__SCAN_IN), .B(n4200), .S(n4558), .Z(U3540) );
  INV_X1 U4761 ( .A(n4143), .ZN(n4144) );
  AOI21_X1 U4762 ( .B1(n4145), .B2(n4534), .A(n4144), .ZN(n4201) );
  MUX2_X1 U4763 ( .A(n4146), .B(n4201), .S(n4558), .Z(n4147) );
  OAI21_X1 U4764 ( .B1(n4168), .B2(n4204), .A(n4147), .ZN(U3539) );
  INV_X1 U4765 ( .A(n4148), .ZN(n4149) );
  AOI21_X1 U4766 ( .B1(n4150), .B2(n4534), .A(n4149), .ZN(n4205) );
  MUX2_X1 U4767 ( .A(n4151), .B(n4205), .S(n4558), .Z(n4152) );
  OAI21_X1 U4768 ( .B1(n4168), .B2(n4208), .A(n4152), .ZN(U3538) );
  AOI21_X1 U4769 ( .B1(n4154), .B2(n4534), .A(n4153), .ZN(n4209) );
  MUX2_X1 U4770 ( .A(n4155), .B(n4209), .S(n4558), .Z(n4156) );
  OAI21_X1 U4771 ( .B1(n4168), .B2(n4212), .A(n4156), .ZN(U3537) );
  OAI211_X1 U4772 ( .C1(n4159), .C2(n4520), .A(n4158), .B(n4157), .ZN(n4213)
         );
  MUX2_X1 U4773 ( .A(REG1_REG_18__SCAN_IN), .B(n4213), .S(n4558), .Z(U3536) );
  AOI21_X1 U4774 ( .B1(n4161), .B2(n4534), .A(n4160), .ZN(n4214) );
  MUX2_X1 U4775 ( .A(n4162), .B(n4214), .S(n4558), .Z(n4163) );
  OAI21_X1 U4776 ( .B1(n4168), .B2(n4217), .A(n4163), .ZN(U3535) );
  AOI21_X1 U4777 ( .B1(n4165), .B2(n4534), .A(n4164), .ZN(n4218) );
  MUX2_X1 U4778 ( .A(n4166), .B(n4218), .S(n4558), .Z(n4167) );
  OAI21_X1 U4779 ( .B1(n4168), .B2(n4222), .A(n4167), .ZN(U3534) );
  INV_X1 U4780 ( .A(n4169), .ZN(n4174) );
  NAND3_X1 U4781 ( .A1(n4171), .A2(n4537), .A3(n4170), .ZN(n4172) );
  OAI211_X1 U4782 ( .C1(n4174), .C2(n4498), .A(n4173), .B(n4172), .ZN(n4223)
         );
  MUX2_X1 U4783 ( .A(REG1_REG_14__SCAN_IN), .B(n4223), .S(n4558), .Z(U3532) );
  NAND2_X1 U4784 ( .A1(n4175), .A2(n4534), .ZN(n4177) );
  OAI211_X1 U4785 ( .C1(n3992), .C2(n4178), .A(n4177), .B(n4176), .ZN(n4224)
         );
  MUX2_X1 U4786 ( .A(REG1_REG_13__SCAN_IN), .B(n4224), .S(n4558), .Z(U3531) );
  INV_X1 U4787 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4179) );
  MUX2_X1 U4788 ( .A(n4179), .B(n4237), .S(n4544), .Z(n4180) );
  OAI21_X1 U4789 ( .B1(n4181), .B2(n4221), .A(n4180), .ZN(U3517) );
  INV_X1 U4790 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4182) );
  MUX2_X1 U4791 ( .A(n4182), .B(n4240), .S(n4544), .Z(n4183) );
  OAI21_X1 U4792 ( .B1(n4184), .B2(n4221), .A(n4183), .ZN(U3516) );
  MUX2_X1 U4793 ( .A(REG0_REG_29__SCAN_IN), .B(n4185), .S(n4544), .Z(U3515) );
  MUX2_X1 U4794 ( .A(REG0_REG_27__SCAN_IN), .B(n4186), .S(n4544), .Z(U3513) );
  INV_X1 U4795 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4188) );
  MUX2_X1 U4796 ( .A(n4188), .B(n4187), .S(n4544), .Z(n4189) );
  OAI21_X1 U4797 ( .B1(n4190), .B2(n4221), .A(n4189), .ZN(U3512) );
  MUX2_X1 U4798 ( .A(REG0_REG_25__SCAN_IN), .B(n4191), .S(n4544), .Z(U3511) );
  MUX2_X1 U4799 ( .A(n4193), .B(n4192), .S(n4544), .Z(n4194) );
  OAI21_X1 U4800 ( .B1(n4195), .B2(n4221), .A(n4194), .ZN(U3510) );
  INV_X1 U4801 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4197) );
  MUX2_X1 U4802 ( .A(n4197), .B(n4196), .S(n4544), .Z(n4198) );
  OAI21_X1 U4803 ( .B1(n4199), .B2(n4221), .A(n4198), .ZN(U3509) );
  MUX2_X1 U4804 ( .A(REG0_REG_22__SCAN_IN), .B(n4200), .S(n4544), .Z(U3508) );
  INV_X1 U4805 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4202) );
  MUX2_X1 U4806 ( .A(n4202), .B(n4201), .S(n4544), .Z(n4203) );
  OAI21_X1 U4807 ( .B1(n4204), .B2(n4221), .A(n4203), .ZN(U3507) );
  INV_X1 U4808 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4206) );
  MUX2_X1 U4809 ( .A(n4206), .B(n4205), .S(n4544), .Z(n4207) );
  OAI21_X1 U4810 ( .B1(n4208), .B2(n4221), .A(n4207), .ZN(U3506) );
  MUX2_X1 U4811 ( .A(n4210), .B(n4209), .S(n4544), .Z(n4211) );
  OAI21_X1 U4812 ( .B1(n4212), .B2(n4221), .A(n4211), .ZN(U3505) );
  MUX2_X1 U4813 ( .A(REG0_REG_18__SCAN_IN), .B(n4213), .S(n4544), .Z(U3503) );
  INV_X1 U4814 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4215) );
  MUX2_X1 U4815 ( .A(n4215), .B(n4214), .S(n4544), .Z(n4216) );
  OAI21_X1 U4816 ( .B1(n4217), .B2(n4221), .A(n4216), .ZN(U3501) );
  INV_X1 U4817 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4219) );
  MUX2_X1 U4818 ( .A(n4219), .B(n4218), .S(n4544), .Z(n4220) );
  OAI21_X1 U4819 ( .B1(n4222), .B2(n4221), .A(n4220), .ZN(U3499) );
  MUX2_X1 U4820 ( .A(REG0_REG_14__SCAN_IN), .B(n4223), .S(n4544), .Z(U3495) );
  MUX2_X1 U4821 ( .A(REG0_REG_13__SCAN_IN), .B(n4224), .S(n4544), .Z(U3493) );
  MUX2_X1 U4822 ( .A(DATAI_30_), .B(n4225), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4823 ( .A(DATAI_29_), .B(n4226), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4824 ( .A(DATAI_27_), .B(n4242), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4825 ( .A(DATAI_25_), .B(n4227), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  INV_X1 U4826 ( .A(n2721), .ZN(n4228) );
  MUX2_X1 U4827 ( .A(n4228), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4828 ( .A(n4229), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4829 ( .A(n4230), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4830 ( .A(DATAI_4_), .B(n4231), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4831 ( .A(n4232), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U4832 ( .A1(STATE_REG_SCAN_IN), .A2(n4234), .B1(n4233), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4833 ( .A1(n4235), .A2(n4438), .B1(n4442), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4236) );
  OAI21_X1 U4834 ( .B1(n4442), .B2(n4237), .A(n4236), .ZN(U3260) );
  AOI22_X1 U4835 ( .A1(n4238), .A2(n4438), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4442), .ZN(n4239) );
  OAI21_X1 U4836 ( .B1(n4442), .B2(n4240), .A(n4239), .ZN(U3261) );
  OAI21_X1 U4837 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4242), .A(n4241), .ZN(n4243)
         );
  XOR2_X1 U4838 ( .A(n4243), .B(IR_REG_0__SCAN_IN), .Z(n4246) );
  AOI22_X1 U4839 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4378), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4244) );
  OAI21_X1 U4840 ( .B1(n4246), .B2(n4245), .A(n4244), .ZN(U3240) );
  AOI211_X1 U4841 ( .C1(n2053), .C2(n4248), .A(n4247), .B(n4354), .ZN(n4250)
         );
  AOI211_X1 U4842 ( .C1(n4378), .C2(ADDR_REG_5__SCAN_IN), .A(n4250), .B(n4249), 
        .ZN(n4255) );
  OAI211_X1 U4843 ( .C1(n4253), .C2(n4252), .A(n4358), .B(n4251), .ZN(n4254)
         );
  OAI211_X1 U4844 ( .C1(n4385), .C2(n4489), .A(n4255), .B(n4254), .ZN(U3245)
         );
  AOI211_X1 U4845 ( .C1(n2374), .C2(n4257), .A(n4256), .B(n4354), .ZN(n4258)
         );
  AOI211_X1 U4846 ( .C1(n4378), .C2(ADDR_REG_6__SCAN_IN), .A(n4259), .B(n4258), 
        .ZN(n4263) );
  OAI211_X1 U4847 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4261), .A(n4358), .B(n4260), 
        .ZN(n4262) );
  OAI211_X1 U4848 ( .C1(n4385), .C2(n4264), .A(n4263), .B(n4262), .ZN(U3246)
         );
  INV_X1 U4849 ( .A(n4265), .ZN(n4485) );
  OAI211_X1 U4850 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4267), .A(n4358), .B(n4266), 
        .ZN(n4269) );
  NAND2_X1 U4851 ( .A1(n4269), .A2(n4268), .ZN(n4270) );
  AOI21_X1 U4852 ( .B1(n4378), .B2(ADDR_REG_8__SCAN_IN), .A(n4270), .ZN(n4274)
         );
  OAI211_X1 U4853 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4272), .A(n4380), .B(n4271), 
        .ZN(n4273) );
  OAI211_X1 U4854 ( .C1(n4385), .C2(n4485), .A(n4274), .B(n4273), .ZN(U3248)
         );
  OAI211_X1 U4855 ( .C1(n4277), .C2(n4276), .A(n4380), .B(n4275), .ZN(n4282)
         );
  OAI211_X1 U4856 ( .C1(n4280), .C2(n4279), .A(n4358), .B(n4278), .ZN(n4281)
         );
  OAI211_X1 U4857 ( .C1(n4385), .C2(n4283), .A(n4282), .B(n4281), .ZN(n4284)
         );
  AOI211_X1 U4858 ( .C1(n4378), .C2(ADDR_REG_9__SCAN_IN), .A(n4285), .B(n4284), 
        .ZN(n4286) );
  INV_X1 U4859 ( .A(n4286), .ZN(U3249) );
  OAI211_X1 U4860 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4289), .A(n4380), .B(n4288), .ZN(n4293) );
  OAI211_X1 U4861 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4291), .A(n4358), .B(n4290), .ZN(n4292) );
  OAI211_X1 U4862 ( .C1(n4385), .C2(n3716), .A(n4293), .B(n4292), .ZN(n4294)
         );
  AOI211_X1 U4863 ( .C1(n4378), .C2(ADDR_REG_10__SCAN_IN), .A(n4295), .B(n4294), .ZN(n4296) );
  INV_X1 U4864 ( .A(n4296), .ZN(U3250) );
  OAI211_X1 U4865 ( .C1(n4299), .C2(n4298), .A(n4380), .B(n4297), .ZN(n4304)
         );
  OAI211_X1 U4866 ( .C1(n4302), .C2(n4301), .A(n4358), .B(n4300), .ZN(n4303)
         );
  OAI211_X1 U4867 ( .C1(n4385), .C2(n4480), .A(n4304), .B(n4303), .ZN(n4305)
         );
  AOI211_X1 U4868 ( .C1(n4378), .C2(ADDR_REG_11__SCAN_IN), .A(n4306), .B(n4305), .ZN(n4307) );
  INV_X1 U4869 ( .A(n4307), .ZN(U3251) );
  OAI211_X1 U4870 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4309), .A(n4358), .B(n4308), .ZN(n4311) );
  NAND2_X1 U4871 ( .A1(n4311), .A2(n4310), .ZN(n4312) );
  AOI21_X1 U4872 ( .B1(n4378), .B2(ADDR_REG_12__SCAN_IN), .A(n4312), .ZN(n4316) );
  OAI211_X1 U4873 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4314), .A(n4380), .B(n4313), .ZN(n4315) );
  OAI211_X1 U4874 ( .C1(n4385), .C2(n4478), .A(n4316), .B(n4315), .ZN(U3252)
         );
  AOI21_X1 U4875 ( .B1(n4477), .B2(n3291), .A(n4317), .ZN(n4320) );
  OAI21_X1 U4876 ( .B1(n4320), .B2(n4319), .A(n4358), .ZN(n4318) );
  AOI21_X1 U4877 ( .B1(n4320), .B2(n4319), .A(n4318), .ZN(n4321) );
  AOI211_X1 U4878 ( .C1(n4378), .C2(ADDR_REG_13__SCAN_IN), .A(n4322), .B(n4321), .ZN(n4327) );
  OAI211_X1 U4879 ( .C1(n4325), .C2(n4324), .A(n4380), .B(n4323), .ZN(n4326)
         );
  OAI211_X1 U4880 ( .C1(n4385), .C2(n4477), .A(n4327), .B(n4326), .ZN(U3253)
         );
  INV_X1 U4881 ( .A(n4328), .ZN(n4333) );
  INV_X1 U4882 ( .A(n4358), .ZN(n4372) );
  AOI211_X1 U4883 ( .C1(n4331), .C2(n4330), .A(n4329), .B(n4372), .ZN(n4332)
         );
  AOI211_X1 U4884 ( .C1(n4378), .C2(ADDR_REG_14__SCAN_IN), .A(n4333), .B(n4332), .ZN(n4337) );
  OAI211_X1 U4885 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4335), .A(n4380), .B(n4334), .ZN(n4336) );
  OAI211_X1 U4886 ( .C1(n4385), .C2(n4475), .A(n4337), .B(n4336), .ZN(U3254)
         );
  INV_X1 U4887 ( .A(n4338), .ZN(n4342) );
  AOI211_X1 U4888 ( .C1(n2041), .C2(n4340), .A(n4339), .B(n4372), .ZN(n4341)
         );
  AOI211_X1 U4889 ( .C1(n4378), .C2(ADDR_REG_15__SCAN_IN), .A(n4342), .B(n4341), .ZN(n4347) );
  OAI211_X1 U4890 ( .C1(n4345), .C2(n4344), .A(n4380), .B(n4343), .ZN(n4346)
         );
  OAI211_X1 U4891 ( .C1(n4385), .C2(n4348), .A(n4347), .B(n4346), .ZN(U3255)
         );
  INV_X1 U4892 ( .A(n4378), .ZN(n4361) );
  OAI21_X1 U4893 ( .B1(n4350), .B2(n2553), .A(n4349), .ZN(n4357) );
  AOI21_X1 U4894 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4352), .A(n4351), .ZN(n4355) );
  OAI22_X1 U4895 ( .A1(n4355), .A2(n4354), .B1(n4353), .B2(n4385), .ZN(n4356)
         );
  AOI21_X1 U4896 ( .B1(n4358), .B2(n4357), .A(n4356), .ZN(n4360) );
  OAI211_X1 U4897 ( .C1(n4362), .C2(n4361), .A(n4360), .B(n4359), .ZN(U3256)
         );
  AOI221_X1 U4898 ( .B1(n4365), .B2(n4364), .C1(n4363), .C2(n4364), .A(n4372), 
        .ZN(n4366) );
  AOI211_X1 U4899 ( .C1(n4378), .C2(ADDR_REG_17__SCAN_IN), .A(n4367), .B(n4366), .ZN(n4371) );
  OAI221_X1 U4900 ( .B1(n4369), .B2(n2034), .C1(n4369), .C2(n4368), .A(n4380), 
        .ZN(n4370) );
  OAI211_X1 U4901 ( .C1(n4385), .C2(n4469), .A(n4371), .B(n4370), .ZN(U3257)
         );
  AOI211_X1 U4902 ( .C1(n4375), .C2(n4374), .A(n4373), .B(n4372), .ZN(n4376)
         );
  AOI211_X1 U4903 ( .C1(n4378), .C2(ADDR_REG_18__SCAN_IN), .A(n4377), .B(n4376), .ZN(n4384) );
  OAI211_X1 U4904 ( .C1(n4382), .C2(n4381), .A(n4380), .B(n4379), .ZN(n4383)
         );
  XNOR2_X1 U4905 ( .A(n4386), .B(n4387), .ZN(n4539) );
  XNOR2_X1 U4906 ( .A(n4388), .B(n4387), .ZN(n4397) );
  OAI22_X1 U4907 ( .A1(n4391), .A2(n4447), .B1(n4390), .B2(n4389), .ZN(n4392)
         );
  AOI21_X1 U4908 ( .B1(n4394), .B2(n4393), .A(n4392), .ZN(n4395) );
  OAI21_X1 U4909 ( .B1(n4397), .B2(n4396), .A(n4395), .ZN(n4398) );
  AOI21_X1 U4910 ( .B1(n4445), .B2(n4539), .A(n4398), .ZN(n4541) );
  AOI22_X1 U4911 ( .A1(n4399), .A2(n4434), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4442), .ZN(n4404) );
  AOI21_X1 U4912 ( .B1(n4402), .B2(n4401), .A(n4400), .ZN(n4536) );
  AOI22_X1 U4913 ( .A1(n4539), .A2(n4443), .B1(n4438), .B2(n4536), .ZN(n4403)
         );
  OAI211_X1 U4914 ( .C1(n4442), .C2(n4541), .A(n4404), .B(n4403), .ZN(U3279)
         );
  OAI22_X1 U4915 ( .A1(n4405), .A2(n4457), .B1(n2447), .B2(n4453), .ZN(n4406)
         );
  INV_X1 U4916 ( .A(n4406), .ZN(n4411) );
  INV_X1 U4917 ( .A(n4407), .ZN(n4408) );
  AOI22_X1 U4918 ( .A1(n4409), .A2(n4443), .B1(n4438), .B2(n4408), .ZN(n4410)
         );
  OAI211_X1 U4919 ( .C1(n4442), .C2(n4412), .A(n4411), .B(n4410), .ZN(U3280)
         );
  AOI22_X1 U4920 ( .A1(n4413), .A2(n4434), .B1(REG2_REG_8__SCAN_IN), .B2(n4442), .ZN(n4418) );
  INV_X1 U4921 ( .A(n4414), .ZN(n4415) );
  AOI22_X1 U4922 ( .A1(n4416), .A2(n4443), .B1(n4438), .B2(n4415), .ZN(n4417)
         );
  OAI211_X1 U4923 ( .C1(n4442), .C2(n4419), .A(n4418), .B(n4417), .ZN(U3282)
         );
  INV_X1 U4924 ( .A(n2841), .ZN(n4420) );
  AOI22_X1 U4925 ( .A1(n4424), .A2(n4423), .B1(n4422), .B2(n4421), .ZN(n4425)
         );
  OAI21_X1 U4926 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n4432) );
  OAI21_X1 U4927 ( .B1(n2841), .B2(n4429), .A(n4428), .ZN(n4499) );
  NOR2_X1 U4928 ( .A1(n4499), .A2(n4430), .ZN(n4431) );
  AOI211_X1 U4929 ( .C1(n4444), .C2(n4433), .A(n4432), .B(n4431), .ZN(n4496)
         );
  AOI22_X1 U4930 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4434), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4442), .ZN(n4441) );
  INV_X1 U4931 ( .A(n4499), .ZN(n4439) );
  OAI21_X1 U4932 ( .B1(n4436), .B2(n4450), .A(n4435), .ZN(n4497) );
  INV_X1 U4933 ( .A(n4497), .ZN(n4437) );
  AOI22_X1 U4934 ( .A1(n4439), .A2(n4443), .B1(n4438), .B2(n4437), .ZN(n4440)
         );
  OAI211_X1 U4935 ( .C1(n4442), .C2(n4496), .A(n4441), .B(n4440), .ZN(U3289)
         );
  AOI22_X1 U4936 ( .A1(n4443), .A2(n4494), .B1(REG2_REG_0__SCAN_IN), .B2(n4442), .ZN(n4456) );
  OAI21_X1 U4937 ( .B1(n4445), .B2(n4444), .A(n4494), .ZN(n4446) );
  OAI21_X1 U4938 ( .B1(n2993), .B2(n4447), .A(n4446), .ZN(n4492) );
  INV_X1 U4939 ( .A(n4448), .ZN(n4449) );
  NOR2_X1 U4940 ( .A1(n4450), .A2(n4449), .ZN(n4493) );
  INV_X1 U4941 ( .A(n4493), .ZN(n4452) );
  NOR2_X1 U4942 ( .A1(n4452), .A2(n4451), .ZN(n4454) );
  OAI21_X1 U4943 ( .B1(n4492), .B2(n4454), .A(n4453), .ZN(n4455) );
  OAI211_X1 U4944 ( .C1(n4457), .C2(n2276), .A(n4456), .B(n4455), .ZN(U3290)
         );
  INV_X1 U4945 ( .A(n4460), .ZN(n4463) );
  NOR2_X1 U4946 ( .A1(n4463), .A2(n4458), .ZN(U3291) );
  AND2_X1 U4947 ( .A1(D_REG_30__SCAN_IN), .A2(n4460), .ZN(U3292) );
  AND2_X1 U4948 ( .A1(D_REG_29__SCAN_IN), .A2(n4460), .ZN(U3293) );
  AND2_X1 U4949 ( .A1(D_REG_28__SCAN_IN), .A2(n4460), .ZN(U3294) );
  AND2_X1 U4950 ( .A1(D_REG_27__SCAN_IN), .A2(n4460), .ZN(U3295) );
  AND2_X1 U4951 ( .A1(D_REG_26__SCAN_IN), .A2(n4460), .ZN(U3296) );
  AND2_X1 U4952 ( .A1(D_REG_25__SCAN_IN), .A2(n4460), .ZN(U3297) );
  AND2_X1 U4953 ( .A1(D_REG_24__SCAN_IN), .A2(n4460), .ZN(U3298) );
  AND2_X1 U4954 ( .A1(D_REG_23__SCAN_IN), .A2(n4460), .ZN(U3299) );
  AND2_X1 U4955 ( .A1(D_REG_22__SCAN_IN), .A2(n4460), .ZN(U3300) );
  AND2_X1 U4956 ( .A1(D_REG_21__SCAN_IN), .A2(n4460), .ZN(U3301) );
  AND2_X1 U4957 ( .A1(D_REG_20__SCAN_IN), .A2(n4460), .ZN(U3302) );
  AND2_X1 U4958 ( .A1(D_REG_19__SCAN_IN), .A2(n4460), .ZN(U3303) );
  AND2_X1 U4959 ( .A1(D_REG_18__SCAN_IN), .A2(n4460), .ZN(U3304) );
  AND2_X1 U4960 ( .A1(D_REG_17__SCAN_IN), .A2(n4460), .ZN(U3305) );
  AND2_X1 U4961 ( .A1(D_REG_16__SCAN_IN), .A2(n4460), .ZN(U3306) );
  AND2_X1 U4962 ( .A1(D_REG_15__SCAN_IN), .A2(n4460), .ZN(U3307) );
  AND2_X1 U4963 ( .A1(D_REG_14__SCAN_IN), .A2(n4460), .ZN(U3308) );
  AND2_X1 U4964 ( .A1(D_REG_13__SCAN_IN), .A2(n4460), .ZN(U3309) );
  NOR2_X1 U4965 ( .A1(n4463), .A2(n4459), .ZN(U3310) );
  AND2_X1 U4966 ( .A1(D_REG_11__SCAN_IN), .A2(n4460), .ZN(U3311) );
  AND2_X1 U4967 ( .A1(D_REG_10__SCAN_IN), .A2(n4460), .ZN(U3312) );
  AND2_X1 U4968 ( .A1(n4460), .A2(D_REG_9__SCAN_IN), .ZN(U3313) );
  AND2_X1 U4969 ( .A1(D_REG_8__SCAN_IN), .A2(n4460), .ZN(U3314) );
  AND2_X1 U4970 ( .A1(D_REG_7__SCAN_IN), .A2(n4460), .ZN(U3315) );
  AND2_X1 U4971 ( .A1(D_REG_6__SCAN_IN), .A2(n4460), .ZN(U3316) );
  AND2_X1 U4972 ( .A1(D_REG_5__SCAN_IN), .A2(n4460), .ZN(U3317) );
  AND2_X1 U4973 ( .A1(D_REG_4__SCAN_IN), .A2(n4460), .ZN(U3318) );
  NOR2_X1 U4974 ( .A1(n4463), .A2(n4461), .ZN(U3319) );
  NOR2_X1 U4975 ( .A1(n4463), .A2(n4462), .ZN(U3320) );
  OAI21_X1 U4976 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4464), .ZN(
        n4465) );
  INV_X1 U4977 ( .A(n4465), .ZN(U3329) );
  INV_X1 U4978 ( .A(DATAI_18_), .ZN(n4466) );
  AOI22_X1 U4979 ( .A1(STATE_REG_SCAN_IN), .A2(n4467), .B1(n4466), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U4980 ( .A(DATAI_17_), .ZN(n4468) );
  AOI22_X1 U4981 ( .A1(STATE_REG_SCAN_IN), .A2(n4469), .B1(n4468), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U4982 ( .A1(U3149), .A2(n4470), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4471) );
  INV_X1 U4983 ( .A(n4471), .ZN(U3336) );
  OAI22_X1 U4984 ( .A1(U3149), .A2(n4472), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4473) );
  INV_X1 U4985 ( .A(n4473), .ZN(U3337) );
  INV_X1 U4986 ( .A(DATAI_14_), .ZN(n4474) );
  AOI22_X1 U4987 ( .A1(STATE_REG_SCAN_IN), .A2(n4475), .B1(n4474), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U4988 ( .A1(STATE_REG_SCAN_IN), .A2(n4477), .B1(n4476), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U4989 ( .A1(STATE_REG_SCAN_IN), .A2(n4478), .B1(n2493), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U4990 ( .A(DATAI_11_), .ZN(n4479) );
  AOI22_X1 U4991 ( .A1(STATE_REG_SCAN_IN), .A2(n4480), .B1(n4479), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U4992 ( .A(DATAI_10_), .ZN(n4481) );
  AOI22_X1 U4993 ( .A1(STATE_REG_SCAN_IN), .A2(n3716), .B1(n4481), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U4994 ( .A1(U3149), .A2(n4482), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4483) );
  INV_X1 U4995 ( .A(n4483), .ZN(U3343) );
  INV_X1 U4996 ( .A(DATAI_8_), .ZN(n4484) );
  AOI22_X1 U4997 ( .A1(STATE_REG_SCAN_IN), .A2(n4485), .B1(n4484), .B2(U3149), 
        .ZN(U3344) );
  OAI22_X1 U4998 ( .A1(U3149), .A2(n4486), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4487) );
  INV_X1 U4999 ( .A(n4487), .ZN(U3346) );
  AOI22_X1 U5000 ( .A1(STATE_REG_SCAN_IN), .A2(n4489), .B1(n4488), .B2(U3149), 
        .ZN(U3347) );
  INV_X1 U5001 ( .A(DATAI_0_), .ZN(n4490) );
  AOI22_X1 U5002 ( .A1(STATE_REG_SCAN_IN), .A2(n2015), .B1(n4490), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5003 ( .C1(n4538), .C2(n4494), .A(n4493), .B(n4492), .ZN(n4545)
         );
  AOI22_X1 U5004 ( .A1(n4544), .A2(n4545), .B1(n4495), .B2(n4542), .ZN(U3467)
         );
  INV_X1 U5005 ( .A(n4496), .ZN(n4501) );
  OAI22_X1 U5006 ( .A1(n4499), .A2(n4498), .B1(n3992), .B2(n4497), .ZN(n4500)
         );
  NOR2_X1 U5007 ( .A1(n4501), .A2(n4500), .ZN(n4547) );
  INV_X1 U5008 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U5009 ( .A1(n4544), .A2(n4547), .B1(n4502), .B2(n4542), .ZN(U3469)
         );
  AND3_X1 U5010 ( .A1(n4504), .A2(n4537), .A3(n4503), .ZN(n4506) );
  AOI211_X1 U5011 ( .C1(n4538), .C2(n4507), .A(n4506), .B(n4505), .ZN(n4549)
         );
  AOI22_X1 U5012 ( .A1(n4544), .A2(n4549), .B1(n4508), .B2(n4542), .ZN(U3471)
         );
  AOI22_X1 U5013 ( .A1(n4510), .A2(n4538), .B1(n4537), .B2(n4509), .ZN(n4511)
         );
  AND2_X1 U5014 ( .A1(n4512), .A2(n4511), .ZN(n4551) );
  INV_X1 U5015 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4513) );
  AOI22_X1 U5016 ( .A1(n4544), .A2(n4551), .B1(n4513), .B2(n4542), .ZN(U3473)
         );
  NAND2_X1 U5017 ( .A1(n4514), .A2(n4538), .ZN(n4516) );
  NAND2_X1 U5018 ( .A1(n4516), .A2(n4515), .ZN(n4517) );
  NOR2_X1 U5019 ( .A1(n4518), .A2(n4517), .ZN(n4552) );
  INV_X1 U5020 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5021 ( .A1(n4544), .A2(n4552), .B1(n4519), .B2(n4542), .ZN(U3475)
         );
  NOR2_X1 U5022 ( .A1(n4521), .A2(n4520), .ZN(n4523) );
  AOI211_X1 U5023 ( .C1(n4537), .C2(n4524), .A(n4523), .B(n4522), .ZN(n4553)
         );
  INV_X1 U5024 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5025 ( .A1(n4544), .A2(n4553), .B1(n4525), .B2(n4542), .ZN(U3477)
         );
  AOI211_X1 U5026 ( .C1(n4528), .C2(n4534), .A(n4527), .B(n4526), .ZN(n4554)
         );
  INV_X1 U5027 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4529) );
  AOI22_X1 U5028 ( .A1(n4544), .A2(n4554), .B1(n4529), .B2(n4542), .ZN(U3481)
         );
  OAI21_X1 U5029 ( .B1(n3992), .B2(n4531), .A(n4530), .ZN(n4532) );
  AOI21_X1 U5030 ( .B1(n4534), .B2(n4533), .A(n4532), .ZN(n4555) );
  INV_X1 U5031 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5032 ( .A1(n4544), .A2(n4555), .B1(n4535), .B2(n4542), .ZN(U3485)
         );
  AOI22_X1 U5033 ( .A1(n4539), .A2(n4538), .B1(n4537), .B2(n4536), .ZN(n4540)
         );
  AND2_X1 U5034 ( .A1(n4541), .A2(n4540), .ZN(n4557) );
  INV_X1 U5035 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5036 ( .A1(n4544), .A2(n4557), .B1(n4543), .B2(n4542), .ZN(U3489)
         );
  AOI22_X1 U5037 ( .A1(n4558), .A2(n4545), .B1(n2283), .B2(n4556), .ZN(U3518)
         );
  AOI22_X1 U5038 ( .A1(n4558), .A2(n4547), .B1(n4546), .B2(n4556), .ZN(U3519)
         );
  AOI22_X1 U5039 ( .A1(n4558), .A2(n4549), .B1(n4548), .B2(n4556), .ZN(U3520)
         );
  AOI22_X1 U5040 ( .A1(n4558), .A2(n4551), .B1(n4550), .B2(n4556), .ZN(U3521)
         );
  AOI22_X1 U5041 ( .A1(n4558), .A2(n4552), .B1(n2330), .B2(n4556), .ZN(U3522)
         );
  AOI22_X1 U5042 ( .A1(n4558), .A2(n4553), .B1(n2355), .B2(n4556), .ZN(U3523)
         );
  AOI22_X1 U5043 ( .A1(n4558), .A2(n4554), .B1(n3004), .B2(n4556), .ZN(U3525)
         );
  AOI22_X1 U5044 ( .A1(n4558), .A2(n4555), .B1(n2430), .B2(n4556), .ZN(U3527)
         );
  AOI22_X1 U5045 ( .A1(n4558), .A2(n4557), .B1(n2466), .B2(n4556), .ZN(U3529)
         );
  CLKBUF_X1 U2262 ( .A(n2319), .Z(n2955) );
  CLKBUF_X1 U2382 ( .A(n2354), .Z(n2953) );
endmodule

