

module b22_C_SARLock_k_128_9 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6558, n6559, n6560, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15407;

  NOR2_X1 U7307 ( .A1(n9285), .A2(n9284), .ZN(n12440) );
  AND2_X1 U7308 ( .A1(n12715), .A2(n12699), .ZN(n6786) );
  INV_X1 U7309 ( .A(n13429), .ZN(n13721) );
  XNOR2_X1 U7310 ( .A(n9190), .B(n9189), .ZN(n11584) );
  NAND2_X1 U7311 ( .A1(n11642), .A2(n11641), .ZN(n11640) );
  CLKBUF_X2 U7312 ( .A(n9963), .Z(n11559) );
  NAND2_X1 U7313 ( .A1(n9680), .A2(n10126), .ZN(n11563) );
  INV_X2 U7314 ( .A(n8901), .ZN(n8849) );
  NAND2_X2 U7315 ( .A1(n9680), .A2(n13307), .ZN(n11564) );
  CLKBUF_X2 U7316 ( .A(n8237), .Z(n8307) );
  CLKBUF_X2 U7317 ( .A(n8270), .Z(n10661) );
  CLKBUF_X2 U7318 ( .A(n8650), .Z(n8671) );
  CLKBUF_X2 U7319 ( .A(n8264), .Z(n8651) );
  NAND2_X1 U7320 ( .A1(n8062), .A2(n8124), .ZN(n8127) );
  INV_X2 U7322 ( .A(n12661), .ZN(n12684) );
  NAND3_X1 U7324 ( .A1(n6750), .A2(n8874), .A3(n8873), .ZN(n12805) );
  AND2_X1 U7325 ( .A1(n12710), .A2(n12693), .ZN(n12715) );
  NOR2_X1 U7326 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7563) );
  NOR2_X1 U7327 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7281) );
  NAND2_X1 U7328 ( .A1(n8748), .A2(n11809), .ZN(n10388) );
  AND2_X1 U7329 ( .A1(n9536), .A2(n9469), .ZN(n8896) );
  INV_X1 U7330 ( .A(n13072), .ZN(n12888) );
  NAND2_X1 U7331 ( .A1(n11149), .A2(n11148), .ZN(n11152) );
  INV_X2 U7332 ( .A(n11476), .ZN(n9952) );
  OR2_X1 U7333 ( .A1(n13830), .A2(n13950), .ZN(n6607) );
  INV_X2 U7334 ( .A(n13444), .ZN(n13472) );
  INV_X1 U7335 ( .A(n13477), .ZN(n13483) );
  AND2_X1 U7336 ( .A1(n7551), .A2(n7501), .ZN(n7362) );
  AND2_X1 U7337 ( .A1(n8176), .A2(n11118), .ZN(n8264) );
  INV_X2 U7339 ( .A(n11911), .ZN(n11948) );
  NAND2_X1 U7340 ( .A1(n8497), .A2(n8496), .ZN(n8517) );
  INV_X2 U7341 ( .A(n12913), .ZN(n9183) );
  INV_X1 U7342 ( .A(n12514), .ZN(n12512) );
  NAND2_X1 U7343 ( .A1(n8808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8809) );
  INV_X2 U7344 ( .A(n9506), .ZN(n7894) );
  INV_X1 U7345 ( .A(n13442), .ZN(n13434) );
  OAI22_X1 U7346 ( .A1(n14117), .A2(n14064), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14063), .ZN(n14065) );
  OAI21_X1 U7347 ( .B1(n12440), .B2(n7024), .A(n12442), .ZN(n6728) );
  NAND2_X1 U7348 ( .A1(n7031), .A2(n12464), .ZN(n12498) );
  AOI21_X1 U7349 ( .B1(n11299), .B2(n6873), .A(n6872), .ZN(n12488) );
  CLKBUF_X3 U7350 ( .A(n8872), .Z(n9239) );
  NAND2_X1 U7351 ( .A1(n7704), .A2(n7703), .ZN(n14578) );
  XNOR2_X1 U7352 ( .A(n14571), .B(n13570), .ZN(n13497) );
  NAND2_X1 U7353 ( .A1(n7717), .A2(n7716), .ZN(n13345) );
  OR2_X1 U7354 ( .A1(n8127), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n8129) );
  NOR2_X1 U7355 ( .A1(n14850), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n14100) );
  INV_X1 U7356 ( .A(n8176), .ZN(n8179) );
  INV_X1 U7357 ( .A(n11962), .ZN(n10182) );
  NAND4_X1 U7358 ( .A1(n8922), .A2(n8921), .A3(n8920), .A4(n8919), .ZN(n12800)
         );
  OR2_X1 U7360 ( .A1(n13886), .A2(n13873), .ZN(n6558) );
  INV_X2 U7361 ( .A(n14550), .ZN(n10480) );
  INV_X2 U7362 ( .A(n7611), .ZN(n13573) );
  NAND2_X1 U7363 ( .A1(n7407), .A2(n7402), .ZN(n8832) );
  NOR2_X2 U7364 ( .A1(n14370), .A2(n11189), .ZN(n11188) );
  XNOR2_X2 U7365 ( .A(n14123), .B(n14124), .ZN(n15393) );
  NAND2_X2 U7366 ( .A1(n14120), .A2(n14119), .ZN(n14123) );
  XNOR2_X2 U7367 ( .A(n8711), .B(n8710), .ZN(n8721) );
  XNOR2_X2 U7368 ( .A(n8809), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U7370 ( .A1(n13449), .A2(n13483), .ZN(n6970) );
  INV_X1 U7372 ( .A(n12512), .ZN(n6560) );
  INV_X2 U7373 ( .A(n7132), .ZN(n10343) );
  AOI211_X2 U7374 ( .C1(n12060), .C2(n14929), .A(n12059), .B(n12058), .ZN(
        n12061) );
  AOI22_X2 U7375 ( .A1(n14089), .A2(n14080), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n14937), .ZN(n14141) );
  AND2_X4 U7376 ( .A1(n8179), .A2(n8175), .ZN(n8298) );
  AOI21_X2 U7377 ( .B1(n10454), .B2(n10451), .A(n10450), .ZN(n10207) );
  AOI21_X2 U7378 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(n10454) );
  INV_X4 U7380 ( .A(n15407), .ZN(n6562) );
  NOR3_X2 U7382 ( .A1(n8837), .A2(n7409), .A3(P2_IR_REG_20__SCAN_IN), .ZN(
        n7401) );
  XNOR2_X2 U7383 ( .A(n8687), .B(P3_IR_REG_20__SCAN_IN), .ZN(n11962) );
  OAI21_X2 U7384 ( .B1(n8276), .B2(n8189), .A(n8190), .ZN(n8289) );
  NAND2_X4 U7385 ( .A1(n6879), .A2(n6878), .ZN(n9469) );
  NAND4_X2 U7386 ( .A1(n12845), .A2(n13681), .A3(n7214), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6879) );
  NAND4_X2 U7387 ( .A1(n7212), .A2(n7213), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6878) );
  XNOR2_X2 U7388 ( .A(n12683), .B(n12682), .ZN(n13473) );
  NOR2_X2 U7389 ( .A1(n7220), .A2(n14171), .ZN(n14395) );
  NOR2_X2 U7390 ( .A1(n14170), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7220) );
  OAI21_X2 U7391 ( .B1(n8674), .B2(n8673), .A(n8675), .ZN(n11752) );
  NAND2_X2 U7392 ( .A1(n8661), .A2(n8660), .ZN(n8674) );
  NOR2_X2 U7393 ( .A1(n14062), .A2(n14061), .ZN(n14117) );
  AOI22_X2 U7394 ( .A1(n10565), .A2(n10566), .B1(n10308), .B2(n10304), .ZN(
        n10551) );
  XNOR2_X2 U7395 ( .A(n12800), .B(n14769), .ZN(n12730) );
  OAI21_X2 U7396 ( .B1(n14137), .B2(n14396), .A(n14393), .ZN(n14400) );
  AND2_X1 U7397 ( .A1(n9393), .A2(n11686), .ZN(n11655) );
  XNOR2_X1 U7398 ( .A(n7023), .B(n12760), .ZN(n13063) );
  AND2_X1 U7399 ( .A1(n11398), .A2(n11397), .ZN(n13065) );
  OAI21_X1 U7400 ( .B1(n11505), .B2(n11504), .A(n13197), .ZN(n13243) );
  AOI21_X1 U7401 ( .B1(n11152), .B2(n7459), .A(n6790), .ZN(n11413) );
  OAI21_X1 U7402 ( .B1(n8517), .B2(n8516), .A(n8518), .ZN(n8538) );
  NAND2_X1 U7403 ( .A1(n8314), .A2(n8313), .ZN(n10619) );
  INV_X1 U7404 ( .A(n13498), .ZN(n10228) );
  NAND2_X1 U7405 ( .A1(n13318), .A2(n13319), .ZN(n14502) );
  OAI21_X2 U7406 ( .B1(n13493), .B2(n10459), .A(n13313), .ZN(n10483) );
  INV_X2 U7407 ( .A(n12536), .ZN(n14769) );
  INV_X4 U7408 ( .A(n13485), .ZN(n6563) );
  NAND2_X1 U7409 ( .A1(n10182), .A2(n12057), .ZN(n9311) );
  NAND2_X1 U7410 ( .A1(n13450), .A2(n13477), .ZN(n13307) );
  NAND2_X1 U7411 ( .A1(n9477), .A2(n12684), .ZN(n8916) );
  CLKBUF_X2 U7412 ( .A(n8902), .Z(n11403) );
  INV_X4 U7413 ( .A(n8877), .ZN(n12913) );
  INV_X1 U7414 ( .A(n14040), .ZN(n7488) );
  AND2_X1 U7415 ( .A1(n7064), .A2(n7437), .ZN(n7062) );
  AND2_X1 U7416 ( .A1(n8802), .A2(n8796), .ZN(n7064) );
  INV_X1 U7417 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n6581) );
  OAI21_X1 U7418 ( .B1(n11728), .B2(n9400), .A(n7515), .ZN(n11604) );
  XNOR2_X1 U7419 ( .A(n11728), .B(n11729), .ZN(n6571) );
  AND2_X1 U7420 ( .A1(n6968), .A2(n11803), .ZN(n7246) );
  NAND2_X2 U7421 ( .A1(n11659), .A2(n9398), .ZN(n11728) );
  NAND2_X1 U7422 ( .A1(n12865), .A2(n11400), .ZN(n7023) );
  NAND2_X1 U7423 ( .A1(n13054), .A2(n12688), .ZN(n12722) );
  NAND2_X1 U7424 ( .A1(n6573), .A2(n9387), .ZN(n11685) );
  CLKBUF_X1 U7425 ( .A(n12851), .Z(n6764) );
  NAND2_X1 U7426 ( .A1(n12663), .A2(n12662), .ZN(n12853) );
  NAND3_X1 U7427 ( .A1(n12498), .A2(n9228), .A3(n12504), .ZN(n12497) );
  NAND2_X1 U7428 ( .A1(n13447), .A2(n13446), .ZN(n13997) );
  NAND2_X1 U7429 ( .A1(n9381), .A2(n9380), .ZN(n9384) );
  AOI21_X1 U7430 ( .B1(n12115), .B2(n12114), .A(n7096), .ZN(n12104) );
  OAI21_X1 U7431 ( .B1(n11752), .B2(n11751), .A(n11753), .ZN(n11758) );
  NAND2_X1 U7432 ( .A1(n12882), .A2(n13065), .ZN(n12868) );
  NAND2_X1 U7433 ( .A1(n13065), .A2(n11425), .ZN(n11426) );
  CLKBUF_X1 U7434 ( .A(n11696), .Z(n6585) );
  NAND2_X1 U7435 ( .A1(n7034), .A2(n7033), .ZN(n7032) );
  OR2_X1 U7436 ( .A1(n12962), .A2(n12961), .ZN(n12964) );
  AND2_X1 U7437 ( .A1(n8047), .A2(n8046), .ZN(n13429) );
  NAND2_X1 U7438 ( .A1(n8102), .A2(n8101), .ZN(n11335) );
  AOI21_X1 U7439 ( .B1(n11353), .B2(n11352), .A(n11351), .ZN(n11358) );
  NAND2_X1 U7440 ( .A1(n6570), .A2(n9371), .ZN(n11634) );
  AND2_X1 U7441 ( .A1(n9231), .A2(n9230), .ZN(n13072) );
  OAI21_X1 U7442 ( .B1(n11332), .B2(n11331), .A(n11330), .ZN(n11353) );
  CLKBUF_X1 U7443 ( .A(n12975), .Z(n6776) );
  XNOR2_X1 U7444 ( .A(n11332), .B(n11331), .ZN(n13165) );
  NAND2_X1 U7445 ( .A1(n11710), .A2(n9370), .ZN(n6570) );
  NAND2_X1 U7446 ( .A1(n6567), .A2(n7558), .ZN(n11710) );
  XNOR2_X1 U7447 ( .A(n8037), .B(n8024), .ZN(n13169) );
  NAND2_X1 U7448 ( .A1(n9365), .A2(n6568), .ZN(n6567) );
  NAND2_X1 U7449 ( .A1(n8766), .A2(n7268), .ZN(n12205) );
  OR2_X1 U7450 ( .A1(n12457), .A2(n6863), .ZN(n6858) );
  AND2_X1 U7451 ( .A1(n12915), .A2(n12914), .ZN(n12917) );
  NAND2_X1 U7452 ( .A1(n7131), .A2(n6639), .ZN(n12206) );
  AND2_X1 U7453 ( .A1(n14145), .A2(n14146), .ZN(n14414) );
  NAND2_X1 U7454 ( .A1(n13288), .A2(n6817), .ZN(n14357) );
  NOR2_X1 U7455 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  NAND2_X1 U7456 ( .A1(n8555), .A2(n8554), .ZN(n12289) );
  AND2_X1 U7457 ( .A1(n11420), .A2(n11394), .ZN(n12961) );
  NOR2_X1 U7458 ( .A1(n14412), .A2(n14411), .ZN(n14410) );
  NAND2_X1 U7459 ( .A1(n8543), .A2(n8542), .ZN(n12293) );
  NOR2_X1 U7460 ( .A1(n9369), .A2(n6569), .ZN(n6568) );
  OAI21_X1 U7461 ( .B1(n14256), .B2(n8435), .A(n8434), .ZN(n11244) );
  NAND2_X1 U7462 ( .A1(n11121), .A2(n9347), .ZN(n11624) );
  NAND2_X1 U7463 ( .A1(n14402), .A2(n7216), .ZN(n14407) );
  NAND2_X1 U7464 ( .A1(n11640), .A2(n6689), .ZN(n11121) );
  NAND2_X1 U7465 ( .A1(n7884), .A2(n7883), .ZN(n13873) );
  NAND2_X1 U7466 ( .A1(n8840), .A2(n8839), .ZN(n13045) );
  NAND2_X1 U7467 ( .A1(n11077), .A2(n7798), .ZN(n11185) );
  AOI22_X1 U7468 ( .A1(n11044), .A2(n11043), .B1(n10949), .B2(n10948), .ZN(
        n10956) );
  NAND2_X1 U7469 ( .A1(n7896), .A2(n7895), .ZN(n14022) );
  OR2_X1 U7470 ( .A1(n10895), .A2(n8757), .ZN(n8759) );
  OAI21_X1 U7471 ( .B1(n14865), .B2(n15070), .A(n14854), .ZN(n12001) );
  NAND2_X1 U7472 ( .A1(n11676), .A2(n6594), .ZN(n7519) );
  OAI21_X1 U7473 ( .B1(n7911), .B2(n7910), .A(n7909), .ZN(n7915) );
  AND3_X1 U7474 ( .A1(n10399), .A2(n6572), .A3(n9329), .ZN(n10518) );
  NAND2_X1 U7475 ( .A1(n9087), .A2(n9086), .ZN(n12599) );
  NAND2_X1 U7476 ( .A1(n7805), .A2(n7804), .ZN(n14370) );
  AOI21_X1 U7477 ( .B1(n14132), .B2(n14131), .A(n14166), .ZN(n14133) );
  AOI22_X1 U7478 ( .A1(n10216), .A2(n10217), .B1(n9327), .B2(n10402), .ZN(
        n10401) );
  NAND2_X1 U7479 ( .A1(n6574), .A2(n9325), .ZN(n10216) );
  OAI21_X1 U7480 ( .B1(n10677), .B2(n15066), .A(n10676), .ZN(n11998) );
  INV_X1 U7481 ( .A(n10519), .ZN(n6572) );
  NAND2_X1 U7482 ( .A1(n9747), .A2(n9748), .ZN(n9881) );
  NAND2_X1 U7483 ( .A1(n9001), .A2(n9000), .ZN(n14803) );
  AND2_X2 U7484 ( .A1(n13707), .A2(n14508), .ZN(n14521) );
  NAND2_X2 U7485 ( .A1(n9847), .A2(n13041), .ZN(n12979) );
  OAI21_X2 U7486 ( .B1(n9692), .B2(n10089), .A(n14508), .ZN(n9693) );
  AOI21_X1 U7487 ( .B1(n13574), .B2(n9685), .A(n9684), .ZN(n9706) );
  AND2_X1 U7488 ( .A1(n10048), .A2(n7267), .ZN(n12342) );
  NAND2_X1 U7489 ( .A1(n7711), .A2(n7710), .ZN(n7325) );
  NAND4_X2 U7490 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(n14978)
         );
  INV_X1 U7491 ( .A(n9308), .ZN(n6564) );
  NAND2_X4 U7492 ( .A1(n11554), .A2(n13884), .ZN(n9958) );
  XNOR2_X1 U7493 ( .A(n10309), .B(n10308), .ZN(n10558) );
  NAND2_X1 U7494 ( .A1(n10307), .A2(n10306), .ZN(n10309) );
  OAI211_X1 U7495 ( .C1(n8277), .C2(n9463), .A(n8247), .B(n8246), .ZN(n10048)
         );
  OAI211_X1 U7496 ( .C1(n8277), .C2(n9452), .A(n8240), .B(n8239), .ZN(n10393)
         );
  NAND2_X1 U7497 ( .A1(n8268), .A2(n6617), .ZN(n14979) );
  NAND2_X2 U7498 ( .A1(n7656), .A2(n7655), .ZN(n14571) );
  NAND2_X1 U7499 ( .A1(n13573), .A2(n10480), .ZN(n13299) );
  NAND4_X1 U7500 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n12329)
         );
  OR2_X2 U7501 ( .A1(n9985), .A2(n13483), .ZN(n13884) );
  NAND2_X1 U7502 ( .A1(n8245), .A2(n12680), .ZN(n8277) );
  BUF_X2 U7503 ( .A(n8245), .Z(n8698) );
  AND2_X1 U7504 ( .A1(n8245), .A2(n9469), .ZN(n8237) );
  NAND2_X1 U7505 ( .A1(n11329), .A2(n12037), .ZN(n8245) );
  CLKBUF_X3 U7506 ( .A(n8904), .Z(n12668) );
  INV_X1 U7508 ( .A(n12011), .ZN(n12057) );
  AOI21_X1 U7509 ( .B1(n7741), .B2(n7333), .A(n7331), .ZN(n7330) );
  NAND2_X1 U7510 ( .A1(n8179), .A2(n11118), .ZN(n8270) );
  NAND2_X1 U7511 ( .A1(n9733), .A2(n9732), .ZN(n13026) );
  BUF_X4 U7512 ( .A(n12037), .Z(n6590) );
  AND2_X1 U7513 ( .A1(n8523), .A2(n8686), .ZN(n12011) );
  NAND2_X1 U7514 ( .A1(n6822), .A2(n6819), .ZN(n14044) );
  CLKBUF_X3 U7515 ( .A(n8896), .Z(n12685) );
  NAND2_X1 U7516 ( .A1(n8066), .A2(n8065), .ZN(n13477) );
  NAND2_X1 U7517 ( .A1(n8128), .A2(n8129), .ZN(n14048) );
  NAND2_X1 U7518 ( .A1(n8712), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8711) );
  OR2_X1 U7519 ( .A1(n13438), .A2(n10468), .ZN(n7588) );
  AND2_X1 U7520 ( .A1(n8176), .A2(n8175), .ZN(n8650) );
  XNOR2_X1 U7521 ( .A(n8685), .B(P3_IR_REG_21__SCAN_IN), .ZN(n11772) );
  OAI21_X1 U7522 ( .B1(n8686), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8685) );
  NAND2_X2 U7523 ( .A1(n9536), .A2(n12680), .ZN(n12661) );
  NAND2_X1 U7524 ( .A1(n8129), .A2(n6741), .ZN(n6822) );
  AND2_X1 U7525 ( .A1(n11334), .A2(n11576), .ZN(n8917) );
  AND2_X1 U7526 ( .A1(n8125), .A2(n8127), .ZN(n9482) );
  NAND2_X2 U7527 ( .A1(n11360), .A2(n7488), .ZN(n13442) );
  NAND2_X1 U7528 ( .A1(n6580), .A2(n6581), .ZN(n8738) );
  NAND2_X1 U7529 ( .A1(n8225), .A2(n8224), .ZN(n12037) );
  NAND2_X1 U7530 ( .A1(n10284), .A2(n10283), .ZN(n10286) );
  AOI21_X1 U7531 ( .B1(n6593), .B2(n6923), .A(n6667), .ZN(n6922) );
  INV_X1 U7532 ( .A(n6593), .ZN(n6924) );
  NAND2_X1 U7533 ( .A1(n8807), .A2(n8808), .ZN(n11334) );
  MUX2_X1 U7534 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8223), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8225) );
  XNOR2_X1 U7535 ( .A(n8220), .B(n8219), .ZN(n11329) );
  NOR2_X1 U7536 ( .A1(n8719), .A2(n8718), .ZN(n8736) );
  OR2_X1 U7537 ( .A1(n8522), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8686) );
  NOR2_X1 U7538 ( .A1(n14055), .A2(n14056), .ZN(n14058) );
  XNOR2_X1 U7539 ( .A(n7571), .B(n7570), .ZN(n14040) );
  NAND2_X1 U7540 ( .A1(n8224), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8220) );
  NOR2_X1 U7541 ( .A1(n6821), .A2(n6820), .ZN(n6819) );
  MUX2_X1 U7542 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8806), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n8807) );
  NAND2_X1 U7543 ( .A1(n14032), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7568) );
  NAND2_X2 U7544 ( .A1(n8042), .A2(P1_U3086), .ZN(n14047) );
  AOI21_X1 U7545 ( .B1(n8837), .B2(n7406), .A(n7403), .ZN(n7402) );
  XNOR2_X1 U7546 ( .A(n8828), .B(n8827), .ZN(n9539) );
  INV_X1 U7547 ( .A(n8689), .ZN(n7533) );
  NAND2_X1 U7548 ( .A1(n8826), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8828) );
  NAND2_X2 U7549 ( .A1(n9474), .A2(P1_U3086), .ZN(n14043) );
  XNOR2_X1 U7550 ( .A(n8825), .B(P2_IR_REG_21__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U7551 ( .A1(n8821), .A2(n8820), .ZN(n8837) );
  INV_X1 U7552 ( .A(n9111), .ZN(n8821) );
  INV_X1 U7553 ( .A(n12680), .ZN(n9474) );
  AOI21_X1 U7554 ( .B1(n14097), .B2(n14098), .A(n7222), .ZN(n14054) );
  NAND2_X2 U7555 ( .A1(n9469), .A2(P2_U3088), .ZN(n13160) );
  NAND2_X1 U7556 ( .A1(n8818), .A2(n6599), .ZN(n9111) );
  INV_X1 U7557 ( .A(n7136), .ZN(n7082) );
  AND2_X1 U7558 ( .A1(n9050), .A2(n7436), .ZN(n7435) );
  AND2_X1 U7559 ( .A1(n6566), .A2(n6565), .ZN(n7507) );
  AND2_X1 U7560 ( .A1(n8161), .A2(n8162), .ZN(n7506) );
  AND4_X1 U7561 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n7542)
         );
  AND2_X1 U7562 ( .A1(n8793), .A2(n8792), .ZN(n9049) );
  AND2_X1 U7563 ( .A1(n6739), .A2(n8794), .ZN(n9050) );
  AND2_X1 U7564 ( .A1(n8397), .A2(n7504), .ZN(n7265) );
  INV_X1 U7565 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9277) );
  INV_X1 U7566 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7567) );
  NOR2_X1 U7567 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8792) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8793) );
  INV_X1 U7569 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7213) );
  INV_X1 U7570 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7212) );
  INV_X4 U7571 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7572 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7573 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7283) );
  NOR2_X1 U7574 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n7276) );
  NOR2_X1 U7575 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7277) );
  NOR2_X1 U7576 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7278) );
  NOR2_X1 U7577 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6820) );
  NOR2_X1 U7578 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6739) );
  INV_X1 U7579 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9244) );
  INV_X1 U7580 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8397) );
  XNOR2_X1 U7581 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14099) );
  NOR2_X1 U7582 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n6566) );
  INV_X1 U7583 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8739) );
  NOR2_X1 U7584 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n6565) );
  INV_X1 U7585 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8710) );
  INV_X1 U7586 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n15181) );
  INV_X1 U7587 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8161) );
  INV_X1 U7588 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7083) );
  INV_X4 U7589 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7590 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8422) );
  INV_X1 U7591 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8437) );
  NOR2_X1 U7592 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8163) );
  INV_X1 U7593 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8500) );
  INV_X1 U7594 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U7595 ( .A1(n9365), .A2(n9364), .ZN(n11361) );
  INV_X1 U7596 ( .A(n9364), .ZN(n6569) );
  NAND2_X1 U7597 ( .A1(n6571), .A2(n11730), .ZN(n11736) );
  NOR2_X2 U7598 ( .A1(n10518), .A2(n9333), .ZN(n11676) );
  NAND2_X1 U7599 ( .A1(n11702), .A2(n9385), .ZN(n6573) );
  NAND3_X1 U7600 ( .A1(n9384), .A2(n12165), .A3(n9385), .ZN(n11702) );
  NAND2_X1 U7601 ( .A1(n9383), .A2(n9382), .ZN(n9385) );
  OAI211_X1 U7602 ( .C1(n10391), .C2(n12336), .A(n6574), .B(n10390), .ZN(
        n10392) );
  NAND2_X1 U7603 ( .A1(n9323), .A2(n10391), .ZN(n6574) );
  NAND2_X1 U7604 ( .A1(n11606), .A2(n9339), .ZN(n11642) );
  XNOR2_X2 U7605 ( .A(n6575), .B(n8172), .ZN(n8176) );
  NOR2_X1 U7606 ( .A1(n12407), .A2(n8716), .ZN(n6575) );
  NOR2_X2 U7607 ( .A1(n8173), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n12407) );
  AOI21_X1 U7608 ( .B1(n7624), .B2(n7625), .A(n7623), .ZN(n7641) );
  OAI21_X2 U7609 ( .B1(n8003), .B2(n8002), .A(n8001), .ZN(n8020) );
  AND2_X2 U7610 ( .A1(n12900), .A2(n12917), .ZN(n12895) );
  OR2_X1 U7611 ( .A1(n10438), .A2(n12545), .ZN(n10509) );
  AND2_X2 U7612 ( .A1(n7219), .A2(n7218), .ZN(n14174) );
  NOR2_X2 U7613 ( .A1(n14113), .A2(n14114), .ZN(n14115) );
  XNOR2_X1 U7614 ( .A(n10343), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U7615 ( .A1(n9393), .A2(n6579), .ZN(n6576) );
  AND2_X2 U7616 ( .A1(n6576), .A2(n6577), .ZN(n11659) );
  OR2_X1 U7617 ( .A1(n6578), .A2(n11656), .ZN(n6577) );
  INV_X1 U7618 ( .A(n11657), .ZN(n6578) );
  AND2_X1 U7619 ( .A1(n11686), .A2(n11657), .ZN(n6579) );
  AND2_X1 U7620 ( .A1(n8739), .A2(n6581), .ZN(n6582) );
  INV_X1 U7621 ( .A(n8709), .ZN(n6580) );
  NAND2_X4 U7622 ( .A1(n8836), .A2(n12762), .ZN(n9731) );
  XNOR2_X2 U7623 ( .A(n12765), .B(n12778), .ZN(n8836) );
  AND2_X2 U7624 ( .A1(n6772), .A2(n6773), .ZN(n14412) );
  AND2_X1 U7625 ( .A1(n11702), .A2(n9385), .ZN(n6583) );
  NAND2_X1 U7626 ( .A1(n10399), .A2(n9329), .ZN(n6584) );
  NAND2_X1 U7627 ( .A1(n9313), .A2(n9312), .ZN(n6586) );
  NAND2_X1 U7629 ( .A1(n10401), .A2(n10400), .ZN(n10399) );
  NAND2_X1 U7630 ( .A1(n9374), .A2(n9373), .ZN(n11696) );
  NAND2_X1 U7631 ( .A1(n9313), .A2(n9312), .ZN(n9326) );
  NAND2_X2 U7632 ( .A1(n9319), .A2(n9317), .ZN(n8748) );
  INV_X2 U7633 ( .A(n8254), .ZN(n9319) );
  NOR2_X2 U7634 ( .A1(n13114), .A2(n13039), .ZN(n13013) );
  OR2_X2 U7635 ( .A1(n13045), .A2(n13038), .ZN(n13039) );
  NOR2_X1 U7636 ( .A1(n8689), .A2(n8501), .ZN(n8505) );
  OAI22_X2 U7637 ( .A1(n12127), .A2(n12126), .B1(n12139), .B2(n12279), .ZN(
        n12115) );
  OAI211_X1 U7638 ( .C1(n12661), .C2(n9525), .A(n8860), .B(n7543), .ZN(n12514)
         );
  CLKBUF_X1 U7639 ( .A(n8896), .Z(n6588) );
  CLKBUF_X2 U7640 ( .A(n12531), .Z(n6589) );
  OAI211_X1 U7641 ( .C1(n12661), .C2(n9501), .A(n8886), .B(n8885), .ZN(n12531)
         );
  OAI21_X1 U7642 ( .B1(n8712), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8713) );
  OR2_X1 U7643 ( .A1(n10106), .A2(n12531), .ZN(n10531) );
  NAND2_X2 U7644 ( .A1(n11625), .A2(n9353), .ZN(n11304) );
  AOI21_X1 U7645 ( .B1(n11809), .B2(n9318), .A(n9320), .ZN(n9324) );
  INV_X1 U7646 ( .A(n9389), .ZN(n9394) );
  OAI21_X2 U7647 ( .B1(n11696), .B2(n7527), .A(n7523), .ZN(n9383) );
  OR2_X1 U7648 ( .A1(n12273), .A2(n12125), .ZN(n11932) );
  AND2_X1 U7649 ( .A1(n11892), .A2(n11891), .ZN(n12218) );
  NOR2_X1 U7650 ( .A1(n13795), .A2(n7318), .ZN(n7317) );
  INV_X1 U7651 ( .A(n8096), .ZN(n7318) );
  NAND2_X1 U7652 ( .A1(n10337), .A2(n10336), .ZN(n10335) );
  NAND2_X1 U7653 ( .A1(n7146), .A2(n10285), .ZN(n10274) );
  NAND2_X1 U7654 ( .A1(n10335), .A2(n10273), .ZN(n7146) );
  OR2_X1 U7655 ( .A1(n12281), .A2(n12154), .ZN(n11924) );
  OR2_X1 U7656 ( .A1(n12300), .A2(n11711), .ZN(n11895) );
  NAND2_X1 U7657 ( .A1(n8810), .A2(n8811), .ZN(n8902) );
  INV_X1 U7658 ( .A(n11334), .ZN(n8810) );
  AND2_X1 U7659 ( .A1(n9731), .A2(n14822), .ZN(n13140) );
  NAND2_X1 U7660 ( .A1(n7932), .A2(n7931), .ZN(n7943) );
  OR2_X1 U7661 ( .A1(n12526), .A2(n12527), .ZN(n7174) );
  AND2_X1 U7662 ( .A1(n12592), .A2(n7182), .ZN(n7181) );
  INV_X1 U7663 ( .A(n12590), .ZN(n7182) );
  NAND2_X1 U7664 ( .A1(n12593), .A2(n12590), .ZN(n7180) );
  NAND2_X1 U7665 ( .A1(n7198), .A2(n7197), .ZN(n12621) );
  NAND2_X1 U7666 ( .A1(n12615), .A2(n12617), .ZN(n7197) );
  NAND2_X1 U7667 ( .A1(n7205), .A2(n12627), .ZN(n7204) );
  INV_X1 U7668 ( .A(n12628), .ZN(n7205) );
  NOR2_X1 U7669 ( .A1(n7372), .A2(n7370), .ZN(n7369) );
  NOR2_X1 U7670 ( .A1(n7007), .A2(n13427), .ZN(n7006) );
  NAND2_X1 U7671 ( .A1(n6922), .A2(n6924), .ZN(n6921) );
  NAND3_X1 U7672 ( .A1(n7265), .A2(n7082), .A3(n7534), .ZN(n7262) );
  NAND2_X1 U7673 ( .A1(n12666), .A2(n12665), .ZN(n12707) );
  NAND2_X1 U7674 ( .A1(n12853), .A2(n12664), .ZN(n12666) );
  INV_X1 U7675 ( .A(n11456), .ZN(n6836) );
  XNOR2_X1 U7676 ( .A(n13297), .B(n13525), .ZN(n13449) );
  NAND2_X1 U7677 ( .A1(n7846), .A2(n8484), .ZN(n7862) );
  OR2_X1 U7678 ( .A1(n7800), .A2(SI_14_), .ZN(n7056) );
  NOR2_X1 U7679 ( .A1(n7762), .A2(n7334), .ZN(n7333) );
  INV_X1 U7680 ( .A(n7745), .ZN(n7334) );
  OAI21_X1 U7681 ( .B1(n7159), .B2(n7158), .A(n7156), .ZN(n11982) );
  INV_X1 U7682 ( .A(n7161), .ZN(n7158) );
  AOI21_X1 U7683 ( .B1(n6591), .B2(n6632), .A(n7157), .ZN(n7156) );
  NAND2_X1 U7684 ( .A1(n10351), .A2(n6591), .ZN(n7159) );
  NOR2_X1 U7685 ( .A1(n12266), .A2(n12079), .ZN(n7098) );
  NAND2_X1 U7686 ( .A1(n12110), .A2(n12117), .ZN(n7099) );
  NAND2_X1 U7687 ( .A1(n6672), .A2(n7100), .ZN(n7097) );
  NAND2_X1 U7688 ( .A1(n12273), .A2(n11970), .ZN(n7100) );
  INV_X1 U7689 ( .A(n11792), .ZN(n7110) );
  INV_X1 U7690 ( .A(n7115), .ZN(n7114) );
  OAI21_X1 U7691 ( .B1(n11788), .B2(n7116), .A(n8479), .ZN(n7115) );
  OR2_X1 U7692 ( .A1(n12279), .A2(n11971), .ZN(n11927) );
  NAND2_X1 U7693 ( .A1(n12176), .A2(n11907), .ZN(n7240) );
  INV_X1 U7694 ( .A(n6955), .ZN(n6954) );
  OAI21_X1 U7695 ( .B1(n8550), .B2(n6956), .A(n8561), .ZN(n6955) );
  NAND2_X1 U7696 ( .A1(n7084), .A2(n7083), .ZN(n7136) );
  INV_X1 U7697 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7084) );
  AND2_X1 U7698 ( .A1(n13078), .A2(n12785), .ZN(n11396) );
  NOR2_X1 U7699 ( .A1(n7339), .A2(n7072), .ZN(n7071) );
  INV_X1 U7700 ( .A(n12755), .ZN(n7072) );
  INV_X1 U7701 ( .A(n9958), .ZN(n11558) );
  INV_X1 U7702 ( .A(n7358), .ZN(n7357) );
  AND2_X1 U7703 ( .A1(n8067), .A2(n13307), .ZN(n11476) );
  INV_X1 U7704 ( .A(n9481), .ZN(n8145) );
  OR2_X1 U7705 ( .A1(n13297), .A2(n13450), .ZN(n9985) );
  OAI21_X1 U7706 ( .B1(n7325), .B2(n6924), .A(n6922), .ZN(n7743) );
  NAND2_X1 U7707 ( .A1(n7346), .A2(n7652), .ZN(n7665) );
  AND2_X1 U7708 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  INV_X1 U7709 ( .A(n12329), .ZN(n10520) );
  OR2_X1 U7710 ( .A1(n10374), .A2(n10273), .ZN(n7147) );
  OR2_X1 U7711 ( .A1(n14871), .A2(n7153), .ZN(n7150) );
  OR2_X1 U7712 ( .A1(n14888), .A2(n14872), .ZN(n7153) );
  NAND2_X1 U7713 ( .A1(n11986), .A2(n7152), .ZN(n7151) );
  INV_X1 U7714 ( .A(n14888), .ZN(n7152) );
  OR2_X1 U7715 ( .A1(n12113), .A2(n8768), .ZN(n8769) );
  AND2_X1 U7716 ( .A1(n12126), .A2(n11924), .ZN(n7274) );
  NAND2_X1 U7717 ( .A1(n7104), .A2(n7106), .ZN(n7101) );
  AND2_X1 U7718 ( .A1(n11895), .A2(n11897), .ZN(n12208) );
  NOR2_X1 U7719 ( .A1(n12218), .A2(n7129), .ZN(n7128) );
  INV_X1 U7720 ( .A(n12236), .ZN(n7129) );
  NAND2_X1 U7721 ( .A1(n11234), .A2(n11788), .ZN(n11233) );
  NAND2_X1 U7722 ( .A1(n10778), .A2(n6631), .ZN(n14948) );
  NAND2_X1 U7723 ( .A1(n11924), .A2(n8596), .ZN(n12140) );
  NAND2_X1 U7724 ( .A1(n12205), .A2(n6650), .ZN(n12186) );
  INV_X1 U7725 ( .A(n12190), .ZN(n7270) );
  INV_X1 U7726 ( .A(n12208), .ZN(n12202) );
  AOI21_X1 U7727 ( .B1(n12235), .B2(n7232), .A(n7231), .ZN(n7230) );
  INV_X1 U7728 ( .A(n11886), .ZN(n7232) );
  XNOR2_X1 U7729 ( .A(n8174), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U7730 ( .A1(n8173), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8174) );
  INV_X1 U7731 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U7732 ( .A1(n6967), .A2(n8210), .ZN(n8467) );
  NAND2_X1 U7733 ( .A1(n8451), .A2(n8449), .ZN(n6967) );
  NAND2_X1 U7734 ( .A1(n12497), .A2(n7025), .ZN(n9285) );
  NAND2_X1 U7735 ( .A1(n9227), .A2(n7026), .ZN(n7025) );
  INV_X1 U7736 ( .A(n9229), .ZN(n7026) );
  AND2_X1 U7737 ( .A1(n9201), .A2(n9200), .ZN(n7035) );
  INV_X1 U7738 ( .A(n12796), .ZN(n10686) );
  INV_X1 U7739 ( .A(n8861), .ZN(n8904) );
  OR2_X1 U7740 ( .A1(n14686), .A2(n14685), .ZN(n14683) );
  NAND2_X1 U7741 ( .A1(n13009), .A2(n11388), .ZN(n7053) );
  NOR2_X1 U7742 ( .A1(n13005), .A2(n13045), .ZN(n11414) );
  INV_X1 U7743 ( .A(n7049), .ZN(n7046) );
  NOR2_X1 U7744 ( .A1(n12746), .A2(n7037), .ZN(n7041) );
  INV_X1 U7745 ( .A(n7043), .ZN(n7037) );
  OR2_X1 U7746 ( .A1(n12594), .A2(n14305), .ZN(n7049) );
  INV_X2 U7747 ( .A(n9536), .ZN(n9135) );
  NAND2_X1 U7748 ( .A1(n8803), .A2(n8827), .ZN(n7470) );
  NAND2_X1 U7749 ( .A1(n15197), .A2(n7410), .ZN(n7409) );
  NAND2_X1 U7750 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n7410) );
  NAND2_X1 U7751 ( .A1(n14040), .A2(n11360), .ZN(n7980) );
  NAND2_X1 U7752 ( .A1(n13747), .A2(n6597), .ZN(n8102) );
  NAND2_X1 U7753 ( .A1(n7315), .A2(n6642), .ZN(n7314) );
  OR2_X2 U7754 ( .A1(n13268), .A2(n13554), .ZN(n8097) );
  NAND2_X1 U7755 ( .A1(n13810), .A2(n7317), .ZN(n13792) );
  NAND2_X1 U7756 ( .A1(n13818), .A2(n7941), .ZN(n13791) );
  NAND2_X1 U7757 ( .A1(n13958), .A2(n6936), .ZN(n13818) );
  AND2_X1 U7758 ( .A1(n13808), .A2(n7926), .ZN(n6936) );
  NAND2_X1 U7759 ( .A1(n6881), .A2(n6880), .ZN(n13886) );
  INV_X1 U7760 ( .A(n10082), .ZN(n7352) );
  INV_X1 U7761 ( .A(n10084), .ZN(n7354) );
  NAND2_X1 U7762 ( .A1(n8107), .A2(n8106), .ZN(n14585) );
  XNOR2_X1 U7763 ( .A(n8020), .B(n8004), .ZN(n13173) );
  INV_X1 U7764 ( .A(n7973), .ZN(n6765) );
  NOR2_X1 U7765 ( .A1(n7343), .A2(n7916), .ZN(n7340) );
  OAI21_X1 U7766 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14898), .A(n14078), .ZN(
        n14090) );
  OR2_X1 U7767 ( .A1(n11712), .A2(n12224), .ZN(n9370) );
  INV_X1 U7768 ( .A(n11974), .ZN(n12179) );
  NOR2_X1 U7769 ( .A1(n8452), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8468) );
  AND2_X1 U7770 ( .A1(n14322), .A2(n9125), .ZN(n9126) );
  NOR2_X1 U7771 ( .A1(n12761), .A2(n12767), .ZN(n6789) );
  XNOR2_X1 U7772 ( .A(n6766), .B(n12762), .ZN(n12761) );
  OAI21_X1 U7773 ( .B1(n12840), .B2(n14695), .A(n6911), .ZN(n6910) );
  AOI21_X1 U7774 ( .B1(n12841), .B2(n14655), .A(n14719), .ZN(n6911) );
  NAND2_X1 U7775 ( .A1(n8026), .A2(n8025), .ZN(n13915) );
  INV_X1 U7776 ( .A(n13321), .ZN(n13571) );
  XNOR2_X1 U7777 ( .A(n13662), .B(n13661), .ZN(n13676) );
  AND2_X1 U7778 ( .A1(n9609), .A2(n14041), .ZN(n14483) );
  NAND2_X1 U7779 ( .A1(n14404), .A2(n14403), .ZN(n14402) );
  OR2_X1 U7780 ( .A1(n12535), .A2(n12534), .ZN(n6787) );
  OR2_X1 U7781 ( .A1(n12546), .A2(n12548), .ZN(n6732) );
  NAND2_X1 U7782 ( .A1(n12560), .A2(n7194), .ZN(n7193) );
  INV_X1 U7783 ( .A(n12559), .ZN(n7194) );
  AND2_X1 U7784 ( .A1(n6986), .A2(n13303), .ZN(n6985) );
  AND2_X1 U7785 ( .A1(n13305), .A2(n13306), .ZN(n7376) );
  NAND2_X1 U7786 ( .A1(n12580), .A2(n12579), .ZN(n12583) );
  OR2_X1 U7787 ( .A1(n12591), .A2(n7181), .ZN(n7176) );
  AND2_X1 U7788 ( .A1(n7180), .A2(n7178), .ZN(n6743) );
  NAND2_X1 U7789 ( .A1(n7179), .A2(n7177), .ZN(n12596) );
  AOI21_X1 U7790 ( .B1(n7181), .B2(n7180), .A(n7178), .ZN(n7177) );
  NAND2_X1 U7791 ( .A1(n6973), .A2(n6972), .ZN(n13347) );
  NAND2_X1 U7792 ( .A1(n13342), .A2(n13344), .ZN(n6972) );
  NAND2_X1 U7793 ( .A1(n13347), .A2(n13348), .ZN(n6971) );
  NAND2_X1 U7794 ( .A1(n13365), .A2(n7384), .ZN(n7383) );
  INV_X1 U7795 ( .A(n13367), .ZN(n6982) );
  AND2_X1 U7796 ( .A1(n6980), .A2(n6983), .ZN(n6978) );
  NAND2_X1 U7797 ( .A1(n7203), .A2(n7201), .ZN(n12631) );
  AOI21_X1 U7798 ( .B1(n7206), .B2(n7204), .A(n7202), .ZN(n7201) );
  NAND2_X1 U7799 ( .A1(n6730), .A2(n6729), .ZN(n7200) );
  INV_X1 U7800 ( .A(n7206), .ZN(n6729) );
  INV_X1 U7801 ( .A(n12629), .ZN(n6730) );
  NAND2_X1 U7802 ( .A1(n7013), .A2(n6645), .ZN(n7012) );
  INV_X1 U7803 ( .A(n7016), .ZN(n7013) );
  AOI21_X1 U7804 ( .B1(n13401), .B2(n13402), .A(n7374), .ZN(n7373) );
  INV_X1 U7805 ( .A(n13399), .ZN(n7374) );
  AND2_X1 U7806 ( .A1(n13384), .A2(n13383), .ZN(n7554) );
  NAND2_X1 U7807 ( .A1(n7015), .A2(n13513), .ZN(n7014) );
  NAND2_X1 U7808 ( .A1(n7016), .A2(n7889), .ZN(n7015) );
  NAND2_X1 U7809 ( .A1(n13406), .A2(n6991), .ZN(n6989) );
  NAND2_X1 U7810 ( .A1(n13408), .A2(n6992), .ZN(n6991) );
  INV_X1 U7811 ( .A(n7372), .ZN(n7368) );
  NAND2_X1 U7812 ( .A1(n13407), .A2(n13409), .ZN(n6990) );
  INV_X1 U7813 ( .A(n13410), .ZN(n7367) );
  NAND2_X1 U7814 ( .A1(n13414), .A2(n13417), .ZN(n6975) );
  INV_X1 U7815 ( .A(n12646), .ZN(n6744) );
  NOR2_X1 U7816 ( .A1(n6598), .A2(n7006), .ZN(n7003) );
  INV_X1 U7817 ( .A(n13425), .ZN(n7363) );
  INV_X1 U7818 ( .A(n7006), .ZN(n7005) );
  NOR2_X1 U7819 ( .A1(n11772), .A2(n10182), .ZN(n9309) );
  NOR2_X1 U7820 ( .A1(n10779), .A2(n8337), .ZN(n7242) );
  INV_X1 U7821 ( .A(n11841), .ZN(n7244) );
  OAI21_X1 U7822 ( .B1(n8090), .B2(n7301), .A(n7298), .ZN(n13860) );
  INV_X1 U7823 ( .A(n13387), .ZN(n7301) );
  AND2_X1 U7824 ( .A1(n13862), .A2(n7299), .ZN(n7298) );
  NAND2_X1 U7825 ( .A1(n7300), .A2(n13387), .ZN(n7299) );
  INV_X1 U7826 ( .A(n7780), .ZN(n6928) );
  OR2_X1 U7827 ( .A1(n7060), .A2(n7816), .ZN(n7057) );
  NAND2_X1 U7828 ( .A1(n7818), .A2(n9824), .ZN(n7844) );
  INV_X1 U7829 ( .A(SI_13_), .ZN(n7782) );
  AOI21_X1 U7830 ( .B1(n7330), .B2(n7332), .A(n7329), .ZN(n7328) );
  INV_X1 U7831 ( .A(n7545), .ZN(n7329) );
  AOI21_X1 U7832 ( .B1(n7663), .B2(n7667), .A(n7680), .ZN(n6869) );
  INV_X1 U7833 ( .A(n7667), .ZN(n6870) );
  INV_X1 U7834 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14057) );
  AND3_X1 U7835 ( .A1(n8296), .A2(n8295), .A3(n8294), .ZN(n9330) );
  INV_X1 U7836 ( .A(n11956), .ZN(n11775) );
  INV_X1 U7837 ( .A(n14285), .ZN(n11771) );
  NOR2_X1 U7838 ( .A1(n8771), .A2(n11944), .ZN(n7250) );
  NAND2_X1 U7839 ( .A1(n11775), .A2(n11774), .ZN(n11804) );
  AOI21_X1 U7840 ( .B1(n11773), .B2(n11799), .A(n11801), .ZN(n11774) );
  NOR2_X1 U7841 ( .A1(n14285), .A2(n11766), .ZN(n11799) );
  INV_X1 U7842 ( .A(n10315), .ZN(n7144) );
  AOI21_X1 U7843 ( .B1(n7143), .B2(n10315), .A(n10308), .ZN(n7142) );
  AND2_X1 U7844 ( .A1(n7105), .A2(n6685), .ZN(n7104) );
  OR2_X1 U7845 ( .A1(n6614), .A2(n7106), .ZN(n7105) );
  INV_X1 U7846 ( .A(n8464), .ZN(n7116) );
  NAND2_X1 U7847 ( .A1(n10520), .A2(n9315), .ZN(n11819) );
  NAND2_X1 U7848 ( .A1(n8748), .A2(n12342), .ZN(n9322) );
  OR2_X1 U7849 ( .A1(n8672), .A2(n12093), .ZN(n7552) );
  OR2_X1 U7850 ( .A1(n12266), .A2(n12102), .ZN(n11941) );
  INV_X1 U7851 ( .A(n11907), .ZN(n7237) );
  OR2_X1 U7852 ( .A1(n12196), .A2(n11975), .ZN(n11902) );
  AND2_X1 U7853 ( .A1(n8219), .A2(n8218), .ZN(n8171) );
  INV_X1 U7854 ( .A(n8552), .ZN(n6956) );
  INV_X1 U7855 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U7856 ( .A1(n9186), .A2(n9185), .ZN(n6864) );
  INV_X1 U7857 ( .A(n9170), .ZN(n6862) );
  NAND2_X1 U7858 ( .A1(n12722), .A2(n12689), .ZN(n6769) );
  INV_X1 U7859 ( .A(n12760), .ZN(n6767) );
  NAND2_X1 U7860 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  NAND2_X1 U7861 ( .A1(n14665), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6897) );
  AND2_X1 U7862 ( .A1(n6896), .A2(n12820), .ZN(n12828) );
  OR2_X1 U7863 ( .A1(n7460), .A2(n7458), .ZN(n7457) );
  INV_X1 U7864 ( .A(n11282), .ZN(n7458) );
  INV_X1 U7865 ( .A(n7045), .ZN(n7039) );
  NOR2_X1 U7866 ( .A1(n11217), .A2(n7464), .ZN(n7463) );
  INV_X1 U7867 ( .A(n11151), .ZN(n7464) );
  NOR2_X1 U7868 ( .A1(n11252), .A2(n7461), .ZN(n7460) );
  INV_X1 U7869 ( .A(n11216), .ZN(n7461) );
  INV_X1 U7870 ( .A(n7444), .ZN(n7439) );
  NAND2_X1 U7871 ( .A1(n6883), .A2(n6882), .ZN(n10852) );
  INV_X1 U7872 ( .A(n14811), .ZN(n6882) );
  INV_X1 U7873 ( .A(n9730), .ZN(n9279) );
  INV_X1 U7874 ( .A(n12727), .ZN(n10098) );
  INV_X1 U7875 ( .A(n11516), .ZN(n6830) );
  AND2_X1 U7876 ( .A1(n13217), .A2(n6845), .ZN(n6844) );
  OR2_X1 U7877 ( .A1(n13234), .A2(n6846), .ZN(n6845) );
  INV_X1 U7878 ( .A(n11538), .ZN(n6846) );
  OR2_X1 U7879 ( .A1(n14384), .A2(n11478), .ZN(n13378) );
  NOR2_X1 U7880 ( .A1(n11101), .A2(n7361), .ZN(n7360) );
  INV_X1 U7881 ( .A(n7815), .ZN(n7361) );
  AOI21_X1 U7882 ( .B1(n7294), .B2(n13508), .A(n7293), .ZN(n7292) );
  INV_X1 U7883 ( .A(n8086), .ZN(n7294) );
  INV_X1 U7884 ( .A(n11190), .ZN(n7293) );
  NOR2_X1 U7885 ( .A1(n13355), .A2(n13352), .ZN(n6877) );
  NOR2_X1 U7886 ( .A1(n8073), .A2(n7311), .ZN(n7310) );
  INV_X1 U7887 ( .A(n13318), .ZN(n7311) );
  NAND2_X1 U7888 ( .A1(n7943), .A2(n6918), .ZN(n6917) );
  NOR2_X1 U7889 ( .A1(n6919), .A2(n7956), .ZN(n6918) );
  INV_X1 U7890 ( .A(n7942), .ZN(n6919) );
  INV_X1 U7891 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7008) );
  INV_X1 U7892 ( .A(n7908), .ZN(n7079) );
  NAND2_X1 U7893 ( .A1(n7876), .A2(n7905), .ZN(n7081) );
  OAI21_X1 U7894 ( .B1(n7874), .B2(n9866), .A(n7873), .ZN(n6914) );
  NAND2_X1 U7895 ( .A1(n7801), .A2(n7800), .ZN(n7054) );
  NAND2_X1 U7896 ( .A1(n7799), .A2(n7550), .ZN(n7801) );
  AND2_X1 U7897 ( .A1(n7800), .A2(SI_14_), .ZN(n7060) );
  INV_X1 U7898 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n15289) );
  NOR2_X1 U7899 ( .A1(n7730), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U7900 ( .A1(n7700), .A2(n7699), .ZN(n7711) );
  AND2_X1 U7901 ( .A1(n14053), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7222) );
  XNOR2_X1 U7902 ( .A(n14058), .B(n14057), .ZN(n14095) );
  AOI21_X1 U7903 ( .B1(n7515), .B2(n9400), .A(n6661), .ZN(n7512) );
  NAND2_X1 U7904 ( .A1(n7517), .A2(n9401), .ZN(n7513) );
  AND2_X1 U7905 ( .A1(n9402), .A2(n7516), .ZN(n7515) );
  NAND2_X1 U7906 ( .A1(n7517), .A2(n9401), .ZN(n7516) );
  AND2_X1 U7907 ( .A1(n11656), .A2(n9392), .ZN(n11686) );
  INV_X1 U7908 ( .A(n11850), .ZN(n11125) );
  INV_X1 U7909 ( .A(n11979), .ZN(n11126) );
  INV_X1 U7910 ( .A(n11719), .ZN(n7520) );
  NAND2_X1 U7911 ( .A1(n9335), .A2(n9334), .ZN(n7521) );
  OR2_X1 U7912 ( .A1(n11676), .A2(n11675), .ZN(n7522) );
  OR2_X1 U7913 ( .A1(n8707), .A2(n12082), .ZN(n11953) );
  OR2_X1 U7914 ( .A1(n10836), .A2(n8737), .ZN(n9446) );
  AND2_X1 U7915 ( .A1(n10273), .A2(n10374), .ZN(n7148) );
  AOI22_X1 U7916 ( .A1(n7145), .A2(n7143), .B1(n7142), .B2(n7144), .ZN(n7141)
         );
  NAND2_X1 U7917 ( .A1(n7138), .A2(n7145), .ZN(n7140) );
  OR2_X1 U7918 ( .A1(n6610), .A2(n14852), .ZN(n7170) );
  OR2_X1 U7919 ( .A1(n11984), .A2(n6711), .ZN(n7168) );
  AND3_X1 U7920 ( .A1(n7150), .A2(n7151), .A3(n6717), .ZN(n11987) );
  NAND2_X1 U7921 ( .A1(n14243), .A2(n14244), .ZN(n14242) );
  OAI21_X1 U7922 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n7089) );
  INV_X1 U7923 ( .A(n7098), .ZN(n7090) );
  OAI21_X1 U7924 ( .B1(n7097), .B2(n12114), .A(n7099), .ZN(n7087) );
  INV_X1 U7925 ( .A(n7100), .ZN(n7096) );
  NAND2_X1 U7926 ( .A1(n8601), .A2(n11690), .ZN(n8617) );
  INV_X1 U7927 ( .A(n8602), .ZN(n8601) );
  OR2_X1 U7928 ( .A1(n11916), .A2(n11917), .ZN(n12151) );
  NAND2_X1 U7929 ( .A1(n6678), .A2(n7110), .ZN(n7107) );
  NAND2_X1 U7930 ( .A1(n8535), .A2(n11975), .ZN(n8536) );
  NAND2_X1 U7931 ( .A1(n8493), .A2(n8765), .ZN(n12233) );
  OR2_X1 U7932 ( .A1(n12309), .A2(n12223), .ZN(n12236) );
  NAND2_X1 U7933 ( .A1(n8702), .A2(n11948), .ZN(n12252) );
  INV_X1 U7934 ( .A(n14977), .ZN(n12254) );
  AND2_X1 U7935 ( .A1(n8418), .A2(n7120), .ZN(n7119) );
  AOI21_X1 U7936 ( .B1(n11784), .B2(n7261), .A(n7260), .ZN(n7259) );
  INV_X1 U7937 ( .A(n11857), .ZN(n7260) );
  INV_X1 U7938 ( .A(n8758), .ZN(n7261) );
  NAND2_X1 U7939 ( .A1(n10972), .A2(n11854), .ZN(n10971) );
  NAND2_X1 U7940 ( .A1(n14963), .A2(n14966), .ZN(n14962) );
  NAND2_X1 U7941 ( .A1(n10585), .A2(n10584), .ZN(n10588) );
  NOR2_X1 U7942 ( .A1(n7127), .A2(n7126), .ZN(n7125) );
  INV_X1 U7943 ( .A(n8705), .ZN(n7126) );
  INV_X1 U7944 ( .A(n6633), .ZN(n7127) );
  AOI21_X1 U7945 ( .B1(n7274), .B2(n12140), .A(n7272), .ZN(n7271) );
  INV_X1 U7946 ( .A(n11927), .ZN(n7272) );
  OR2_X1 U7947 ( .A1(n12141), .A2(n12140), .ZN(n12143) );
  OR2_X1 U7948 ( .A1(n11792), .A2(n6625), .ZN(n12162) );
  OR2_X1 U7949 ( .A1(n12173), .A2(n12176), .ZN(n12175) );
  NOR2_X1 U7950 ( .A1(n12202), .A2(n7269), .ZN(n7268) );
  AND2_X1 U7951 ( .A1(n8463), .A2(n8464), .ZN(n11788) );
  AND2_X1 U7952 ( .A1(n9446), .A2(n15075), .ZN(n10238) );
  OR2_X1 U7953 ( .A1(n9404), .A2(n10581), .ZN(n9432) );
  AND2_X1 U7954 ( .A1(n8563), .A2(n8553), .ZN(n8561) );
  AND2_X1 U7955 ( .A1(n8552), .A2(n8541), .ZN(n8550) );
  NAND2_X1 U7956 ( .A1(n8540), .A2(n8539), .ZN(n8551) );
  AND2_X1 U7957 ( .A1(n7265), .A2(n8163), .ZN(n7264) );
  NAND2_X1 U7958 ( .A1(n8204), .A2(n8203), .ZN(n8413) );
  AND2_X1 U7959 ( .A1(n7507), .A2(n7506), .ZN(n7503) );
  NOR2_X1 U7960 ( .A1(n8346), .A2(n6965), .ZN(n6964) );
  INV_X1 U7961 ( .A(n8198), .ZN(n6965) );
  NAND2_X1 U7962 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n6963), .ZN(n6962) );
  INV_X1 U7963 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8194) );
  XNOR2_X1 U7964 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8305) );
  OR2_X1 U7965 ( .A1(n9116), .A2(n9115), .ZN(n9118) );
  INV_X1 U7966 ( .A(n12479), .ZN(n7033) );
  NAND2_X1 U7967 ( .A1(n10894), .A2(n9067), .ZN(n10986) );
  XNOR2_X1 U7968 ( .A(n14819), .B(n12433), .ZN(n10888) );
  AND2_X1 U7969 ( .A1(n12778), .A2(n12767), .ZN(n9534) );
  NAND2_X1 U7970 ( .A1(n6908), .A2(n6907), .ZN(n6906) );
  NAND2_X1 U7971 ( .A1(n9567), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6907) );
  AND2_X1 U7972 ( .A1(n6906), .A2(n9568), .ZN(n9585) );
  NAND2_X1 U7973 ( .A1(n14644), .A2(n14645), .ZN(n14643) );
  OR2_X1 U7974 ( .A1(n14661), .A2(n14662), .ZN(n6898) );
  NAND2_X1 U7975 ( .A1(n14683), .A2(n12832), .ZN(n14693) );
  NOR2_X1 U7976 ( .A1(n14694), .A2(n6893), .ZN(n12836) );
  NOR2_X1 U7977 ( .A1(n6894), .A2(n11291), .ZN(n6893) );
  INV_X1 U7978 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12845) );
  NAND2_X1 U7979 ( .A1(n6734), .A2(n12684), .ZN(n12663) );
  AND2_X1 U7980 ( .A1(n12882), .A2(n6890), .ZN(n12855) );
  NOR2_X1 U7981 ( .A1(n12853), .A2(n6891), .ZN(n6890) );
  OR2_X1 U7982 ( .A1(n13059), .A2(n12872), .ZN(n6891) );
  NAND2_X1 U7983 ( .A1(n7051), .A2(n7050), .ZN(n12867) );
  AOI21_X1 U7984 ( .B1(n6609), .B2(n11396), .A(n6592), .ZN(n7050) );
  NAND2_X1 U7985 ( .A1(n11400), .A2(n11399), .ZN(n12861) );
  NAND2_X1 U7986 ( .A1(n13065), .A2(n12692), .ZN(n11399) );
  INV_X1 U7987 ( .A(n7456), .ZN(n7449) );
  NAND2_X1 U7988 ( .A1(n7448), .A2(n7456), .ZN(n7447) );
  INV_X1 U7989 ( .A(n7452), .ZN(n7451) );
  XNOR2_X1 U7990 ( .A(n12888), .B(n12894), .ZN(n12877) );
  OAI22_X1 U7991 ( .A1(n11424), .A2(n7454), .B1(n12785), .B2(n12900), .ZN(
        n7453) );
  INV_X1 U7992 ( .A(n11424), .ZN(n7455) );
  AND2_X1 U7993 ( .A1(n8817), .A2(n8816), .ZN(n12912) );
  NOR2_X2 U7994 ( .A1(n12909), .A2(n12908), .ZN(n12907) );
  NOR2_X1 U7995 ( .A1(n7067), .A2(n7337), .ZN(n7066) );
  NAND2_X1 U7996 ( .A1(n12964), .A2(n7071), .ZN(n7070) );
  NAND2_X1 U7997 ( .A1(n6776), .A2(n11419), .ZN(n7434) );
  NAND2_X1 U7998 ( .A1(n7434), .A2(n7433), .ZN(n12957) );
  AND2_X1 U7999 ( .A1(n12961), .A2(n6612), .ZN(n7433) );
  NAND2_X1 U8000 ( .A1(n11391), .A2(n11390), .ZN(n12973) );
  AND2_X1 U8001 ( .A1(n11418), .A2(n11417), .ZN(n12996) );
  OR2_X1 U8002 ( .A1(n10723), .A2(n12661), .ZN(n8840) );
  AOI21_X1 U8003 ( .B1(n7045), .B2(n7044), .A(n6640), .ZN(n7043) );
  INV_X1 U8004 ( .A(n6615), .ZN(n7044) );
  NAND2_X1 U8005 ( .A1(n11152), .A2(n7463), .ZN(n7462) );
  NAND2_X1 U8006 ( .A1(n7462), .A2(n7460), .ZN(n11283) );
  NAND2_X1 U8007 ( .A1(n9071), .A2(n9070), .ZN(n12594) );
  NAND2_X1 U8008 ( .A1(n11021), .A2(n11020), .ZN(n11149) );
  NAND2_X1 U8009 ( .A1(n11000), .A2(n7465), .ZN(n11021) );
  NOR2_X1 U8010 ( .A1(n7467), .A2(n7466), .ZN(n7465) );
  INV_X1 U8011 ( .A(n10999), .ZN(n7466) );
  OR2_X1 U8012 ( .A1(n10845), .A2(n12742), .ZN(n11000) );
  OAI21_X1 U8013 ( .B1(n10607), .B2(n7440), .A(n7438), .ZN(n10691) );
  INV_X1 U8014 ( .A(n7441), .ZN(n7440) );
  AOI21_X1 U8015 ( .B1(n7441), .B2(n7439), .A(n6647), .ZN(n7438) );
  NOR2_X1 U8016 ( .A1(n10687), .A2(n7442), .ZN(n7441) );
  AND2_X1 U8017 ( .A1(n12737), .A2(n10600), .ZN(n7073) );
  NAND2_X1 U8018 ( .A1(n10634), .A2(n10633), .ZN(n7074) );
  NAND2_X1 U8019 ( .A1(n6559), .A2(n9279), .ZN(n8877) );
  NAND2_X1 U8020 ( .A1(n10423), .A2(n12730), .ZN(n10432) );
  XNOR2_X1 U8021 ( .A(n12801), .B(n12511), .ZN(n12529) );
  INV_X1 U8022 ( .A(n13006), .ZN(n13030) );
  XNOR2_X1 U8023 ( .A(n12802), .B(n6589), .ZN(n12727) );
  OR2_X1 U8024 ( .A1(n12778), .A2(n12767), .ZN(n9730) );
  NAND2_X1 U8025 ( .A1(n9157), .A2(n9156), .ZN(n13105) );
  NAND2_X1 U8026 ( .A1(n12764), .A2(n9279), .ZN(n14797) );
  INV_X1 U8027 ( .A(n7470), .ZN(n7468) );
  NOR2_X1 U8028 ( .A1(n9248), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U8029 ( .A1(n7406), .A2(n7409), .ZN(n7405) );
  NAND2_X1 U8030 ( .A1(n8822), .A2(n8805), .ZN(n7404) );
  NOR2_X1 U8031 ( .A1(n8822), .A2(n8805), .ZN(n7406) );
  AND2_X1 U8032 ( .A1(n8797), .A2(n7417), .ZN(n7416) );
  NAND2_X1 U8033 ( .A1(n6844), .A2(n6846), .ZN(n6840) );
  NOR2_X1 U8034 ( .A1(n6842), .A2(n7484), .ZN(n6841) );
  INV_X1 U8035 ( .A(n6844), .ZN(n6842) );
  NAND2_X1 U8036 ( .A1(n6848), .A2(n6622), .ZN(n6847) );
  INV_X1 U8037 ( .A(n6851), .ZN(n6848) );
  NAND2_X1 U8038 ( .A1(n9881), .A2(n6616), .ZN(n9957) );
  INV_X1 U8039 ( .A(n9885), .ZN(n9882) );
  NAND2_X1 U8040 ( .A1(n13280), .A2(n7483), .ZN(n7482) );
  NAND2_X1 U8041 ( .A1(n10792), .A2(n6854), .ZN(n6853) );
  INV_X1 U8042 ( .A(n10794), .ZN(n6854) );
  NAND2_X1 U8043 ( .A1(n14357), .A2(n11489), .ZN(n13225) );
  NAND2_X1 U8044 ( .A1(n13241), .A2(n6644), .ZN(n13206) );
  AND2_X1 U8045 ( .A1(n6834), .A2(n7496), .ZN(n6833) );
  OR2_X1 U8046 ( .A1(n11470), .A2(n7544), .ZN(n7496) );
  AND4_X1 U8047 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n13430)
         );
  AND4_X1 U8048 ( .A1(n7618), .A2(n7617), .A3(n7616), .A4(n7615), .ZN(n9877)
         );
  OR2_X1 U8049 ( .A1(n13442), .A2(n7586), .ZN(n7589) );
  NAND2_X1 U8050 ( .A1(n6815), .A2(n6814), .ZN(n6813) );
  NAND2_X1 U8051 ( .A1(n13626), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8052 ( .A1(n6813), .A2(n6812), .ZN(n6811) );
  INV_X1 U8053 ( .A(n9636), .ZN(n6812) );
  NOR2_X1 U8054 ( .A1(n14420), .A2(n6706), .ZN(n14435) );
  NOR2_X1 U8055 ( .A1(n14433), .A2(n6809), .ZN(n13668) );
  AND2_X1 U8056 ( .A1(n13667), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6809) );
  INV_X1 U8057 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13681) );
  NAND2_X1 U8058 ( .A1(n13759), .A2(n7319), .ZN(n13747) );
  NOR2_X1 U8059 ( .A1(n13744), .A2(n7320), .ZN(n7319) );
  INV_X1 U8060 ( .A(n8099), .ZN(n7320) );
  INV_X1 U8061 ( .A(n13516), .ZN(n13744) );
  NAND2_X1 U8062 ( .A1(n8097), .A2(n7951), .ZN(n13795) );
  AOI21_X1 U8063 ( .B1(n7323), .B2(n13840), .A(n7322), .ZN(n7321) );
  INV_X1 U8064 ( .A(n13807), .ZN(n7322) );
  NAND2_X1 U8065 ( .A1(n6945), .A2(n7357), .ZN(n6941) );
  NAND2_X1 U8066 ( .A1(n6984), .A2(n7843), .ZN(n6945) );
  NAND2_X1 U8067 ( .A1(n11185), .A2(n7357), .ZN(n6942) );
  NAND2_X1 U8068 ( .A1(n11187), .A2(n7360), .ZN(n11093) );
  NAND2_X1 U8069 ( .A1(n6944), .A2(n6984), .ZN(n11187) );
  INV_X1 U8070 ( .A(n11185), .ZN(n6944) );
  NAND2_X1 U8071 ( .A1(n7313), .A2(n7312), .ZN(n10801) );
  AOI21_X1 U8072 ( .B1(n13504), .B2(n8083), .A(n10813), .ZN(n7312) );
  NAND2_X1 U8073 ( .A1(n10166), .A2(n13500), .ZN(n7295) );
  NAND2_X1 U8074 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  NAND2_X1 U8075 ( .A1(n8072), .A2(n7310), .ZN(n7309) );
  OR2_X1 U8076 ( .A1(n10080), .A2(n10079), .ZN(n13707) );
  NAND2_X1 U8077 ( .A1(n13456), .A2(n13455), .ZN(n13905) );
  AND2_X1 U8078 ( .A1(n14050), .A2(n9506), .ZN(n13946) );
  NAND2_X1 U8079 ( .A1(n7853), .A2(n7852), .ZN(n13988) );
  NAND2_X1 U8080 ( .A1(n10089), .A2(n8151), .ZN(n14549) );
  AND2_X1 U8081 ( .A1(n11340), .A2(n14553), .ZN(n13991) );
  NOR2_X1 U8082 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7502) );
  NAND2_X1 U8083 ( .A1(n6917), .A2(n6915), .ZN(n7969) );
  NOR2_X1 U8084 ( .A1(n6916), .A2(n7958), .ZN(n6915) );
  INV_X1 U8085 ( .A(n7955), .ZN(n6916) );
  NAND2_X1 U8086 ( .A1(n7566), .A2(n6618), .ZN(n8066) );
  NOR2_X1 U8087 ( .A1(n8057), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n8062) );
  INV_X1 U8088 ( .A(n7081), .ZN(n7076) );
  OR2_X1 U8089 ( .A1(n7911), .A2(n9972), .ZN(n7891) );
  NAND2_X1 U8090 ( .A1(n7327), .A2(n7330), .ZN(n7779) );
  OR2_X1 U8091 ( .A1(n7743), .A2(n7332), .ZN(n7327) );
  NAND2_X1 U8092 ( .A1(n6871), .A2(n7745), .ZN(n7763) );
  NAND2_X1 U8093 ( .A1(n7743), .A2(n7742), .ZN(n6871) );
  XNOR2_X1 U8094 ( .A(n7681), .B(n7680), .ZN(n9494) );
  NAND2_X1 U8095 ( .A1(n6868), .A2(n7667), .ZN(n7681) );
  NAND2_X1 U8096 ( .A1(n7665), .A2(n7664), .ZN(n6868) );
  NAND2_X1 U8097 ( .A1(n7175), .A2(n7607), .ZN(n7624) );
  NOR2_X1 U8098 ( .A1(n14070), .A2(n14069), .ZN(n14129) );
  NOR2_X1 U8099 ( .A1(n15151), .A2(n14094), .ZN(n14069) );
  AOI21_X1 U8100 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14075), .A(n14074), .ZN(
        n14136) );
  AOI22_X1 U8101 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14428), .B1(n14090), 
        .B2(n14079), .ZN(n14089) );
  OAI21_X1 U8102 ( .B1(n14174), .B2(n14175), .A(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n7217) );
  NAND2_X1 U8103 ( .A1(n8588), .A2(n8587), .ZN(n12281) );
  OR2_X1 U8104 ( .A1(n11764), .A2(n15288), .ZN(n8587) );
  AND3_X1 U8105 ( .A1(n8403), .A2(n8402), .A3(n8401), .ZN(n11627) );
  AND3_X1 U8106 ( .A1(n8549), .A2(n8548), .A3(n8547), .ZN(n12166) );
  OR2_X1 U8107 ( .A1(n9328), .A2(n10520), .ZN(n9329) );
  OR2_X1 U8108 ( .A1(n8277), .A2(SI_2_), .ZN(n8260) );
  OR2_X1 U8109 ( .A1(n8698), .A2(n10343), .ZN(n8261) );
  INV_X1 U8110 ( .A(n11976), .ZN(n12240) );
  NAND2_X1 U8111 ( .A1(n8336), .A2(n8335), .ZN(n14960) );
  INV_X1 U8112 ( .A(n8334), .ZN(n8335) );
  OAI21_X1 U8113 ( .B1(n8277), .B2(n9460), .A(n8333), .ZN(n8334) );
  INV_X1 U8114 ( .A(n11733), .ZN(n11740) );
  INV_X1 U8115 ( .A(n12252), .ZN(n14980) );
  OAI211_X1 U8116 ( .C1(n10661), .C2(n12372), .A(n8560), .B(n8559), .ZN(n11974) );
  INV_X1 U8117 ( .A(n12166), .ZN(n12192) );
  OR2_X1 U8118 ( .A1(n11764), .A2(n10410), .ZN(n8554) );
  NAND2_X1 U8119 ( .A1(n8509), .A2(n8508), .ZN(n12300) );
  NAND2_X1 U8120 ( .A1(n8230), .A2(n8229), .ZN(n12303) );
  NAND2_X1 U8121 ( .A1(n8472), .A2(n8471), .ZN(n12313) );
  AND3_X1 U8122 ( .A1(n8351), .A2(n8350), .A3(n8349), .ZN(n15042) );
  NAND2_X1 U8123 ( .A1(n9188), .A2(n9187), .ZN(n13094) );
  NAND2_X1 U8124 ( .A1(n9137), .A2(n9136), .ZN(n13114) );
  NAND2_X1 U8125 ( .A1(n8848), .A2(n8847), .ZN(n12618) );
  NAND2_X1 U8126 ( .A1(n9203), .A2(n9202), .ZN(n13089) );
  AOI21_X1 U8127 ( .B1(n7413), .B2(n7415), .A(n6724), .ZN(n7411) );
  INV_X1 U8128 ( .A(n8995), .ZN(n7415) );
  NAND2_X1 U8129 ( .A1(n7020), .A2(n7392), .ZN(n6872) );
  AND2_X1 U8130 ( .A1(n11298), .A2(n12420), .ZN(n6873) );
  INV_X1 U8131 ( .A(n12422), .ZN(n7392) );
  NAND2_X1 U8132 ( .A1(n9098), .A2(n9097), .ZN(n13137) );
  INV_X1 U8133 ( .A(n12912), .ZN(n12785) );
  NAND2_X1 U8134 ( .A1(n9211), .A2(n9210), .ZN(n12944) );
  OR2_X1 U8135 ( .A1(n8872), .A2(n9850), .ZN(n8873) );
  AND2_X1 U8136 ( .A1(n8875), .A2(n8876), .ZN(n6750) );
  AND2_X1 U8137 ( .A1(n9543), .A2(n6777), .ZN(n14655) );
  INV_X1 U8138 ( .A(n12853), .ZN(n13057) );
  NAND2_X1 U8139 ( .A1(n9114), .A2(n9113), .ZN(n14327) );
  INV_X1 U8140 ( .A(n6780), .ZN(n6779) );
  OAI21_X1 U8141 ( .B1(n13063), .B2(n13140), .A(n6925), .ZN(n6780) );
  NOR2_X1 U8142 ( .A1(n7470), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7469) );
  INV_X1 U8143 ( .A(n7408), .ZN(n8833) );
  AOI21_X1 U8144 ( .B1(n8837), .B2(P2_IR_REG_31__SCAN_IN), .A(n7409), .ZN(
        n7408) );
  INV_X1 U8145 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10713) );
  NOR2_X1 U8146 ( .A1(n14044), .A2(n14048), .ZN(n6818) );
  NAND2_X1 U8147 ( .A1(n7962), .A2(n7961), .ZN(n13939) );
  NAND2_X1 U8148 ( .A1(n6816), .A2(n7471), .ZN(n13197) );
  AOI21_X1 U8149 ( .B1(n7473), .B2(n7474), .A(n7472), .ZN(n7471) );
  NAND2_X1 U8150 ( .A1(n13225), .A2(n7473), .ZN(n6816) );
  INV_X1 U8151 ( .A(n13198), .ZN(n7472) );
  OR2_X1 U8152 ( .A1(n13444), .A2(n9525), .ZN(n7597) );
  NAND2_X1 U8153 ( .A1(n7935), .A2(n7934), .ZN(n13950) );
  AND2_X1 U8154 ( .A1(n7920), .A2(n7919), .ZN(n13831) );
  OR2_X1 U8155 ( .A1(n11592), .A2(n13444), .ZN(n7920) );
  INV_X1 U8156 ( .A(n13946), .ZN(n13268) );
  OR2_X1 U8157 ( .A1(n10723), .A2(n13444), .ZN(n7884) );
  NAND2_X1 U8158 ( .A1(n8006), .A2(n8005), .ZN(n13729) );
  INV_X1 U8159 ( .A(n14384), .ZN(n13296) );
  NAND2_X1 U8160 ( .A1(n13491), .A2(n13490), .ZN(n13540) );
  OR2_X1 U8161 ( .A1(n13491), .A2(n13488), .ZN(n13541) );
  NAND2_X1 U8162 ( .A1(n9691), .A2(n9868), .ZN(n13543) );
  INV_X1 U8163 ( .A(n9877), .ZN(n13572) );
  INV_X1 U8164 ( .A(n9750), .ZN(n7486) );
  AOI21_X1 U8165 ( .B1(n14425), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14417), .ZN(
        n14431) );
  AOI21_X1 U8166 ( .B1(n13676), .B2(n14483), .A(n14493), .ZN(n6799) );
  OAI21_X1 U8167 ( .B1(n13681), .B2(n14499), .A(n13680), .ZN(n6797) );
  OR2_X1 U8168 ( .A1(n8056), .A2(n13695), .ZN(n13724) );
  AOI21_X1 U8169 ( .B1(n8118), .B2(n14585), .A(n11570), .ZN(n13715) );
  AND2_X1 U8170 ( .A1(n6693), .A2(n11337), .ZN(n13918) );
  NAND2_X1 U8171 ( .A1(n7353), .A2(n10082), .ZN(n10125) );
  NAND2_X1 U8172 ( .A1(n7354), .A2(n10083), .ZN(n7353) );
  NAND2_X1 U8173 ( .A1(n7583), .A2(n6760), .ZN(n7288) );
  NOR2_X1 U8174 ( .A1(n7501), .A2(n14033), .ZN(n6760) );
  NAND2_X1 U8175 ( .A1(n8122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8060) );
  INV_X1 U8176 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10724) );
  OAI21_X1 U8177 ( .B1(n14404), .B2(n14403), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n7216) );
  NOR2_X1 U8178 ( .A1(n14407), .A2(n14408), .ZN(n14406) );
  NAND2_X1 U8179 ( .A1(n6731), .A2(n7192), .ZN(n12552) );
  NAND2_X1 U8180 ( .A1(n12548), .A2(n12546), .ZN(n7192) );
  NAND2_X1 U8181 ( .A1(n7196), .A2(n12559), .ZN(n7195) );
  INV_X1 U8182 ( .A(n12570), .ZN(n7211) );
  NAND2_X1 U8183 ( .A1(n6673), .A2(n6563), .ZN(n6988) );
  NAND2_X1 U8184 ( .A1(n13310), .A2(n13485), .ZN(n6987) );
  NAND2_X1 U8185 ( .A1(n6999), .A2(n6998), .ZN(n6997) );
  INV_X1 U8186 ( .A(n13324), .ZN(n6998) );
  NAND2_X1 U8187 ( .A1(n7375), .A2(n13320), .ZN(n13325) );
  NAND2_X1 U8188 ( .A1(n13323), .A2(n13324), .ZN(n7001) );
  AND2_X1 U8189 ( .A1(n6997), .A2(n13327), .ZN(n6996) );
  NAND2_X1 U8190 ( .A1(n13332), .A2(n7381), .ZN(n7380) );
  NAND2_X1 U8191 ( .A1(n6996), .A2(n7000), .ZN(n6993) );
  INV_X1 U8192 ( .A(n7001), .ZN(n7000) );
  NAND2_X1 U8193 ( .A1(n13343), .A2(n7378), .ZN(n7377) );
  NAND2_X1 U8194 ( .A1(n7176), .A2(n6743), .ZN(n6742) );
  NAND2_X1 U8195 ( .A1(n13354), .A2(n7387), .ZN(n7386) );
  NAND2_X1 U8196 ( .A1(n12626), .A2(n12625), .ZN(n12629) );
  AND2_X1 U8197 ( .A1(n7207), .A2(n12628), .ZN(n7206) );
  INV_X1 U8198 ( .A(n12627), .ZN(n7207) );
  AND2_X1 U8199 ( .A1(n6979), .A2(n6977), .ZN(n13385) );
  AOI22_X1 U8200 ( .A1(n13371), .A2(n6978), .B1(n13376), .B2(n6983), .ZN(n6977) );
  NOR2_X1 U8201 ( .A1(n6984), .A2(n6982), .ZN(n6981) );
  AND2_X1 U8202 ( .A1(n7018), .A2(n7017), .ZN(n7016) );
  NAND2_X1 U8203 ( .A1(n13396), .A2(n6630), .ZN(n7017) );
  INV_X1 U8204 ( .A(n13395), .ZN(n7018) );
  NAND2_X1 U8205 ( .A1(n7200), .A2(n6637), .ZN(n12633) );
  NOR2_X1 U8206 ( .A1(n13401), .A2(n13402), .ZN(n7372) );
  INV_X1 U8207 ( .A(n7011), .ZN(n7010) );
  OAI21_X1 U8208 ( .B1(n7014), .B2(n7012), .A(n7373), .ZN(n7011) );
  OAI21_X1 U8209 ( .B1(n13411), .B2(n7366), .A(n7365), .ZN(n13415) );
  NAND2_X1 U8210 ( .A1(n13413), .A2(n13410), .ZN(n7365) );
  AND2_X1 U8211 ( .A1(n13412), .A2(n7367), .ZN(n7366) );
  INV_X1 U8212 ( .A(n13414), .ZN(n6976) );
  INV_X1 U8213 ( .A(n7302), .ZN(n7300) );
  AND2_X1 U8214 ( .A1(n10673), .A2(n7161), .ZN(n7157) );
  NAND2_X1 U8215 ( .A1(n10675), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7161) );
  INV_X1 U8216 ( .A(n14960), .ZN(n9314) );
  INV_X1 U8217 ( .A(n10393), .ZN(n9317) );
  NOR2_X1 U8218 ( .A1(n12653), .A2(n7184), .ZN(n7183) );
  NAND2_X1 U8219 ( .A1(n6679), .A2(n7189), .ZN(n7187) );
  NAND2_X1 U8220 ( .A1(n12656), .A2(n12657), .ZN(n7191) );
  NOR2_X1 U8221 ( .A1(n7184), .A2(n7186), .ZN(n7185) );
  INV_X1 U8222 ( .A(n12650), .ZN(n7186) );
  NOR2_X1 U8223 ( .A1(n10699), .A2(n14803), .ZN(n6883) );
  AOI22_X1 U8224 ( .A1(n7005), .A2(n6596), .B1(n7007), .B2(n13427), .ZN(n7004)
         );
  INV_X1 U8225 ( .A(n7713), .ZN(n6923) );
  INV_X1 U8226 ( .A(n9377), .ZN(n7528) );
  AOI21_X1 U8227 ( .B1(n7526), .B2(n7525), .A(n7524), .ZN(n7523) );
  INV_X1 U8228 ( .A(n9379), .ZN(n7524) );
  INV_X1 U8229 ( .A(n11695), .ZN(n7525) );
  NAND2_X1 U8230 ( .A1(n11772), .A2(n10182), .ZN(n9310) );
  OAI21_X1 U8231 ( .B1(n12027), .B2(n15274), .A(n14889), .ZN(n12003) );
  OAI21_X1 U8232 ( .B1(n12045), .B2(n12310), .A(n14202), .ZN(n12009) );
  NOR2_X1 U8233 ( .A1(n7098), .A2(n7095), .ZN(n7094) );
  NAND2_X1 U8234 ( .A1(n7099), .A2(n12114), .ZN(n7095) );
  AND2_X1 U8235 ( .A1(n7097), .A2(n7099), .ZN(n7091) );
  NAND2_X1 U8236 ( .A1(n8647), .A2(n8646), .ZN(n8666) );
  INV_X1 U8237 ( .A(n7107), .ZN(n7106) );
  NAND2_X1 U8238 ( .A1(n8557), .A2(n8556), .ZN(n8572) );
  AND2_X1 U8239 ( .A1(n8545), .A2(n8544), .ZN(n8557) );
  AND2_X1 U8240 ( .A1(n8488), .A2(n11669), .ZN(n8177) );
  NAND2_X1 U8241 ( .A1(n8177), .A2(n11368), .ZN(n8510) );
  NOR2_X1 U8242 ( .A1(n8473), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8488) );
  OR2_X1 U8243 ( .A1(n8457), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U8244 ( .A1(n8442), .A2(n11273), .ZN(n8457) );
  NOR2_X1 U8245 ( .A1(n7122), .A2(n11784), .ZN(n7118) );
  INV_X1 U8246 ( .A(n8417), .ZN(n7122) );
  NAND2_X1 U8247 ( .A1(n8417), .A2(n7121), .ZN(n7120) );
  INV_X1 U8248 ( .A(n8404), .ZN(n7121) );
  AND3_X1 U8249 ( .A1(n8384), .A2(n8383), .A3(n8382), .ZN(n11850) );
  AOI21_X1 U8250 ( .B1(n11836), .B2(n7245), .A(n7244), .ZN(n7243) );
  INV_X1 U8251 ( .A(n11834), .ZN(n7245) );
  NAND2_X1 U8252 ( .A1(n10393), .A2(n8254), .ZN(n11809) );
  NAND2_X1 U8253 ( .A1(n11772), .A2(n11966), .ZN(n11911) );
  NOR2_X1 U8254 ( .A1(n7233), .A2(n7229), .ZN(n7228) );
  AND2_X1 U8255 ( .A1(n8170), .A2(n8221), .ZN(n8218) );
  INV_X1 U8256 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U8257 ( .A1(n8419), .A2(n8206), .ZN(n8207) );
  NAND2_X1 U8258 ( .A1(n8207), .A2(n9828), .ZN(n8208) );
  INV_X1 U8259 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U8260 ( .A1(n6769), .A2(n12706), .ZN(n12709) );
  INV_X1 U8261 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7436) );
  OR2_X1 U8262 ( .A1(n8872), .A2(n9551), .ZN(n8862) );
  AND2_X1 U8263 ( .A1(n9232), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9292) );
  OAI21_X1 U8264 ( .B1(n7453), .B2(n7455), .A(n12877), .ZN(n7452) );
  INV_X1 U8265 ( .A(n7453), .ZN(n7448) );
  AND2_X1 U8266 ( .A1(n13084), .A2(n12928), .ZN(n11423) );
  INV_X1 U8267 ( .A(n7071), .ZN(n7067) );
  AND2_X1 U8268 ( .A1(n13089), .A2(n12944), .ZN(n7337) );
  NAND2_X1 U8269 ( .A1(n13094), .A2(n12927), .ZN(n11421) );
  NAND2_X1 U8270 ( .A1(n11420), .A2(n7429), .ZN(n7428) );
  INV_X1 U8271 ( .A(n6612), .ZN(n7429) );
  NOR2_X1 U8272 ( .A1(n7432), .A2(n7431), .ZN(n7430) );
  INV_X1 U8273 ( .A(n11419), .ZN(n7431) );
  NOR2_X1 U8274 ( .A1(n12990), .A2(n13105), .ZN(n6886) );
  NOR2_X1 U8275 ( .A1(n6888), .A2(n14327), .ZN(n6887) );
  INV_X1 U8276 ( .A(n6889), .ZN(n6888) );
  NOR2_X1 U8277 ( .A1(n12599), .A2(n13137), .ZN(n6889) );
  AND2_X1 U8278 ( .A1(n9002), .A2(n8780), .ZN(n9037) );
  NOR2_X1 U8279 ( .A1(n9004), .A2(n9003), .ZN(n9002) );
  INV_X1 U8280 ( .A(n7446), .ZN(n7442) );
  NOR2_X1 U8281 ( .A1(n10609), .A2(n7445), .ZN(n7444) );
  INV_X1 U8282 ( .A(n10606), .ZN(n7445) );
  NAND2_X1 U8283 ( .A1(n12805), .A2(n10025), .ZN(n12520) );
  NAND2_X1 U8284 ( .A1(n10020), .A2(n10024), .ZN(n12515) );
  NAND2_X1 U8285 ( .A1(n12900), .A2(n12912), .ZN(n7335) );
  NOR2_X1 U8286 ( .A1(n12937), .A2(n7069), .ZN(n7068) );
  INV_X1 U8287 ( .A(n12756), .ZN(n7069) );
  INV_X1 U8288 ( .A(n6883), .ZN(n10767) );
  OR2_X1 U8289 ( .A1(n8998), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9014) );
  AND2_X1 U8290 ( .A1(n6622), .A2(n10206), .ZN(n6850) );
  INV_X1 U8291 ( .A(n11545), .ZN(n7483) );
  NOR2_X1 U8292 ( .A1(n7544), .A2(n7498), .ZN(n7497) );
  OR2_X1 U8293 ( .A1(n7490), .A2(n6836), .ZN(n6835) );
  INV_X1 U8294 ( .A(n13250), .ZN(n7498) );
  NAND2_X1 U8295 ( .A1(n6623), .A2(n6836), .ZN(n6834) );
  OR2_X1 U8296 ( .A1(n13449), .A2(n13450), .ZN(n6969) );
  NAND2_X1 U8297 ( .A1(n13778), .A2(n7316), .ZN(n7315) );
  INV_X1 U8298 ( .A(n8097), .ZN(n7316) );
  NOR2_X1 U8299 ( .A1(n13392), .A2(n6943), .ZN(n6940) );
  INV_X1 U8300 ( .A(n8074), .ZN(n7308) );
  INV_X1 U8301 ( .A(n7310), .ZN(n7305) );
  AND2_X1 U8302 ( .A1(n9750), .A2(n13311), .ZN(n13300) );
  NAND2_X1 U8303 ( .A1(n13981), .A2(n13387), .ZN(n13861) );
  AOI21_X1 U8304 ( .B1(n8145), .B2(n9487), .A(n9485), .ZN(n10078) );
  AND2_X1 U8305 ( .A1(n7862), .A2(n7848), .ZN(n7860) );
  AND2_X1 U8306 ( .A1(n6927), .A2(n7055), .ZN(n6926) );
  AND2_X1 U8307 ( .A1(n7057), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U8308 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  AND2_X1 U8309 ( .A1(n7844), .A2(n7820), .ZN(n7821) );
  INV_X1 U8310 ( .A(n7761), .ZN(n7331) );
  INV_X1 U8311 ( .A(n7333), .ZN(n7332) );
  AOI21_X1 U8312 ( .B1(n6869), .B2(n6870), .A(n6666), .ZN(n6866) );
  OAI21_X1 U8313 ( .B1(n7641), .B2(n7640), .A(n7643), .ZN(n7650) );
  NAND2_X1 U8314 ( .A1(n9469), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7536) );
  INV_X1 U8315 ( .A(n7215), .ZN(n14060) );
  OAI21_X1 U8316 ( .B1(n14095), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6620), .ZN(
        n7215) );
  NOR2_X1 U8317 ( .A1(n14066), .A2(n14067), .ZN(n14068) );
  NOR2_X1 U8318 ( .A1(n14121), .A2(n14122), .ZN(n14066) );
  XNOR2_X1 U8319 ( .A(n14068), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n14094) );
  OAI21_X1 U8320 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14072), .A(n14071), .ZN(
        n14092) );
  AND3_X1 U8321 ( .A1(n8281), .A2(n8280), .A3(n8279), .ZN(n9315) );
  NAND2_X1 U8322 ( .A1(n6585), .A2(n11695), .ZN(n7529) );
  AND2_X1 U8323 ( .A1(n9398), .A2(n9397), .ZN(n11657) );
  NAND2_X1 U8324 ( .A1(n8369), .A2(n15364), .ZN(n8387) );
  INV_X1 U8325 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15364) );
  AOI21_X1 U8326 ( .B1(n9322), .B2(n9394), .A(n6752), .ZN(n9323) );
  INV_X1 U8327 ( .A(n12336), .ZN(n6752) );
  OR2_X1 U8328 ( .A1(n7248), .A2(n11804), .ZN(n6968) );
  AND2_X1 U8329 ( .A1(n7253), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U8330 ( .A1(n11953), .A2(n7250), .ZN(n7249) );
  INV_X1 U8331 ( .A(n11804), .ZN(n7252) );
  AND2_X1 U8332 ( .A1(n11773), .A2(n11769), .ZN(n11956) );
  OAI21_X1 U8333 ( .B1(n10276), .B2(n7144), .A(n7142), .ZN(n10318) );
  AND2_X1 U8334 ( .A1(n7141), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7137) );
  OAI21_X1 U8335 ( .B1(n10312), .B2(n15062), .A(n10541), .ZN(n10353) );
  NAND2_X1 U8336 ( .A1(n6591), .A2(n10322), .ZN(n10351) );
  NAND2_X1 U8337 ( .A1(n11999), .A2(n12000), .ZN(n14856) );
  AND2_X1 U8338 ( .A1(n7168), .A2(n7167), .ZN(n11985) );
  AND2_X1 U8339 ( .A1(n7170), .A2(n6712), .ZN(n7167) );
  INV_X1 U8340 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14898) );
  INV_X1 U8341 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11273) );
  OR2_X1 U8342 ( .A1(n14912), .A2(n14911), .ZN(n14914) );
  OR2_X1 U8343 ( .A1(n14934), .A2(n14935), .ZN(n14931) );
  NOR2_X1 U8344 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  OR2_X1 U8345 ( .A1(n8666), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U8346 ( .A1(n11946), .A2(n11944), .ZN(n12077) );
  OR2_X1 U8347 ( .A1(n11937), .A2(n11936), .ZN(n12100) );
  AND2_X1 U8348 ( .A1(n8623), .A2(n8622), .ZN(n12125) );
  NAND2_X1 U8349 ( .A1(n8526), .A2(n8525), .ZN(n12196) );
  NAND2_X1 U8350 ( .A1(n12303), .A2(n11976), .ZN(n7130) );
  NAND2_X1 U8351 ( .A1(n12233), .A2(n12236), .ZN(n12219) );
  AOI21_X1 U8352 ( .B1(n7114), .B2(n7116), .A(n6651), .ZN(n7113) );
  AOI21_X1 U8353 ( .B1(n6595), .B2(n11854), .A(n7255), .ZN(n7254) );
  INV_X1 U8354 ( .A(n11861), .ZN(n7255) );
  AND2_X1 U8355 ( .A1(n11871), .A2(n11865), .ZN(n14264) );
  OR2_X1 U8356 ( .A1(n8387), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8405) );
  OR2_X1 U8357 ( .A1(n8405), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U8358 ( .A1(n14948), .A2(n6643), .ZN(n10896) );
  INV_X1 U8359 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8354) );
  AND2_X1 U8360 ( .A1(n8355), .A2(n8354), .ZN(n8369) );
  NOR2_X1 U8361 ( .A1(n8339), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U8362 ( .A1(n14967), .A2(n8338), .ZN(n10780) );
  NAND2_X1 U8363 ( .A1(n7085), .A2(n10619), .ZN(n14967) );
  AND2_X1 U8364 ( .A1(n8337), .A2(n8315), .ZN(n7085) );
  NOR2_X1 U8365 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8299) );
  NAND2_X1 U8366 ( .A1(n14976), .A2(n8753), .ZN(n14975) );
  NAND2_X1 U8367 ( .A1(n11819), .A2(n11818), .ZN(n14983) );
  NAND2_X1 U8368 ( .A1(n10048), .A2(n12337), .ZN(n12336) );
  AND2_X1 U8369 ( .A1(n10238), .A2(n15043), .ZN(n10586) );
  AND2_X1 U8370 ( .A1(n8742), .A2(n8741), .ZN(n10585) );
  AOI21_X1 U8371 ( .B1(n7238), .B2(n7237), .A(n6657), .ZN(n7236) );
  OR2_X1 U8372 ( .A1(n12173), .A2(n7239), .ZN(n7235) );
  INV_X1 U8373 ( .A(n14988), .ZN(n15043) );
  NAND2_X1 U8374 ( .A1(n11801), .A2(n11805), .ZN(n14988) );
  INV_X1 U8375 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U8376 ( .A1(n8222), .A2(n8218), .ZN(n8224) );
  NAND2_X1 U8377 ( .A1(n8222), .A2(n8221), .ZN(n8717) );
  NAND2_X1 U8378 ( .A1(n8628), .A2(n8627), .ZN(n8641) );
  NAND2_X1 U8379 ( .A1(n8626), .A2(n8625), .ZN(n8628) );
  NAND2_X1 U8380 ( .A1(n8598), .A2(n8597), .ZN(n8611) );
  XNOR2_X1 U8381 ( .A(n8740), .B(n8739), .ZN(n10240) );
  NAND2_X1 U8382 ( .A1(n8581), .A2(n8580), .ZN(n8585) );
  NAND2_X1 U8383 ( .A1(n8585), .A2(n8584), .ZN(n8598) );
  AOI21_X1 U8384 ( .B1(n6954), .B2(n6956), .A(n6952), .ZN(n6951) );
  INV_X1 U8385 ( .A(n8563), .ZN(n6952) );
  INV_X1 U8386 ( .A(n8688), .ZN(n7532) );
  AND2_X1 U8387 ( .A1(n8539), .A2(n8519), .ZN(n8537) );
  NAND2_X1 U8388 ( .A1(n8495), .A2(n8494), .ZN(n8497) );
  NAND2_X1 U8389 ( .A1(n8216), .A2(n8215), .ZN(n8495) );
  NAND2_X1 U8390 ( .A1(n8482), .A2(n8480), .ZN(n8216) );
  INV_X1 U8391 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8499) );
  AND2_X1 U8392 ( .A1(n8212), .A2(n8211), .ZN(n8465) );
  AND2_X1 U8393 ( .A1(n8210), .A2(n8209), .ZN(n8449) );
  NAND2_X1 U8394 ( .A1(n8208), .A2(n6753), .ZN(n8436) );
  OR2_X1 U8395 ( .A1(n8207), .A2(n9828), .ZN(n6753) );
  AOI21_X1 U8396 ( .B1(n6966), .B2(n6606), .A(n6709), .ZN(n8421) );
  AND2_X1 U8397 ( .A1(n8206), .A2(n8205), .ZN(n8420) );
  INV_X1 U8398 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8162) );
  OR2_X1 U8399 ( .A1(n8364), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8379) );
  AOI21_X1 U8400 ( .B1(n6957), .B2(n6960), .A(n6958), .ZN(n8378) );
  AND2_X1 U8401 ( .A1(n8201), .A2(n8200), .ZN(n8377) );
  OR2_X1 U8402 ( .A1(n8331), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8364) );
  XNOR2_X1 U8403 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8288) );
  AND2_X1 U8404 ( .A1(n8867), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U8405 ( .A1(n8786), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U8406 ( .A1(n9133), .A2(n7394), .ZN(n7393) );
  INV_X1 U8407 ( .A(n9134), .ZN(n7394) );
  INV_X1 U8408 ( .A(n9139), .ZN(n8784) );
  OR2_X1 U8409 ( .A1(n7420), .A2(n9081), .ZN(n7418) );
  NAND2_X1 U8410 ( .A1(n7391), .A2(n12420), .ZN(n7020) );
  INV_X1 U8411 ( .A(n7393), .ZN(n7391) );
  OR3_X1 U8412 ( .A1(n9160), .A2(n9159), .A3(n9158), .ZN(n9175) );
  NAND2_X1 U8413 ( .A1(n7390), .A2(n9029), .ZN(n10818) );
  INV_X1 U8414 ( .A(n10882), .ZN(n7390) );
  NAND2_X1 U8415 ( .A1(n8783), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8852) );
  OR2_X1 U8416 ( .A1(n8852), .A2(n8841), .ZN(n9139) );
  NAND2_X1 U8417 ( .A1(n6674), .A2(n6726), .ZN(n6766) );
  AND2_X1 U8418 ( .A1(n6769), .A2(n6677), .ZN(n6726) );
  AND4_X1 U8419 ( .A1(n12861), .A2(n12759), .A3(n12877), .A4(n12901), .ZN(
        n6768) );
  INV_X1 U8420 ( .A(n8917), .ZN(n12670) );
  OR2_X1 U8421 ( .A1(n8902), .A2(n9849), .ZN(n8875) );
  NOR2_X1 U8422 ( .A1(n9718), .A2(n6902), .ZN(n9720) );
  AND2_X1 U8423 ( .A1(n9723), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U8424 ( .A1(n9720), .A2(n9719), .ZN(n9796) );
  NOR2_X1 U8425 ( .A1(n9796), .A2(n6901), .ZN(n9801) );
  AND2_X1 U8426 ( .A1(n9797), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8427 ( .A1(n9801), .A2(n9800), .ZN(n9931) );
  NOR2_X1 U8428 ( .A1(n10928), .A2(n6900), .ZN(n12808) );
  AND2_X1 U8429 ( .A1(n10929), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U8430 ( .A1(n12808), .A2(n12807), .ZN(n12806) );
  NAND2_X1 U8431 ( .A1(n12806), .A2(n6899), .ZN(n14644) );
  OR2_X1 U8432 ( .A1(n12812), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U8433 ( .A1(n6896), .A2(n12820), .ZN(n6895) );
  XNOR2_X1 U8434 ( .A(n12836), .B(n14718), .ZN(n14713) );
  NAND2_X1 U8435 ( .A1(n12687), .A2(n12686), .ZN(n12851) );
  NAND2_X1 U8436 ( .A1(n13084), .A2(n12893), .ZN(n7336) );
  NOR2_X1 U8437 ( .A1(n12946), .A2(n13089), .ZN(n12914) );
  NAND2_X1 U8438 ( .A1(n6886), .A2(n6885), .ZN(n12965) );
  INV_X1 U8439 ( .A(n6884), .ZN(n12946) );
  NOR2_X1 U8440 ( .A1(n12965), .A2(n13094), .ZN(n6884) );
  INV_X1 U8441 ( .A(n6886), .ZN(n12980) );
  AND2_X1 U8442 ( .A1(n11282), .A2(n7463), .ZN(n7459) );
  NAND2_X1 U8443 ( .A1(n7457), .A2(n6641), .ZN(n6790) );
  OAI21_X1 U8444 ( .B1(n11154), .B2(n7040), .A(n7038), .ZN(n11289) );
  INV_X1 U8445 ( .A(n7041), .ZN(n7040) );
  AOI21_X1 U8446 ( .B1(n7041), .B2(n7039), .A(n6653), .ZN(n7038) );
  NAND2_X1 U8447 ( .A1(n11155), .A2(n6889), .ZN(n11256) );
  NAND2_X1 U8448 ( .A1(n11155), .A2(n14333), .ZN(n11258) );
  AND2_X1 U8449 ( .A1(n11030), .A2(n14340), .ZN(n11155) );
  AND2_X1 U8450 ( .A1(n11004), .A2(n11086), .ZN(n11030) );
  NAND2_X1 U8451 ( .A1(n7443), .A2(n7446), .ZN(n10688) );
  NAND2_X1 U8452 ( .A1(n10607), .A2(n7444), .ZN(n7443) );
  NAND2_X1 U8453 ( .A1(n10529), .A2(n10422), .ZN(n10423) );
  INV_X1 U8454 ( .A(n10014), .ZN(n10017) );
  INV_X1 U8455 ( .A(n12805), .ZN(n10020) );
  INV_X1 U8456 ( .A(n13062), .ZN(n6925) );
  NAND2_X1 U8457 ( .A1(n7052), .A2(n6609), .ZN(n13070) );
  AND2_X1 U8458 ( .A1(n7070), .A2(n7068), .ZN(n12936) );
  NAND2_X1 U8459 ( .A1(n9275), .A2(n9277), .ZN(n9248) );
  INV_X1 U8460 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U8461 ( .A1(n7542), .A2(n8818), .ZN(n8824) );
  OAI21_X1 U8462 ( .B1(n8837), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8834) );
  INV_X1 U8463 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n15197) );
  OR2_X1 U8464 ( .A1(n8981), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8998) );
  OR2_X1 U8465 ( .A1(n8946), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8962) );
  OR2_X1 U8466 ( .A1(n9047), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8928) );
  OR2_X1 U8467 ( .A1(n9469), .A2(n6688), .ZN(n8869) );
  OR3_X1 U8468 ( .A1(n7809), .A2(n7808), .A3(n7807), .ZN(n7836) );
  AND2_X1 U8469 ( .A1(n14348), .A2(n14349), .ZN(n11470) );
  AND2_X1 U8470 ( .A1(n6829), .A2(n11523), .ZN(n6828) );
  NAND2_X1 U8471 ( .A1(n13260), .A2(n6830), .ZN(n6829) );
  INV_X1 U8472 ( .A(n13260), .ZN(n6831) );
  NAND2_X1 U8473 ( .A1(n6824), .A2(n9879), .ZN(n9880) );
  OR2_X1 U8474 ( .A1(n7475), .A2(n7555), .ZN(n7473) );
  AND2_X1 U8475 ( .A1(n13270), .A2(n7476), .ZN(n7475) );
  OR2_X1 U8476 ( .A1(n7477), .A2(n13226), .ZN(n7476) );
  NAND2_X1 U8477 ( .A1(n7478), .A2(n11496), .ZN(n7474) );
  INV_X1 U8478 ( .A(n6853), .ZN(n6852) );
  NAND2_X1 U8479 ( .A1(n7772), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7809) );
  NOR2_X1 U8480 ( .A1(n7495), .A2(n7561), .ZN(n7490) );
  INV_X1 U8481 ( .A(n11140), .ZN(n7495) );
  INV_X1 U8482 ( .A(n7992), .ZN(n7993) );
  INV_X1 U8483 ( .A(n7978), .ZN(n7979) );
  AOI21_X1 U8484 ( .B1(n6828), .B2(n6831), .A(n6827), .ZN(n6826) );
  INV_X1 U8485 ( .A(n13190), .ZN(n6827) );
  OR2_X1 U8486 ( .A1(n7721), .A2(n7720), .ZN(n7734) );
  AOI22_X1 U8487 ( .A1(n11554), .A2(n9986), .B1(n9681), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9682) );
  OR2_X1 U8488 ( .A1(n7898), .A2(n7897), .ZN(n7921) );
  NOR2_X1 U8489 ( .A1(n7734), .A2(n7733), .ZN(n7754) );
  NOR2_X1 U8490 ( .A1(n11061), .A2(n7494), .ZN(n7493) );
  INV_X1 U8491 ( .A(n11058), .ZN(n7494) );
  NAND2_X1 U8492 ( .A1(n13225), .A2(n13226), .ZN(n13224) );
  INV_X1 U8493 ( .A(n13542), .ZN(n13864) );
  INV_X1 U8494 ( .A(n13686), .ZN(n13262) );
  AND4_X1 U8495 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n11464)
         );
  AND4_X1 U8496 ( .A1(n7639), .A2(n7638), .A3(n7637), .A4(n7636), .ZN(n13321)
         );
  AND4_X2 U8497 ( .A1(n7603), .A2(n7602), .A3(n7601), .A4(n7600), .ZN(n7611)
         );
  OR2_X1 U8498 ( .A1(n13442), .A2(n7598), .ZN(n7601) );
  OR2_X1 U8499 ( .A1(n9620), .A2(n9619), .ZN(n6803) );
  OR2_X1 U8500 ( .A1(n9675), .A2(n9674), .ZN(n6801) );
  INV_X1 U8501 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15151) );
  AND2_X1 U8502 ( .A1(n6801), .A2(n6800), .ZN(n9818) );
  NAND2_X1 U8503 ( .A1(n9814), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6800) );
  NOR2_X1 U8504 ( .A1(n10066), .A2(n6804), .ZN(n10071) );
  AND2_X1 U8505 ( .A1(n10067), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6804) );
  NOR2_X1 U8506 ( .A1(n10071), .A2(n10070), .ZN(n13633) );
  NAND2_X1 U8507 ( .A1(n13641), .A2(n6746), .ZN(n13643) );
  OR2_X1 U8508 ( .A1(n13642), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6746) );
  NAND2_X1 U8509 ( .A1(n13643), .A2(n13644), .ZN(n13652) );
  NOR2_X1 U8510 ( .A1(n14435), .A2(n14434), .ZN(n14433) );
  NAND2_X1 U8511 ( .A1(n14446), .A2(n6634), .ZN(n6795) );
  AND2_X1 U8512 ( .A1(n14469), .A2(n13672), .ZN(n13673) );
  AND2_X1 U8513 ( .A1(n14465), .A2(n13658), .ZN(n13659) );
  NOR2_X1 U8514 ( .A1(n13701), .A2(n13905), .ZN(n13690) );
  NAND2_X1 U8515 ( .A1(n11342), .A2(n13429), .ZN(n13701) );
  AND2_X1 U8516 ( .A1(n6671), .A2(n7952), .ZN(n7356) );
  INV_X1 U8517 ( .A(n7945), .ZN(n7946) );
  NAND2_X1 U8518 ( .A1(n8093), .A2(n13513), .ZN(n13843) );
  AND2_X1 U8519 ( .A1(n7303), .A2(n8089), .ZN(n7302) );
  INV_X1 U8520 ( .A(n13891), .ZN(n7303) );
  AND2_X1 U8521 ( .A1(n7854), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U8522 ( .A1(n7291), .A2(n7289), .ZN(n11193) );
  AND2_X1 U8523 ( .A1(n13377), .A2(n7290), .ZN(n7289) );
  NAND2_X1 U8524 ( .A1(n7292), .A2(n11078), .ZN(n7290) );
  NAND2_X1 U8525 ( .A1(n10859), .A2(n8086), .ZN(n11068) );
  NAND2_X1 U8526 ( .A1(n11068), .A2(n13508), .ZN(n11191) );
  NAND2_X1 U8527 ( .A1(n10727), .A2(n6761), .ZN(n11189) );
  NOR2_X1 U8528 ( .A1(n6763), .A2(n6762), .ZN(n6761) );
  INV_X1 U8529 ( .A(n6877), .ZN(n6763) );
  NAND2_X1 U8530 ( .A1(n6876), .A2(n6875), .ZN(n6762) );
  NAND2_X1 U8531 ( .A1(n6877), .A2(n6716), .ZN(n11074) );
  NAND2_X1 U8532 ( .A1(n6877), .A2(n10727), .ZN(n10866) );
  NAND2_X1 U8533 ( .A1(n10725), .A2(n7740), .ZN(n10814) );
  AND2_X1 U8534 ( .A1(n10727), .A2(n10967), .ZN(n10807) );
  AND2_X1 U8535 ( .A1(n14586), .A2(n8081), .ZN(n10648) );
  INV_X1 U8536 ( .A(n7694), .ZN(n6934) );
  OAI21_X1 U8537 ( .B1(n8072), .B2(n7306), .A(n7304), .ZN(n10227) );
  INV_X1 U8538 ( .A(n7307), .ZN(n7306) );
  AOI21_X1 U8539 ( .B1(n7307), .B2(n7305), .A(n6658), .ZN(n7304) );
  NOR2_X1 U8540 ( .A1(n8076), .A2(n7308), .ZN(n7307) );
  NAND2_X1 U8541 ( .A1(n6758), .A2(n6874), .ZN(n10226) );
  INV_X1 U8542 ( .A(n10133), .ZN(n6758) );
  NAND2_X1 U8543 ( .A1(n14515), .A2(n14559), .ZN(n14514) );
  NAND2_X1 U8544 ( .A1(n6759), .A2(n14565), .ZN(n10133) );
  INV_X1 U8545 ( .A(n14514), .ZN(n6759) );
  INV_X1 U8546 ( .A(n13495), .ZN(n10484) );
  AOI21_X1 U8547 ( .B1(n8145), .B2(n9484), .A(n8144), .ZN(n10079) );
  NAND2_X1 U8548 ( .A1(n7566), .A2(n7362), .ZN(n7584) );
  NOR2_X1 U8549 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7286) );
  NOR2_X1 U8550 ( .A1(n6823), .A2(n14033), .ZN(n6741) );
  INV_X1 U8551 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6823) );
  INV_X1 U8552 ( .A(n7583), .ZN(n6821) );
  XNOR2_X1 U8553 ( .A(n8147), .B(n8146), .ZN(n9504) );
  INV_X1 U8554 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8146) );
  INV_X1 U8555 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8059) );
  NOR2_X1 U8556 ( .A1(n7345), .A2(n15138), .ZN(n7344) );
  INV_X1 U8557 ( .A(n7914), .ZN(n7345) );
  NAND2_X1 U8558 ( .A1(n7876), .A2(n6605), .ZN(n7077) );
  OR2_X1 U8559 ( .A1(n7850), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n7879) );
  AND2_X1 U8560 ( .A1(n7827), .A2(n7826), .ZN(n7831) );
  XNOR2_X1 U8561 ( .A(n7803), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13667) );
  NAND2_X1 U8562 ( .A1(n7059), .A2(n7061), .ZN(n7817) );
  NAND2_X1 U8563 ( .A1(n7801), .A2(n7060), .ZN(n7061) );
  NAND2_X1 U8564 ( .A1(n7054), .A2(n9784), .ZN(n7059) );
  OR2_X1 U8565 ( .A1(n7827), .A2(n14033), .ZN(n7750) );
  OR2_X1 U8566 ( .A1(n7714), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U8567 ( .A1(n7325), .A2(n7713), .ZN(n7728) );
  OR2_X1 U8568 ( .A1(n7701), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7714) );
  AND2_X1 U8569 ( .A1(n7669), .A2(n7668), .ZN(n7684) );
  INV_X1 U8570 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7668) );
  NOR2_X1 U8571 ( .A1(n7653), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7669) );
  OR2_X1 U8572 ( .A1(n7619), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n7653) );
  INV_X1 U8573 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8574 ( .A1(n7591), .A2(n8869), .ZN(n7605) );
  NAND2_X1 U8575 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7224), .ZN(n7223) );
  XNOR2_X1 U8576 ( .A(n14054), .B(n15220), .ZN(n14106) );
  XNOR2_X1 U8577 ( .A(n14095), .B(n6774), .ZN(n14096) );
  NAND2_X1 U8578 ( .A1(n14125), .A2(n14126), .ZN(n14127) );
  NAND2_X1 U8579 ( .A1(n15393), .A2(n15394), .ZN(n14125) );
  AOI21_X1 U8580 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14879), .A(n14077), .ZN(
        n14138) );
  NOR2_X1 U8581 ( .A1(n14136), .A2(n14135), .ZN(n14077) );
  AND2_X1 U8582 ( .A1(n7512), .A2(n7510), .ZN(n7509) );
  INV_X1 U8583 ( .A(n7515), .ZN(n7510) );
  NAND2_X1 U8584 ( .A1(n7512), .A2(n7514), .ZN(n7511) );
  OR2_X1 U8585 ( .A1(n9402), .A2(n9400), .ZN(n7514) );
  NAND2_X1 U8586 ( .A1(n9388), .A2(n11685), .ZN(n11616) );
  INV_X1 U8587 ( .A(n14979), .ZN(n10402) );
  NAND2_X1 U8588 ( .A1(n7529), .A2(n9377), .ZN(n11648) );
  AND3_X1 U8589 ( .A1(n8312), .A2(n8311), .A3(n8310), .ZN(n11679) );
  NAND2_X1 U8590 ( .A1(n11640), .A2(n7538), .ZN(n11123) );
  AOI21_X1 U8591 ( .B1(n9518), .B2(n8307), .A(n8416), .ZN(n14280) );
  INV_X1 U8592 ( .A(n14259), .ZN(n11305) );
  OR2_X1 U8593 ( .A1(n7547), .A2(n9368), .ZN(n7558) );
  NAND2_X1 U8594 ( .A1(n7522), .A2(n6594), .ZN(n11721) );
  NAND2_X1 U8595 ( .A1(n7522), .A2(n7521), .ZN(n11720) );
  NAND2_X1 U8596 ( .A1(n9420), .A2(n9419), .ZN(n11733) );
  INV_X1 U8597 ( .A(n11731), .ZN(n11744) );
  INV_X1 U8598 ( .A(n11737), .ZN(n11746) );
  INV_X1 U8599 ( .A(n11730), .ZN(n11748) );
  AND2_X1 U8600 ( .A1(n10665), .A2(n8682), .ZN(n12082) );
  INV_X1 U8601 ( .A(n12125), .ZN(n11970) );
  NAND2_X1 U8602 ( .A1(n8609), .A2(n8608), .ZN(n11971) );
  NAND2_X1 U8603 ( .A1(n8671), .A2(n11680), .ZN(n8302) );
  INV_X1 U8604 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14850) );
  NAND2_X1 U8605 ( .A1(n10274), .A2(n7149), .ZN(n10367) );
  NAND2_X1 U8606 ( .A1(n10276), .A2(n10277), .ZN(n10316) );
  AND2_X1 U8607 ( .A1(n8308), .A2(n8293), .ZN(n10297) );
  INV_X1 U8608 ( .A(n7160), .ZN(n10674) );
  OAI21_X1 U8609 ( .B1(n10351), .B2(n10783), .A(n6591), .ZN(n7160) );
  NAND2_X1 U8610 ( .A1(n7168), .A2(n7170), .ZN(n14851) );
  AND2_X1 U8611 ( .A1(n7169), .A2(n6610), .ZN(n14853) );
  OR2_X1 U8612 ( .A1(n11984), .A2(n10901), .ZN(n7169) );
  OR2_X1 U8613 ( .A1(n14871), .A2(n14872), .ZN(n7155) );
  NAND2_X1 U8614 ( .A1(n7151), .A2(n7150), .ZN(n14887) );
  NOR2_X1 U8615 ( .A1(n11988), .A2(n14906), .ZN(n14925) );
  INV_X1 U8616 ( .A(n7165), .ZN(n14195) );
  OR2_X1 U8617 ( .A1(n14193), .A2(n14194), .ZN(n7165) );
  INV_X1 U8618 ( .A(n11990), .ZN(n7164) );
  OAI21_X1 U8619 ( .B1(n14193), .B2(n7163), .A(n7162), .ZN(n14200) );
  NAND2_X1 U8620 ( .A1(n7166), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U8621 ( .A1(n11990), .A2(n7166), .ZN(n7162) );
  INV_X1 U8622 ( .A(n14201), .ZN(n7166) );
  NOR2_X1 U8623 ( .A1(n14218), .A2(n11995), .ZN(n14238) );
  NAND2_X1 U8624 ( .A1(n14242), .A2(n6733), .ZN(n12012) );
  NAND2_X1 U8625 ( .A1(n14239), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6733) );
  AOI21_X1 U8626 ( .B1(n12412), .B2(n8307), .A(n11765), .ZN(n12261) );
  NAND2_X1 U8627 ( .A1(n11756), .A2(n11755), .ZN(n14285) );
  OR2_X1 U8628 ( .A1(n11764), .A2(n11327), .ZN(n8664) );
  NAND2_X1 U8629 ( .A1(n7088), .A2(n7086), .ZN(n12091) );
  INV_X1 U8630 ( .A(n7087), .ZN(n7086) );
  OR2_X1 U8631 ( .A1(n11764), .A2(n11051), .ZN(n8644) );
  NAND2_X1 U8632 ( .A1(n8614), .A2(n8613), .ZN(n12273) );
  OR2_X1 U8633 ( .A1(n11764), .A2(n10835), .ZN(n8613) );
  NAND2_X1 U8634 ( .A1(n12419), .A2(n8698), .ZN(n12279) );
  NAND2_X1 U8635 ( .A1(n12143), .A2(n7274), .ZN(n12124) );
  NAND2_X1 U8636 ( .A1(n7103), .A2(n7107), .ZN(n12152) );
  NAND2_X1 U8637 ( .A1(n12177), .A2(n6614), .ZN(n7103) );
  NAND2_X1 U8638 ( .A1(n8571), .A2(n8570), .ZN(n12285) );
  AND2_X1 U8639 ( .A1(n7108), .A2(n7111), .ZN(n12163) );
  NAND2_X1 U8640 ( .A1(n12177), .A2(n12176), .ZN(n7108) );
  NAND2_X1 U8641 ( .A1(n8487), .A2(n8486), .ZN(n12309) );
  NAND2_X1 U8642 ( .A1(n11233), .A2(n8464), .ZN(n12248) );
  NAND2_X1 U8643 ( .A1(n8456), .A2(n8455), .ZN(n12316) );
  NAND2_X1 U8644 ( .A1(n10971), .A2(n8404), .ZN(n14273) );
  NAND2_X1 U8645 ( .A1(n7258), .A2(n7259), .ZN(n14279) );
  OR2_X1 U8646 ( .A1(n8759), .A2(n11854), .ZN(n7258) );
  NAND2_X1 U8647 ( .A1(n8759), .A2(n8758), .ZN(n10975) );
  NAND2_X1 U8648 ( .A1(n14962), .A2(n11834), .ZN(n10777) );
  AND2_X1 U8649 ( .A1(n10182), .A2(n12011), .ZN(n14999) );
  INV_X1 U8650 ( .A(n10048), .ZN(n10740) );
  NOR2_X1 U8651 ( .A1(n7124), .A2(n15056), .ZN(n7123) );
  INV_X1 U8652 ( .A(n7125), .ZN(n7124) );
  NAND2_X1 U8653 ( .A1(n12175), .A2(n11907), .ZN(n12161) );
  NAND2_X1 U8654 ( .A1(n12205), .A2(n11895), .ZN(n12188) );
  NAND2_X1 U8655 ( .A1(n8766), .A2(n11891), .ZN(n12203) );
  NAND2_X1 U8656 ( .A1(n7234), .A2(n11886), .ZN(n12232) );
  NAND2_X1 U8657 ( .A1(n12246), .A2(n12247), .ZN(n7234) );
  AND2_X1 U8658 ( .A1(n10240), .A2(P3_STATE_REG_SCAN_IN), .ZN(n15075) );
  INV_X1 U8659 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8172) );
  INV_X1 U8660 ( .A(n8175), .ZN(n11118) );
  XNOR2_X1 U8661 ( .A(n8713), .B(n15181), .ZN(n10836) );
  INV_X1 U8662 ( .A(SI_23_), .ZN(n15288) );
  NAND2_X1 U8663 ( .A1(n6953), .A2(n8552), .ZN(n8562) );
  NAND2_X1 U8664 ( .A1(n8551), .A2(n8550), .ZN(n6953) );
  INV_X1 U8665 ( .A(SI_19_), .ZN(n15339) );
  INV_X1 U8666 ( .A(SI_18_), .ZN(n9972) );
  INV_X1 U8667 ( .A(SI_17_), .ZN(n9866) );
  INV_X1 U8668 ( .A(SI_15_), .ZN(n9824) );
  INV_X1 U8669 ( .A(SI_12_), .ZN(n15245) );
  INV_X1 U8670 ( .A(SI_11_), .ZN(n15182) );
  INV_X1 U8671 ( .A(n12016), .ZN(n14880) );
  NAND2_X1 U8672 ( .A1(n6961), .A2(n6962), .ZN(n8363) );
  NAND2_X1 U8673 ( .A1(n8327), .A2(n6964), .ZN(n6961) );
  INV_X1 U8674 ( .A(n10348), .ZN(n10352) );
  NAND2_X1 U8675 ( .A1(n8327), .A2(n8198), .ZN(n8347) );
  INV_X1 U8676 ( .A(n10297), .ZN(n10314) );
  NAND2_X1 U8677 ( .A1(n8716), .A2(n8161), .ZN(n7134) );
  NAND2_X1 U8678 ( .A1(n8980), .A2(n10113), .ZN(n12446) );
  NAND2_X1 U8679 ( .A1(n10987), .A2(n7419), .ZN(n14304) );
  NAND2_X1 U8680 ( .A1(n10987), .A2(n9083), .ZN(n14301) );
  NAND2_X1 U8681 ( .A1(n12786), .A2(n9183), .ZN(n7036) );
  NAND2_X1 U8682 ( .A1(n9019), .A2(n9018), .ZN(n14811) );
  NAND2_X1 U8683 ( .A1(n11297), .A2(n7393), .ZN(n12424) );
  NAND2_X1 U8684 ( .A1(n9054), .A2(n9053), .ZN(n12589) );
  NAND2_X1 U8685 ( .A1(n7032), .A2(n9213), .ZN(n7031) );
  INV_X1 U8686 ( .A(n7032), .ZN(n12478) );
  INV_X1 U8687 ( .A(n7034), .ZN(n12480) );
  NAND2_X1 U8688 ( .A1(n9833), .A2(n9832), .ZN(n10002) );
  NAND2_X1 U8689 ( .A1(n8995), .A2(n12446), .ZN(n12445) );
  NAND2_X1 U8690 ( .A1(n9147), .A2(n9146), .ZN(n13109) );
  NAND2_X1 U8691 ( .A1(n9082), .A2(n9081), .ZN(n10987) );
  AND2_X1 U8692 ( .A1(n6858), .A2(n6859), .ZN(n6855) );
  NOR2_X1 U8693 ( .A1(n6857), .A2(n9184), .ZN(n6856) );
  INV_X1 U8694 ( .A(n6859), .ZN(n6857) );
  XNOR2_X1 U8695 ( .A(n10888), .B(n9045), .ZN(n10828) );
  OR2_X1 U8696 ( .A1(n9863), .A2(n6626), .ZN(n9979) );
  AND2_X1 U8697 ( .A1(n9132), .A2(n9131), .ZN(n7395) );
  XNOR2_X1 U8698 ( .A(n9133), .B(n9134), .ZN(n11298) );
  NAND2_X1 U8699 ( .A1(n11299), .A2(n11298), .ZN(n11297) );
  NOR2_X1 U8700 ( .A1(n10034), .A2(n7400), .ZN(n7399) );
  INV_X1 U8701 ( .A(n8945), .ZN(n7400) );
  NAND2_X1 U8702 ( .A1(n9919), .A2(n8945), .ZN(n10035) );
  NAND2_X1 U8703 ( .A1(n6931), .A2(n8831), .ZN(n13078) );
  NAND2_X1 U8704 ( .A1(n13173), .A2(n12684), .ZN(n6931) );
  NAND2_X1 U8705 ( .A1(n9858), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14331) );
  NAND2_X1 U8706 ( .A1(n9534), .A2(n9541), .ZN(n13004) );
  NAND4_X1 U8707 ( .A1(n8908), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(n12801)
         );
  INV_X1 U8708 ( .A(n10013), .ZN(n12803) );
  INV_X1 U8709 ( .A(n6906), .ZN(n9570) );
  NOR2_X1 U8710 ( .A1(n9585), .A2(n6903), .ZN(n14632) );
  NOR2_X1 U8711 ( .A1(n6905), .A2(n6904), .ZN(n6903) );
  INV_X1 U8712 ( .A(n6898), .ZN(n14660) );
  AND2_X1 U8713 ( .A1(n14693), .A2(n12834), .ZN(n14694) );
  OAI21_X1 U8714 ( .B1(n14722), .B2(n12845), .A(n12844), .ZN(n6913) );
  INV_X1 U8715 ( .A(n12855), .ZN(n12856) );
  AND2_X1 U8716 ( .A1(n12864), .A2(n12863), .ZN(n13068) );
  INV_X1 U8717 ( .A(n7450), .ZN(n12878) );
  AOI21_X1 U8718 ( .B1(n12907), .B2(n7455), .A(n7453), .ZN(n7450) );
  INV_X1 U8719 ( .A(n13078), .ZN(n12900) );
  AOI21_X1 U8720 ( .B1(n6793), .B2(n13026), .A(n6791), .ZN(n13080) );
  INV_X1 U8721 ( .A(n6792), .ZN(n6791) );
  XNOR2_X1 U8722 ( .A(n6624), .B(n12901), .ZN(n6793) );
  AOI22_X1 U8723 ( .A1(n12894), .A2(n13030), .B1(n13029), .B2(n12893), .ZN(
        n6792) );
  NAND2_X1 U8724 ( .A1(n7070), .A2(n12756), .ZN(n12938) );
  NAND2_X1 U8725 ( .A1(n12964), .A2(n7338), .ZN(n12952) );
  NAND2_X1 U8726 ( .A1(n12957), .A2(n11420), .ZN(n12942) );
  AND2_X1 U8727 ( .A1(n12960), .A2(n12959), .ZN(n13101) );
  AND2_X1 U8728 ( .A1(n7434), .A2(n6612), .ZN(n12958) );
  NAND2_X1 U8729 ( .A1(n7053), .A2(n11389), .ZN(n12988) );
  NAND2_X1 U8730 ( .A1(n7042), .A2(n7043), .ZN(n11263) );
  NAND2_X1 U8731 ( .A1(n11154), .A2(n7045), .ZN(n7042) );
  NAND2_X1 U8732 ( .A1(n7462), .A2(n11216), .ZN(n11253) );
  NAND2_X1 U8733 ( .A1(n11152), .A2(n11151), .ZN(n11218) );
  NAND2_X1 U8734 ( .A1(n7047), .A2(n7049), .ZN(n11225) );
  NAND2_X1 U8735 ( .A1(n7048), .A2(n6615), .ZN(n7047) );
  INV_X1 U8736 ( .A(n11154), .ZN(n7048) );
  NAND2_X1 U8737 ( .A1(n11000), .A2(n10999), .ZN(n11001) );
  NAND2_X1 U8738 ( .A1(n9033), .A2(n9032), .ZN(n14819) );
  NAND2_X1 U8739 ( .A1(n7074), .A2(n10600), .ZN(n10602) );
  NAND2_X1 U8740 ( .A1(n8984), .A2(n8983), .ZN(n12561) );
  NAND2_X1 U8741 ( .A1(n12979), .A2(n10425), .ZN(n13002) );
  NAND2_X1 U8742 ( .A1(n10432), .A2(n10431), .ZN(n10499) );
  INV_X1 U8743 ( .A(n13002), .ZN(n13049) );
  NAND2_X1 U8744 ( .A1(n6588), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U8745 ( .A1(n12979), .A2(n12762), .ZN(n13047) );
  AND2_X1 U8746 ( .A1(n12979), .A2(n10051), .ZN(n13044) );
  NOR2_X1 U8747 ( .A1(n13083), .A2(n6736), .ZN(n13085) );
  NAND2_X1 U8748 ( .A1(n13082), .A2(n6737), .ZN(n6736) );
  NAND2_X1 U8749 ( .A1(n13084), .A2(n14818), .ZN(n6737) );
  OR3_X1 U8750 ( .A1(n13129), .A2(n13128), .A3(n13127), .ZN(n13156) );
  NOR2_X1 U8751 ( .A1(n14724), .A2(n14753), .ZN(n14746) );
  CLKBUF_X1 U8752 ( .A(n14746), .Z(n14749) );
  AND2_X1 U8753 ( .A1(n9289), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14751) );
  INV_X1 U8754 ( .A(n8811), .ZN(n11576) );
  NAND2_X1 U8755 ( .A1(n6738), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U8756 ( .A1(n8804), .A2(n7468), .ZN(n6738) );
  CLKBUF_X1 U8757 ( .A(n13170), .Z(n6777) );
  AND2_X1 U8758 ( .A1(n9247), .A2(n8829), .ZN(n13174) );
  INV_X1 U8759 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U8760 ( .A1(n7405), .A2(n7404), .ZN(n7403) );
  INV_X1 U8761 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10412) );
  INV_X1 U8762 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10185) );
  AND2_X1 U8763 ( .A1(n9112), .A2(n9111), .ZN(n14689) );
  INV_X1 U8764 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U8765 ( .A1(n8797), .A2(n8818), .ZN(n9095) );
  INV_X1 U8766 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9831) );
  INV_X1 U8767 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9790) );
  INV_X1 U8768 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9655) );
  INV_X1 U8769 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9558) );
  INV_X1 U8770 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9533) );
  INV_X1 U8771 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9496) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U8773 ( .A1(n10207), .A2(n10206), .ZN(n10793) );
  NOR2_X1 U8774 ( .A1(n6669), .A2(n6839), .ZN(n6838) );
  NOR2_X1 U8775 ( .A1(n6840), .A2(n7484), .ZN(n6839) );
  NAND2_X1 U8776 ( .A1(n9881), .A2(n9880), .ZN(n9884) );
  INV_X1 U8777 ( .A(n7479), .ZN(n11569) );
  OAI21_X1 U8778 ( .B1(n11546), .B2(n7481), .A(n7480), .ZN(n7479) );
  AOI21_X1 U8779 ( .B1(n6669), .B2(n13182), .A(n7537), .ZN(n7480) );
  NAND2_X1 U8780 ( .A1(n13182), .A2(n13280), .ZN(n7481) );
  NAND2_X1 U8781 ( .A1(n13241), .A2(n11511), .ZN(n13208) );
  NAND2_X1 U8782 ( .A1(n7491), .A2(n7490), .ZN(n11457) );
  NAND2_X1 U8783 ( .A1(n6843), .A2(n11538), .ZN(n13216) );
  AND2_X1 U8784 ( .A1(n14356), .A2(n14358), .ZN(n6817) );
  INV_X1 U8785 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U8786 ( .A1(n13251), .A2(n13250), .ZN(n14350) );
  NAND2_X1 U8787 ( .A1(n11457), .A2(n11456), .ZN(n13251) );
  NAND2_X1 U8788 ( .A1(n13259), .A2(n13260), .ZN(n13258) );
  NAND2_X1 U8789 ( .A1(n13206), .A2(n11516), .ZN(n13259) );
  INV_X1 U8790 ( .A(n7491), .ZN(n11136) );
  NAND2_X1 U8791 ( .A1(n11059), .A2(n11058), .ZN(n11060) );
  INV_X1 U8792 ( .A(n14360), .ZN(n14353) );
  NAND2_X1 U8793 ( .A1(n13224), .A2(n11496), .ZN(n13269) );
  NAND2_X1 U8794 ( .A1(n9494), .A2(n13472), .ZN(n6947) );
  OR2_X1 U8795 ( .A1(n9692), .A2(n9687), .ZN(n13286) );
  INV_X1 U8796 ( .A(n13286), .ZN(n14365) );
  INV_X1 U8797 ( .A(n10462), .ZN(n13574) );
  INV_X1 U8798 ( .A(n6811), .ZN(n9635) );
  INV_X1 U8799 ( .A(n6813), .ZN(n9637) );
  NOR2_X1 U8800 ( .A1(n13624), .A2(n6748), .ZN(n9631) );
  NOR2_X1 U8801 ( .A1(n6749), .A2(n7635), .ZN(n6748) );
  NAND2_X1 U8802 ( .A1(n9631), .A2(n9632), .ZN(n9630) );
  NAND2_X1 U8803 ( .A1(n9633), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6810) );
  AOI21_X1 U8804 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9622), .A(n9621), .ZN(
        n9625) );
  INV_X1 U8805 ( .A(n6803), .ZN(n9671) );
  AND2_X1 U8806 ( .A1(n6803), .A2(n6802), .ZN(n9675) );
  NAND2_X1 U8807 ( .A1(n9672), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6802) );
  INV_X1 U8808 ( .A(n6801), .ZN(n9813) );
  NOR2_X1 U8809 ( .A1(n9891), .A2(n9890), .ZN(n10066) );
  NOR2_X1 U8810 ( .A1(n9889), .A2(n6805), .ZN(n9891) );
  AND2_X1 U8811 ( .A1(n9894), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6805) );
  AOI21_X1 U8812 ( .B1(n10067), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10060), .ZN(
        n10063) );
  XNOR2_X1 U8813 ( .A(n13668), .B(n6747), .ZN(n14447) );
  XNOR2_X1 U8814 ( .A(n13654), .B(n6747), .ZN(n14444) );
  NAND2_X1 U8815 ( .A1(n14444), .A2(n14443), .ZN(n14442) );
  INV_X1 U8816 ( .A(n6795), .ZN(n14456) );
  AND2_X1 U8817 ( .A1(n6949), .A2(n6948), .ZN(n13917) );
  AOI21_X1 U8818 ( .B1(n11341), .B2(n14585), .A(n13183), .ZN(n6948) );
  OR2_X1 U8819 ( .A1(n13918), .A2(n11340), .ZN(n6949) );
  NAND2_X1 U8820 ( .A1(n13747), .A2(n8100), .ZN(n13735) );
  NAND2_X1 U8821 ( .A1(n13759), .A2(n8099), .ZN(n13745) );
  NAND2_X1 U8822 ( .A1(n13792), .A2(n8097), .ZN(n13779) );
  NAND2_X1 U8823 ( .A1(n7953), .A2(n7952), .ZN(n13777) );
  NAND2_X1 U8824 ( .A1(n13810), .A2(n8096), .ZN(n13794) );
  NAND2_X1 U8825 ( .A1(n13958), .A2(n7926), .ZN(n13820) );
  NAND2_X1 U8826 ( .A1(n13843), .A2(n7323), .ZN(n13806) );
  NAND2_X1 U8827 ( .A1(n8090), .A2(n7302), .ZN(n13981) );
  NAND2_X1 U8828 ( .A1(n8090), .A2(n8089), .ZN(n13892) );
  NAND2_X1 U8829 ( .A1(n6942), .A2(n6938), .ZN(n13879) );
  AND2_X1 U8830 ( .A1(n6941), .A2(n7859), .ZN(n6938) );
  NAND2_X1 U8831 ( .A1(n11093), .A2(n7843), .ZN(n11176) );
  NAND2_X1 U8832 ( .A1(n7835), .A2(n7834), .ZN(n14384) );
  INV_X1 U8833 ( .A(n14512), .ZN(n14376) );
  NAND2_X1 U8834 ( .A1(n10744), .A2(n8083), .ZN(n10802) );
  OR2_X1 U8835 ( .A1(n10731), .A2(n13504), .ZN(n10744) );
  NAND2_X1 U8836 ( .A1(n7295), .A2(n7296), .ZN(n14586) );
  NOR2_X1 U8837 ( .A1(n13502), .A2(n7297), .ZN(n7296) );
  INV_X1 U8838 ( .A(n8079), .ZN(n7297) );
  NAND2_X1 U8839 ( .A1(n7295), .A2(n8079), .ZN(n10148) );
  NAND2_X1 U8840 ( .A1(n10140), .A2(n13502), .ZN(n10139) );
  NAND2_X1 U8841 ( .A1(n10155), .A2(n7694), .ZN(n10140) );
  OAI21_X1 U8842 ( .B1(n7354), .B2(n7348), .A(n7349), .ZN(n10224) );
  AOI21_X1 U8843 ( .B1(n7351), .B2(n7647), .A(n7350), .ZN(n7349) );
  NAND2_X1 U8844 ( .A1(n7309), .A2(n8074), .ZN(n10127) );
  NAND2_X1 U8845 ( .A1(n8072), .A2(n13318), .ZN(n10085) );
  NAND2_X1 U8846 ( .A1(n14536), .A2(n10081), .ZN(n13895) );
  AND2_X1 U8847 ( .A1(n14536), .A2(n14522), .ZN(n14512) );
  NAND2_X1 U8848 ( .A1(n9691), .A2(n9690), .ZN(n14508) );
  INV_X1 U8849 ( .A(n9986), .ZN(n14526) );
  AND2_X1 U8850 ( .A1(n14536), .A2(n14585), .ZN(n14532) );
  INV_X1 U8851 ( .A(n13976), .ZN(n13969) );
  CLKBUF_X1 U8852 ( .A(n14597), .Z(n14600) );
  AOI21_X1 U8853 ( .B1(n13911), .B2(n14585), .A(n13910), .ZN(n13912) );
  INV_X1 U8854 ( .A(n13729), .ZN(n14004) );
  NAND2_X1 U8855 ( .A1(n7990), .A2(n7989), .ZN(n14007) );
  NAND2_X1 U8856 ( .A1(n7977), .A2(n7976), .ZN(n14011) );
  INV_X1 U8857 ( .A(n13831), .ZN(n14018) );
  AND2_X1 U8858 ( .A1(n14044), .A2(n14048), .ZN(n9485) );
  AND2_X1 U8859 ( .A1(n9504), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9486) );
  AND2_X1 U8860 ( .A1(n7551), .A2(n7500), .ZN(n7499) );
  AND2_X1 U8861 ( .A1(n7502), .A2(n7570), .ZN(n7500) );
  XNOR2_X1 U8862 ( .A(n7960), .B(SI_23_), .ZN(n11171) );
  XNOR2_X1 U8863 ( .A(n7944), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14050) );
  INV_X1 U8864 ( .A(n8062), .ZN(n8063) );
  NAND2_X1 U8865 ( .A1(n7892), .A2(n7878), .ZN(n10723) );
  INV_X1 U8866 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n15334) );
  INV_X1 U8867 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10154) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10045) );
  INV_X1 U8869 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9930) );
  INV_X1 U8870 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9828) );
  AND2_X1 U8871 ( .A1(n7789), .A2(n7802), .ZN(n14425) );
  INV_X1 U8872 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9788) );
  INV_X1 U8873 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9701) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9658) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9530) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9499) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9476) );
  XNOR2_X1 U8878 ( .A(n6807), .B(n6806), .ZN(n13596) );
  NOR2_X1 U8879 ( .A1(n7608), .A2(n14033), .ZN(n6807) );
  XNOR2_X1 U8880 ( .A(n7594), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13577) );
  XNOR2_X1 U8881 ( .A(n14115), .B(n14638), .ZN(n14160) );
  XNOR2_X1 U8882 ( .A(n14127), .B(n14128), .ZN(n14165) );
  AND2_X1 U8883 ( .A1(n14133), .A2(n14134), .ZN(n14170) );
  NAND2_X1 U8884 ( .A1(n14398), .A2(n6775), .ZN(n14404) );
  OAI21_X1 U8885 ( .B1(n14400), .B2(n14399), .A(P2_ADDR_REG_12__SCAN_IN), .ZN(
        n6775) );
  NAND2_X1 U8886 ( .A1(n6740), .A2(n14692), .ZN(n7219) );
  INV_X1 U8887 ( .A(n14415), .ZN(n7218) );
  NAND2_X1 U8888 ( .A1(n14174), .A2(n14175), .ZN(n14173) );
  CLKBUF_X1 U8889 ( .A(n11973), .Z(P3_U3897) );
  NAND2_X1 U8890 ( .A1(n7560), .A2(n6646), .ZN(P3_U3488) );
  NAND2_X1 U8891 ( .A1(n9283), .A2(n9282), .ZN(n9307) );
  OAI211_X1 U8892 ( .C1(n12843), .C2(n12842), .A(n6912), .B(n6909), .ZN(
        P2_U3233) );
  INV_X1 U8893 ( .A(n6913), .ZN(n6912) );
  NAND2_X1 U8894 ( .A1(n6910), .A2(n12842), .ZN(n6909) );
  NAND2_X1 U8895 ( .A1(n14827), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8896 ( .A1(n13144), .A2(n14829), .ZN(n7022) );
  AND3_X1 U8897 ( .A1(n13541), .A2(n13540), .A3(n13539), .ZN(n13547) );
  NAND2_X1 U8898 ( .A1(n7487), .A2(n7485), .ZN(P1_U3561) );
  OR2_X1 U8899 ( .A1(n13591), .A2(n9526), .ZN(n7487) );
  AND3_X1 U8900 ( .A1(n14496), .A2(n14495), .A3(n14494), .ZN(n14498) );
  AOI21_X1 U8901 ( .B1(n6798), .B2(n13525), .A(n6797), .ZN(n6796) );
  INV_X1 U8902 ( .A(n13676), .ZN(n13678) );
  OAI21_X1 U8903 ( .B1(n13429), .B2(n13976), .A(n8157), .ZN(n8158) );
  AOI21_X1 U8904 ( .B1(n13526), .B2(n14023), .A(n6756), .ZN(n6755) );
  NOR2_X1 U8905 ( .A1(n8150), .A2(n13993), .ZN(n6756) );
  NAND2_X1 U8906 ( .A1(n8156), .A2(n8150), .ZN(n8153) );
  XNOR2_X1 U8907 ( .A(n14184), .B(n6725), .ZN(n7225) );
  NAND2_X1 U8908 ( .A1(n10321), .A2(n10352), .ZN(n6591) );
  AND2_X1 U8909 ( .A1(n12888), .A2(n12894), .ZN(n6592) );
  XOR2_X1 U8910 ( .A(n7729), .B(SI_9_), .Z(n6593) );
  AND2_X1 U8911 ( .A1(n7520), .A2(n7521), .ZN(n6594) );
  AND2_X1 U8912 ( .A1(n7259), .A2(n7257), .ZN(n6595) );
  NAND4_X1 U8913 ( .A1(n8304), .A2(n8303), .A3(n8302), .A4(n8301), .ZN(n14965)
         );
  INV_X1 U8914 ( .A(n7566), .ZN(n8057) );
  NAND2_X1 U8915 ( .A1(n12660), .A2(n7190), .ZN(n7189) );
  INV_X1 U8916 ( .A(n7189), .ZN(n7184) );
  NAND2_X1 U8917 ( .A1(n7732), .A2(n7731), .ZN(n13352) );
  AND2_X1 U8918 ( .A1(n7364), .A2(n13425), .ZN(n6596) );
  INV_X1 U8919 ( .A(n12117), .ZN(n10445) );
  AND2_X1 U8920 ( .A1(n8638), .A2(n8637), .ZN(n12117) );
  NAND2_X1 U8921 ( .A1(n8645), .A2(n8644), .ZN(n12266) );
  AND2_X1 U8922 ( .A1(n6676), .A2(n8100), .ZN(n6597) );
  AND2_X1 U8923 ( .A1(n13426), .A2(n7363), .ZN(n6598) );
  INV_X1 U8924 ( .A(n7843), .ZN(n7359) );
  INV_X1 U8925 ( .A(n6960), .ZN(n6959) );
  AND2_X1 U8926 ( .A1(n6694), .A2(n6962), .ZN(n6960) );
  AND2_X1 U8927 ( .A1(n7416), .A2(n8819), .ZN(n6599) );
  INV_X1 U8928 ( .A(n13526), .ZN(n13994) );
  NAND2_X1 U8929 ( .A1(n13476), .A2(n13475), .ZN(n13526) );
  AND2_X1 U8930 ( .A1(n9046), .A2(n9045), .ZN(n6600) );
  AND2_X1 U8931 ( .A1(n10382), .A2(n8997), .ZN(n6601) );
  AND2_X1 U8932 ( .A1(n9215), .A2(n9214), .ZN(n12915) );
  INV_X1 U8933 ( .A(n12915), .ZN(n13084) );
  INV_X1 U8934 ( .A(n13405), .ZN(n7370) );
  OR2_X1 U8935 ( .A1(n8579), .A2(n12165), .ZN(n6602) );
  AND2_X1 U8936 ( .A1(n7418), .A2(n9109), .ZN(n6603) );
  AND2_X1 U8937 ( .A1(n7147), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6604) );
  AND2_X2 U8938 ( .A1(n12516), .A2(n12509), .ZN(n12528) );
  NAND2_X1 U8939 ( .A1(n6708), .A2(n7503), .ZN(n8399) );
  AND2_X1 U8940 ( .A1(n7908), .A2(n7905), .ZN(n6605) );
  NAND2_X1 U8941 ( .A1(n9701), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6606) );
  INV_X1 U8942 ( .A(n12247), .ZN(n7229) );
  NAND2_X1 U8943 ( .A1(n7771), .A2(n7770), .ZN(n13363) );
  INV_X1 U8944 ( .A(n13363), .ZN(n6876) );
  NAND2_X1 U8945 ( .A1(n11059), .A2(n7493), .ZN(n7491) );
  INV_X1 U8946 ( .A(n9326), .ZN(n9316) );
  OR2_X1 U8947 ( .A1(n10163), .A2(n14578), .ZN(n6608) );
  INV_X1 U8948 ( .A(n11729), .ZN(n7517) );
  AND2_X1 U8949 ( .A1(n12883), .A2(n7335), .ZN(n6609) );
  OR2_X1 U8950 ( .A1(n11983), .A2(n11982), .ZN(n6610) );
  OR2_X1 U8951 ( .A1(n12828), .A2(n6895), .ZN(n6611) );
  NAND2_X1 U8952 ( .A1(n13105), .A2(n12492), .ZN(n6612) );
  OR3_X1 U8953 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        n10253), .ZN(n6613) );
  AND2_X1 U8954 ( .A1(n7110), .A2(n12176), .ZN(n6614) );
  NAND2_X1 U8955 ( .A1(n12594), .A2(n14305), .ZN(n6615) );
  NOR2_X1 U8956 ( .A1(n11224), .A2(n7046), .ZN(n7045) );
  AND2_X1 U8957 ( .A1(n9882), .A2(n9880), .ZN(n6616) );
  AND3_X1 U8958 ( .A1(n8267), .A2(n8266), .A3(n8265), .ZN(n6617) );
  AND2_X1 U8959 ( .A1(n8058), .A2(n7008), .ZN(n6618) );
  AND4_X1 U8960 ( .A1(n7437), .A2(n7435), .A3(n7542), .A4(n8796), .ZN(n6619)
         );
  OR2_X1 U8961 ( .A1(n14058), .A2(n14057), .ZN(n6620) );
  AND2_X1 U8962 ( .A1(n13939), .A2(n13553), .ZN(n6621) );
  OAI21_X1 U8963 ( .B1(n13206), .B2(n6831), .A(n6828), .ZN(n13189) );
  NAND2_X1 U8964 ( .A1(n10944), .A2(n10943), .ZN(n6622) );
  INV_X1 U8965 ( .A(n10308), .ZN(n10564) );
  AND2_X1 U8966 ( .A1(n7497), .A2(n6835), .ZN(n6623) );
  INV_X1 U8967 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8913) );
  INV_X1 U8968 ( .A(n13280), .ZN(n7484) );
  INV_X1 U8969 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15220) );
  INV_X1 U8970 ( .A(n11891), .ZN(n7269) );
  NAND2_X1 U8971 ( .A1(n7646), .A2(n7645), .ZN(n13322) );
  INV_X1 U8972 ( .A(n13322), .ZN(n14565) );
  INV_X1 U8973 ( .A(n10277), .ZN(n7143) );
  OR2_X1 U8974 ( .A1(n12907), .A2(n11423), .ZN(n6624) );
  NAND2_X1 U8975 ( .A1(n8804), .A2(n7469), .ZN(n8808) );
  AND2_X1 U8976 ( .A1(n12289), .A2(n11974), .ZN(n6625) );
  XNOR2_X1 U8977 ( .A(n14578), .B(n8080), .ZN(n13502) );
  INV_X1 U8978 ( .A(n13502), .ZN(n6935) );
  NAND2_X1 U8979 ( .A1(n9174), .A2(n9173), .ZN(n13099) );
  INV_X1 U8980 ( .A(n13099), .ZN(n6885) );
  INV_X1 U8981 ( .A(n11887), .ZN(n7231) );
  OR2_X1 U8982 ( .A1(n9856), .A2(n9901), .ZN(n6626) );
  AND2_X1 U8983 ( .A1(n6811), .A2(n6810), .ZN(n6627) );
  AND2_X1 U8984 ( .A1(n7330), .A2(n6921), .ZN(n6628) );
  INV_X1 U8985 ( .A(n12632), .ZN(n7202) );
  OR2_X1 U8986 ( .A1(n7058), .A2(n9784), .ZN(n6629) );
  NOR2_X1 U8987 ( .A1(n13392), .A2(n13391), .ZN(n6630) );
  AND2_X1 U8988 ( .A1(n13397), .A2(n13398), .ZN(n13513) );
  INV_X1 U8989 ( .A(n12599), .ZN(n14333) );
  NAND2_X1 U8990 ( .A1(n7753), .A2(n7752), .ZN(n13355) );
  AND2_X1 U8991 ( .A1(n14949), .A2(n8353), .ZN(n6631) );
  AND2_X1 U8992 ( .A1(n7161), .A2(n10783), .ZN(n6632) );
  OR2_X1 U8993 ( .A1(n8708), .A2(n14988), .ZN(n6633) );
  OAI22_X1 U8994 ( .A1(n12658), .A2(n12659), .B1(n12656), .B2(n12657), .ZN(
        n7190) );
  AND2_X1 U8995 ( .A1(n13669), .A2(n6794), .ZN(n6634) );
  AND2_X1 U8996 ( .A1(n12651), .A2(n7185), .ZN(n6635) );
  AND2_X1 U8997 ( .A1(n12143), .A2(n11924), .ZN(n6636) );
  NAND2_X1 U8998 ( .A1(n11941), .A2(n11943), .ZN(n12089) );
  INV_X1 U8999 ( .A(n12089), .ZN(n7092) );
  NAND2_X1 U9000 ( .A1(n11834), .A2(n11833), .ZN(n8337) );
  OR2_X1 U9001 ( .A1(n12263), .A2(n12093), .ZN(n11946) );
  AND2_X1 U9002 ( .A1(n7204), .A2(n7202), .ZN(n6637) );
  AND2_X1 U9003 ( .A1(n11953), .A2(n11946), .ZN(n6638) );
  AND2_X1 U9004 ( .A1(n12202), .A2(n7130), .ZN(n6639) );
  AND2_X1 U9005 ( .A1(n12599), .A2(n12790), .ZN(n6640) );
  NAND2_X1 U9006 ( .A1(n14327), .A2(n11281), .ZN(n6641) );
  NAND2_X1 U9007 ( .A1(n13939), .A2(n8098), .ZN(n6642) );
  AND2_X1 U9008 ( .A1(n8385), .A2(n8368), .ZN(n6643) );
  AND2_X1 U9009 ( .A1(n11513), .A2(n11511), .ZN(n6644) );
  OR2_X1 U9010 ( .A1(n13394), .A2(n6630), .ZN(n6645) );
  AND2_X1 U9011 ( .A1(n8779), .A2(n8778), .ZN(n6646) );
  AND2_X1 U9012 ( .A1(n12561), .A2(n10686), .ZN(n6647) );
  AND3_X1 U9013 ( .A1(n6994), .A2(n13326), .A3(n6993), .ZN(n6648) );
  AND2_X1 U9014 ( .A1(n7165), .A2(n7164), .ZN(n6649) );
  AND2_X1 U9015 ( .A1(n8656), .A2(n8655), .ZN(n12102) );
  AND2_X1 U9016 ( .A1(n7270), .A2(n11895), .ZN(n6650) );
  AND2_X1 U9017 ( .A1(n12313), .A2(n11977), .ZN(n6651) );
  INV_X1 U9018 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8716) );
  INV_X1 U9019 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8827) );
  AND2_X1 U9020 ( .A1(n7211), .A2(n12571), .ZN(n6652) );
  NOR2_X1 U9021 ( .A1(n13137), .A2(n14307), .ZN(n6653) );
  AND2_X1 U9022 ( .A1(n7529), .A2(n7526), .ZN(n6654) );
  AND2_X1 U9023 ( .A1(n13721), .A2(n13708), .ZN(n6655) );
  AND2_X1 U9024 ( .A1(n8164), .A2(n7531), .ZN(n6656) );
  NOR2_X1 U9025 ( .A1(n12289), .A2(n12179), .ZN(n6657) );
  AND2_X1 U9026 ( .A1(n13372), .A2(n13373), .ZN(n13377) );
  INV_X1 U9027 ( .A(n13377), .ZN(n6984) );
  AND2_X1 U9028 ( .A1(n14571), .A2(n8075), .ZN(n6658) );
  AND2_X1 U9029 ( .A1(n10308), .A2(n10315), .ZN(n7145) );
  AND2_X1 U9030 ( .A1(n13357), .A2(n13356), .ZN(n6659) );
  INV_X1 U9031 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8822) );
  INV_X1 U9032 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U9033 ( .A1(n7371), .A2(n7368), .ZN(n6660) );
  INV_X1 U9034 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14033) );
  NOR2_X1 U9035 ( .A1(n9402), .A2(n7513), .ZN(n6661) );
  AND2_X1 U9036 ( .A1(n6995), .A2(n7001), .ZN(n6662) );
  AND2_X1 U9037 ( .A1(n6971), .A2(n13346), .ZN(n6663) );
  INV_X1 U9038 ( .A(n7561), .ZN(n7492) );
  AND2_X1 U9039 ( .A1(n7317), .A2(n13778), .ZN(n6664) );
  NAND2_X1 U9040 ( .A1(n13843), .A2(n13398), .ZN(n6665) );
  AND2_X1 U9041 ( .A1(n7682), .A2(SI_6_), .ZN(n6666) );
  AND2_X1 U9042 ( .A1(n7729), .A2(SI_9_), .ZN(n6667) );
  AND2_X1 U9043 ( .A1(n13419), .A2(n13418), .ZN(n6668) );
  NAND2_X1 U9044 ( .A1(n7482), .A2(n11553), .ZN(n6669) );
  AND2_X1 U9045 ( .A1(n6660), .A2(n7370), .ZN(n6670) );
  INV_X1 U9046 ( .A(n7527), .ZN(n7526) );
  OR2_X1 U9047 ( .A1(n11649), .A2(n7528), .ZN(n7527) );
  OR2_X1 U9048 ( .A1(n13939), .A2(n13553), .ZN(n6671) );
  INV_X1 U9049 ( .A(n12110), .ZN(n12268) );
  AND2_X1 U9050 ( .A1(n8630), .A2(n8629), .ZN(n12110) );
  OAI21_X1 U9051 ( .B1(n6964), .B2(n6959), .A(n8199), .ZN(n6958) );
  OR2_X1 U9052 ( .A1(n12110), .A2(n12117), .ZN(n6672) );
  AND2_X1 U9053 ( .A1(n13309), .A2(n13308), .ZN(n6673) );
  NAND2_X1 U9054 ( .A1(n12333), .A2(n10402), .ZN(n8751) );
  AND2_X1 U9055 ( .A1(n6768), .A2(n6767), .ZN(n6674) );
  INV_X1 U9056 ( .A(n6892), .ZN(n12854) );
  AND2_X1 U9057 ( .A1(n9336), .A2(n11980), .ZN(n6675) );
  NAND2_X1 U9058 ( .A1(n13729), .A2(n11336), .ZN(n6676) );
  INV_X1 U9059 ( .A(n11420), .ZN(n7432) );
  OR2_X1 U9060 ( .A1(n13099), .A2(n12978), .ZN(n11420) );
  NAND2_X1 U9061 ( .A1(n10462), .A2(n9986), .ZN(n13310) );
  XOR2_X1 U9062 ( .A(n12853), .B(n12726), .Z(n6677) );
  OR2_X1 U9063 ( .A1(n6625), .A2(n7109), .ZN(n6678) );
  INV_X1 U9064 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9524) );
  INV_X1 U9065 ( .A(n12560), .ZN(n7196) );
  INV_X1 U9066 ( .A(n13426), .ZN(n7364) );
  NAND2_X1 U9067 ( .A1(n12660), .A2(n7191), .ZN(n6679) );
  INV_X1 U9068 ( .A(n12597), .ZN(n7178) );
  XNOR2_X1 U9069 ( .A(n8061), .B(P1_IR_REG_21__SCAN_IN), .ZN(n13450) );
  OR2_X1 U9070 ( .A1(n14128), .A2(n14127), .ZN(n6680) );
  AND3_X1 U9071 ( .A1(n8802), .A2(n8803), .A3(n8796), .ZN(n6681) );
  OR2_X1 U9072 ( .A1(n14178), .A2(n14177), .ZN(n6682) );
  AND2_X1 U9073 ( .A1(n10828), .A2(n9044), .ZN(n6683) );
  NOR2_X1 U9074 ( .A1(n14578), .A2(n13567), .ZN(n6684) );
  INV_X1 U9075 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6963) );
  OR2_X1 U9076 ( .A1(n12285), .A2(n11972), .ZN(n6685) );
  AND2_X1 U9077 ( .A1(n6887), .A2(n13126), .ZN(n6686) );
  AND2_X1 U9078 ( .A1(n11389), .A2(n7535), .ZN(n6687) );
  NAND2_X1 U9079 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6688) );
  AND2_X1 U9080 ( .A1(n11927), .A2(n11925), .ZN(n12126) );
  INV_X1 U9081 ( .A(n7816), .ZN(n7058) );
  AND2_X1 U9082 ( .A1(n9343), .A2(n7538), .ZN(n6689) );
  OR2_X1 U9083 ( .A1(n7068), .A2(n7337), .ZN(n6690) );
  INV_X1 U9084 ( .A(n10431), .ZN(n7030) );
  NAND2_X1 U9085 ( .A1(n13045), .A2(n13005), .ZN(n6691) );
  INV_X1 U9086 ( .A(n7339), .ZN(n7338) );
  NOR2_X1 U9087 ( .A1(n6885), .A2(n12978), .ZN(n7339) );
  AND2_X1 U9088 ( .A1(n6618), .A2(n8059), .ZN(n6692) );
  NAND2_X1 U9089 ( .A1(n11339), .A2(n11338), .ZN(n6693) );
  NAND2_X1 U9090 ( .A1(n9530), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6694) );
  INV_X1 U9091 ( .A(n7662), .ZN(n7350) );
  INV_X1 U9092 ( .A(n14543), .ZN(n13311) );
  INV_X1 U9093 ( .A(n7555), .ZN(n7478) );
  INV_X1 U9094 ( .A(n7239), .ZN(n7238) );
  NAND2_X1 U9095 ( .A1(n7240), .A2(n8767), .ZN(n7239) );
  INV_X1 U9096 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7570) );
  OR2_X1 U9097 ( .A1(n7647), .A2(n7350), .ZN(n6695) );
  INV_X1 U9098 ( .A(n7324), .ZN(n7323) );
  NAND2_X1 U9099 ( .A1(n13834), .A2(n13398), .ZN(n7324) );
  INV_X1 U9100 ( .A(n7420), .ZN(n7419) );
  NAND2_X1 U9101 ( .A1(n7421), .A2(n9083), .ZN(n7420) );
  INV_X1 U9102 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9502) );
  INV_X1 U9103 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6806) );
  INV_X1 U9104 ( .A(n6930), .ZN(n6929) );
  NAND2_X1 U9105 ( .A1(n7550), .A2(n6629), .ZN(n6930) );
  INV_X1 U9106 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9470) );
  AND2_X1 U9107 ( .A1(n7052), .A2(n7335), .ZN(n6696) );
  AND2_X1 U9108 ( .A1(n14350), .A2(n11470), .ZN(n6697) );
  AND2_X1 U9109 ( .A1(n13416), .A2(n6976), .ZN(n6698) );
  INV_X1 U9110 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7501) );
  NAND3_X1 U9111 ( .A1(n7266), .A2(n7264), .A3(n7507), .ZN(n6699) );
  NAND2_X1 U9112 ( .A1(n12233), .A2(n7128), .ZN(n7131) );
  OR2_X1 U9113 ( .A1(n8259), .A2(n7133), .ZN(n7132) );
  AND2_X1 U9114 ( .A1(n11155), .A2(n6887), .ZN(n6700) );
  INV_X1 U9115 ( .A(n14278), .ZN(n7257) );
  INV_X1 U9116 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7417) );
  INV_X1 U9117 ( .A(n11972), .ZN(n12165) );
  INV_X1 U9118 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6904) );
  AND2_X1 U9119 ( .A1(n9222), .A2(n9221), .ZN(n12928) );
  INV_X1 U9120 ( .A(n12928), .ZN(n12893) );
  AND2_X1 U9121 ( .A1(n9242), .A2(n9241), .ZN(n12695) );
  INV_X1 U9122 ( .A(n12695), .ZN(n12894) );
  INV_X1 U9123 ( .A(n6881), .ZN(n13885) );
  AND2_X1 U9124 ( .A1(n10793), .A2(n6851), .ZN(n6701) );
  NAND2_X1 U9125 ( .A1(n7131), .A2(n7130), .ZN(n6702) );
  AND2_X1 U9126 ( .A1(n6855), .A2(n6860), .ZN(n6703) );
  AND2_X1 U9127 ( .A1(n11187), .A2(n7815), .ZN(n6704) );
  AND2_X1 U9128 ( .A1(n7491), .A2(n7492), .ZN(n6705) );
  INV_X1 U9129 ( .A(n12154), .ZN(n11617) );
  AND2_X1 U9130 ( .A1(n8595), .A2(n8594), .ZN(n12154) );
  AND2_X1 U9131 ( .A1(n14425), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6706) );
  AND2_X1 U9132 ( .A1(n7042), .A2(n7041), .ZN(n6707) );
  AND3_X1 U9133 ( .A1(n7082), .A2(n8163), .A3(n8397), .ZN(n6708) );
  INV_X1 U9134 ( .A(n11496), .ZN(n7477) );
  INV_X1 U9135 ( .A(n7343), .ZN(n7342) );
  NOR2_X1 U9136 ( .A1(n7914), .A2(SI_20_), .ZN(n7343) );
  AND2_X1 U9137 ( .A1(n9698), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U9138 ( .A1(n8818), .A2(n7416), .ZN(n6710) );
  OR2_X1 U9139 ( .A1(n14852), .A2(n10901), .ZN(n6711) );
  NAND2_X1 U9140 ( .A1(n12018), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6712) );
  INV_X1 U9141 ( .A(n7111), .ZN(n7109) );
  NAND2_X1 U9142 ( .A1(n12293), .A2(n12192), .ZN(n7111) );
  NAND2_X1 U9143 ( .A1(n12616), .A2(n7199), .ZN(n6713) );
  AND2_X1 U9144 ( .A1(n7505), .A2(n7506), .ZN(n6714) );
  INV_X1 U9145 ( .A(n14028), .ZN(n14023) );
  INV_X1 U9146 ( .A(n12743), .ZN(n7467) );
  AND2_X1 U9147 ( .A1(n10818), .A2(n6683), .ZN(n6715) );
  INV_X1 U9148 ( .A(n8316), .ZN(n10658) );
  INV_X1 U9149 ( .A(n8298), .ZN(n8316) );
  INV_X1 U9150 ( .A(n12235), .ZN(n7233) );
  NAND2_X1 U9151 ( .A1(n7117), .A2(n7119), .ZN(n14256) );
  AND2_X1 U9152 ( .A1(n11829), .A2(n11828), .ZN(n11825) );
  INV_X1 U9153 ( .A(n11825), .ZN(n8313) );
  INV_X1 U9154 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U9155 ( .A1(n7867), .A2(n7866), .ZN(n13979) );
  INV_X1 U9156 ( .A(n13979), .ZN(n6880) );
  OR2_X1 U9157 ( .A1(n13497), .A2(n7352), .ZN(n7348) );
  AND2_X1 U9158 ( .A1(n10727), .A2(n6876), .ZN(n6716) );
  INV_X2 U9159 ( .A(n15056), .ZN(n15055) );
  AND2_X1 U9160 ( .A1(n9438), .A2(n9437), .ZN(n15056) );
  NAND2_X1 U9161 ( .A1(n14899), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6717) );
  AND2_X1 U9162 ( .A1(n7353), .A2(n7351), .ZN(n6718) );
  AND2_X1 U9163 ( .A1(n10778), .A2(n8353), .ZN(n6719) );
  AND2_X1 U9164 ( .A1(n10619), .A2(n8315), .ZN(n6720) );
  AND2_X1 U9165 ( .A1(n14948), .A2(n8368), .ZN(n6721) );
  INV_X1 U9166 ( .A(n7859), .ZN(n6943) );
  AND2_X1 U9167 ( .A1(n7155), .A2(n7154), .ZN(n6722) );
  NAND2_X1 U9168 ( .A1(n7793), .A2(n7792), .ZN(n13366) );
  INV_X1 U9169 ( .A(n13366), .ZN(n6875) );
  AND2_X2 U9170 ( .A1(n10030), .A2(n14750), .ZN(n14829) );
  INV_X1 U9171 ( .A(n14445), .ZN(n6747) );
  OR2_X1 U9172 ( .A1(n12045), .A2(n11991), .ZN(n6723) );
  AND2_X1 U9173 ( .A1(n8691), .A2(n9405), .ZN(n12249) );
  INV_X1 U9174 ( .A(n12249), .ZN(n14982) );
  XOR2_X1 U9175 ( .A(n9010), .B(n9011), .Z(n6724) );
  NAND3_X1 U9176 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(n12337) );
  INV_X1 U9177 ( .A(n12337), .ZN(n7267) );
  INV_X1 U9178 ( .A(n14571), .ZN(n6874) );
  INV_X1 U9179 ( .A(n10113), .ZN(n7414) );
  INV_X1 U9180 ( .A(n9590), .ZN(n6905) );
  INV_X1 U9181 ( .A(n13525), .ZN(n14523) );
  NAND2_X1 U9182 ( .A1(n6559), .A2(n12842), .ZN(n12725) );
  INV_X1 U9183 ( .A(n14703), .ZN(n6894) );
  NAND2_X1 U9184 ( .A1(n7499), .A2(n7566), .ZN(n14032) );
  NAND2_X1 U9185 ( .A1(n13627), .A2(n13628), .ZN(n6815) );
  NAND2_X1 U9186 ( .A1(n14613), .A2(n14614), .ZN(n6908) );
  XOR2_X1 U9187 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n6725) );
  INV_X1 U9188 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7224) );
  INV_X1 U9189 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6774) );
  INV_X1 U9190 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U9191 ( .A1(n13019), .A2(n13031), .ZN(n7423) );
  NAND2_X1 U9192 ( .A1(n7019), .A2(n7862), .ZN(n7874) );
  OAI21_X1 U9193 ( .B1(n7781), .B2(n6930), .A(n6926), .ZN(n7822) );
  NAND2_X1 U9194 ( .A1(n12679), .A2(n12678), .ZN(n12683) );
  OAI21_X1 U9195 ( .B1(n12444), .B2(n12443), .A(n6727), .ZN(P2_U3192) );
  INV_X1 U9196 ( .A(n6728), .ZN(n6727) );
  NAND2_X1 U9197 ( .A1(n7412), .A2(n7411), .ZN(n10386) );
  OAI21_X1 U9198 ( .B1(n12488), .B2(n12484), .A(n12485), .ZN(n12459) );
  NAND2_X1 U9199 ( .A1(n7273), .A2(n7271), .ZN(n12113) );
  NAND2_X1 U9200 ( .A1(n7227), .A2(n7230), .ZN(n12217) );
  NAND2_X1 U9201 ( .A1(n7241), .A2(n7243), .ZN(n14947) );
  NAND2_X1 U9202 ( .A1(n7256), .A2(n7254), .ZN(n14266) );
  OAI21_X1 U9203 ( .B1(n12150), .B2(n11916), .A(n11793), .ZN(n12141) );
  OAI21_X1 U9204 ( .B1(n12101), .B2(n11937), .A(n11791), .ZN(n12090) );
  NAND2_X1 U9205 ( .A1(n12539), .A2(n12540), .ZN(n12538) );
  NAND2_X1 U9206 ( .A1(n12533), .A2(n6787), .ZN(n12539) );
  NAND2_X1 U9207 ( .A1(n6745), .A2(n6744), .ZN(n12648) );
  NAND3_X1 U9208 ( .A1(n12544), .A2(n12543), .A3(n6732), .ZN(n6731) );
  NAND2_X1 U9209 ( .A1(n12598), .A2(n6742), .ZN(n12603) );
  NAND2_X1 U9210 ( .A1(n7208), .A2(n7210), .ZN(n12647) );
  OAI21_X1 U9211 ( .B1(n6935), .B2(n10155), .A(n6933), .ZN(n10645) );
  OAI21_X2 U9213 ( .B1(n13859), .B2(n7890), .A(n7889), .ZN(n13839) );
  NAND2_X2 U9214 ( .A1(n13743), .A2(n13744), .ZN(n13742) );
  AND3_X4 U9215 ( .A1(n7284), .A2(n7279), .A3(n7280), .ZN(n7566) );
  NAND2_X1 U9216 ( .A1(n13314), .A2(n13299), .ZN(n13495) );
  INV_X2 U9217 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9683) );
  NOR2_X2 U9218 ( .A1(n13695), .A2(n6655), .ZN(n13696) );
  NAND2_X1 U9219 ( .A1(n13791), .A2(n13795), .ZN(n7953) );
  INV_X4 U9220 ( .A(n13438), .ZN(n7991) );
  OAI211_X1 U9221 ( .C1(n10084), .C2(n6695), .A(n10228), .B(n7347), .ZN(n10223) );
  NAND2_X1 U9222 ( .A1(n7355), .A2(n13518), .ZN(n11337) );
  NAND2_X1 U9223 ( .A1(n6946), .A2(n7872), .ZN(n13859) );
  NAND2_X1 U9224 ( .A1(n10645), .A2(n13503), .ZN(n10644) );
  NAND2_X1 U9225 ( .A1(n6942), .A2(n6939), .ZN(n6946) );
  NAND2_X1 U9226 ( .A1(n7613), .A2(n7612), .ZN(n14501) );
  NAND2_X1 U9227 ( .A1(n10870), .A2(n7778), .ZN(n11079) );
  NAND2_X1 U9228 ( .A1(n7904), .A2(n7903), .ZN(n13835) );
  NAND2_X2 U9229 ( .A1(n6937), .A2(n13825), .ZN(n13958) );
  XNOR2_X2 U9230 ( .A(n7568), .B(n7567), .ZN(n11360) );
  NAND2_X1 U9231 ( .A1(n7135), .A2(n7134), .ZN(n7133) );
  NAND2_X1 U9232 ( .A1(n8041), .A2(n8040), .ZN(n11332) );
  NAND2_X1 U9233 ( .A1(n7988), .A2(n7987), .ZN(n8003) );
  INV_X1 U9234 ( .A(n13445), .ZN(n6734) );
  NAND2_X1 U9235 ( .A1(n11359), .A2(n12679), .ZN(n13445) );
  OAI211_X1 U9236 ( .C1(n11604), .C2(n11605), .A(n6735), .B(n11603), .ZN(
        P3_U3160) );
  NAND4_X1 U9237 ( .A1(n11604), .A2(n11600), .A3(n11596), .A4(n11730), .ZN(
        n6735) );
  NAND2_X1 U9238 ( .A1(n7519), .A2(n7518), .ZN(n11608) );
  NAND2_X1 U9239 ( .A1(n11608), .A2(n11607), .ZN(n11606) );
  INV_X1 U9240 ( .A(n7530), .ZN(n8689) );
  NAND2_X2 U9241 ( .A1(n13170), .A2(n9539), .ZN(n9536) );
  XNOR2_X2 U9242 ( .A(n8830), .B(n8803), .ZN(n13170) );
  NOR2_X2 U9243 ( .A1(n12924), .A2(n12925), .ZN(n12923) );
  AOI21_X2 U9244 ( .B1(n11413), .B2(n11412), .A(n11411), .ZN(n13025) );
  NAND2_X1 U9245 ( .A1(n10506), .A2(n10505), .ZN(n10604) );
  NAND2_X1 U9246 ( .A1(n10526), .A2(n10415), .ZN(n10417) );
  NAND2_X1 U9247 ( .A1(n12994), .A2(n11418), .ZN(n12975) );
  NAND2_X1 U9248 ( .A1(n10690), .A2(n10689), .ZN(n10757) );
  AOI21_X1 U9249 ( .B1(n7424), .B2(n6691), .A(n11414), .ZN(n13003) );
  NOR2_X1 U9250 ( .A1(n8902), .A2(n10052), .ZN(n8865) );
  NAND2_X1 U9251 ( .A1(n12521), .A2(n12517), .ZN(n10015) );
  INV_X1 U9252 ( .A(n10015), .ZN(n10018) );
  NAND2_X1 U9253 ( .A1(n10414), .A2(n10413), .ZN(n10527) );
  NAND2_X1 U9254 ( .A1(n10530), .A2(n12731), .ZN(n10529) );
  OAI21_X1 U9255 ( .B1(n12973), .B2(n11393), .A(n11392), .ZN(n12962) );
  NOR2_X2 U9256 ( .A1(n11334), .A2(n8811), .ZN(n8861) );
  OAI21_X2 U9257 ( .B1(n12906), .B2(n11395), .A(n7336), .ZN(n12902) );
  INV_X1 U9258 ( .A(n14414), .ZN(n6740) );
  OAI21_X1 U9259 ( .B1(n14165), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6680), .ZN(
        n7221) );
  AOI21_X2 U9260 ( .B1(n14679), .B2(n14143), .A(n14410), .ZN(n14145) );
  NOR2_X1 U9261 ( .A1(n14395), .A2(n14394), .ZN(n14137) );
  NAND2_X2 U9262 ( .A1(n6818), .A2(n9482), .ZN(n9680) );
  NAND2_X1 U9263 ( .A1(n7608), .A2(n6806), .ZN(n7619) );
  NAND2_X1 U9264 ( .A1(n6849), .A2(n6847), .ZN(n10947) );
  NAND2_X1 U9265 ( .A1(n14052), .A2(n7223), .ZN(n14097) );
  NAND2_X1 U9266 ( .A1(n7217), .A2(n14173), .ZN(n14177) );
  INV_X1 U9267 ( .A(n7221), .ZN(n14168) );
  OAI21_X1 U9268 ( .B1(n14179), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6682), .ZN(
        n7226) );
  OAI21_X2 U9269 ( .B1(n13233), .B2(n6846), .A(n6844), .ZN(n11546) );
  NAND2_X1 U9270 ( .A1(n9712), .A2(n9711), .ZN(n9746) );
  INV_X1 U9271 ( .A(n12647), .ZN(n6745) );
  INV_X2 U9272 ( .A(n12691), .ZN(n12606) );
  OAI21_X1 U9273 ( .B1(n13677), .B2(n14488), .A(n6799), .ZN(n6798) );
  OAI21_X1 U9274 ( .B1(n13679), .B2(n13525), .A(n6796), .ZN(P1_U3262) );
  INV_X1 U9275 ( .A(n13626), .ZN(n6749) );
  NAND2_X1 U9276 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NAND2_X1 U9277 ( .A1(n8023), .A2(n8022), .ZN(n8037) );
  NAND2_X1 U9278 ( .A1(n6751), .A2(n7605), .ZN(n7175) );
  NAND2_X1 U9279 ( .A1(n7604), .A2(n7536), .ZN(n6751) );
  NAND2_X1 U9280 ( .A1(n8213), .A2(n8212), .ZN(n8482) );
  NAND2_X1 U9281 ( .A1(n8421), .A2(n8420), .ZN(n8419) );
  INV_X1 U9282 ( .A(n8327), .ZN(n6957) );
  NAND2_X1 U9283 ( .A1(n8567), .A2(n8566), .ZN(n8581) );
  INV_X1 U9284 ( .A(n8413), .ZN(n6966) );
  NAND2_X1 U9285 ( .A1(n8188), .A2(n8187), .ZN(n8276) );
  NAND2_X1 U9286 ( .A1(n8717), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U9287 ( .A1(n8643), .A2(n8642), .ZN(n8659) );
  NAND2_X1 U9288 ( .A1(n8378), .A2(n8377), .ZN(n8376) );
  OAI21_X2 U9289 ( .B1(n8436), .B2(n9831), .A(n8208), .ZN(n8451) );
  NAND2_X1 U9290 ( .A1(n8538), .A2(n8537), .ZN(n8540) );
  NAND2_X1 U9291 ( .A1(n8289), .A2(n8288), .ZN(n8193) );
  NAND2_X1 U9292 ( .A1(n11802), .A2(n11801), .ZN(n11803) );
  XNOR2_X1 U9293 ( .A(n7251), .B(n12057), .ZN(n11963) );
  INV_X1 U9294 ( .A(n13058), .ZN(n6781) );
  NAND2_X1 U9295 ( .A1(n6781), .A2(n6779), .ZN(n13144) );
  NAND2_X1 U9296 ( .A1(n7022), .A2(n7021), .ZN(P2_U3496) );
  NAND2_X1 U9297 ( .A1(n6754), .A2(n6765), .ZN(n7988) );
  NAND2_X1 U9298 ( .A1(n7969), .A2(n15288), .ZN(n7971) );
  INV_X1 U9299 ( .A(n7974), .ZN(n6754) );
  NAND2_X1 U9300 ( .A1(n7971), .A2(n7970), .ZN(n7974) );
  INV_X4 U9301 ( .A(n9469), .ZN(n12680) );
  MUX2_X1 U9302 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n9469), .Z(n7642) );
  NAND3_X1 U9303 ( .A1(n7341), .A2(n7927), .A3(n7340), .ZN(n7928) );
  AND2_X1 U9304 ( .A1(n12716), .A2(n12717), .ZN(n6778) );
  INV_X1 U9305 ( .A(n13835), .ZN(n6937) );
  AOI21_X1 U9306 ( .B1(n13502), .B2(n6934), .A(n6684), .ZN(n6933) );
  NAND2_X1 U9307 ( .A1(n7533), .A2(n7532), .ZN(n8709) );
  NAND2_X1 U9308 ( .A1(n8720), .A2(n8736), .ZN(n8723) );
  NAND2_X1 U9309 ( .A1(n11615), .A2(n11685), .ZN(n9393) );
  NAND2_X1 U9310 ( .A1(n6757), .A2(n6755), .ZN(P1_U3527) );
  OR2_X1 U9311 ( .A1(n13992), .A2(n14577), .ZN(n6757) );
  NAND2_X2 U9312 ( .A1(n9506), .A2(n9469), .ZN(n13444) );
  INV_X1 U9313 ( .A(n13690), .ZN(n13703) );
  NAND2_X1 U9314 ( .A1(n6770), .A2(n15138), .ZN(n7341) );
  NAND2_X1 U9315 ( .A1(n6914), .A2(n7875), .ZN(n7911) );
  NAND2_X1 U9316 ( .A1(n7845), .A2(n7844), .ZN(n7861) );
  INV_X1 U9317 ( .A(n7915), .ZN(n6770) );
  OAI21_X1 U9318 ( .B1(n12774), .B2(n12725), .A(n6789), .ZN(n6788) );
  NAND2_X1 U9319 ( .A1(n7861), .A2(n7860), .ZN(n7019) );
  NAND2_X1 U9320 ( .A1(n7822), .A2(n7821), .ZN(n7845) );
  NAND2_X1 U9321 ( .A1(n6867), .A2(n6866), .ZN(n7697) );
  NAND2_X1 U9322 ( .A1(n6771), .A2(n14109), .ZN(n14112) );
  NAND2_X1 U9323 ( .A1(n15389), .A2(n15388), .ZN(n6771) );
  NAND2_X1 U9324 ( .A1(n14140), .A2(n10937), .ZN(n6772) );
  INV_X1 U9325 ( .A(n14406), .ZN(n6773) );
  NOR2_X1 U9326 ( .A1(n14106), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n14055) );
  XNOR2_X1 U9327 ( .A(n7226), .B(n7225), .ZN(SUB_1596_U4) );
  NAND2_X1 U9328 ( .A1(n10019), .A2(n10018), .ZN(n10100) );
  AND2_X2 U9329 ( .A1(n9049), .A2(n8795), .ZN(n7437) );
  INV_X1 U9330 ( .A(n8804), .ZN(n8829) );
  NAND2_X1 U9331 ( .A1(n11439), .A2(n11438), .ZN(n13058) );
  NAND2_X1 U9332 ( .A1(n12718), .A2(n6778), .ZN(n12724) );
  AND2_X2 U9333 ( .A1(n7062), .A2(n7063), .ZN(n8804) );
  NAND2_X1 U9334 ( .A1(n10604), .A2(n12734), .ZN(n10607) );
  INV_X1 U9335 ( .A(n7422), .ZN(n12995) );
  NOR2_X1 U9336 ( .A1(n8055), .A2(n8103), .ZN(n13695) );
  NAND2_X1 U9337 ( .A1(n12724), .A2(n12723), .ZN(n12774) );
  OAI21_X1 U9338 ( .B1(n6635), .B2(n6782), .A(n6786), .ZN(n12718) );
  NAND2_X1 U9339 ( .A1(n7188), .A2(n7187), .ZN(n6782) );
  NAND2_X1 U9340 ( .A1(n12648), .A2(n12649), .ZN(n12652) );
  INV_X1 U9341 ( .A(n6788), .ZN(n12776) );
  OAI22_X1 U9342 ( .A1(n12572), .A2(n6652), .B1(n12571), .B2(n7211), .ZN(
        n12575) );
  NAND3_X1 U9343 ( .A1(n6784), .A2(n6783), .A3(n7209), .ZN(n7208) );
  NAND2_X1 U9344 ( .A1(n12640), .A2(n12639), .ZN(n6783) );
  NAND2_X1 U9345 ( .A1(n12636), .A2(n12635), .ZN(n6784) );
  NAND2_X1 U9346 ( .A1(n6785), .A2(n7195), .ZN(n12564) );
  NAND3_X1 U9347 ( .A1(n12557), .A2(n12556), .A3(n7193), .ZN(n6785) );
  OR2_X1 U9348 ( .A1(n12603), .A2(n12602), .ZN(n12604) );
  AND2_X2 U9349 ( .A1(n8883), .A2(n9048), .ZN(n8796) );
  OAI21_X1 U9350 ( .B1(n13003), .B2(n11416), .A(n7423), .ZN(n7422) );
  INV_X1 U9351 ( .A(n13025), .ZN(n7424) );
  NOR2_X2 U9352 ( .A1(n8866), .A2(n8865), .ZN(n10013) );
  NAND2_X1 U9353 ( .A1(n6795), .A2(n13670), .ZN(n14470) );
  NAND2_X1 U9354 ( .A1(n14446), .A2(n13669), .ZN(n14458) );
  INV_X1 U9355 ( .A(n14457), .ZN(n6794) );
  AND2_X2 U9356 ( .A1(n9683), .A2(n6808), .ZN(n7608) );
  INV_X1 U9357 ( .A(n9878), .ZN(n6824) );
  NAND2_X1 U9358 ( .A1(n13206), .A2(n6828), .ZN(n6825) );
  NAND2_X1 U9359 ( .A1(n6825), .A2(n6826), .ZN(n11531) );
  NAND2_X1 U9360 ( .A1(n7491), .A2(n6623), .ZN(n6832) );
  NAND2_X1 U9361 ( .A1(n6832), .A2(n6833), .ZN(n11485) );
  NAND2_X1 U9362 ( .A1(n13233), .A2(n6841), .ZN(n6837) );
  NAND2_X1 U9363 ( .A1(n6837), .A2(n6838), .ZN(n13181) );
  NAND2_X1 U9364 ( .A1(n13233), .A2(n13234), .ZN(n6843) );
  NAND2_X1 U9365 ( .A1(n10207), .A2(n6850), .ZN(n6849) );
  NAND2_X1 U9366 ( .A1(n10793), .A2(n6853), .ZN(n10795) );
  NOR2_X1 U9367 ( .A1(n10796), .A2(n6852), .ZN(n6851) );
  NAND3_X1 U9368 ( .A1(n6858), .A2(n6860), .A3(n6856), .ZN(n6865) );
  NAND2_X1 U9369 ( .A1(n12457), .A2(n6861), .ZN(n6860) );
  NAND2_X1 U9370 ( .A1(n12457), .A2(n9170), .ZN(n9186) );
  NAND2_X1 U9371 ( .A1(n9185), .A2(n6862), .ZN(n6859) );
  NOR2_X1 U9372 ( .A1(n9185), .A2(n6862), .ZN(n6861) );
  INV_X1 U9373 ( .A(n9185), .ZN(n6863) );
  INV_X1 U9374 ( .A(n6865), .ZN(n11583) );
  AND2_X2 U9375 ( .A1(n6865), .A2(n6864), .ZN(n9190) );
  NAND2_X1 U9376 ( .A1(n7665), .A2(n6869), .ZN(n6867) );
  NOR2_X1 U9378 ( .A1(n11584), .A2(n7036), .ZN(n11591) );
  INV_X2 U9379 ( .A(n14511), .ZN(n14559) );
  NOR2_X2 U9380 ( .A1(n10476), .A2(n14550), .ZN(n14515) );
  NOR2_X2 U9381 ( .A1(n6558), .A2(n14022), .ZN(n13849) );
  NOR2_X2 U9382 ( .A1(n11179), .A2(n13988), .ZN(n6881) );
  NOR2_X2 U9383 ( .A1(n13727), .A2(n13915), .ZN(n11342) );
  NOR2_X2 U9384 ( .A1(n10852), .A2(n14819), .ZN(n11004) );
  NAND2_X1 U9385 ( .A1(n6686), .A2(n11155), .ZN(n13038) );
  NAND2_X2 U9386 ( .A1(n8829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8830) );
  NOR2_X2 U9387 ( .A1(n12868), .A2(n13059), .ZN(n6892) );
  NOR2_X2 U9388 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8883) );
  NAND2_X1 U9389 ( .A1(n6917), .A2(n7955), .ZN(n7959) );
  NAND2_X1 U9390 ( .A1(n7943), .A2(n7942), .ZN(n7957) );
  NAND2_X1 U9391 ( .A1(n7325), .A2(n6922), .ZN(n6920) );
  NAND2_X1 U9392 ( .A1(n6920), .A2(n6628), .ZN(n7326) );
  NAND2_X1 U9393 ( .A1(n7781), .A2(n7780), .ZN(n7799) );
  NAND2_X1 U9394 ( .A1(n9469), .A2(n9502), .ZN(n6932) );
  OAI21_X1 U9395 ( .B1(n9469), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n6932), .ZN(
        n7622) );
  AND2_X1 U9396 ( .A1(n6941), .A2(n6940), .ZN(n6939) );
  NAND2_X2 U9397 ( .A1(n6947), .A2(n7671), .ZN(n13330) );
  NAND2_X1 U9398 ( .A1(n8551), .A2(n6954), .ZN(n6950) );
  NAND2_X1 U9399 ( .A1(n6950), .A2(n6951), .ZN(n8567) );
  OAI21_X2 U9400 ( .B1(n8611), .B2(n8610), .A(n8612), .ZN(n8626) );
  XNOR2_X2 U9401 ( .A(n8060), .B(P1_IR_REG_22__SCAN_IN), .ZN(n13297) );
  NAND3_X1 U9402 ( .A1(n13341), .A2(n7377), .A3(n13340), .ZN(n6973) );
  OR2_X1 U9403 ( .A1(n13415), .A2(n6698), .ZN(n6974) );
  NAND2_X1 U9404 ( .A1(n6974), .A2(n6975), .ZN(n13420) );
  INV_X1 U9405 ( .A(n13420), .ZN(n13423) );
  NAND3_X1 U9406 ( .A1(n13368), .A2(n6981), .A3(n6983), .ZN(n6979) );
  NOR2_X1 U9407 ( .A1(n6984), .A2(n13370), .ZN(n6980) );
  INV_X1 U9408 ( .A(n13382), .ZN(n6983) );
  NAND4_X1 U9409 ( .A1(n13317), .A2(n7376), .A3(n13304), .A4(n6985), .ZN(n7375) );
  NAND3_X1 U9410 ( .A1(n13316), .A2(n6988), .A3(n6987), .ZN(n6986) );
  OAI21_X1 U9411 ( .B1(n6989), .B2(n6670), .A(n6990), .ZN(n13411) );
  INV_X1 U9412 ( .A(n13407), .ZN(n6992) );
  NAND2_X1 U9413 ( .A1(n13325), .A2(n6996), .ZN(n6994) );
  NAND2_X1 U9414 ( .A1(n13325), .A2(n6997), .ZN(n6995) );
  INV_X1 U9415 ( .A(n13323), .ZN(n6999) );
  NAND2_X1 U9416 ( .A1(n13424), .A2(n7003), .ZN(n7002) );
  OAI21_X1 U9417 ( .B1(n7002), .B2(n6668), .A(n7004), .ZN(n13433) );
  INV_X1 U9418 ( .A(n13428), .ZN(n7007) );
  NAND2_X1 U9419 ( .A1(n7566), .A2(n6692), .ZN(n8122) );
  OR2_X1 U9420 ( .A1(n13393), .A2(n7014), .ZN(n7009) );
  NAND2_X1 U9421 ( .A1(n7009), .A2(n7010), .ZN(n7371) );
  NAND3_X1 U9422 ( .A1(n12443), .A2(n12441), .A3(n9282), .ZN(n7024) );
  NAND2_X1 U9423 ( .A1(n7029), .A2(n7027), .ZN(n10501) );
  INV_X1 U9424 ( .A(n7028), .ZN(n7027) );
  OAI21_X1 U9425 ( .B1(n7030), .B2(n12730), .A(n10498), .ZN(n7028) );
  NAND3_X1 U9426 ( .A1(n10431), .A2(n10422), .A3(n10529), .ZN(n7029) );
  NAND2_X1 U9427 ( .A1(n12902), .A2(n6609), .ZN(n7051) );
  OR2_X1 U9428 ( .A1(n12902), .A2(n11396), .ZN(n7052) );
  NAND2_X1 U9429 ( .A1(n7053), .A2(n6687), .ZN(n11391) );
  NAND3_X1 U9430 ( .A1(n7063), .A2(n7437), .A3(n6681), .ZN(n8826) );
  AND2_X2 U9431 ( .A1(n7435), .A2(n7542), .ZN(n7063) );
  NAND2_X1 U9432 ( .A1(n12964), .A2(n7066), .ZN(n7065) );
  NAND2_X1 U9433 ( .A1(n6690), .A2(n7065), .ZN(n12906) );
  NAND2_X1 U9434 ( .A1(n7074), .A2(n7073), .ZN(n10696) );
  INV_X1 U9435 ( .A(n7891), .ZN(n7075) );
  NAND2_X1 U9436 ( .A1(n7075), .A2(n7908), .ZN(n7080) );
  NAND2_X1 U9437 ( .A1(n7076), .A2(n7891), .ZN(n7892) );
  NAND2_X1 U9438 ( .A1(n7891), .A2(n7876), .ZN(n7877) );
  NAND3_X1 U9439 ( .A1(n7080), .A2(n7078), .A3(n7077), .ZN(n10831) );
  NAND3_X1 U9440 ( .A1(n7891), .A2(n7079), .A3(n7081), .ZN(n7078) );
  NAND2_X1 U9441 ( .A1(n7082), .A2(n8161), .ZN(n8290) );
  AND2_X1 U9442 ( .A1(n7506), .A2(n7082), .ZN(n7266) );
  AND2_X1 U9443 ( .A1(n7082), .A2(n8163), .ZN(n7505) );
  INV_X1 U9444 ( .A(n8337), .ZN(n14966) );
  AND2_X2 U9445 ( .A1(n7530), .A2(n8169), .ZN(n8222) );
  OR2_X1 U9446 ( .A1(n12115), .A2(n7097), .ZN(n7088) );
  NAND2_X1 U9447 ( .A1(n7093), .A2(n7089), .ZN(n12078) );
  NAND2_X1 U9448 ( .A1(n12115), .A2(n7094), .ZN(n7093) );
  NAND2_X1 U9449 ( .A1(n12177), .A2(n7104), .ZN(n7102) );
  NAND3_X1 U9450 ( .A1(n7102), .A2(n7101), .A3(n6602), .ZN(n12137) );
  NAND2_X1 U9451 ( .A1(n7112), .A2(n7113), .ZN(n12234) );
  NAND2_X1 U9452 ( .A1(n11234), .A2(n7114), .ZN(n7112) );
  NAND2_X1 U9453 ( .A1(n10972), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U9454 ( .A1(n8706), .A2(n7125), .ZN(n9429) );
  NAND2_X1 U9455 ( .A1(n8706), .A2(n7123), .ZN(n9441) );
  NAND2_X1 U9456 ( .A1(n8706), .A2(n8705), .ZN(n12068) );
  INV_X1 U9457 ( .A(n7131), .ZN(n12222) );
  MUX2_X1 U9458 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n15005), .S(n7132), .Z(n10337) );
  NAND3_X1 U9459 ( .A1(n7136), .A2(P3_IR_REG_2__SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U9460 ( .A1(n10276), .A2(n7142), .ZN(n7139) );
  NAND3_X1 U9461 ( .A1(n7140), .A2(n7137), .A3(n7139), .ZN(n10319) );
  INV_X1 U9462 ( .A(n10276), .ZN(n7138) );
  NAND3_X1 U9463 ( .A1(n7140), .A2(n7141), .A3(n7139), .ZN(n10560) );
  NAND2_X1 U9464 ( .A1(n10335), .A2(n7148), .ZN(n7149) );
  OAI211_X1 U9465 ( .C1(n10335), .C2(n10374), .A(n6604), .B(n7149), .ZN(n10275) );
  INV_X1 U9466 ( .A(n7155), .ZN(n14870) );
  INV_X1 U9467 ( .A(n11986), .ZN(n7154) );
  XNOR2_X1 U9468 ( .A(n11989), .B(n14185), .ZN(n14193) );
  NAND2_X1 U9469 ( .A1(n7650), .A2(n7649), .ZN(n7346) );
  AND3_X4 U9470 ( .A1(n7595), .A2(n7596), .A3(n7597), .ZN(n14543) );
  NOR2_X2 U9471 ( .A1(n10226), .A2(n13330), .ZN(n10225) );
  AND2_X2 U9472 ( .A1(n8124), .A2(n7565), .ZN(n7551) );
  NOR2_X1 U9473 ( .A1(n7287), .A2(n7286), .ZN(n7285) );
  OAI21_X1 U9474 ( .B1(n11289), .B2(n11288), .A(n11287), .ZN(n11383) );
  NAND2_X1 U9475 ( .A1(n10997), .A2(n10996), .ZN(n11027) );
  NAND2_X1 U9476 ( .A1(n11386), .A2(n12752), .ZN(n13037) );
  OAI211_X2 U9477 ( .C1(n12661), .C2(n9475), .A(n8900), .B(n8899), .ZN(n12511)
         );
  NOR2_X2 U9478 ( .A1(n10509), .A2(n12549), .ZN(n10635) );
  NOR2_X2 U9479 ( .A1(n10531), .A2(n12511), .ZN(n10533) );
  NAND2_X1 U9480 ( .A1(n10099), .A2(n10098), .ZN(n10421) );
  NAND2_X1 U9481 ( .A1(n11992), .A2(n6723), .ZN(n11993) );
  OAI211_X1 U9482 ( .C1(n12530), .C2(n7173), .A(n7171), .B(n12529), .ZN(n12533) );
  NAND2_X1 U9483 ( .A1(n7172), .A2(n12532), .ZN(n7171) );
  NAND2_X1 U9484 ( .A1(n7173), .A2(n12530), .ZN(n7172) );
  NAND2_X1 U9485 ( .A1(n12525), .A2(n7174), .ZN(n7173) );
  NAND2_X1 U9486 ( .A1(n12591), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U9487 ( .A1(n12654), .A2(n7183), .ZN(n7188) );
  NAND3_X1 U9488 ( .A1(n12614), .A2(n12613), .A3(n6713), .ZN(n7198) );
  INV_X1 U9489 ( .A(n12615), .ZN(n7199) );
  NAND2_X1 U9490 ( .A1(n12629), .A2(n7204), .ZN(n7203) );
  OR2_X1 U9491 ( .A1(n12643), .A2(n12641), .ZN(n7209) );
  NAND2_X1 U9492 ( .A1(n12643), .A2(n12641), .ZN(n7210) );
  NAND2_X1 U9493 ( .A1(n12575), .A2(n12576), .ZN(n12574) );
  INV_X1 U9494 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7214) );
  NAND2_X1 U9495 ( .A1(n12246), .A2(n7228), .ZN(n7227) );
  NAND2_X1 U9496 ( .A1(n7235), .A2(n7236), .ZN(n12150) );
  NAND2_X1 U9497 ( .A1(n14963), .A2(n7242), .ZN(n7241) );
  OAI21_X1 U9498 ( .B1(n12075), .B2(n7247), .A(n7246), .ZN(n7251) );
  NAND2_X1 U9499 ( .A1(n7252), .A2(n6638), .ZN(n7247) );
  AOI21_X1 U9500 ( .B1(n12075), .B2(n11944), .A(n8771), .ZN(n11768) );
  INV_X1 U9501 ( .A(n11767), .ZN(n7253) );
  NAND2_X1 U9502 ( .A1(n8759), .A2(n6595), .ZN(n7256) );
  NOR2_X2 U9503 ( .A1(n7263), .A2(n7262), .ZN(n7530) );
  NAND4_X1 U9504 ( .A1(n7507), .A2(n7506), .A3(n8163), .A4(n6656), .ZN(n7263)
         );
  NAND4_X1 U9505 ( .A1(n6714), .A2(n7265), .A3(n7507), .A4(n7534), .ZN(n8452)
         );
  NAND2_X1 U9506 ( .A1(n12141), .A2(n7274), .ZN(n7273) );
  NOR2_X2 U9508 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7275) );
  NOR2_X2 U9509 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7825) );
  AND4_X2 U9510 ( .A1(n7825), .A2(n7283), .A3(n7282), .A4(n7281), .ZN(n7280)
         );
  INV_X1 U9512 ( .A(n7619), .ZN(n7284) );
  NAND2_X2 U9513 ( .A1(n7285), .A2(n7288), .ZN(n14041) );
  INV_X1 U9514 ( .A(n7584), .ZN(n7287) );
  NAND2_X1 U9515 ( .A1(n10859), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U9516 ( .A1(n10731), .A2(n8083), .ZN(n7313) );
  AOI21_X1 U9517 ( .B1(n13810), .B2(n6664), .A(n7314), .ZN(n13761) );
  OAI21_X1 U9518 ( .B1(n8093), .B2(n7324), .A(n7321), .ZN(n8094) );
  NAND2_X1 U9519 ( .A1(n7326), .A2(n7328), .ZN(n7781) );
  NAND2_X1 U9520 ( .A1(n7915), .A2(n7344), .ZN(n7927) );
  NAND3_X1 U9521 ( .A1(n7341), .A2(n7342), .A3(n7927), .ZN(n7917) );
  NAND2_X1 U9522 ( .A1(n7348), .A2(n7662), .ZN(n7347) );
  INV_X1 U9523 ( .A(n7348), .ZN(n7351) );
  NAND2_X1 U9524 ( .A1(n11337), .A2(n8035), .ZN(n8055) );
  INV_X1 U9525 ( .A(n11339), .ZN(n7355) );
  NAND2_X1 U9526 ( .A1(n13766), .A2(n13767), .ZN(n13765) );
  AOI21_X2 U9527 ( .B1(n7953), .B2(n7356), .A(n6621), .ZN(n13767) );
  OAI21_X1 U9528 ( .B1(n7360), .B2(n7359), .A(n7858), .ZN(n7358) );
  XNOR2_X2 U9529 ( .A(n14543), .B(n9750), .ZN(n13493) );
  NAND2_X1 U9530 ( .A1(n7371), .A2(n7369), .ZN(n13404) );
  INV_X1 U9531 ( .A(n13342), .ZN(n7378) );
  OAI22_X1 U9532 ( .A1(n7379), .A2(n6648), .B1(n7381), .B2(n13332), .ZN(n13336) );
  NAND2_X1 U9533 ( .A1(n13329), .A2(n7380), .ZN(n7379) );
  INV_X1 U9534 ( .A(n13331), .ZN(n7381) );
  OAI22_X1 U9535 ( .A1(n7382), .A2(n6659), .B1(n7384), .B2(n13365), .ZN(n13369) );
  NAND2_X1 U9536 ( .A1(n13362), .A2(n7383), .ZN(n7382) );
  INV_X1 U9537 ( .A(n13364), .ZN(n7384) );
  NAND2_X1 U9538 ( .A1(n13351), .A2(n7386), .ZN(n7385) );
  OAI22_X1 U9539 ( .A1(n7385), .A2(n6663), .B1(n7387), .B2(n13354), .ZN(n13358) );
  INV_X1 U9540 ( .A(n13353), .ZN(n7387) );
  NAND2_X1 U9541 ( .A1(n7388), .A2(n7389), .ZN(n9063) );
  NAND2_X1 U9542 ( .A1(n10882), .A2(n6683), .ZN(n7388) );
  AOI21_X1 U9543 ( .B1(n6683), .B2(n10883), .A(n6600), .ZN(n7389) );
  NOR2_X2 U9544 ( .A1(n11161), .A2(n7395), .ZN(n11299) );
  NAND2_X1 U9545 ( .A1(n8882), .A2(n9863), .ZN(n7398) );
  XNOR2_X1 U9546 ( .A(n8878), .B(n8879), .ZN(n9863) );
  NAND2_X1 U9547 ( .A1(n8882), .A2(n6626), .ZN(n7397) );
  NAND2_X1 U9548 ( .A1(n7398), .A2(n7396), .ZN(n9982) );
  AND2_X1 U9549 ( .A1(n7397), .A2(n9974), .ZN(n7396) );
  NAND2_X1 U9550 ( .A1(n9919), .A2(n7399), .ZN(n10036) );
  NAND2_X1 U9551 ( .A1(n8941), .A2(n9913), .ZN(n9919) );
  INV_X1 U9552 ( .A(n7401), .ZN(n7407) );
  NAND2_X1 U9553 ( .A1(n8980), .A2(n7413), .ZN(n7412) );
  AOI21_X1 U9554 ( .B1(n8995), .B2(n7414), .A(n6601), .ZN(n7413) );
  INV_X1 U9555 ( .A(n14300), .ZN(n7421) );
  OAI21_X1 U9556 ( .B1(n9082), .B2(n7420), .A(n6603), .ZN(n9127) );
  NAND2_X1 U9557 ( .A1(n8861), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8863) );
  OAI211_X1 U9558 ( .C1(n12961), .C2(n7432), .A(n7428), .B(n11421), .ZN(n7426)
         );
  NAND2_X1 U9559 ( .A1(n7427), .A2(n7425), .ZN(n11422) );
  INV_X1 U9560 ( .A(n7426), .ZN(n7425) );
  NAND2_X1 U9561 ( .A1(n12975), .A2(n7430), .ZN(n7427) );
  AND4_X2 U9562 ( .A1(n9050), .A2(n8796), .A3(n8795), .A4(n9049), .ZN(n8818)
         );
  INV_X1 U9563 ( .A(n8818), .ZN(n9084) );
  NAND2_X1 U9564 ( .A1(n10607), .A2(n10606), .ZN(n10629) );
  INV_X1 U9565 ( .A(n10691), .ZN(n10690) );
  OR2_X1 U9566 ( .A1(n10608), .A2(n12558), .ZN(n7446) );
  OAI22_X1 U9567 ( .A1(n7451), .A2(n7449), .B1(n12907), .B2(n7447), .ZN(n12862) );
  INV_X1 U9568 ( .A(n11423), .ZN(n7454) );
  NAND2_X1 U9569 ( .A1(n12862), .A2(n12861), .ZN(n12860) );
  NAND2_X1 U9570 ( .A1(n12888), .A2(n12695), .ZN(n7456) );
  OAI21_X1 U9571 ( .B1(n13225), .B2(n7474), .A(n7473), .ZN(n13199) );
  NAND2_X1 U9572 ( .A1(n11546), .A2(n11545), .ZN(n13279) );
  AND4_X4 U9573 ( .A1(n7587), .A2(n7589), .A3(n7588), .A4(n7590), .ZN(n9750)
         );
  NOR2_X1 U9574 ( .A1(n9750), .A2(n13311), .ZN(n13301) );
  NAND2_X1 U9575 ( .A1(n7486), .A2(n13311), .ZN(n13312) );
  XNOR2_X1 U9576 ( .A(n10465), .B(n7486), .ZN(n10460) );
  NAND2_X1 U9577 ( .A1(n13591), .A2(n7486), .ZN(n7485) );
  OR2_X2 U9578 ( .A1(n11360), .A2(n7488), .ZN(n13438) );
  INV_X1 U9579 ( .A(n11360), .ZN(n7489) );
  XNOR2_X1 U9580 ( .A(n11485), .B(n11483), .ZN(n13290) );
  NAND2_X1 U9581 ( .A1(n7566), .A2(n7551), .ZN(n7583) );
  NAND3_X1 U9582 ( .A1(n7566), .A2(n7551), .A3(n7502), .ZN(n7569) );
  AND3_X1 U9583 ( .A1(n7507), .A2(n7506), .A3(n7505), .ZN(n8396) );
  NAND2_X1 U9584 ( .A1(n11728), .A2(n7509), .ZN(n7508) );
  OAI211_X1 U9585 ( .C1(n11728), .C2(n7511), .A(n7508), .B(n11730), .ZN(n9428)
         );
  AOI21_X1 U9586 ( .B1(n6594), .B2(n11675), .A(n6675), .ZN(n7518) );
  NAND3_X1 U9587 ( .A1(n9388), .A2(n12154), .A3(n11685), .ZN(n11615) );
  OAI21_X2 U9588 ( .B1(n11271), .B2(n11267), .A(n11268), .ZN(n11375) );
  OAI21_X2 U9589 ( .B1(n11304), .B2(n9359), .A(n9358), .ZN(n11271) );
  OAI21_X2 U9590 ( .B1(n8723), .B2(P3_D_REG_0__SCAN_IN), .A(n8722), .ZN(n9308)
         );
  NAND2_X1 U9591 ( .A1(n9384), .A2(n9385), .ZN(n11704) );
  NAND2_X1 U9592 ( .A1(n9429), .A2(n15072), .ZN(n8779) );
  NAND2_X1 U9593 ( .A1(n10896), .A2(n8386), .ZN(n10972) );
  NAND2_X1 U9594 ( .A1(n12774), .A2(n12771), .ZN(n12772) );
  XNOR2_X1 U9595 ( .A(n11353), .B(n11352), .ZN(n13454) );
  OAI21_X1 U9596 ( .B1(n9307), .B2(n12440), .A(n9306), .ZN(P2_U3186) );
  OAI21_X1 U9597 ( .B1(n6636), .B2(n12126), .A(n12124), .ZN(n12276) );
  XNOR2_X1 U9598 ( .A(n9031), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12812) );
  CLKBUF_X1 U9599 ( .A(n10018), .Z(n12728) );
  NAND2_X1 U9600 ( .A1(n8087), .A2(n13511), .ZN(n8090) );
  AND4_X2 U9601 ( .A1(n7578), .A2(n7577), .A3(n7576), .A4(n7575), .ZN(n10462)
         );
  INV_X1 U9602 ( .A(n8717), .ZN(n8718) );
  NAND2_X1 U9603 ( .A1(n9285), .A2(n9284), .ZN(n9283) );
  NAND2_X1 U9604 ( .A1(n6564), .A2(n9309), .ZN(n9313) );
  XNOR2_X1 U9605 ( .A(n9705), .B(n11476), .ZN(n9744) );
  OR2_X1 U9606 ( .A1(n6562), .A2(n13575), .ZN(n7587) );
  AOI22_X2 U9607 ( .A1(n12137), .A2(n12140), .B1(n12281), .B2(n11617), .ZN(
        n12127) );
  AND2_X1 U9608 ( .A1(n10259), .A2(n6590), .ZN(n14929) );
  INV_X1 U9609 ( .A(n13513), .ZN(n13840) );
  AND2_X1 U9610 ( .A1(n8422), .A2(n8437), .ZN(n7534) );
  AND2_X2 U9611 ( .A1(n10585), .A2(n8747), .ZN(n15072) );
  OR2_X1 U9612 ( .A1(n13109), .A2(n12787), .ZN(n7535) );
  INV_X1 U9613 ( .A(n12752), .ZN(n13034) );
  AND2_X1 U9614 ( .A1(n11562), .A2(n11561), .ZN(n7537) );
  OR2_X1 U9615 ( .A1(n9342), .A2(n11126), .ZN(n7538) );
  AND2_X1 U9616 ( .A1(n12714), .A2(n12713), .ZN(n7539) );
  AND2_X1 U9617 ( .A1(n7556), .A2(n8152), .ZN(n7540) );
  AND2_X1 U9618 ( .A1(n13470), .A2(n7553), .ZN(n7541) );
  OR2_X1 U9619 ( .A1(n9536), .A2(n8859), .ZN(n7543) );
  AND2_X1 U9620 ( .A1(n11473), .A2(n11472), .ZN(n7544) );
  AND2_X1 U9621 ( .A1(n7780), .A2(n7766), .ZN(n7545) );
  OR2_X1 U9622 ( .A1(n8122), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n7546) );
  OR2_X1 U9623 ( .A1(n9302), .A2(n9281), .ZN(n14302) );
  INV_X1 U9624 ( .A(n14302), .ZN(n9282) );
  AND2_X1 U9625 ( .A1(n9366), .A2(n12240), .ZN(n7547) );
  AND2_X1 U9626 ( .A1(n8234), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7548) );
  INV_X1 U9627 ( .A(n12196), .ZN(n8535) );
  INV_X1 U9628 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13159) );
  AND2_X1 U9629 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7549) );
  INV_X1 U9630 ( .A(n12945), .ZN(n12978) );
  AND2_X1 U9631 ( .A1(n7800), .A2(n7785), .ZN(n7550) );
  INV_X2 U9632 ( .A(n14521), .ZN(n14536) );
  AND2_X1 U9633 ( .A1(n9300), .A2(n9299), .ZN(n12692) );
  INV_X2 U9634 ( .A(n14600), .ZN(n14598) );
  NOR2_X2 U9635 ( .A1(n8155), .A2(n8154), .ZN(n14597) );
  NOR2_X1 U9636 ( .A1(n9961), .A2(n9960), .ZN(n9990) );
  INV_X1 U9637 ( .A(n12719), .ZN(n12664) );
  OR2_X1 U9638 ( .A1(n13469), .A2(n13468), .ZN(n7553) );
  AND2_X1 U9639 ( .A1(n11502), .A2(n11501), .ZN(n7555) );
  INV_X1 U9640 ( .A(n13065), .ZN(n12872) );
  OR2_X1 U9641 ( .A1(n13429), .A2(n14028), .ZN(n7556) );
  AND2_X1 U9642 ( .A1(n10402), .A2(n10219), .ZN(n7557) );
  XNOR2_X1 U9643 ( .A(n8901), .B(n6560), .ZN(n8878) );
  INV_X1 U9644 ( .A(n14983), .ZN(n8753) );
  OR2_X1 U9645 ( .A1(n12073), .A2(n12405), .ZN(n7559) );
  OR2_X1 U9646 ( .A1(n12073), .A2(n12325), .ZN(n7560) );
  INV_X1 U9647 ( .A(n11772), .ZN(n11801) );
  AND2_X1 U9648 ( .A1(n11135), .A2(n11134), .ZN(n7561) );
  INV_X1 U9649 ( .A(n12520), .ZN(n12518) );
  AND3_X1 U9650 ( .A1(n13315), .A2(n13314), .A3(n13299), .ZN(n13316) );
  NAND2_X1 U9651 ( .A1(n12569), .A2(n12568), .ZN(n12572) );
  OAI21_X1 U9652 ( .B1(n7554), .B2(n13390), .A(n13389), .ZN(n13393) );
  INV_X1 U9653 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U9654 ( .A1(n12783), .A2(n12719), .ZN(n12665) );
  INV_X1 U9655 ( .A(n12692), .ZN(n11425) );
  INV_X1 U9656 ( .A(n9171), .ZN(n7954) );
  INV_X1 U9657 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8544) );
  INV_X1 U9658 ( .A(n11797), .ZN(n8683) );
  INV_X1 U9659 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8164) );
  AND2_X1 U9660 ( .A1(n13114), .A2(n11415), .ZN(n11416) );
  INV_X1 U9661 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8794) );
  AND2_X1 U9662 ( .A1(n13520), .A2(n13699), .ZN(n13521) );
  INV_X1 U9663 ( .A(n14951), .ZN(n9345) );
  AND2_X1 U9664 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  NOR2_X1 U9665 ( .A1(n11766), .A2(n12063), .ZN(n8704) );
  OR2_X1 U9666 ( .A1(n8723), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8725) );
  INV_X1 U9667 ( .A(n9168), .ZN(n9169) );
  NAND2_X1 U9668 ( .A1(n12715), .A2(n7539), .ZN(n12716) );
  INV_X1 U9669 ( .A(n9292), .ZN(n9294) );
  INV_X1 U9670 ( .A(n9118), .ZN(n8783) );
  INV_X1 U9671 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8986) );
  INV_X1 U9672 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8897) );
  INV_X1 U9673 ( .A(n11563), .ZN(n9963) );
  INV_X1 U9674 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7733) );
  INV_X1 U9675 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7672) );
  INV_X1 U9676 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7562) );
  INV_X1 U9677 ( .A(SI_16_), .ZN(n8484) );
  INV_X1 U9678 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7683) );
  NAND2_X1 U9679 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  INV_X1 U9680 ( .A(n8617), .ZN(n8616) );
  OR2_X1 U9681 ( .A1(n8589), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8602) );
  OR2_X1 U9682 ( .A1(n8572), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8589) );
  OR2_X1 U9683 ( .A1(n8510), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8527) );
  INV_X1 U9684 ( .A(SI_22_), .ZN(n8569) );
  NOR2_X1 U9685 ( .A1(n8427), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U9686 ( .A1(n9314), .A2(n11980), .ZN(n11833) );
  AND2_X1 U9687 ( .A1(n8725), .A2(n8724), .ZN(n10581) );
  INV_X1 U9688 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8221) );
  AND2_X1 U9689 ( .A1(n8215), .A2(n8214), .ZN(n8480) );
  AND2_X1 U9690 ( .A1(n9471), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8189) );
  OR2_X1 U9691 ( .A1(n14317), .A2(n11207), .ZN(n9125) );
  NAND2_X1 U9692 ( .A1(n9167), .A2(n9169), .ZN(n9170) );
  AND2_X1 U9693 ( .A1(n9294), .A2(n9235), .ZN(n12884) );
  NAND2_X1 U9694 ( .A1(n8784), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9160) );
  OR2_X1 U9695 ( .A1(n8970), .A2(n10121), .ZN(n8987) );
  AND2_X1 U9696 ( .A1(n14649), .A2(n10918), .ZN(n14658) );
  OAI21_X1 U9697 ( .B1(n12692), .B2(n13004), .A(n11436), .ZN(n11437) );
  OR2_X1 U9698 ( .A1(n8987), .A2(n8986), .ZN(n9004) );
  AND2_X1 U9699 ( .A1(n6619), .A2(n9244), .ZN(n9275) );
  INV_X1 U9700 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8819) );
  NOR2_X1 U9701 ( .A1(n10187), .A2(n10186), .ZN(n10189) );
  NAND2_X1 U9702 ( .A1(n9708), .A2(n9952), .ZN(n9709) );
  INV_X1 U9703 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n15166) );
  INV_X1 U9704 ( .A(n11056), .ZN(n11057) );
  INV_X1 U9705 ( .A(n7963), .ZN(n7964) );
  INV_X1 U9706 ( .A(n13939), .ZN(n8119) );
  AND2_X1 U9707 ( .A1(n7754), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U9708 ( .A1(n7959), .A2(n7958), .ZN(n7970) );
  INV_X1 U9709 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n15352) );
  INV_X1 U9710 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14059) );
  NOR2_X1 U9711 ( .A1(n14092), .A2(n14093), .ZN(n14074) );
  AND2_X1 U9712 ( .A1(n10242), .A2(n8698), .ZN(n10248) );
  NOR2_X1 U9713 ( .A1(n8527), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8545) );
  OR2_X1 U9714 ( .A1(n11607), .A2(n9338), .ZN(n9339) );
  NAND2_X1 U9715 ( .A1(n8616), .A2(n8615), .ZN(n8631) );
  INV_X1 U9716 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10559) );
  INV_X1 U9717 ( .A(n12224), .ZN(n11711) );
  OR2_X1 U9718 ( .A1(n8631), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8648) );
  INV_X1 U9719 ( .A(n9311), .ZN(n11960) );
  INV_X1 U9720 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11669) );
  INV_X1 U9721 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n11368) );
  AND2_X1 U9722 ( .A1(n10250), .A2(n10248), .ZN(n10259) );
  INV_X1 U9723 ( .A(n11971), .ZN(n12139) );
  INV_X1 U9724 ( .A(n11977), .ZN(n12239) );
  INV_X1 U9725 ( .A(n11978), .ZN(n12251) );
  OR2_X1 U9726 ( .A1(n8317), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8339) );
  INV_X1 U9727 ( .A(n15072), .ZN(n8777) );
  INV_X1 U9728 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9439) );
  AND2_X1 U9729 ( .A1(n11881), .A2(n11886), .ZN(n12247) );
  OR2_X1 U9730 ( .A1(n14267), .A2(n14274), .ZN(n11871) );
  INV_X1 U9731 ( .A(n12131), .ZN(n15038) );
  INV_X1 U9732 ( .A(n11966), .ZN(n11805) );
  AND2_X1 U9733 ( .A1(n9037), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9055) );
  OR2_X1 U9734 ( .A1(n9204), .A2(n12474), .ZN(n9216) );
  INV_X1 U9735 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9909) );
  INV_X1 U9736 ( .A(n10985), .ZN(n9081) );
  OR2_X1 U9737 ( .A1(n12870), .A2(n11403), .ZN(n9300) );
  INV_X1 U9738 ( .A(n11403), .ZN(n9236) );
  OR2_X1 U9739 ( .A1(n14647), .A2(n14646), .ZN(n14649) );
  INV_X1 U9740 ( .A(n13044), .ZN(n13018) );
  NAND2_X1 U9741 ( .A1(n14751), .A2(n9287), .ZN(n13041) );
  INV_X1 U9742 ( .A(n14797), .ZN(n14818) );
  INV_X1 U9743 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9245) );
  NOR2_X1 U9744 ( .A1(n7836), .A2(n15166), .ZN(n7854) );
  NOR2_X1 U9745 ( .A1(n13246), .A2(n7921), .ZN(n7936) );
  NAND2_X1 U9746 ( .A1(n11055), .A2(n11057), .ZN(n11058) );
  OR2_X1 U9747 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  OR2_X1 U9748 ( .A1(n9688), .A2(n13543), .ZN(n14360) );
  NAND2_X1 U9749 ( .A1(n7885), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7898) );
  AND2_X1 U9750 ( .A1(n7868), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7885) );
  OR2_X1 U9751 ( .A1(n9612), .A2(n13589), .ZN(n14475) );
  INV_X1 U9752 ( .A(n13519), .ZN(n8103) );
  INV_X1 U9753 ( .A(n13726), .ZN(n13751) );
  NAND2_X1 U9754 ( .A1(n13780), .A2(n8119), .ZN(n13781) );
  INV_X1 U9755 ( .A(n13780), .ZN(n13798) );
  INV_X1 U9756 ( .A(n13825), .ZN(n13834) );
  INV_X1 U9757 ( .A(n9689), .ZN(n9690) );
  INV_X1 U9758 ( .A(n13543), .ZN(n10077) );
  NAND2_X1 U9759 ( .A1(n14577), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8152) );
  INV_X1 U9760 ( .A(n13808), .ZN(n13821) );
  OR2_X1 U9761 ( .A1(n9985), .A2(n13477), .ZN(n10089) );
  INV_X1 U9762 ( .A(n14585), .ZN(n14505) );
  INV_X1 U9763 ( .A(n14549), .ZN(n14582) );
  INV_X1 U9764 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8058) );
  NOR2_X1 U9765 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14110), .ZN(n14061) );
  AND2_X1 U9766 ( .A1(n9408), .A2(n10238), .ZN(n11730) );
  INV_X1 U9767 ( .A(n15075), .ZN(n9756) );
  NOR2_X1 U9768 ( .A1(n14219), .A2(n14220), .ZN(n14218) );
  OR2_X1 U9769 ( .A1(n10588), .A2(n14999), .ZN(n14268) );
  AND2_X1 U9770 ( .A1(n11948), .A2(n8701), .ZN(n14977) );
  INV_X1 U9771 ( .A(n12134), .ZN(n14253) );
  INV_X1 U9772 ( .A(n15010), .ZN(n14991) );
  NAND2_X1 U9773 ( .A1(n10586), .A2(n14999), .ZN(n15010) );
  AND2_X1 U9774 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  OR2_X1 U9775 ( .A1(n12131), .A2(n15049), .ZN(n15054) );
  AND2_X1 U9776 ( .A1(n14999), .A2(n11805), .ZN(n15049) );
  OR2_X1 U9777 ( .A1(n9436), .A2(n9435), .ZN(n9437) );
  NOR2_X1 U9778 ( .A1(n9757), .A2(n9756), .ZN(n9759) );
  XNOR2_X1 U9779 ( .A(n8690), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U9780 ( .A1(n8376), .A2(n8201), .ZN(n8395) );
  NAND2_X1 U9781 ( .A1(n9055), .A2(n8781), .ZN(n9100) );
  NAND2_X1 U9782 ( .A1(n12459), .A2(n12458), .ZN(n12457) );
  NAND2_X1 U9783 ( .A1(n9288), .A2(n13041), .ZN(n14328) );
  OR2_X1 U9784 ( .A1(n9552), .A2(n6777), .ZN(n14695) );
  INV_X1 U9785 ( .A(n14695), .ZN(n14715) );
  AND2_X1 U9786 ( .A1(n14639), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14719) );
  INV_X1 U9787 ( .A(n12762), .ZN(n12842) );
  XNOR2_X1 U9788 ( .A(n13059), .B(n11409), .ZN(n12760) );
  INV_X1 U9789 ( .A(n13047), .ZN(n13023) );
  INV_X1 U9790 ( .A(n13004), .ZN(n13029) );
  INV_X1 U9791 ( .A(n14750), .ZN(n9739) );
  OR2_X1 U9792 ( .A1(n12882), .A2(n12881), .ZN(n13075) );
  OR2_X1 U9793 ( .A1(n12725), .A2(n12778), .ZN(n14822) );
  INV_X1 U9794 ( .A(n13140), .ZN(n14787) );
  AND2_X1 U9795 ( .A1(n14752), .A2(n9738), .ZN(n10030) );
  AND2_X1 U9796 ( .A1(n13174), .A2(n9257), .ZN(n14724) );
  OR2_X1 U9797 ( .A1(n13174), .A2(n9258), .ZN(n9259) );
  XNOR2_X1 U9798 ( .A(n9278), .B(n9277), .ZN(n11172) );
  INV_X1 U9799 ( .A(n14369), .ZN(n13293) );
  INV_X1 U9800 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14116) );
  OR2_X1 U9801 ( .A1(n9612), .A2(n9601), .ZN(n14488) );
  INV_X1 U9802 ( .A(n14488), .ZN(n14468) );
  INV_X1 U9803 ( .A(n13884), .ZN(n14513) );
  INV_X1 U9804 ( .A(n13888), .ZN(n14517) );
  INV_X1 U9805 ( .A(n13991), .ZN(n14590) );
  OR2_X1 U9806 ( .A1(n10078), .A2(n8142), .ZN(n8155) );
  AND2_X1 U9807 ( .A1(n9680), .A2(n9486), .ZN(n9691) );
  XNOR2_X1 U9808 ( .A(n7642), .B(SI_3_), .ZN(n7640) );
  INV_X1 U9809 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14122) );
  AND2_X1 U9810 ( .A1(n10250), .A2(n10249), .ZN(n14860) );
  INV_X1 U9811 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U9812 ( .A1(n9409), .A2(n10586), .ZN(n11737) );
  INV_X1 U9813 ( .A(n12102), .ZN(n12079) );
  NOR2_X1 U9814 ( .A1(n9446), .A2(n9756), .ZN(n11973) );
  INV_X1 U9815 ( .A(n14860), .ZN(n14936) );
  INV_X1 U9816 ( .A(n14192), .ZN(n14945) );
  OR2_X1 U9817 ( .A1(n14268), .A2(n14988), .ZN(n12134) );
  AND2_X1 U9818 ( .A1(n15013), .A2(n10776), .ZN(n14269) );
  NAND2_X2 U9819 ( .A1(n10588), .A2(n15010), .ZN(n14995) );
  NAND2_X1 U9820 ( .A1(n15072), .A2(n15054), .ZN(n12325) );
  OR2_X1 U9821 ( .A1(n15056), .A2(n14288), .ZN(n12405) );
  INV_X1 U9822 ( .A(SI_25_), .ZN(n10835) );
  INV_X1 U9823 ( .A(SI_20_), .ZN(n15138) );
  INV_X1 U9824 ( .A(SI_14_), .ZN(n9784) );
  INV_X1 U9825 ( .A(n10677), .ZN(n10675) );
  OR2_X1 U9826 ( .A1(n9302), .A2(n12777), .ZN(n12438) );
  INV_X1 U9827 ( .A(n12594), .ZN(n14340) );
  INV_X1 U9828 ( .A(n14328), .ZN(n14310) );
  INV_X1 U9829 ( .A(P2_U3947), .ZN(n12795) );
  INV_X1 U9830 ( .A(P2_U3947), .ZN(n12804) );
  INV_X1 U9831 ( .A(n14719), .ZN(n14621) );
  AND2_X1 U9832 ( .A1(n10927), .A2(n10926), .ZN(n12819) );
  OR2_X1 U9833 ( .A1(n9546), .A2(P2_U3088), .ZN(n14722) );
  AND2_X2 U9834 ( .A1(n10030), .A2(n9739), .ZN(n14842) );
  OR3_X1 U9835 ( .A1(n13123), .A2(n13122), .A3(n13121), .ZN(n13155) );
  INV_X1 U9836 ( .A(n14829), .ZN(n14827) );
  INV_X1 U9837 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15260) );
  XNOR2_X1 U9838 ( .A(n9250), .B(n9249), .ZN(n11175) );
  INV_X1 U9839 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10832) );
  INV_X1 U9840 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9698) );
  INV_X1 U9841 ( .A(n13352), .ZN(n10967) );
  AND2_X1 U9842 ( .A1(n9871), .A2(n13546), .ZN(n14369) );
  NAND2_X1 U9843 ( .A1(n9510), .A2(n9508), .ZN(n14499) );
  OR2_X1 U9844 ( .A1(n14521), .A2(n13481), .ZN(n13877) );
  NAND2_X1 U9845 ( .A1(n8150), .A2(n14549), .ZN(n14028) );
  OR2_X1 U9846 ( .A1(n8155), .A2(n8149), .ZN(n14577) );
  INV_X1 U9847 ( .A(n14537), .ZN(n14538) );
  INV_X1 U9848 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9561) );
  AND2_X1 U9849 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9538), .ZN(P2_U3947) );
  NOR2_X1 U9850 ( .A1(n9680), .A2(n9445), .ZN(P1_U4016) );
  NAND2_X1 U9851 ( .A1(n8153), .A2(n7540), .ZN(P1_U3524) );
  NOR2_X1 U9852 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7564) );
  NOR3_X1 U9854 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U9855 ( .A1(n7569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7571) );
  NAND2_X1 U9856 ( .A1(n13439), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7578) );
  INV_X1 U9857 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7572) );
  OR2_X1 U9858 ( .A1(n6562), .A2(n7572), .ZN(n7577) );
  INV_X1 U9859 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7573) );
  OR2_X1 U9860 ( .A1(n13442), .A2(n7573), .ZN(n7576) );
  INV_X1 U9861 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7574) );
  OR2_X1 U9862 ( .A1(n13438), .A2(n7574), .ZN(n7575) );
  AND2_X1 U9863 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7579) );
  NAND2_X1 U9864 ( .A1(n9469), .A2(n7579), .ZN(n7591) );
  INV_X1 U9865 ( .A(SI_0_), .ZN(n9463) );
  INV_X1 U9866 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8242) );
  OAI21_X1 U9867 ( .B1(n12680), .B2(n9463), .A(n8242), .ZN(n7580) );
  AND2_X1 U9868 ( .A1(n7591), .A2(n7580), .ZN(n14051) );
  XNOR2_X2 U9869 ( .A(n7582), .B(n7581), .ZN(n8115) );
  MUX2_X1 U9870 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14051), .S(n9506), .Z(n9986)
         );
  NOR2_X1 U9871 ( .A1(n10462), .A2(n14526), .ZN(n10459) );
  INV_X1 U9872 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7585) );
  OR2_X1 U9873 ( .A1(n7980), .A2(n7585), .ZN(n7590) );
  INV_X1 U9874 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7586) );
  INV_X1 U9875 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13575) );
  XNOR2_X1 U9876 ( .A(n7605), .B(SI_1_), .ZN(n7593) );
  INV_X1 U9877 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9520) );
  MUX2_X1 U9878 ( .A(n9520), .B(n9526), .S(n12680), .Z(n7592) );
  XNOR2_X1 U9879 ( .A(n7593), .B(n7592), .ZN(n9525) );
  AND2_X4 U9880 ( .A1(n9506), .A2(n12680), .ZN(n13474) );
  NAND2_X1 U9881 ( .A1(n13474), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9882 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7594) );
  NAND2_X1 U9883 ( .A1(n7894), .A2(n13577), .ZN(n7595) );
  NAND2_X1 U9884 ( .A1(n9750), .A2(n14543), .ZN(n13313) );
  NAND2_X1 U9885 ( .A1(n7991), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7603) );
  INV_X1 U9886 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13594) );
  OR2_X1 U9887 ( .A1(n6562), .A2(n13594), .ZN(n7602) );
  INV_X1 U9888 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7598) );
  INV_X1 U9889 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7599) );
  OR2_X1 U9890 ( .A1(n7980), .A2(n7599), .ZN(n7600) );
  XNOR2_X1 U9891 ( .A(n7622), .B(SI_2_), .ZN(n7625) );
  AOI21_X1 U9892 ( .B1(n12680), .B2(P1_DATAO_REG_1__SCAN_IN), .A(SI_1_), .ZN(
        n7604) );
  NAND2_X1 U9893 ( .A1(n12680), .A2(n9526), .ZN(n7606) );
  OAI211_X1 U9894 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n12680), .A(n7606), .B(
        SI_1_), .ZN(n7607) );
  XNOR2_X1 U9895 ( .A(n7625), .B(n7624), .ZN(n9501) );
  NAND2_X1 U9896 ( .A1(n13474), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7610) );
  NAND2_X1 U9897 ( .A1(n7894), .A2(n13596), .ZN(n7609) );
  OAI211_X2 U9898 ( .C1(n13444), .C2(n9501), .A(n7610), .B(n7609), .ZN(n14550)
         );
  NAND2_X1 U9899 ( .A1(n7611), .A2(n14550), .ZN(n13314) );
  NAND2_X1 U9900 ( .A1(n10483), .A2(n13495), .ZN(n7613) );
  NAND2_X1 U9901 ( .A1(n7611), .A2(n10480), .ZN(n7612) );
  NAND2_X1 U9902 ( .A1(n13434), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7618) );
  INV_X1 U9903 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14509) );
  OR2_X1 U9904 ( .A1(n13438), .A2(n14509), .ZN(n7617) );
  OR2_X1 U9905 ( .A1(n6562), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7616) );
  INV_X1 U9906 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7614) );
  OR2_X1 U9907 ( .A1(n7980), .A2(n7614), .ZN(n7615) );
  NAND2_X1 U9908 ( .A1(n7619), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7621) );
  INV_X1 U9909 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7620) );
  XNOR2_X1 U9910 ( .A(n7621), .B(n7620), .ZN(n13606) );
  OAI22_X1 U9911 ( .A1(n7790), .A2(n9476), .B1(n9506), .B2(n13606), .ZN(n7627)
         );
  INV_X1 U9912 ( .A(SI_2_), .ZN(n9467) );
  NOR2_X1 U9913 ( .A1(n7622), .A2(n9467), .ZN(n7623) );
  XNOR2_X1 U9914 ( .A(n7641), .B(n7640), .ZN(n9475) );
  NOR2_X1 U9915 ( .A1(n9475), .A2(n13444), .ZN(n7626) );
  OR2_X2 U9916 ( .A1(n7627), .A2(n7626), .ZN(n14511) );
  NAND2_X1 U9917 ( .A1(n9877), .A2(n14511), .ZN(n13318) );
  NAND2_X1 U9918 ( .A1(n14559), .A2(n13572), .ZN(n13319) );
  NAND2_X1 U9919 ( .A1(n14501), .A2(n14502), .ZN(n7629) );
  NAND2_X1 U9920 ( .A1(n9877), .A2(n14559), .ZN(n7628) );
  NAND2_X1 U9921 ( .A1(n7629), .A2(n7628), .ZN(n10084) );
  NAND2_X1 U9922 ( .A1(n13439), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7639) );
  INV_X1 U9923 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7630) );
  OR2_X1 U9924 ( .A1(n13438), .A2(n7630), .ZN(n7638) );
  AND2_X1 U9925 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7657) );
  INV_X1 U9926 ( .A(n7657), .ZN(n7634) );
  INV_X1 U9927 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7632) );
  INV_X1 U9928 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U9929 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  NAND2_X1 U9930 ( .A1(n7634), .A2(n7633), .ZN(n10090) );
  OR2_X1 U9931 ( .A1(n6562), .A2(n10090), .ZN(n7637) );
  INV_X1 U9932 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7635) );
  OR2_X1 U9933 ( .A1(n13442), .A2(n7635), .ZN(n7636) );
  NAND2_X1 U9934 ( .A1(n7642), .A2(SI_3_), .ZN(n7643) );
  MUX2_X1 U9935 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n12680), .Z(n7651) );
  XNOR2_X1 U9936 ( .A(n7651), .B(SI_4_), .ZN(n7648) );
  XNOR2_X1 U9937 ( .A(n7650), .B(n7648), .ZN(n9477) );
  NAND2_X1 U9938 ( .A1(n9477), .A2(n13472), .ZN(n7646) );
  NAND2_X1 U9939 ( .A1(n7653), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7644) );
  XNOR2_X1 U9940 ( .A(n7644), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U9941 ( .A1(n13474), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7894), .B2(
        n13626), .ZN(n7645) );
  OR2_X1 U9942 ( .A1(n13571), .A2(n13322), .ZN(n10083) );
  INV_X1 U9943 ( .A(n10083), .ZN(n7647) );
  NAND2_X1 U9944 ( .A1(n13322), .A2(n13571), .ZN(n10082) );
  INV_X1 U9945 ( .A(n7648), .ZN(n7649) );
  NAND2_X1 U9946 ( .A1(n7651), .A2(SI_4_), .ZN(n7652) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n12680), .Z(n7666) );
  XNOR2_X1 U9948 ( .A(n7666), .B(SI_5_), .ZN(n7663) );
  XNOR2_X1 U9949 ( .A(n7665), .B(n7663), .ZN(n9488) );
  NAND2_X1 U9950 ( .A1(n9488), .A2(n13472), .ZN(n7656) );
  OR2_X1 U9951 ( .A1(n7669), .A2(n14033), .ZN(n7654) );
  XNOR2_X1 U9952 ( .A(n7654), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9633) );
  AOI22_X1 U9953 ( .A1(n13474), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7894), .B2(
        n9633), .ZN(n7655) );
  NAND2_X1 U9954 ( .A1(n13439), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9955 ( .A1(n7991), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9956 ( .A1(n7657), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7673) );
  OAI21_X1 U9957 ( .B1(n7657), .B2(P1_REG3_REG_5__SCAN_IN), .A(n7673), .ZN(
        n10131) );
  OR2_X1 U9958 ( .A1(n6562), .A2(n10131), .ZN(n7659) );
  INV_X1 U9959 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9608) );
  OR2_X1 U9960 ( .A1(n13442), .A2(n9608), .ZN(n7658) );
  NAND4_X1 U9961 ( .A1(n7661), .A2(n7660), .A3(n7659), .A4(n7658), .ZN(n13570)
         );
  OR2_X1 U9962 ( .A1(n14571), .A2(n13570), .ZN(n7662) );
  INV_X1 U9963 ( .A(n7663), .ZN(n7664) );
  NAND2_X1 U9964 ( .A1(n7666), .A2(SI_5_), .ZN(n7667) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n12680), .Z(n7682) );
  XNOR2_X1 U9966 ( .A(n7682), .B(SI_6_), .ZN(n7680) );
  OR2_X1 U9967 ( .A1(n7684), .A2(n14033), .ZN(n7670) );
  XNOR2_X1 U9968 ( .A(n7670), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9622) );
  AOI22_X1 U9969 ( .A1(n13474), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7894), .B2(
        n9622), .ZN(n7671) );
  NAND2_X1 U9970 ( .A1(n7991), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U9971 ( .A1(n13434), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U9972 ( .A1(n13439), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7676) );
  AND2_X1 U9973 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  NOR2_X1 U9974 ( .A1(n7673), .A2(n7672), .ZN(n7688) );
  OR2_X1 U9975 ( .A1(n7674), .A2(n7688), .ZN(n10490) );
  OR2_X1 U9976 ( .A1(n6562), .A2(n10490), .ZN(n7675) );
  NAND4_X1 U9977 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), .ZN(n13569)
         );
  XNOR2_X1 U9978 ( .A(n13330), .B(n13569), .ZN(n13498) );
  OR2_X1 U9979 ( .A1(n13330), .A2(n13569), .ZN(n7679) );
  NAND2_X1 U9980 ( .A1(n10223), .A2(n7679), .ZN(n10157) );
  MUX2_X1 U9981 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n12680), .Z(n7698) );
  XNOR2_X1 U9982 ( .A(n7698), .B(SI_7_), .ZN(n7695) );
  XNOR2_X1 U9983 ( .A(n7697), .B(n7695), .ZN(n9516) );
  NAND2_X1 U9984 ( .A1(n9516), .A2(n13472), .ZN(n7687) );
  NAND2_X1 U9985 ( .A1(n7684), .A2(n7683), .ZN(n7701) );
  NAND2_X1 U9986 ( .A1(n7701), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7685) );
  XNOR2_X1 U9987 ( .A(n7685), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U9988 ( .A1(n13474), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7894), .B2(
        n9672), .ZN(n7686) );
  NAND2_X1 U9989 ( .A1(n7687), .A2(n7686), .ZN(n13333) );
  NAND2_X1 U9990 ( .A1(n13439), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9991 ( .A1(n7991), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9992 ( .A1(n13434), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9993 ( .A1(n7688), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7721) );
  OR2_X1 U9994 ( .A1(n7688), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9995 ( .A1(n7721), .A2(n7689), .ZN(n10211) );
  OR2_X1 U9996 ( .A1(n6562), .A2(n10211), .ZN(n7690) );
  NAND4_X1 U9997 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n13568)
         );
  XNOR2_X1 U9998 ( .A(n13333), .B(n13568), .ZN(n13500) );
  INV_X1 U9999 ( .A(n13500), .ZN(n10156) );
  OR2_X1 U10000 ( .A1(n13333), .A2(n13568), .ZN(n7694) );
  INV_X1 U10001 ( .A(n7695), .ZN(n7696) );
  NAND2_X1 U10002 ( .A1(n7697), .A2(n7696), .ZN(n7700) );
  NAND2_X1 U10003 ( .A1(n7698), .A2(SI_7_), .ZN(n7699) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n12680), .Z(n7712) );
  XNOR2_X1 U10005 ( .A(n7712), .B(SI_8_), .ZN(n7709) );
  XNOR2_X1 U10006 ( .A(n7711), .B(n7709), .ZN(n9528) );
  NAND2_X1 U10007 ( .A1(n9528), .A2(n13472), .ZN(n7704) );
  NAND2_X1 U10008 ( .A1(n7714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U10009 ( .A(n7702), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10010 ( .A1(n13474), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7894), 
        .B2(n9814), .ZN(n7703) );
  NAND2_X1 U10011 ( .A1(n13439), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U10012 ( .A1(n7991), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7707) );
  INV_X1 U10013 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7719) );
  XNOR2_X1 U10014 ( .A(n7721), .B(n7719), .ZN(n10788) );
  OR2_X1 U10015 ( .A1(n6562), .A2(n10788), .ZN(n7706) );
  INV_X1 U10016 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9667) );
  OR2_X1 U10017 ( .A1(n13442), .A2(n9667), .ZN(n7705) );
  NAND4_X1 U10018 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n13567) );
  INV_X1 U10019 ( .A(n13567), .ZN(n8080) );
  INV_X1 U10020 ( .A(n7709), .ZN(n7710) );
  NAND2_X1 U10021 ( .A1(n7712), .A2(SI_8_), .ZN(n7713) );
  INV_X4 U10022 ( .A(n9474), .ZN(n8042) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8042), .Z(n7729) );
  XNOR2_X1 U10024 ( .A(n7728), .B(n6924), .ZN(n9557) );
  NAND2_X1 U10025 ( .A1(n9557), .A2(n13472), .ZN(n7717) );
  NAND2_X1 U10026 ( .A1(n7730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7715) );
  XNOR2_X1 U10027 ( .A(n7715), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9894) );
  AOI22_X1 U10028 ( .A1(n7894), .A2(n9894), .B1(n13474), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U10029 ( .A1(n13439), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10030 ( .A1(n7991), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7725) );
  INV_X1 U10031 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7718) );
  OAI21_X1 U10032 ( .B1(n7721), .B2(n7719), .A(n7718), .ZN(n7722) );
  NAND2_X1 U10033 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n7720) );
  NAND2_X1 U10034 ( .A1(n7722), .A2(n7734), .ZN(n11042) );
  OR2_X1 U10035 ( .A1(n6562), .A2(n11042), .ZN(n7724) );
  INV_X1 U10036 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9807) );
  OR2_X1 U10037 ( .A1(n13442), .A2(n9807), .ZN(n7723) );
  NAND4_X1 U10038 ( .A1(n7726), .A2(n7725), .A3(n7724), .A4(n7723), .ZN(n13566) );
  INV_X1 U10039 ( .A(n13566), .ZN(n10962) );
  XNOR2_X1 U10040 ( .A(n13345), .B(n10962), .ZN(n13503) );
  OR2_X1 U10041 ( .A1(n13345), .A2(n13566), .ZN(n7727) );
  NAND2_X1 U10042 ( .A1(n10644), .A2(n7727), .ZN(n10726) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8042), .Z(n7744) );
  XNOR2_X1 U10044 ( .A(n7744), .B(SI_10_), .ZN(n7741) );
  XNOR2_X1 U10045 ( .A(n7743), .B(n7741), .ZN(n9654) );
  NAND2_X1 U10046 ( .A1(n9654), .A2(n13472), .ZN(n7732) );
  XNOR2_X1 U10047 ( .A(n7750), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U10048 ( .A1(n10067), .A2(n7894), .B1(n13474), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10049 ( .A1(n13439), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U10050 ( .A1(n7991), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10051 ( .A1(n13434), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7737) );
  AND2_X1 U10052 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  OR2_X1 U10053 ( .A1(n7735), .A2(n7754), .ZN(n10957) );
  OR2_X1 U10054 ( .A1(n6562), .A2(n10957), .ZN(n7736) );
  NAND4_X1 U10055 ( .A1(n7739), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n13565) );
  INV_X1 U10056 ( .A(n13565), .ZN(n10953) );
  XNOR2_X1 U10057 ( .A(n13352), .B(n10953), .ZN(n13504) );
  NAND2_X1 U10058 ( .A1(n10726), .A2(n13504), .ZN(n10725) );
  OR2_X1 U10059 ( .A1(n13352), .A2(n13565), .ZN(n7740) );
  INV_X1 U10060 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U10061 ( .A1(n7744), .A2(SI_10_), .ZN(n7745) );
  MUX2_X1 U10062 ( .A(n9701), .B(n9698), .S(n8042), .Z(n7746) );
  NAND2_X1 U10063 ( .A1(n7746), .A2(n15182), .ZN(n7761) );
  INV_X1 U10064 ( .A(n7746), .ZN(n7747) );
  NAND2_X1 U10065 ( .A1(n7747), .A2(SI_11_), .ZN(n7748) );
  NAND2_X1 U10066 ( .A1(n7761), .A2(n7748), .ZN(n7762) );
  XNOR2_X1 U10067 ( .A(n7763), .B(n7762), .ZN(n9696) );
  NAND2_X1 U10068 ( .A1(n9696), .A2(n13472), .ZN(n7753) );
  INV_X1 U10069 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U10070 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  NAND2_X1 U10071 ( .A1(n7751), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7768) );
  XNOR2_X1 U10072 ( .A(n7768), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U10073 ( .A1(n13642), .A2(n7894), .B1(n13474), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n7752) );
  NAND2_X1 U10074 ( .A1(n13439), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10075 ( .A1(n7991), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7758) );
  NOR2_X1 U10076 ( .A1(n7754), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7755) );
  OR2_X1 U10077 ( .A1(n7772), .A2(n7755), .ZN(n11064) );
  OR2_X1 U10078 ( .A1(n6562), .A2(n11064), .ZN(n7757) );
  INV_X1 U10079 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10061) );
  OR2_X1 U10080 ( .A1(n13442), .A2(n10061), .ZN(n7756) );
  NAND4_X1 U10081 ( .A1(n7759), .A2(n7758), .A3(n7757), .A4(n7756), .ZN(n13564) );
  XNOR2_X1 U10082 ( .A(n13355), .B(n13564), .ZN(n13505) );
  INV_X1 U10083 ( .A(n13505), .ZN(n10813) );
  NAND2_X1 U10084 ( .A1(n10814), .A2(n10813), .ZN(n10812) );
  OR2_X1 U10085 ( .A1(n13355), .A2(n13564), .ZN(n7760) );
  NAND2_X1 U10086 ( .A1(n10812), .A2(n7760), .ZN(n10872) );
  MUX2_X1 U10087 ( .A(n9788), .B(n9790), .S(n8042), .Z(n7764) );
  NAND2_X1 U10088 ( .A1(n7764), .A2(n15245), .ZN(n7780) );
  INV_X1 U10089 ( .A(n7764), .ZN(n7765) );
  NAND2_X1 U10090 ( .A1(n7765), .A2(SI_12_), .ZN(n7766) );
  XNOR2_X1 U10091 ( .A(n7779), .B(n7545), .ZN(n9786) );
  NAND2_X1 U10092 ( .A1(n9786), .A2(n13472), .ZN(n7771) );
  INV_X1 U10093 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U10094 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  NAND2_X1 U10095 ( .A1(n7769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7786) );
  XNOR2_X1 U10096 ( .A(n7786), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U10097 ( .A1(n13666), .A2(n7894), .B1(n13474), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U10098 ( .A1(n13439), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7777) );
  INV_X1 U10099 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10867) );
  OR2_X1 U10100 ( .A1(n13438), .A2(n10867), .ZN(n7776) );
  OR2_X1 U10101 ( .A1(n7772), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10102 ( .A1(n7809), .A2(n7773), .ZN(n11141) );
  OR2_X1 U10103 ( .A1(n6562), .A2(n11141), .ZN(n7775) );
  INV_X1 U10104 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n13640) );
  OR2_X1 U10105 ( .A1(n13442), .A2(n13640), .ZN(n7774) );
  NAND4_X1 U10106 ( .A1(n7777), .A2(n7776), .A3(n7775), .A4(n7774), .ZN(n13563) );
  XNOR2_X1 U10107 ( .A(n13363), .B(n13563), .ZN(n13506) );
  INV_X1 U10108 ( .A(n13506), .ZN(n10871) );
  NAND2_X1 U10109 ( .A1(n10872), .A2(n10871), .ZN(n10870) );
  OR2_X1 U10110 ( .A1(n13363), .A2(n13563), .ZN(n7778) );
  MUX2_X1 U10111 ( .A(n9828), .B(n9831), .S(n8042), .Z(n7783) );
  NAND2_X1 U10112 ( .A1(n7783), .A2(n7782), .ZN(n7800) );
  INV_X1 U10113 ( .A(n7783), .ZN(n7784) );
  NAND2_X1 U10114 ( .A1(n7784), .A2(SI_13_), .ZN(n7785) );
  XNOR2_X1 U10115 ( .A(n7799), .B(n7550), .ZN(n9826) );
  NAND2_X1 U10116 ( .A1(n9826), .A2(n13472), .ZN(n7793) );
  AOI21_X1 U10117 ( .B1(n7786), .B2(n15289), .A(n14033), .ZN(n7787) );
  NAND2_X1 U10118 ( .A1(n7787), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n7789) );
  INV_X1 U10119 ( .A(n7787), .ZN(n7788) );
  NAND2_X1 U10120 ( .A1(n7788), .A2(n15352), .ZN(n7802) );
  NOR2_X1 U10121 ( .A1(n7790), .A2(n9828), .ZN(n7791) );
  AOI21_X1 U10122 ( .B1(n14425), .B2(n7894), .A(n7791), .ZN(n7792) );
  NAND2_X1 U10123 ( .A1(n7991), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U10124 ( .A1(n13434), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U10125 ( .A1(n13439), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7795) );
  INV_X1 U10126 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U10127 ( .A(n7809), .B(n7808), .ZN(n13252) );
  OR2_X1 U10128 ( .A1(n6562), .A2(n13252), .ZN(n7794) );
  NAND4_X1 U10129 ( .A1(n7797), .A2(n7796), .A3(n7795), .A4(n7794), .ZN(n13562) );
  XNOR2_X1 U10130 ( .A(n13366), .B(n13562), .ZN(n13508) );
  INV_X1 U10131 ( .A(n13508), .ZN(n11078) );
  NAND2_X1 U10132 ( .A1(n11079), .A2(n11078), .ZN(n11077) );
  OR2_X1 U10133 ( .A1(n13366), .A2(n13562), .ZN(n7798) );
  MUX2_X1 U10134 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8042), .Z(n7816) );
  XNOR2_X1 U10135 ( .A(n7817), .B(n7816), .ZN(n9927) );
  NAND2_X1 U10136 ( .A1(n9927), .A2(n13472), .ZN(n7805) );
  NAND2_X1 U10137 ( .A1(n7802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7803) );
  AOI22_X1 U10138 ( .A1(n13667), .A2(n7894), .B1(n13474), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U10139 ( .A1(n13439), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7814) );
  INV_X1 U10140 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7806) );
  OR2_X1 U10141 ( .A1(n13438), .A2(n7806), .ZN(n7813) );
  INV_X1 U10142 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7807) );
  OAI21_X1 U10143 ( .B1(n7809), .B2(n7808), .A(n7807), .ZN(n7810) );
  NAND2_X1 U10144 ( .A1(n7810), .A2(n7836), .ZN(n14372) );
  OR2_X1 U10145 ( .A1(n14372), .A2(n6562), .ZN(n7812) );
  INV_X1 U10146 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13651) );
  OR2_X1 U10147 ( .A1(n13442), .A2(n13651), .ZN(n7811) );
  OR2_X1 U10148 ( .A1(n14370), .A2(n11464), .ZN(n13372) );
  NAND2_X1 U10149 ( .A1(n14370), .A2(n11464), .ZN(n13373) );
  INV_X1 U10150 ( .A(n11464), .ZN(n13561) );
  NAND2_X1 U10151 ( .A1(n14370), .A2(n13561), .ZN(n7815) );
  MUX2_X1 U10152 ( .A(n10045), .B(n10047), .S(n8042), .Z(n7818) );
  INV_X1 U10153 ( .A(n7818), .ZN(n7819) );
  NAND2_X1 U10154 ( .A1(n7819), .A2(SI_15_), .ZN(n7820) );
  OR2_X1 U10155 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NAND2_X1 U10156 ( .A1(n7845), .A2(n7823), .ZN(n10044) );
  NAND2_X1 U10157 ( .A1(n10044), .A2(n13472), .ZN(n7835) );
  INV_X1 U10158 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7824) );
  AND4_X1 U10159 ( .A1(n7825), .A2(n15289), .A3(n15352), .A4(n7824), .ZN(n7826) );
  INV_X1 U10160 ( .A(n7831), .ZN(n7828) );
  NAND2_X1 U10161 ( .A1(n7828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7829) );
  MUX2_X1 U10162 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7829), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n7832) );
  INV_X1 U10163 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10164 ( .A1(n7831), .A2(n7830), .ZN(n7850) );
  NAND2_X1 U10165 ( .A1(n7832), .A2(n7850), .ZN(n14445) );
  OAI22_X1 U10166 ( .A1(n14445), .A2(n9506), .B1(n7790), .B2(n10045), .ZN(
        n7833) );
  INV_X1 U10167 ( .A(n7833), .ZN(n7834) );
  AND2_X1 U10168 ( .A1(n7836), .A2(n15166), .ZN(n7837) );
  OR2_X1 U10169 ( .A1(n7837), .A2(n7854), .ZN(n11096) );
  NAND2_X1 U10170 ( .A1(n13434), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7838) );
  OAI21_X1 U10171 ( .B1(n11096), .B2(n6562), .A(n7838), .ZN(n7842) );
  INV_X1 U10172 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10173 ( .A1(n13439), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7839) );
  OAI21_X1 U10174 ( .B1(n7840), .B2(n13438), .A(n7839), .ZN(n7841) );
  NOR2_X1 U10175 ( .A1(n7842), .A2(n7841), .ZN(n11478) );
  NAND2_X1 U10176 ( .A1(n14384), .A2(n11478), .ZN(n13379) );
  NAND2_X1 U10177 ( .A1(n13378), .A2(n13379), .ZN(n13510) );
  INV_X1 U10178 ( .A(n13510), .ZN(n11101) );
  INV_X1 U10179 ( .A(n11478), .ZN(n13560) );
  OR2_X1 U10180 ( .A1(n14384), .A2(n13560), .ZN(n7843) );
  MUX2_X1 U10181 ( .A(n10154), .B(n10185), .S(n8042), .Z(n7846) );
  INV_X1 U10182 ( .A(n7846), .ZN(n7847) );
  NAND2_X1 U10183 ( .A1(n7847), .A2(SI_16_), .ZN(n7848) );
  XNOR2_X1 U10184 ( .A(n7861), .B(n7860), .ZN(n10152) );
  NAND2_X1 U10185 ( .A1(n10152), .A2(n13472), .ZN(n7853) );
  NAND2_X1 U10186 ( .A1(n7850), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7849) );
  MUX2_X1 U10187 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7849), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n7851) );
  AND2_X1 U10188 ( .A1(n7851), .A2(n7879), .ZN(n14461) );
  AOI22_X1 U10189 ( .A1(n14461), .A2(n7894), .B1(n13474), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n7852) );
  NOR2_X1 U10190 ( .A1(n7854), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7855) );
  OR2_X1 U10191 ( .A1(n7868), .A2(n7855), .ZN(n14368) );
  AOI22_X1 U10192 ( .A1(n13434), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n13439), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U10193 ( .A1(n7991), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7856) );
  OAI211_X1 U10194 ( .C1(n14368), .C2(n6562), .A(n7857), .B(n7856), .ZN(n13559) );
  NAND2_X1 U10195 ( .A1(n13988), .A2(n13559), .ZN(n7858) );
  OR2_X1 U10196 ( .A1(n13988), .A2(n13559), .ZN(n7859) );
  MUX2_X1 U10197 ( .A(n15334), .B(n10412), .S(n8042), .Z(n7873) );
  XNOR2_X1 U10198 ( .A(n7873), .B(SI_17_), .ZN(n7863) );
  XNOR2_X1 U10199 ( .A(n7874), .B(n7863), .ZN(n10398) );
  NAND2_X1 U10200 ( .A1(n10398), .A2(n13472), .ZN(n7867) );
  NAND2_X1 U10201 ( .A1(n7879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7864) );
  XNOR2_X1 U10202 ( .A(n7864), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13671) );
  NOR2_X1 U10203 ( .A1(n7790), .A2(n15334), .ZN(n7865) );
  AOI21_X1 U10204 ( .B1(n13671), .B2(n7894), .A(n7865), .ZN(n7866) );
  NOR2_X1 U10205 ( .A1(n7868), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7869) );
  OR2_X1 U10206 ( .A1(n7885), .A2(n7869), .ZN(n13228) );
  AOI22_X1 U10207 ( .A1(n7991), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13434), 
        .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10208 ( .A1(n13439), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7870) );
  OAI211_X1 U10209 ( .C1(n13228), .C2(n6562), .A(n7871), .B(n7870), .ZN(n13865) );
  NOR2_X1 U10210 ( .A1(n13979), .A2(n13865), .ZN(n13392) );
  NAND2_X1 U10211 ( .A1(n13979), .A2(n13865), .ZN(n7872) );
  NAND2_X1 U10212 ( .A1(n7874), .A2(n9866), .ZN(n7875) );
  NAND2_X1 U10213 ( .A1(n7911), .A2(n9972), .ZN(n7876) );
  MUX2_X1 U10214 ( .A(n10724), .B(n10713), .S(n8042), .Z(n7906) );
  NAND2_X1 U10215 ( .A1(n7877), .A2(n7906), .ZN(n7878) );
  OAI21_X1 U10216 ( .B1(n7879), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7881) );
  INV_X1 U10217 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7880) );
  XNOR2_X1 U10218 ( .A(n7881), .B(n7880), .ZN(n14491) );
  OAI22_X1 U10219 ( .A1(n14491), .A2(n9506), .B1(n7790), .B2(n10724), .ZN(
        n7882) );
  INV_X1 U10220 ( .A(n7882), .ZN(n7883) );
  OR2_X1 U10221 ( .A1(n7885), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10222 ( .A1(n7898), .A2(n7886), .ZN(n13870) );
  AOI22_X1 U10223 ( .A1(n7991), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13439), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n7888) );
  INV_X1 U10224 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14479) );
  OR2_X1 U10225 ( .A1(n13442), .A2(n14479), .ZN(n7887) );
  OAI211_X1 U10226 ( .C1(n13870), .C2(n6562), .A(n7888), .B(n7887), .ZN(n13558) );
  NAND2_X1 U10227 ( .A1(n13873), .A2(n13558), .ZN(n13394) );
  INV_X1 U10228 ( .A(n13394), .ZN(n7890) );
  NOR2_X1 U10229 ( .A1(n13873), .A2(n13558), .ZN(n13396) );
  INV_X1 U10230 ( .A(n13396), .ZN(n7889) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8042), .Z(n7912) );
  XNOR2_X1 U10232 ( .A(n7912), .B(SI_19_), .ZN(n7908) );
  NAND2_X1 U10233 ( .A1(n10831), .A2(n13472), .ZN(n7896) );
  NAND2_X1 U10234 ( .A1(n8057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7893) );
  XNOR2_X2 U10235 ( .A(n7893), .B(P1_IR_REG_19__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U10236 ( .A1(n13474), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13525), 
        .B2(n7894), .ZN(n7895) );
  INV_X1 U10237 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10238 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  AND2_X1 U10239 ( .A1(n7921), .A2(n7899), .ZN(n13850) );
  INV_X1 U10240 ( .A(n6562), .ZN(n7925) );
  INV_X1 U10241 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13661) );
  NAND2_X1 U10242 ( .A1(n13439), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10243 ( .A1(n7991), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7900) );
  OAI211_X1 U10244 ( .C1(n13661), .C2(n13442), .A(n7901), .B(n7900), .ZN(n7902) );
  AOI21_X1 U10245 ( .B1(n13850), .B2(n7925), .A(n7902), .ZN(n13271) );
  OR2_X1 U10246 ( .A1(n14022), .A2(n13271), .ZN(n13397) );
  NAND2_X1 U10247 ( .A1(n14022), .A2(n13271), .ZN(n13398) );
  NAND2_X1 U10248 ( .A1(n13839), .A2(n13840), .ZN(n7904) );
  INV_X1 U10249 ( .A(n13271), .ZN(n13557) );
  OR2_X1 U10250 ( .A1(n14022), .A2(n13557), .ZN(n7903) );
  INV_X1 U10251 ( .A(n7906), .ZN(n7905) );
  NOR2_X1 U10252 ( .A1(n7905), .A2(SI_18_), .ZN(n7910) );
  NOR2_X1 U10253 ( .A1(n7906), .A2(n9972), .ZN(n7907) );
  NOR2_X1 U10254 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  INV_X1 U10255 ( .A(n7912), .ZN(n7913) );
  NAND2_X1 U10256 ( .A1(n7913), .A2(n15339), .ZN(n7914) );
  INV_X1 U10257 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10830) );
  MUX2_X1 U10258 ( .A(n10830), .B(n15175), .S(n8042), .Z(n7916) );
  NAND2_X1 U10259 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  NAND2_X1 U10260 ( .A1(n7928), .A2(n7918), .ZN(n11592) );
  NAND2_X1 U10261 ( .A1(n13474), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7919) );
  AOI21_X1 U10262 ( .B1(n7921), .B2(n13246), .A(n7936), .ZN(n13826) );
  INV_X1 U10263 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U10264 ( .A1(n13439), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10265 ( .A1(n13434), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7922) );
  OAI211_X1 U10266 ( .C1(n13438), .C2(n13829), .A(n7923), .B(n7922), .ZN(n7924) );
  AOI21_X1 U10267 ( .B1(n13826), .B2(n7925), .A(n7924), .ZN(n13400) );
  XNOR2_X1 U10268 ( .A(n14018), .B(n13400), .ZN(n13825) );
  OR2_X1 U10269 ( .A1(n13831), .A2(n13400), .ZN(n7926) );
  NAND2_X1 U10270 ( .A1(n7928), .A2(n7927), .ZN(n7932) );
  MUX2_X1 U10271 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n12680), .Z(n7929) );
  NAND2_X1 U10272 ( .A1(n7929), .A2(SI_21_), .ZN(n7942) );
  OAI21_X1 U10273 ( .B1(SI_21_), .B2(n7929), .A(n7942), .ZN(n7930) );
  INV_X1 U10274 ( .A(n7930), .ZN(n7931) );
  OR2_X1 U10275 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U10276 ( .A1(n7943), .A2(n7933), .ZN(n10970) );
  OR2_X1 U10277 ( .A1(n10970), .A2(n13444), .ZN(n7935) );
  NAND2_X1 U10278 ( .A1(n13474), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10279 ( .A1(n7991), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7940) );
  NAND2_X1 U10280 ( .A1(n13439), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10281 ( .A1(n13434), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U10282 ( .A1(n7936), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7945) );
  OAI21_X1 U10283 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n7936), .A(n7945), .ZN(
        n13814) );
  OR2_X1 U10284 ( .A1(n6562), .A2(n13814), .ZN(n7937) );
  NAND4_X1 U10285 ( .A1(n7940), .A2(n7939), .A3(n7938), .A4(n7937), .ZN(n13555) );
  INV_X1 U10286 ( .A(n13555), .ZN(n8095) );
  XNOR2_X1 U10287 ( .A(n13950), .B(n8095), .ZN(n13808) );
  OR2_X1 U10288 ( .A1(n13950), .A2(n13555), .ZN(n7941) );
  XNOR2_X1 U10289 ( .A(n7957), .B(SI_22_), .ZN(n9172) );
  OR2_X1 U10290 ( .A1(n9172), .A2(n12680), .ZN(n7944) );
  NAND2_X1 U10291 ( .A1(n7991), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10292 ( .A1(n13434), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10293 ( .A1(n13439), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10294 ( .A1(n7946), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7963) );
  OAI21_X1 U10295 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n7946), .A(n7963), .ZN(
        n13802) );
  OR2_X1 U10296 ( .A1(n6562), .A2(n13802), .ZN(n7947) );
  NAND4_X1 U10297 ( .A1(n7950), .A2(n7949), .A3(n7948), .A4(n7947), .ZN(n13554) );
  NAND2_X1 U10298 ( .A1(n13268), .A2(n13554), .ZN(n7951) );
  OR2_X1 U10299 ( .A1(n13946), .A2(n13554), .ZN(n7952) );
  MUX2_X1 U10300 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n12680), .Z(n9171) );
  NOR2_X1 U10301 ( .A1(n7954), .A2(n8569), .ZN(n7956) );
  NAND2_X1 U10302 ( .A1(n7954), .A2(n8569), .ZN(n7955) );
  INV_X1 U10303 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8582) );
  INV_X1 U10304 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n15285) );
  MUX2_X1 U10305 ( .A(n8582), .B(n15285), .S(n12680), .Z(n7958) );
  NAND2_X1 U10306 ( .A1(n7969), .A2(n7970), .ZN(n7960) );
  NAND2_X1 U10307 ( .A1(n11171), .A2(n13472), .ZN(n7962) );
  NAND2_X1 U10308 ( .A1(n13474), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10309 ( .A1(n13439), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U10310 ( .A1(n7991), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10311 ( .A1(n7964), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7978) );
  OAI21_X1 U10312 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n7964), .A(n7978), .ZN(
        n13783) );
  OR2_X1 U10313 ( .A1(n6562), .A2(n13783), .ZN(n7966) );
  INV_X1 U10314 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15349) );
  OR2_X1 U10315 ( .A1(n13442), .A2(n15349), .ZN(n7965) );
  NAND4_X1 U10316 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n13553) );
  MUX2_X1 U10317 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8042), .Z(n7972) );
  NAND2_X1 U10318 ( .A1(n7972), .A2(SI_24_), .ZN(n7987) );
  OAI21_X1 U10319 ( .B1(SI_24_), .B2(n7972), .A(n7987), .ZN(n7973) );
  NAND2_X1 U10320 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  NAND2_X1 U10321 ( .A1(n7988), .A2(n7975), .ZN(n11202) );
  OR2_X1 U10322 ( .A1(n11202), .A2(n13444), .ZN(n7977) );
  NAND2_X1 U10323 ( .A1(n13474), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10324 ( .A1(n7991), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10325 ( .A1(n13434), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U10326 ( .A1(n7979), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7992) );
  OAI21_X1 U10327 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7979), .A(n7992), .ZN(
        n13770) );
  OR2_X1 U10328 ( .A1(n6562), .A2(n13770), .ZN(n7982) );
  INV_X1 U10329 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15217) );
  OR2_X1 U10330 ( .A1(n7980), .A2(n15217), .ZN(n7981) );
  NAND4_X1 U10331 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n13552) );
  XNOR2_X1 U10332 ( .A(n14011), .B(n13552), .ZN(n13760) );
  INV_X1 U10333 ( .A(n13760), .ZN(n13766) );
  INV_X1 U10334 ( .A(n14011), .ZN(n8120) );
  INV_X1 U10335 ( .A(n13552), .ZN(n7985) );
  NAND2_X1 U10336 ( .A1(n8120), .A2(n7985), .ZN(n7986) );
  AND2_X2 U10337 ( .A1(n13765), .A2(n7986), .ZN(n13743) );
  MUX2_X1 U10338 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n8042), .Z(n7999) );
  XNOR2_X1 U10339 ( .A(n7999), .B(SI_25_), .ZN(n8002) );
  XNOR2_X1 U10340 ( .A(n8003), .B(n8002), .ZN(n13176) );
  NAND2_X1 U10341 ( .A1(n13176), .A2(n13472), .ZN(n7990) );
  NAND2_X1 U10342 ( .A1(n13474), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10343 ( .A1(n13439), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U10344 ( .A1(n7991), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10345 ( .A1(n13434), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10346 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n7993), .ZN(n8009) );
  OAI21_X1 U10347 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n7993), .A(n8009), .ZN(
        n13752) );
  OR2_X1 U10348 ( .A1(n6562), .A2(n13752), .ZN(n7994) );
  NAND4_X1 U10349 ( .A1(n7997), .A2(n7996), .A3(n7995), .A4(n7994), .ZN(n13551) );
  XNOR2_X1 U10350 ( .A(n14007), .B(n13551), .ZN(n13516) );
  NAND2_X1 U10351 ( .A1(n14007), .A2(n13551), .ZN(n7998) );
  NAND2_X1 U10352 ( .A1(n13742), .A2(n7998), .ZN(n13725) );
  INV_X1 U10353 ( .A(n7999), .ZN(n8000) );
  NAND2_X1 U10354 ( .A1(n8000), .A2(n10835), .ZN(n8001) );
  INV_X1 U10355 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14046) );
  INV_X1 U10356 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15293) );
  MUX2_X1 U10357 ( .A(n14046), .B(n15293), .S(n8042), .Z(n8017) );
  XNOR2_X1 U10358 ( .A(n8017), .B(SI_26_), .ZN(n8004) );
  NAND2_X1 U10359 ( .A1(n13173), .A2(n13472), .ZN(n8006) );
  NAND2_X1 U10360 ( .A1(n13474), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U10361 ( .A1(n13439), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10362 ( .A1(n7991), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10363 ( .A1(n13434), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8012) );
  INV_X1 U10364 ( .A(n8009), .ZN(n8007) );
  NAND2_X1 U10365 ( .A1(n8007), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8029) );
  INV_X1 U10366 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10367 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  NAND2_X1 U10368 ( .A1(n8029), .A2(n8010), .ZN(n13730) );
  OR2_X1 U10369 ( .A1(n6562), .A2(n13730), .ZN(n8011) );
  NAND4_X1 U10370 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n13550) );
  INV_X1 U10371 ( .A(n13550), .ZN(n11336) );
  XNOR2_X1 U10372 ( .A(n13729), .B(n11336), .ZN(n13734) );
  NAND2_X1 U10373 ( .A1(n13725), .A2(n13734), .ZN(n8016) );
  NAND2_X1 U10374 ( .A1(n13729), .A2(n13550), .ZN(n8015) );
  NAND2_X1 U10375 ( .A1(n8016), .A2(n8015), .ZN(n11339) );
  INV_X1 U10376 ( .A(SI_26_), .ZN(n10983) );
  NAND2_X1 U10377 ( .A1(n8020), .A2(n10983), .ZN(n8019) );
  INV_X1 U10378 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U10379 ( .A1(n8019), .A2(n8018), .ZN(n8023) );
  INV_X1 U10380 ( .A(n8020), .ZN(n8021) );
  NAND2_X1 U10381 ( .A1(n8021), .A2(SI_26_), .ZN(n8022) );
  INV_X1 U10382 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15299) );
  INV_X1 U10383 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13172) );
  MUX2_X1 U10384 ( .A(n15299), .B(n13172), .S(n8042), .Z(n8038) );
  XNOR2_X1 U10385 ( .A(n8038), .B(SI_27_), .ZN(n8036) );
  INV_X1 U10386 ( .A(n8036), .ZN(n8024) );
  NAND2_X1 U10387 ( .A1(n13169), .A2(n13472), .ZN(n8026) );
  NAND2_X1 U10388 ( .A1(n13474), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8025) );
  NAND2_X1 U10389 ( .A1(n7991), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8034) );
  NAND2_X1 U10390 ( .A1(n13439), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8033) );
  INV_X1 U10391 ( .A(n8029), .ZN(n8027) );
  NAND2_X1 U10392 ( .A1(n8027), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8108) );
  INV_X1 U10393 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10394 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  NAND2_X1 U10395 ( .A1(n8108), .A2(n8030), .ZN(n13185) );
  OR2_X1 U10396 ( .A1(n6562), .A2(n13185), .ZN(n8032) );
  INV_X1 U10397 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15140) );
  OR2_X1 U10398 ( .A1(n13442), .A2(n15140), .ZN(n8031) );
  NAND4_X1 U10399 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n13549) );
  INV_X1 U10400 ( .A(n13549), .ZN(n13281) );
  XNOR2_X1 U10401 ( .A(n13915), .B(n13281), .ZN(n13518) );
  INV_X1 U10402 ( .A(n13518), .ZN(n11338) );
  OR2_X1 U10403 ( .A1(n13915), .A2(n13549), .ZN(n8035) );
  NAND2_X1 U10404 ( .A1(n8037), .A2(n8036), .ZN(n8041) );
  INV_X1 U10405 ( .A(n8038), .ZN(n8039) );
  NAND2_X1 U10406 ( .A1(n8039), .A2(SI_27_), .ZN(n8040) );
  INV_X1 U10407 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11325) );
  INV_X1 U10408 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13168) );
  MUX2_X1 U10409 ( .A(n11325), .B(n13168), .S(n8042), .Z(n8043) );
  INV_X1 U10410 ( .A(SI_28_), .ZN(n11327) );
  NAND2_X1 U10411 ( .A1(n8043), .A2(n11327), .ZN(n11330) );
  INV_X1 U10412 ( .A(n8043), .ZN(n8044) );
  NAND2_X1 U10413 ( .A1(n8044), .A2(SI_28_), .ZN(n8045) );
  NAND2_X1 U10414 ( .A1(n11330), .A2(n8045), .ZN(n11331) );
  NAND2_X1 U10415 ( .A1(n13165), .A2(n13472), .ZN(n8047) );
  NAND2_X1 U10416 ( .A1(n13474), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10417 ( .A1(n13439), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8053) );
  INV_X1 U10418 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13717) );
  OR2_X1 U10419 ( .A1(n13438), .A2(n13717), .ZN(n8052) );
  INV_X1 U10420 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8048) );
  XNOR2_X1 U10421 ( .A(n8108), .B(n8048), .ZN(n13716) );
  OR2_X1 U10422 ( .A1(n6562), .A2(n13716), .ZN(n8051) );
  INV_X1 U10423 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8049) );
  OR2_X1 U10424 ( .A1(n13442), .A2(n8049), .ZN(n8050) );
  NAND2_X1 U10425 ( .A1(n13721), .A2(n13430), .ZN(n13697) );
  OR2_X1 U10426 ( .A1(n13721), .A2(n13430), .ZN(n8054) );
  NAND2_X1 U10427 ( .A1(n13697), .A2(n8054), .ZN(n13519) );
  AND2_X1 U10428 ( .A1(n8055), .A2(n8103), .ZN(n8056) );
  NAND2_X1 U10429 ( .A1(n13297), .A2(n14523), .ZN(n8067) );
  NAND2_X1 U10430 ( .A1(n8066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10431 ( .A1(n8063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8064) );
  MUX2_X1 U10432 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8064), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8065) );
  INV_X1 U10433 ( .A(n13307), .ZN(n10126) );
  AND2_X1 U10434 ( .A1(n10126), .A2(n13297), .ZN(n8068) );
  NOR2_X1 U10435 ( .A1(n11476), .A2(n8068), .ZN(n10081) );
  NAND2_X1 U10436 ( .A1(n10081), .A2(n14523), .ZN(n11340) );
  NAND2_X1 U10437 ( .A1(n13477), .A2(n13525), .ZN(n8069) );
  OR2_X1 U10438 ( .A1(n8069), .A2(n13297), .ZN(n14553) );
  INV_X1 U10439 ( .A(n13300), .ZN(n8070) );
  OAI21_X1 U10440 ( .B1(n13310), .B2(n13301), .A(n8070), .ZN(n10473) );
  NAND2_X1 U10441 ( .A1(n10473), .A2(n10484), .ZN(n8071) );
  NAND2_X1 U10442 ( .A1(n8071), .A2(n13314), .ZN(n14503) );
  INV_X1 U10443 ( .A(n14502), .ZN(n13317) );
  NAND2_X1 U10444 ( .A1(n14503), .A2(n13317), .ZN(n8072) );
  NOR2_X1 U10445 ( .A1(n13571), .A2(n14565), .ZN(n8073) );
  NAND2_X1 U10446 ( .A1(n13571), .A2(n14565), .ZN(n8074) );
  INV_X1 U10447 ( .A(n13570), .ZN(n8075) );
  NOR2_X1 U10448 ( .A1(n14571), .A2(n8075), .ZN(n8076) );
  NAND2_X1 U10449 ( .A1(n10227), .A2(n13498), .ZN(n8078) );
  INV_X1 U10450 ( .A(n13569), .ZN(n10195) );
  NAND2_X1 U10451 ( .A1(n13330), .A2(n10195), .ZN(n8077) );
  NAND2_X1 U10452 ( .A1(n8078), .A2(n8077), .ZN(n10166) );
  INV_X1 U10453 ( .A(n13568), .ZN(n10204) );
  NAND2_X1 U10454 ( .A1(n13333), .A2(n10204), .ZN(n8079) );
  OR2_X1 U10455 ( .A1(n14578), .A2(n8080), .ZN(n8081) );
  INV_X1 U10456 ( .A(n13503), .ZN(n10647) );
  NAND2_X1 U10457 ( .A1(n10648), .A2(n10647), .ZN(n10646) );
  NAND2_X1 U10458 ( .A1(n13345), .A2(n10962), .ZN(n8082) );
  NAND2_X1 U10459 ( .A1(n10646), .A2(n8082), .ZN(n10731) );
  OR2_X1 U10460 ( .A1(n13352), .A2(n10953), .ZN(n8083) );
  INV_X1 U10461 ( .A(n13564), .ZN(n8084) );
  OR2_X1 U10462 ( .A1(n13355), .A2(n8084), .ZN(n8085) );
  NAND2_X1 U10463 ( .A1(n10801), .A2(n8085), .ZN(n10860) );
  NAND2_X1 U10464 ( .A1(n10860), .A2(n13506), .ZN(n10859) );
  INV_X1 U10465 ( .A(n13563), .ZN(n11137) );
  OR2_X1 U10466 ( .A1(n13363), .A2(n11137), .ZN(n8086) );
  INV_X1 U10467 ( .A(n13562), .ZN(n11458) );
  OR2_X1 U10468 ( .A1(n13366), .A2(n11458), .ZN(n11190) );
  NAND2_X1 U10469 ( .A1(n11193), .A2(n13372), .ZN(n11102) );
  NAND2_X1 U10470 ( .A1(n11102), .A2(n11101), .ZN(n14382) );
  NAND2_X1 U10471 ( .A1(n14382), .A2(n13378), .ZN(n11177) );
  INV_X1 U10472 ( .A(n11177), .ZN(n8087) );
  XNOR2_X1 U10473 ( .A(n13988), .B(n13559), .ZN(n13511) );
  INV_X1 U10474 ( .A(n13559), .ZN(n8088) );
  NAND2_X1 U10475 ( .A1(n13988), .A2(n8088), .ZN(n8089) );
  INV_X1 U10476 ( .A(n13865), .ZN(n13273) );
  OR2_X1 U10477 ( .A1(n13979), .A2(n13273), .ZN(n13387) );
  NAND2_X1 U10478 ( .A1(n13979), .A2(n13273), .ZN(n13388) );
  NAND2_X1 U10479 ( .A1(n13387), .A2(n13388), .ZN(n13891) );
  XNOR2_X1 U10480 ( .A(n13873), .B(n13558), .ZN(n13862) );
  INV_X1 U10481 ( .A(n13558), .ZN(n8091) );
  OR2_X1 U10482 ( .A1(n13873), .A2(n8091), .ZN(n8092) );
  NAND2_X1 U10483 ( .A1(n13860), .A2(n8092), .ZN(n13841) );
  INV_X1 U10484 ( .A(n13841), .ZN(n8093) );
  INV_X1 U10485 ( .A(n13400), .ZN(n13556) );
  NAND2_X1 U10486 ( .A1(n13831), .A2(n13556), .ZN(n13807) );
  NAND2_X1 U10487 ( .A1(n8094), .A2(n13821), .ZN(n13810) );
  OR2_X1 U10488 ( .A1(n13950), .A2(n8095), .ZN(n8096) );
  XNOR2_X1 U10489 ( .A(n13939), .B(n13553), .ZN(n13778) );
  INV_X1 U10490 ( .A(n13553), .ZN(n8098) );
  NAND2_X1 U10491 ( .A1(n13761), .A2(n13760), .ZN(n13759) );
  NAND2_X1 U10492 ( .A1(n8120), .A2(n13552), .ZN(n8099) );
  INV_X1 U10493 ( .A(n13551), .ZN(n13282) );
  NAND2_X1 U10494 ( .A1(n14007), .A2(n13282), .ZN(n8100) );
  OR2_X1 U10495 ( .A1(n13729), .A2(n11336), .ZN(n8101) );
  INV_X1 U10496 ( .A(n13915), .ZN(n11345) );
  OAI22_X1 U10497 ( .A1(n11335), .A2(n13518), .B1(n11345), .B2(n13549), .ZN(
        n8104) );
  NAND2_X1 U10498 ( .A1(n8104), .A2(n8103), .ZN(n13698) );
  OR2_X1 U10499 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  NAND2_X1 U10500 ( .A1(n13698), .A2(n8105), .ZN(n8118) );
  NAND2_X1 U10501 ( .A1(n13297), .A2(n13525), .ZN(n8107) );
  NAND2_X1 U10502 ( .A1(n13450), .A2(n13483), .ZN(n8106) );
  NAND2_X1 U10503 ( .A1(n13439), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10504 ( .A1(n7991), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8113) );
  INV_X1 U10505 ( .A(n8108), .ZN(n8109) );
  NAND2_X1 U10506 ( .A1(n8109), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13706) );
  OR2_X1 U10507 ( .A1(n6562), .A2(n13706), .ZN(n8112) );
  INV_X1 U10508 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15143) );
  OR2_X1 U10509 ( .A1(n13442), .A2(n15143), .ZN(n8111) );
  NAND4_X1 U10510 ( .A1(n8114), .A2(n8113), .A3(n8112), .A4(n8111), .ZN(n13548) );
  NAND2_X1 U10511 ( .A1(n13297), .A2(n13450), .ZN(n13480) );
  INV_X1 U10512 ( .A(n8115), .ZN(n13589) );
  OR2_X1 U10513 ( .A1(n13480), .A2(n13589), .ZN(n13686) );
  NAND2_X1 U10514 ( .A1(n13548), .A2(n13262), .ZN(n8117) );
  OR2_X1 U10515 ( .A1(n13480), .A2(n8115), .ZN(n13542) );
  NAND2_X1 U10516 ( .A1(n13549), .A2(n13864), .ZN(n8116) );
  NAND2_X1 U10517 ( .A1(n8117), .A2(n8116), .ZN(n11570) );
  NAND2_X1 U10518 ( .A1(n14543), .A2(n14526), .ZN(n10476) );
  INV_X1 U10519 ( .A(n13333), .ZN(n10215) );
  NAND2_X1 U10520 ( .A1(n10225), .A2(n10215), .ZN(n10163) );
  NOR2_X2 U10521 ( .A1(n6608), .A2(n13345), .ZN(n10727) );
  INV_X1 U10522 ( .A(n13355), .ZN(n10909) );
  NAND2_X1 U10523 ( .A1(n13296), .A2(n11188), .ZN(n11179) );
  NAND2_X1 U10524 ( .A1(n13849), .A2(n13831), .ZN(n13830) );
  NOR2_X2 U10525 ( .A1(n6607), .A2(n13946), .ZN(n13780) );
  INV_X1 U10526 ( .A(n13781), .ZN(n8121) );
  NAND2_X1 U10527 ( .A1(n8121), .A2(n8120), .ZN(n13769) );
  NOR2_X2 U10528 ( .A1(n13769), .A2(n14007), .ZN(n13726) );
  NAND2_X1 U10529 ( .A1(n14004), .A2(n13726), .ZN(n13727) );
  OAI211_X1 U10530 ( .C1(n13429), .C2(n11342), .A(n14513), .B(n13701), .ZN(
        n13718) );
  OAI211_X1 U10531 ( .C1(n13724), .C2(n13991), .A(n13715), .B(n13718), .ZN(
        n8156) );
  OAI21_X1 U10532 ( .B1(n7546), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8123) );
  MUX2_X1 U10533 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8123), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8125) );
  NAND2_X1 U10534 ( .A1(n8127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8126) );
  MUX2_X1 U10535 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8126), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8128) );
  NAND2_X1 U10536 ( .A1(n14048), .A2(P1_B_REG_SCAN_IN), .ZN(n8131) );
  INV_X1 U10537 ( .A(n14044), .ZN(n8143) );
  INV_X1 U10538 ( .A(P1_B_REG_SCAN_IN), .ZN(n13684) );
  NAND2_X1 U10539 ( .A1(n9482), .A2(n13684), .ZN(n8130) );
  OAI211_X1 U10540 ( .C1(n9482), .C2(n8131), .A(n8143), .B(n8130), .ZN(n9481)
         );
  INV_X1 U10541 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9487) );
  NOR4_X1 U10542 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8140) );
  NOR4_X1 U10543 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n8139) );
  INV_X1 U10544 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15363) );
  INV_X1 U10545 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15360) );
  INV_X1 U10546 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15259) );
  INV_X1 U10547 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15300) );
  NAND4_X1 U10548 ( .A1(n15363), .A2(n15360), .A3(n15259), .A4(n15300), .ZN(
        n8137) );
  NOR4_X1 U10549 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8135) );
  NOR4_X1 U10550 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8134) );
  NOR4_X1 U10551 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8133) );
  NOR4_X1 U10552 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8132) );
  NAND4_X1 U10553 ( .A1(n8135), .A2(n8134), .A3(n8133), .A4(n8132), .ZN(n8136)
         );
  NOR4_X1 U10554 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8137), .A4(n8136), .ZN(n8138) );
  NAND3_X1 U10555 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n8141) );
  NAND2_X1 U10556 ( .A1(n8145), .A2(n8141), .ZN(n10076) );
  NAND2_X1 U10557 ( .A1(n14513), .A2(n13525), .ZN(n9689) );
  NAND2_X1 U10558 ( .A1(n10076), .A2(n9689), .ZN(n8142) );
  INV_X1 U10559 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9484) );
  NOR2_X1 U10560 ( .A1(n9482), .A2(n8143), .ZN(n8144) );
  NAND2_X1 U10561 ( .A1(n7546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8147) );
  AND2_X1 U10562 ( .A1(n13477), .A2(n14523), .ZN(n8148) );
  OR2_X1 U10563 ( .A1(n13480), .A2(n8148), .ZN(n9868) );
  OR2_X1 U10564 ( .A1(n10079), .A2(n13543), .ZN(n8149) );
  INV_X2 U10565 ( .A(n14577), .ZN(n8150) );
  OR2_X1 U10566 ( .A1(n9985), .A2(n14523), .ZN(n8151) );
  NAND2_X1 U10567 ( .A1(n10079), .A2(n10077), .ZN(n8154) );
  NAND2_X1 U10568 ( .A1(n8156), .A2(n14597), .ZN(n8160) );
  NAND2_X1 U10569 ( .A1(n14600), .A2(n14549), .ZN(n13976) );
  NAND2_X1 U10570 ( .A1(n14598), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8157) );
  INV_X1 U10571 ( .A(n8158), .ZN(n8159) );
  NAND2_X1 U10572 ( .A1(n8160), .A2(n8159), .ZN(P1_U3556) );
  NOR2_X1 U10573 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n8167) );
  NOR2_X1 U10574 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8166) );
  NAND4_X1 U10575 ( .A1(n8167), .A2(n8166), .A3(n8165), .A4(n8500), .ZN(n8688)
         );
  NAND4_X1 U10576 ( .A1(n15181), .A2(n8710), .A3(n8739), .A4(n6581), .ZN(n8168) );
  NOR2_X1 U10577 ( .A1(n8688), .A2(n8168), .ZN(n8169) );
  NAND2_X1 U10578 ( .A1(n8222), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U10579 ( .A1(n8651), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10580 ( .A1(n10658), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10581 ( .A1(n8299), .A2(n10559), .ZN(n8317) );
  OR2_X1 U10582 ( .A1(n8177), .A2(n11368), .ZN(n8178) );
  NAND2_X1 U10583 ( .A1(n8510), .A2(n8178), .ZN(n12227) );
  NAND2_X1 U10584 ( .A1(n8671), .A2(n12227), .ZN(n8181) );
  INV_X1 U10585 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12387) );
  OR2_X1 U10586 ( .A1(n10661), .A2(n12387), .ZN(n8180) );
  NAND4_X1 U10587 ( .A1(n8183), .A2(n8182), .A3(n8181), .A4(n8180), .ZN(n11976) );
  XNOR2_X1 U10588 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8236) );
  INV_X1 U10589 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U10590 ( .A1(n8236), .A2(n8241), .ZN(n8185) );
  NAND2_X1 U10591 ( .A1(n9526), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10592 ( .A1(n8185), .A2(n8184), .ZN(n8258) );
  NAND2_X1 U10593 ( .A1(n9502), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U10594 ( .A1(n8258), .A2(n8186), .ZN(n8188) );
  NAND2_X1 U10595 ( .A1(n9470), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10596 ( .A1(n9476), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8190) );
  INV_X1 U10597 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U10598 ( .A1(n8191), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10599 ( .A1(n8193), .A2(n8192), .ZN(n8306) );
  NAND2_X1 U10600 ( .A1(n8306), .A2(n8305), .ZN(n8196) );
  NAND2_X1 U10601 ( .A1(n8194), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10602 ( .A1(n8196), .A2(n8195), .ZN(n8325) );
  NAND2_X1 U10603 ( .A1(n9496), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10604 ( .A1(n9499), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10605 ( .A1(n8198), .A2(n8197), .ZN(n8324) );
  OR2_X2 U10606 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  XNOR2_X1 U10607 ( .A(n6963), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10608 ( .A1(n9533), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U10609 ( .A1(n9561), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10610 ( .A1(n9558), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10611 ( .A1(n9655), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10612 ( .A1(n8395), .A2(n8202), .ZN(n8204) );
  NAND2_X1 U10613 ( .A1(n9658), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10614 ( .A1(n9788), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10615 ( .A1(n9790), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10616 ( .A1(n9930), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8210) );
  INV_X1 U10617 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9928) );
  NAND2_X1 U10618 ( .A1(n9928), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U10619 ( .A1(n10045), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10620 ( .A1(n10047), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U10621 ( .A1(n8467), .A2(n8465), .ZN(n8213) );
  NAND2_X1 U10622 ( .A1(n10154), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U10623 ( .A1(n10185), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8214) );
  AOI22_X1 U10624 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(
        P1_DATAO_REG_17__SCAN_IN), .B1(n10412), .B2(n15334), .ZN(n8217) );
  XNOR2_X1 U10625 ( .A(n8495), .B(n8217), .ZN(n9865) );
  NAND2_X1 U10626 ( .A1(n9865), .A2(n8307), .ZN(n8230) );
  OR2_X1 U10627 ( .A1(n7533), .A2(n8716), .ZN(n8483) );
  NAND2_X1 U10628 ( .A1(n8483), .A2(n8499), .ZN(n8226) );
  NAND2_X1 U10629 ( .A1(n8226), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8227) );
  XNOR2_X1 U10630 ( .A(n8500), .B(n8227), .ZN(n14229) );
  OAI22_X1 U10631 ( .A1(n11764), .A2(n9866), .B1(n8698), .B2(n14229), .ZN(
        n8228) );
  INV_X1 U10632 ( .A(n8228), .ZN(n8229) );
  NAND2_X1 U10633 ( .A1(n8650), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U10634 ( .A1(n8298), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U10635 ( .A1(n8264), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8231) );
  NAND3_X1 U10636 ( .A1(n8233), .A2(n8232), .A3(n8231), .ZN(n8235) );
  INV_X1 U10637 ( .A(n8270), .ZN(n8234) );
  NOR2_X2 U10638 ( .A1(n8235), .A2(n7548), .ZN(n8254) );
  INV_X1 U10639 ( .A(SI_1_), .ZN(n9452) );
  XNOR2_X1 U10640 ( .A(n8236), .B(n8241), .ZN(n9450) );
  NAND2_X1 U10641 ( .A1(n8237), .A2(n9450), .ZN(n8240) );
  NAND2_X1 U10642 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8238) );
  XNOR2_X1 U10643 ( .A(n7083), .B(n8238), .ZN(n10255) );
  OR2_X1 U10644 ( .A1(n8245), .A2(n10255), .ZN(n8239) );
  INV_X1 U10645 ( .A(n8241), .ZN(n8244) );
  NAND2_X1 U10646 ( .A1(n8242), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10647 ( .A1(n8244), .A2(n8243), .ZN(n9462) );
  NAND2_X1 U10648 ( .A1(n8237), .A2(n9462), .ZN(n8247) );
  INV_X1 U10649 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15154) );
  OR2_X1 U10650 ( .A1(n8698), .A2(n15154), .ZN(n8246) );
  NAND2_X1 U10651 ( .A1(n8264), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8253) );
  INV_X1 U10652 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8248) );
  OR2_X1 U10653 ( .A1(n8270), .A2(n8248), .ZN(n8252) );
  NAND2_X1 U10654 ( .A1(n8298), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10655 ( .A1(n8650), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8249) );
  AND2_X1 U10656 ( .A1(n8250), .A2(n8249), .ZN(n8251) );
  NAND2_X1 U10657 ( .A1(n10388), .A2(n12336), .ZN(n8256) );
  NAND2_X1 U10658 ( .A1(n8254), .A2(n9317), .ZN(n8255) );
  NAND2_X1 U10659 ( .A1(n8256), .A2(n8255), .ZN(n12327) );
  XNOR2_X1 U10660 ( .A(n9470), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n8257) );
  XNOR2_X1 U10661 ( .A(n8258), .B(n8257), .ZN(n9468) );
  NAND2_X1 U10662 ( .A1(n8237), .A2(n9468), .ZN(n8262) );
  INV_X1 U10663 ( .A(n8290), .ZN(n8259) );
  NAND3_X1 U10664 ( .A1(n8262), .A2(n8261), .A3(n8260), .ZN(n10219) );
  INV_X1 U10665 ( .A(n10219), .ZN(n12333) );
  INV_X1 U10666 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8263) );
  OR2_X1 U10667 ( .A1(n8270), .A2(n8263), .ZN(n8268) );
  NAND2_X1 U10668 ( .A1(n8650), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U10669 ( .A1(n8298), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10670 ( .A1(n8264), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10671 ( .A1(n14979), .A2(n10219), .ZN(n11812) );
  NAND2_X2 U10672 ( .A1(n8751), .A2(n11812), .ZN(n8749) );
  AOI21_X2 U10673 ( .B1(n12327), .B2(n8749), .A(n7557), .ZN(n14984) );
  INV_X1 U10674 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8269) );
  OR2_X1 U10675 ( .A1(n8270), .A2(n8269), .ZN(n8274) );
  NAND2_X1 U10676 ( .A1(n8298), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8273) );
  INV_X1 U10677 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n14990) );
  NAND2_X1 U10678 ( .A1(n8650), .A2(n14990), .ZN(n8272) );
  NAND2_X1 U10679 ( .A1(n8264), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U10680 ( .A(n9471), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n8275) );
  XNOR2_X1 U10681 ( .A(n8276), .B(n8275), .ZN(n9466) );
  NAND2_X1 U10682 ( .A1(n8237), .A2(n9466), .ZN(n8281) );
  OR2_X1 U10683 ( .A1(n8277), .A2(SI_3_), .ZN(n8280) );
  NAND2_X1 U10684 ( .A1(n8290), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8278) );
  XNOR2_X1 U10685 ( .A(n8278), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10374) );
  OR2_X1 U10686 ( .A1(n8698), .A2(n10374), .ZN(n8279) );
  INV_X1 U10687 ( .A(n9315), .ZN(n14989) );
  NAND2_X1 U10688 ( .A1(n12329), .A2(n14989), .ZN(n11818) );
  NAND2_X1 U10689 ( .A1(n14984), .A2(n14983), .ZN(n14981) );
  NAND2_X1 U10690 ( .A1(n12329), .A2(n9315), .ZN(n8282) );
  NAND2_X1 U10691 ( .A1(n14981), .A2(n8282), .ZN(n10574) );
  NAND2_X1 U10692 ( .A1(n10658), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10693 ( .A1(n8651), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8286) );
  OR2_X1 U10694 ( .A1(n7549), .A2(n8299), .ZN(n10590) );
  NAND2_X1 U10695 ( .A1(n8671), .A2(n10590), .ZN(n8285) );
  INV_X1 U10696 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8283) );
  OR2_X1 U10697 ( .A1(n10661), .A2(n8283), .ZN(n8284) );
  INV_X1 U10698 ( .A(n14978), .ZN(n9331) );
  XNOR2_X1 U10699 ( .A(n8289), .B(n8288), .ZN(n9455) );
  NAND2_X1 U10700 ( .A1(n8307), .A2(n9455), .ZN(n8296) );
  OR2_X1 U10701 ( .A1(n8277), .A2(SI_4_), .ZN(n8295) );
  NOR2_X1 U10702 ( .A1(n8290), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8329) );
  OR2_X1 U10703 ( .A1(n8329), .A2(n8716), .ZN(n8292) );
  INV_X1 U10704 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10705 ( .A1(n8292), .A2(n8291), .ZN(n8308) );
  OR2_X1 U10706 ( .A1(n8292), .A2(n8291), .ZN(n8293) );
  OR2_X1 U10707 ( .A1(n8698), .A2(n10297), .ZN(n8294) );
  NAND2_X1 U10708 ( .A1(n9331), .A2(n9330), .ZN(n11823) );
  INV_X1 U10709 ( .A(n9330), .ZN(n10589) );
  NAND2_X1 U10710 ( .A1(n14978), .A2(n10589), .ZN(n11822) );
  NAND2_X1 U10711 ( .A1(n11823), .A2(n11822), .ZN(n11779) );
  NAND2_X1 U10712 ( .A1(n10574), .A2(n11779), .ZN(n10573) );
  NAND2_X1 U10713 ( .A1(n14978), .A2(n9330), .ZN(n8297) );
  NAND2_X1 U10714 ( .A1(n10573), .A2(n8297), .ZN(n10620) );
  INV_X1 U10715 ( .A(n10620), .ZN(n8314) );
  NAND2_X1 U10716 ( .A1(n8651), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U10717 ( .A1(n8298), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8303) );
  OR2_X1 U10718 ( .A1(n8299), .A2(n10559), .ZN(n8300) );
  NAND2_X1 U10719 ( .A1(n8317), .A2(n8300), .ZN(n11680) );
  OR2_X1 U10720 ( .A1(n10661), .A2(n15032), .ZN(n8301) );
  INV_X1 U10721 ( .A(n14965), .ZN(n9334) );
  XNOR2_X1 U10722 ( .A(n8306), .B(n8305), .ZN(n9454) );
  NAND2_X1 U10723 ( .A1(n8307), .A2(n9454), .ZN(n8312) );
  OR2_X1 U10724 ( .A1(n8277), .A2(SI_5_), .ZN(n8311) );
  NAND2_X1 U10725 ( .A1(n8308), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U10726 ( .A(n8309), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10308) );
  OR2_X1 U10727 ( .A1(n8698), .A2(n10308), .ZN(n8310) );
  NAND2_X1 U10728 ( .A1(n9334), .A2(n11679), .ZN(n11829) );
  INV_X1 U10729 ( .A(n11679), .ZN(n10626) );
  NAND2_X1 U10730 ( .A1(n14965), .A2(n10626), .ZN(n11828) );
  NAND2_X1 U10731 ( .A1(n9334), .A2(n10626), .ZN(n8315) );
  NAND2_X1 U10732 ( .A1(n8651), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10733 ( .A1(n8298), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10734 ( .A1(n8317), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10735 ( .A1(n8339), .A2(n8318), .ZN(n14961) );
  NAND2_X1 U10736 ( .A1(n8671), .A2(n14961), .ZN(n8321) );
  INV_X1 U10737 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10738 ( .A1(n10661), .A2(n8319), .ZN(n8320) );
  NAND4_X1 U10739 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n11980) );
  INV_X1 U10740 ( .A(n11980), .ZN(n9337) );
  NAND2_X1 U10741 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  NAND2_X1 U10742 ( .A1(n8327), .A2(n8326), .ZN(n9459) );
  NAND2_X1 U10743 ( .A1(n8307), .A2(n9459), .ZN(n8336) );
  INV_X1 U10744 ( .A(SI_6_), .ZN(n9460) );
  NOR2_X1 U10745 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8328) );
  NAND2_X1 U10746 ( .A1(n8329), .A2(n8328), .ZN(n8331) );
  NAND2_X1 U10747 ( .A1(n8331), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8330) );
  MUX2_X1 U10748 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8330), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8332) );
  NAND2_X1 U10749 ( .A1(n8332), .A2(n8364), .ZN(n10550) );
  OR2_X1 U10750 ( .A1(n8698), .A2(n10550), .ZN(n8333) );
  NAND2_X1 U10751 ( .A1(n9337), .A2(n14960), .ZN(n11834) );
  NAND2_X1 U10752 ( .A1(n11980), .A2(n14960), .ZN(n8338) );
  NAND2_X1 U10753 ( .A1(n10658), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U10754 ( .A1(n8651), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8344) );
  AND2_X1 U10755 ( .A1(n8339), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8340) );
  OR2_X1 U10756 ( .A1(n8340), .A2(n8355), .ZN(n11610) );
  NAND2_X1 U10757 ( .A1(n8671), .A2(n11610), .ZN(n8343) );
  INV_X1 U10758 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8341) );
  OR2_X1 U10759 ( .A1(n10661), .A2(n8341), .ZN(n8342) );
  NAND4_X1 U10760 ( .A1(n8345), .A2(n8344), .A3(n8343), .A4(n8342), .ZN(n14964) );
  INV_X1 U10761 ( .A(n14964), .ZN(n9338) );
  XNOR2_X1 U10762 ( .A(n8347), .B(n8346), .ZN(n9458) );
  NAND2_X1 U10763 ( .A1(n8307), .A2(n9458), .ZN(n8351) );
  OR2_X1 U10764 ( .A1(n8277), .A2(SI_7_), .ZN(n8350) );
  NAND2_X1 U10765 ( .A1(n8364), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8348) );
  XNOR2_X1 U10766 ( .A(n8348), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10348) );
  OR2_X1 U10767 ( .A1(n8698), .A2(n10348), .ZN(n8349) );
  NAND2_X1 U10768 ( .A1(n9338), .A2(n15042), .ZN(n11841) );
  INV_X1 U10769 ( .A(n15042), .ZN(n8352) );
  NAND2_X1 U10770 ( .A1(n14964), .A2(n8352), .ZN(n11840) );
  NAND2_X1 U10771 ( .A1(n11841), .A2(n11840), .ZN(n10779) );
  NAND2_X1 U10772 ( .A1(n10780), .A2(n10779), .ZN(n10778) );
  NAND2_X1 U10773 ( .A1(n14964), .A2(n15042), .ZN(n8353) );
  NAND2_X1 U10774 ( .A1(n8298), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10775 ( .A1(n8651), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8360) );
  NOR2_X1 U10776 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  OR2_X1 U10777 ( .A1(n8369), .A2(n8356), .ZN(n14956) );
  NAND2_X1 U10778 ( .A1(n8671), .A2(n14956), .ZN(n8359) );
  INV_X1 U10779 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8357) );
  OR2_X1 U10780 ( .A1(n10661), .A2(n8357), .ZN(n8358) );
  NAND4_X1 U10781 ( .A1(n8361), .A2(n8360), .A3(n8359), .A4(n8358), .ZN(n11979) );
  INV_X1 U10782 ( .A(SI_8_), .ZN(n9448) );
  XNOR2_X1 U10783 ( .A(n9533), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10784 ( .A(n8363), .B(n8362), .ZN(n9447) );
  NAND2_X1 U10785 ( .A1(n8307), .A2(n9447), .ZN(n8367) );
  NAND2_X1 U10786 ( .A1(n8379), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8365) );
  XNOR2_X1 U10787 ( .A(n8365), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10677) );
  OR2_X1 U10788 ( .A1(n8698), .A2(n10675), .ZN(n8366) );
  OAI211_X1 U10789 ( .C1(n8277), .C2(n9448), .A(n8367), .B(n8366), .ZN(n14955)
         );
  NAND2_X1 U10790 ( .A1(n11126), .A2(n14955), .ZN(n11845) );
  INV_X1 U10791 ( .A(n14955), .ZN(n9340) );
  NAND2_X1 U10792 ( .A1(n11979), .A2(n9340), .ZN(n11844) );
  NAND2_X1 U10793 ( .A1(n11845), .A2(n11844), .ZN(n14949) );
  NAND2_X1 U10794 ( .A1(n11126), .A2(n9340), .ZN(n8368) );
  NAND2_X1 U10795 ( .A1(n8651), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8375) );
  OR2_X1 U10796 ( .A1(n8369), .A2(n15364), .ZN(n8370) );
  NAND2_X1 U10797 ( .A1(n8387), .A2(n8370), .ZN(n11129) );
  NAND2_X1 U10798 ( .A1(n8671), .A2(n11129), .ZN(n8374) );
  NAND2_X1 U10799 ( .A1(n10658), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8373) );
  INV_X1 U10800 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8371) );
  OR2_X1 U10801 ( .A1(n10661), .A2(n8371), .ZN(n8372) );
  NAND4_X1 U10802 ( .A1(n8375), .A2(n8374), .A3(n8373), .A4(n8372), .ZN(n14951) );
  OAI21_X1 U10803 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n9473) );
  NAND2_X1 U10804 ( .A1(n8307), .A2(n9473), .ZN(n8384) );
  OR2_X1 U10805 ( .A1(n11764), .A2(SI_9_), .ZN(n8383) );
  OAI21_X1 U10806 ( .B1(n8379), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8381) );
  INV_X1 U10807 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8380) );
  XNOR2_X1 U10808 ( .A(n8381), .B(n8380), .ZN(n12020) );
  INV_X1 U10809 ( .A(n12020), .ZN(n11983) );
  OR2_X1 U10810 ( .A1(n8698), .A2(n11983), .ZN(n8382) );
  XNOR2_X1 U10811 ( .A(n14951), .B(n11850), .ZN(n11847) );
  INV_X1 U10812 ( .A(n11847), .ZN(n8385) );
  NAND2_X1 U10813 ( .A1(n14951), .A2(n11850), .ZN(n8386) );
  NAND2_X1 U10814 ( .A1(n8651), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10815 ( .A1(n10658), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10816 ( .A1(n8387), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10817 ( .A1(n8405), .A2(n8388), .ZN(n11628) );
  NAND2_X1 U10818 ( .A1(n8671), .A2(n11628), .ZN(n8391) );
  INV_X1 U10819 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8389) );
  OR2_X1 U10820 ( .A1(n10661), .A2(n8389), .ZN(n8390) );
  NAND4_X1 U10821 ( .A1(n8393), .A2(n8392), .A3(n8391), .A4(n8390), .ZN(n14275) );
  INV_X1 U10822 ( .A(n14275), .ZN(n9348) );
  XNOR2_X1 U10823 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8394) );
  XNOR2_X1 U10824 ( .A(n8395), .B(n8394), .ZN(n9480) );
  NAND2_X1 U10825 ( .A1(n9480), .A2(n8307), .ZN(n8403) );
  OR2_X1 U10826 ( .A1(n8396), .A2(n8716), .ZN(n8398) );
  MUX2_X1 U10827 ( .A(n8398), .B(P3_IR_REG_31__SCAN_IN), .S(n8397), .Z(n8400)
         );
  NAND2_X1 U10828 ( .A1(n8400), .A2(n8399), .ZN(n12018) );
  INV_X1 U10829 ( .A(n12018), .ZN(n14865) );
  OR2_X1 U10830 ( .A1(n8698), .A2(n14865), .ZN(n8402) );
  OR2_X1 U10831 ( .A1(n11764), .A2(SI_10_), .ZN(n8401) );
  NAND2_X1 U10832 ( .A1(n9348), .A2(n11627), .ZN(n11858) );
  INV_X1 U10833 ( .A(n11627), .ZN(n10976) );
  NAND2_X1 U10834 ( .A1(n14275), .A2(n10976), .ZN(n11857) );
  NAND2_X1 U10835 ( .A1(n11858), .A2(n11857), .ZN(n11854) );
  NAND2_X1 U10836 ( .A1(n14275), .A2(n11627), .ZN(n8404) );
  NAND2_X1 U10837 ( .A1(n8405), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10838 ( .A1(n8427), .A2(n8406), .ZN(n14277) );
  NAND2_X1 U10839 ( .A1(n8671), .A2(n14277), .ZN(n8411) );
  NAND2_X1 U10840 ( .A1(n8651), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10841 ( .A1(n10658), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8409) );
  INV_X1 U10842 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8407) );
  OR2_X1 U10843 ( .A1(n10661), .A2(n8407), .ZN(n8408) );
  NAND4_X1 U10844 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n14259) );
  XNOR2_X1 U10845 ( .A(n9698), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8412) );
  XNOR2_X1 U10846 ( .A(n8413), .B(n8412), .ZN(n9518) );
  NAND2_X1 U10847 ( .A1(n8399), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8414) );
  MUX2_X1 U10848 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8414), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8415) );
  AND2_X1 U10849 ( .A1(n8415), .A2(n6699), .ZN(n12016) );
  OAI22_X1 U10850 ( .A1(n11764), .A2(n15182), .B1(n8698), .B2(n14880), .ZN(
        n8416) );
  NAND2_X1 U10851 ( .A1(n11305), .A2(n14280), .ZN(n8417) );
  INV_X1 U10852 ( .A(n14280), .ZN(n8760) );
  NAND2_X1 U10853 ( .A1(n14259), .A2(n8760), .ZN(n8418) );
  OAI21_X1 U10854 ( .B1(n8421), .B2(n8420), .A(n8419), .ZN(n9527) );
  NAND2_X1 U10855 ( .A1(n9527), .A2(n8307), .ZN(n8426) );
  NAND2_X1 U10856 ( .A1(n6699), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8423) );
  XNOR2_X1 U10857 ( .A(n8423), .B(n8422), .ZN(n14899) );
  INV_X1 U10858 ( .A(n14899), .ZN(n12027) );
  OAI22_X1 U10859 ( .A1(n11764), .A2(SI_12_), .B1(n12027), .B2(n8698), .ZN(
        n8424) );
  INV_X1 U10860 ( .A(n8424), .ZN(n8425) );
  NAND2_X1 U10861 ( .A1(n8426), .A2(n8425), .ZN(n14267) );
  AND2_X1 U10862 ( .A1(n8427), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8428) );
  NOR2_X1 U10863 ( .A1(n8442), .A2(n8428), .ZN(n14262) );
  INV_X1 U10864 ( .A(n14262), .ZN(n11321) );
  NAND2_X1 U10865 ( .A1(n8671), .A2(n11321), .ZN(n8433) );
  NAND2_X1 U10866 ( .A1(n10658), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10867 ( .A1(n8651), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8431) );
  INV_X1 U10868 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8429) );
  OR2_X1 U10869 ( .A1(n10661), .A2(n8429), .ZN(n8430) );
  NAND4_X1 U10870 ( .A1(n8433), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(n14274) );
  INV_X1 U10871 ( .A(n14274), .ZN(n11307) );
  NOR2_X1 U10872 ( .A1(n14267), .A2(n11307), .ZN(n8435) );
  NAND2_X1 U10873 ( .A1(n14267), .A2(n11307), .ZN(n8434) );
  XNOR2_X1 U10874 ( .A(n8436), .B(n9831), .ZN(n14155) );
  NAND2_X1 U10875 ( .A1(n14155), .A2(n8307), .ZN(n8441) );
  OAI21_X1 U10876 ( .B1(n6699), .B2(P3_IR_REG_12__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8438) );
  XNOR2_X1 U10877 ( .A(n8438), .B(n8437), .ZN(n14916) );
  INV_X1 U10878 ( .A(n14916), .ZN(n12031) );
  OAI22_X1 U10879 ( .A1(n11764), .A2(SI_13_), .B1(n12031), .B2(n8698), .ZN(
        n8439) );
  INV_X1 U10880 ( .A(n8439), .ZN(n8440) );
  NAND2_X1 U10881 ( .A1(n8441), .A2(n8440), .ZN(n11246) );
  NAND2_X1 U10882 ( .A1(n10658), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10883 ( .A1(n8651), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8446) );
  OR2_X1 U10884 ( .A1(n8442), .A2(n11273), .ZN(n8443) );
  NAND2_X1 U10885 ( .A1(n8457), .A2(n8443), .ZN(n11272) );
  NAND2_X1 U10886 ( .A1(n8671), .A2(n11272), .ZN(n8445) );
  INV_X1 U10887 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12403) );
  OR2_X1 U10888 ( .A1(n10661), .A2(n12403), .ZN(n8444) );
  NAND4_X1 U10889 ( .A1(n8447), .A2(n8446), .A3(n8445), .A4(n8444), .ZN(n14258) );
  OR2_X1 U10890 ( .A1(n11246), .A2(n14258), .ZN(n11873) );
  NAND2_X1 U10891 ( .A1(n11246), .A2(n14258), .ZN(n11872) );
  NAND2_X1 U10892 ( .A1(n11873), .A2(n11872), .ZN(n11787) );
  INV_X1 U10893 ( .A(n14258), .ZN(n11379) );
  AND2_X1 U10894 ( .A1(n11246), .A2(n11379), .ZN(n8448) );
  AOI21_X2 U10895 ( .B1(n11244), .B2(n11787), .A(n8448), .ZN(n11234) );
  INV_X1 U10896 ( .A(n8449), .ZN(n8450) );
  XNOR2_X1 U10897 ( .A(n8451), .B(n8450), .ZN(n9783) );
  NAND2_X1 U10898 ( .A1(n9783), .A2(n8307), .ZN(n8456) );
  NAND2_X1 U10899 ( .A1(n8452), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8453) );
  XNOR2_X1 U10900 ( .A(n8453), .B(n7531), .ZN(n14938) );
  OAI22_X1 U10901 ( .A1(n11764), .A2(n9784), .B1(n8698), .B2(n14938), .ZN(
        n8454) );
  INV_X1 U10902 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U10903 ( .A1(n10658), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10904 ( .A1(n8651), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10905 ( .A1(n8457), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10906 ( .A1(n8473), .A2(n8458), .ZN(n11376) );
  NAND2_X1 U10907 ( .A1(n8671), .A2(n11376), .ZN(n8460) );
  INV_X1 U10908 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12398) );
  OR2_X1 U10909 ( .A1(n10661), .A2(n12398), .ZN(n8459) );
  NAND4_X1 U10910 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(n11978) );
  OR2_X1 U10911 ( .A1(n12316), .A2(n11978), .ZN(n8463) );
  NAND2_X1 U10912 ( .A1(n12316), .A2(n11978), .ZN(n8464) );
  INV_X1 U10913 ( .A(n8465), .ZN(n8466) );
  XNOR2_X1 U10914 ( .A(n8467), .B(n8466), .ZN(n9823) );
  NAND2_X1 U10915 ( .A1(n9823), .A2(n8307), .ZN(n8472) );
  OR2_X1 U10916 ( .A1(n8468), .A2(n8716), .ZN(n8469) );
  XNOR2_X1 U10917 ( .A(n8469), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14185) );
  INV_X1 U10918 ( .A(n14185), .ZN(n12039) );
  OAI22_X1 U10919 ( .A1(n11764), .A2(n9824), .B1(n8698), .B2(n12039), .ZN(
        n8470) );
  INV_X1 U10920 ( .A(n8470), .ZN(n8471) );
  NAND2_X1 U10921 ( .A1(n10658), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10922 ( .A1(n8651), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8477) );
  AND2_X1 U10923 ( .A1(n8473), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8474) );
  OR2_X1 U10924 ( .A1(n8474), .A2(n8488), .ZN(n12255) );
  NAND2_X1 U10925 ( .A1(n8671), .A2(n12255), .ZN(n8476) );
  INV_X1 U10926 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12395) );
  OR2_X1 U10927 ( .A1(n10661), .A2(n12395), .ZN(n8475) );
  NAND4_X1 U10928 ( .A1(n8478), .A2(n8477), .A3(n8476), .A4(n8475), .ZN(n11977) );
  OR2_X1 U10929 ( .A1(n12313), .A2(n11977), .ZN(n8479) );
  INV_X1 U10930 ( .A(n12234), .ZN(n8493) );
  INV_X1 U10931 ( .A(n8480), .ZN(n8481) );
  XNOR2_X1 U10932 ( .A(n8482), .B(n8481), .ZN(n14163) );
  NAND2_X1 U10933 ( .A1(n14163), .A2(n8307), .ZN(n8487) );
  XNOR2_X1 U10934 ( .A(n8483), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12045) );
  INV_X1 U10935 ( .A(n12045), .ZN(n14211) );
  OAI22_X1 U10936 ( .A1(n11764), .A2(n8484), .B1(n8698), .B2(n14211), .ZN(
        n8485) );
  INV_X1 U10937 ( .A(n8485), .ZN(n8486) );
  NAND2_X1 U10938 ( .A1(n8298), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U10939 ( .A1(n8651), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8491) );
  XNOR2_X1 U10940 ( .A(n8488), .B(n11669), .ZN(n12241) );
  NAND2_X1 U10941 ( .A1(n8671), .A2(n12241), .ZN(n8490) );
  INV_X1 U10942 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12391) );
  OR2_X1 U10943 ( .A1(n10661), .A2(n12391), .ZN(n8489) );
  NAND4_X1 U10944 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n12223) );
  NAND2_X1 U10945 ( .A1(n12309), .A2(n12223), .ZN(n8765) );
  OR2_X1 U10946 ( .A1(n12303), .A2(n12240), .ZN(n11892) );
  NAND2_X1 U10947 ( .A1(n12303), .A2(n12240), .ZN(n11891) );
  NAND2_X1 U10948 ( .A1(n10412), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10949 ( .A1(n15334), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10950 ( .A1(n10713), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10951 ( .A1(n10724), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U10952 ( .A1(n8518), .A2(n8498), .ZN(n8516) );
  XNOR2_X1 U10953 ( .A(n8517), .B(n8516), .ZN(n9971) );
  NAND2_X1 U10954 ( .A1(n9971), .A2(n8307), .ZN(n8509) );
  NAND2_X1 U10955 ( .A1(n8500), .A2(n8499), .ZN(n8501) );
  INV_X1 U10956 ( .A(n8505), .ZN(n8502) );
  NAND2_X1 U10957 ( .A1(n8502), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8503) );
  MUX2_X1 U10958 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8503), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8506) );
  NAND2_X1 U10959 ( .A1(n8505), .A2(n8504), .ZN(n8522) );
  NAND2_X1 U10960 ( .A1(n8506), .A2(n8522), .ZN(n14239) );
  OAI22_X1 U10961 ( .A1(n11764), .A2(n9972), .B1(n8698), .B2(n14239), .ZN(
        n8507) );
  INV_X1 U10962 ( .A(n8507), .ZN(n8508) );
  NAND2_X1 U10963 ( .A1(n8651), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10964 ( .A1(n8510), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U10965 ( .A1(n8527), .A2(n8511), .ZN(n12211) );
  NAND2_X1 U10966 ( .A1(n8671), .A2(n12211), .ZN(n8514) );
  NAND2_X1 U10967 ( .A1(n10658), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8513) );
  INV_X1 U10968 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12383) );
  OR2_X1 U10969 ( .A1(n10661), .A2(n12383), .ZN(n8512) );
  NAND4_X1 U10970 ( .A1(n8515), .A2(n8514), .A3(n8513), .A4(n8512), .ZN(n12224) );
  NAND2_X1 U10971 ( .A1(n12300), .A2(n11711), .ZN(n11897) );
  NAND2_X1 U10972 ( .A1(n10832), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8539) );
  INV_X1 U10973 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n15176) );
  NAND2_X1 U10974 ( .A1(n15176), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8519) );
  INV_X1 U10975 ( .A(n8537), .ZN(n8520) );
  XNOR2_X1 U10976 ( .A(n8538), .B(n8520), .ZN(n10012) );
  NAND2_X1 U10977 ( .A1(n10012), .A2(n8307), .ZN(n8526) );
  NAND2_X1 U10978 ( .A1(n8522), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8521) );
  MUX2_X1 U10979 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8521), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8523) );
  OAI22_X1 U10980 ( .A1(n11764), .A2(SI_19_), .B1(n12011), .B2(n8698), .ZN(
        n8524) );
  INV_X1 U10981 ( .A(n8524), .ZN(n8525) );
  INV_X1 U10982 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12379) );
  AND2_X1 U10983 ( .A1(n8527), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8528) );
  OR2_X1 U10984 ( .A1(n8528), .A2(n8545), .ZN(n12197) );
  NAND2_X1 U10985 ( .A1(n12197), .A2(n8671), .ZN(n8532) );
  NAND2_X1 U10986 ( .A1(n8298), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U10987 ( .A1(n8651), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8529) );
  AND2_X1 U10988 ( .A1(n8530), .A2(n8529), .ZN(n8531) );
  OAI211_X1 U10989 ( .C1(n10661), .C2(n12379), .A(n8532), .B(n8531), .ZN(
        n11975) );
  NAND2_X1 U10990 ( .A1(n12196), .A2(n11975), .ZN(n11903) );
  NAND2_X1 U10991 ( .A1(n11902), .A2(n11903), .ZN(n12190) );
  INV_X1 U10992 ( .A(n12300), .ZN(n8533) );
  NAND2_X1 U10993 ( .A1(n8533), .A2(n11711), .ZN(n12191) );
  AND2_X1 U10994 ( .A1(n12190), .A2(n12191), .ZN(n8534) );
  NAND2_X1 U10995 ( .A1(n12206), .A2(n8534), .ZN(n12189) );
  INV_X1 U10996 ( .A(n11975), .ZN(n12210) );
  NAND2_X1 U10997 ( .A1(n12189), .A2(n8536), .ZN(n12177) );
  NAND2_X1 U10998 ( .A1(n15175), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10999 ( .A1(n10830), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8541) );
  XNOR2_X1 U11000 ( .A(n8551), .B(n8550), .ZN(n10180) );
  NAND2_X1 U11001 ( .A1(n10180), .A2(n8307), .ZN(n8543) );
  OR2_X1 U11002 ( .A1(n11764), .A2(n15138), .ZN(n8542) );
  NOR2_X1 U11003 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  OR2_X1 U11004 ( .A1(n8557), .A2(n8546), .ZN(n12180) );
  NAND2_X1 U11005 ( .A1(n12180), .A2(n8671), .ZN(n8549) );
  AOI22_X1 U11006 ( .A1(n8298), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n8651), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n8548) );
  INV_X1 U11007 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n15385) );
  OR2_X1 U11008 ( .A1(n10661), .A2(n15385), .ZN(n8547) );
  XNOR2_X1 U11009 ( .A(n12293), .B(n12166), .ZN(n12176) );
  INV_X1 U11010 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U11011 ( .A1(n10968), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8563) );
  INV_X1 U11012 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n15292) );
  NAND2_X1 U11013 ( .A1(n15292), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8553) );
  XNOR2_X1 U11014 ( .A(n8562), .B(n8561), .ZN(n10408) );
  NAND2_X1 U11015 ( .A1(n10408), .A2(n8307), .ZN(n8555) );
  INV_X1 U11016 ( .A(SI_21_), .ZN(n10410) );
  INV_X1 U11017 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12372) );
  INV_X1 U11018 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8556) );
  OR2_X1 U11019 ( .A1(n8557), .A2(n8556), .ZN(n8558) );
  NAND2_X1 U11020 ( .A1(n8572), .A2(n8558), .ZN(n12167) );
  NAND2_X1 U11021 ( .A1(n12167), .A2(n8671), .ZN(n8560) );
  AOI22_X1 U11022 ( .A1(n8298), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8264), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n8559) );
  NOR2_X1 U11023 ( .A1(n12289), .A2(n11974), .ZN(n11792) );
  INV_X1 U11024 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11108) );
  NAND2_X1 U11025 ( .A1(n11108), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8580) );
  INV_X1 U11026 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U11027 ( .A1(n8564), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8565) );
  AND2_X1 U11028 ( .A1(n8580), .A2(n8565), .ZN(n8566) );
  OR2_X1 U11029 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  NAND2_X1 U11030 ( .A1(n8581), .A2(n8568), .ZN(n10515) );
  NAND2_X1 U11031 ( .A1(n10515), .A2(n8307), .ZN(n8571) );
  OR2_X1 U11032 ( .A1(n11764), .A2(n8569), .ZN(n8570) );
  NAND2_X1 U11033 ( .A1(n8572), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11034 ( .A1(n8589), .A2(n8573), .ZN(n12155) );
  NAND2_X1 U11035 ( .A1(n12155), .A2(n8671), .ZN(n8578) );
  INV_X1 U11036 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U11037 ( .A1(n8298), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U11038 ( .A1(n8651), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8574) );
  OAI211_X1 U11039 ( .C1(n12368), .C2(n10661), .A(n8575), .B(n8574), .ZN(n8576) );
  INV_X1 U11040 ( .A(n8576), .ZN(n8577) );
  NAND2_X1 U11041 ( .A1(n8578), .A2(n8577), .ZN(n11972) );
  INV_X1 U11042 ( .A(n12285), .ZN(n8579) );
  NAND2_X1 U11043 ( .A1(n15285), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11044 ( .A1(n8582), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8583) );
  AND2_X1 U11045 ( .A1(n8597), .A2(n8583), .ZN(n8584) );
  OR2_X1 U11046 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  NAND2_X1 U11047 ( .A1(n8598), .A2(n8586), .ZN(n10708) );
  NAND2_X1 U11048 ( .A1(n10708), .A2(n8307), .ZN(n8588) );
  NAND2_X1 U11049 ( .A1(n8589), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U11050 ( .A1(n8602), .A2(n8590), .ZN(n12144) );
  NAND2_X1 U11051 ( .A1(n12144), .A2(n8671), .ZN(n8595) );
  INV_X1 U11052 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12364) );
  NAND2_X1 U11053 ( .A1(n8298), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11054 ( .A1(n8651), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8591) );
  OAI211_X1 U11055 ( .C1(n12364), .C2(n10661), .A(n8592), .B(n8591), .ZN(n8593) );
  INV_X1 U11056 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U11057 ( .A1(n12281), .A2(n12154), .ZN(n8596) );
  XNOR2_X1 U11058 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .ZN(n8599) );
  XNOR2_X1 U11059 ( .A(n8611), .B(n8599), .ZN(n8600) );
  MUX2_X1 U11060 ( .A(SI_24_), .B(n8600), .S(n9474), .Z(n12419) );
  INV_X1 U11061 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n11690) );
  NAND2_X1 U11062 ( .A1(n8602), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U11063 ( .A1(n8617), .A2(n8603), .ZN(n12132) );
  NAND2_X1 U11064 ( .A1(n12132), .A2(n8671), .ZN(n8609) );
  INV_X1 U11065 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8606) );
  NAND2_X1 U11066 ( .A1(n8298), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U11067 ( .A1(n8651), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8604) );
  OAI211_X1 U11068 ( .C1(n8606), .C2(n10661), .A(n8605), .B(n8604), .ZN(n8607)
         );
  INV_X1 U11069 ( .A(n8607), .ZN(n8608) );
  NAND2_X1 U11070 ( .A1(n12279), .A2(n11971), .ZN(n11925) );
  INV_X1 U11071 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11174) );
  AND2_X1 U11072 ( .A1(n11174), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8610) );
  INV_X1 U11073 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11203) );
  NAND2_X1 U11074 ( .A1(n11203), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8612) );
  INV_X1 U11075 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15366) );
  XNOR2_X1 U11076 ( .A(n15366), .B(P1_DATAO_REG_25__SCAN_IN), .ZN(n8624) );
  XNOR2_X1 U11077 ( .A(n8626), .B(n8624), .ZN(n10834) );
  NAND2_X1 U11078 ( .A1(n10834), .A2(n8307), .ZN(n8614) );
  INV_X1 U11079 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11080 ( .A1(n8617), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11081 ( .A1(n8631), .A2(n8618), .ZN(n12118) );
  NAND2_X1 U11082 ( .A1(n12118), .A2(n8671), .ZN(n8623) );
  INV_X1 U11083 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U11084 ( .A1(n8298), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U11085 ( .A1(n8651), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8619) );
  OAI211_X1 U11086 ( .C1(n12359), .C2(n10661), .A(n8620), .B(n8619), .ZN(n8621) );
  INV_X1 U11087 ( .A(n8621), .ZN(n8622) );
  NAND2_X1 U11088 ( .A1(n12273), .A2(n12125), .ZN(n11933) );
  NAND2_X1 U11089 ( .A1(n11932), .A2(n11933), .ZN(n12114) );
  INV_X1 U11090 ( .A(n8624), .ZN(n8625) );
  NAND2_X1 U11091 ( .A1(n15366), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U11092 ( .A(n14046), .B(P1_DATAO_REG_26__SCAN_IN), .ZN(n8639) );
  XNOR2_X1 U11093 ( .A(n8641), .B(n8639), .ZN(n10981) );
  NAND2_X1 U11094 ( .A1(n10981), .A2(n8307), .ZN(n8630) );
  OR2_X1 U11095 ( .A1(n11764), .A2(n10983), .ZN(n8629) );
  NAND2_X1 U11096 ( .A1(n8631), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11097 ( .A1(n8648), .A2(n8632), .ZN(n12108) );
  NAND2_X1 U11098 ( .A1(n12108), .A2(n8671), .ZN(n8638) );
  INV_X1 U11099 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U11100 ( .A1(n8298), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U11101 ( .A1(n8651), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8633) );
  OAI211_X1 U11102 ( .C1(n8635), .C2(n10661), .A(n8634), .B(n8633), .ZN(n8636)
         );
  INV_X1 U11103 ( .A(n8636), .ZN(n8637) );
  INV_X1 U11104 ( .A(n8639), .ZN(n8640) );
  NAND2_X1 U11105 ( .A1(n8641), .A2(n8640), .ZN(n8643) );
  NAND2_X1 U11106 ( .A1(n14046), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8642) );
  XNOR2_X1 U11107 ( .A(n15299), .B(P1_DATAO_REG_27__SCAN_IN), .ZN(n8657) );
  XNOR2_X1 U11108 ( .A(n8659), .B(n8657), .ZN(n11049) );
  NAND2_X1 U11109 ( .A1(n11049), .A2(n8307), .ZN(n8645) );
  INV_X1 U11110 ( .A(SI_27_), .ZN(n11051) );
  INV_X1 U11111 ( .A(n8648), .ZN(n8647) );
  INV_X1 U11112 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11113 ( .A1(n8648), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U11114 ( .A1(n8666), .A2(n8649), .ZN(n12094) );
  NAND2_X1 U11115 ( .A1(n12094), .A2(n8650), .ZN(n8656) );
  INV_X1 U11116 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U11117 ( .A1(n8651), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11118 ( .A1(n8234), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8652) );
  OAI211_X1 U11119 ( .C1(n8316), .C2(n15246), .A(n8653), .B(n8652), .ZN(n8654)
         );
  INV_X1 U11120 ( .A(n8654), .ZN(n8655) );
  NAND2_X1 U11121 ( .A1(n12266), .A2(n12102), .ZN(n11943) );
  INV_X1 U11122 ( .A(n12266), .ZN(n9425) );
  INV_X1 U11123 ( .A(n8657), .ZN(n8658) );
  NAND2_X1 U11124 ( .A1(n8659), .A2(n8658), .ZN(n8661) );
  NAND2_X1 U11125 ( .A1(n15299), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8660) );
  AOI22_X1 U11126 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13168), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11325), .ZN(n8662) );
  INV_X1 U11127 ( .A(n8662), .ZN(n8663) );
  XNOR2_X1 U11128 ( .A(n8674), .B(n8663), .ZN(n11326) );
  NAND2_X1 U11129 ( .A1(n11326), .A2(n8307), .ZN(n8665) );
  NAND2_X2 U11130 ( .A1(n8665), .A2(n8664), .ZN(n12263) );
  NAND2_X1 U11131 ( .A1(n8666), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11132 ( .A1(n12066), .A2(n8667), .ZN(n12083) );
  INV_X1 U11133 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n15276) );
  NAND2_X1 U11134 ( .A1(n8234), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11135 ( .A1(n8264), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U11136 ( .C1(n8316), .C2(n15276), .A(n8669), .B(n8668), .ZN(n8670)
         );
  AOI21_X1 U11137 ( .B1(n12083), .B2(n8671), .A(n8670), .ZN(n12093) );
  NAND2_X1 U11138 ( .A1(n12263), .A2(n12093), .ZN(n11944) );
  NAND2_X1 U11139 ( .A1(n12078), .A2(n12077), .ZN(n12076) );
  INV_X1 U11140 ( .A(n12263), .ZN(n8672) );
  NAND2_X1 U11141 ( .A1(n12076), .A2(n7552), .ZN(n8684) );
  NOR2_X1 U11142 ( .A1(n13168), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U11143 ( .A1(n13168), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8675) );
  XNOR2_X1 U11144 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11750) );
  XNOR2_X1 U11145 ( .A(n11752), .B(n11750), .ZN(n11117) );
  NAND2_X1 U11146 ( .A1(n11117), .A2(n8307), .ZN(n8677) );
  INV_X1 U11147 ( .A(SI_29_), .ZN(n11120) );
  OR2_X1 U11148 ( .A1(n11764), .A2(n11120), .ZN(n8676) );
  NAND2_X1 U11149 ( .A1(n8677), .A2(n8676), .ZN(n8707) );
  INV_X1 U11150 ( .A(n12066), .ZN(n8678) );
  NAND2_X1 U11151 ( .A1(n8678), .A2(n8671), .ZN(n10665) );
  NAND2_X1 U11152 ( .A1(n8264), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11153 ( .A1(n10658), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U11154 ( .C1(n10661), .C2(n9439), .A(n8680), .B(n8679), .ZN(n8681)
         );
  INV_X1 U11155 ( .A(n8681), .ZN(n8682) );
  NAND2_X1 U11156 ( .A1(n8707), .A2(n12082), .ZN(n11951) );
  NAND2_X1 U11157 ( .A1(n11953), .A2(n11951), .ZN(n11797) );
  XNOR2_X1 U11158 ( .A(n8684), .B(n8683), .ZN(n8692) );
  NAND2_X1 U11159 ( .A1(n8686), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11160 ( .A1(n11772), .A2(n11962), .ZN(n8691) );
  NAND2_X1 U11161 ( .A1(n8709), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U11162 ( .A1(n12011), .A2(n11966), .ZN(n9405) );
  NAND2_X1 U11163 ( .A1(n8692), .A2(n14982), .ZN(n8706) );
  INV_X1 U11164 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U11165 ( .A1(n10658), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U11166 ( .A1(n8651), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8693) );
  OAI211_X1 U11167 ( .C1(n8695), .C2(n10661), .A(n8694), .B(n8693), .ZN(n8696)
         );
  INV_X1 U11168 ( .A(n8696), .ZN(n8697) );
  AND2_X1 U11169 ( .A1(n10665), .A2(n8697), .ZN(n11766) );
  OR2_X1 U11170 ( .A1(n11329), .A2(n6590), .ZN(n10257) );
  NAND2_X1 U11171 ( .A1(n8698), .A2(n10257), .ZN(n8701) );
  INV_X1 U11172 ( .A(P3_B_REG_SCAN_IN), .ZN(n8699) );
  OR2_X1 U11173 ( .A1(n11329), .A2(n8699), .ZN(n8700) );
  NAND2_X1 U11174 ( .A1(n14977), .A2(n8700), .ZN(n12063) );
  INV_X1 U11175 ( .A(n8701), .ZN(n8702) );
  NOR2_X1 U11176 ( .A1(n12093), .A2(n12252), .ZN(n8703) );
  INV_X1 U11177 ( .A(n8707), .ZN(n8708) );
  NAND2_X1 U11178 ( .A1(n6582), .A2(n6580), .ZN(n8712) );
  XNOR2_X1 U11179 ( .A(n8721), .B(P3_B_REG_SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11180 ( .A1(n8714), .A2(n10836), .ZN(n8720) );
  NOR2_X1 U11181 ( .A1(n8222), .A2(n8716), .ZN(n8715) );
  MUX2_X1 U11182 ( .A(n8716), .B(n8715), .S(P3_IR_REG_26__SCAN_IN), .Z(n8719)
         );
  INV_X1 U11183 ( .A(n8736), .ZN(n10984) );
  NAND2_X1 U11184 ( .A1(n8721), .A2(n10984), .ZN(n8722) );
  NAND2_X1 U11185 ( .A1(n10836), .A2(n10984), .ZN(n8724) );
  XNOR2_X1 U11186 ( .A(n9308), .B(n10581), .ZN(n8742) );
  NOR4_X1 U11187 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8734) );
  INV_X1 U11188 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n15336) );
  INV_X1 U11189 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15303) );
  INV_X1 U11190 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n15178) );
  INV_X1 U11191 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15219) );
  NAND4_X1 U11192 ( .A1(n15336), .A2(n15303), .A3(n15178), .A4(n15219), .ZN(
        n8731) );
  NOR4_X1 U11193 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8729) );
  NOR4_X1 U11194 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8728) );
  NOR4_X1 U11195 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8727) );
  NOR4_X1 U11196 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8726) );
  NAND4_X1 U11197 ( .A1(n8729), .A2(n8728), .A3(n8727), .A4(n8726), .ZN(n8730)
         );
  NOR4_X1 U11198 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8731), .A4(n8730), .ZN(n8733) );
  NOR4_X1 U11199 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8732) );
  AND3_X1 U11200 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8735) );
  OR2_X1 U11201 ( .A1(n8723), .A2(n8735), .ZN(n9403) );
  INV_X1 U11202 ( .A(n8721), .ZN(n12418) );
  NAND2_X1 U11203 ( .A1(n12418), .A2(n8736), .ZN(n8737) );
  NAND2_X1 U11204 ( .A1(n8738), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8740) );
  AND2_X1 U11205 ( .A1(n9403), .A2(n10238), .ZN(n8741) );
  NAND3_X1 U11206 ( .A1(n12057), .A2(n11962), .A3(n11966), .ZN(n10578) );
  MUX2_X1 U11207 ( .A(n9311), .B(n10578), .S(n11911), .Z(n10577) );
  NAND2_X1 U11208 ( .A1(n10581), .A2(n10577), .ZN(n8746) );
  NAND2_X1 U11209 ( .A1(n11801), .A2(n10182), .ZN(n8772) );
  NAND2_X1 U11210 ( .A1(n9311), .A2(n9405), .ZN(n8743) );
  AOI21_X1 U11211 ( .B1(n11805), .B2(n8772), .A(n8743), .ZN(n8744) );
  INV_X1 U11212 ( .A(n10581), .ZN(n15073) );
  OAI21_X1 U11213 ( .B1(n11948), .B2(n8744), .A(n15073), .ZN(n8745) );
  NAND2_X1 U11214 ( .A1(n9322), .A2(n11809), .ZN(n12326) );
  INV_X1 U11215 ( .A(n8749), .ZN(n8750) );
  NAND2_X1 U11216 ( .A1(n12326), .A2(n8750), .ZN(n8752) );
  NAND2_X1 U11217 ( .A1(n8752), .A2(n8751), .ZN(n14976) );
  NAND2_X1 U11218 ( .A1(n14975), .A2(n11819), .ZN(n10572) );
  INV_X1 U11219 ( .A(n11779), .ZN(n11821) );
  NAND2_X1 U11220 ( .A1(n10572), .A2(n11821), .ZN(n8754) );
  NAND2_X1 U11221 ( .A1(n8754), .A2(n11823), .ZN(n10618) );
  NAND2_X1 U11222 ( .A1(n10618), .A2(n11825), .ZN(n8755) );
  NAND2_X1 U11223 ( .A1(n8755), .A2(n11829), .ZN(n14963) );
  INV_X1 U11224 ( .A(n10779), .ZN(n11836) );
  INV_X1 U11225 ( .A(n14949), .ZN(n11843) );
  NAND2_X1 U11226 ( .A1(n14947), .A2(n11843), .ZN(n8756) );
  NAND2_X1 U11227 ( .A1(n8756), .A2(n11845), .ZN(n10895) );
  NOR2_X1 U11228 ( .A1(n14951), .A2(n11125), .ZN(n8757) );
  NAND2_X1 U11229 ( .A1(n14951), .A2(n11125), .ZN(n8758) );
  INV_X1 U11230 ( .A(n11854), .ZN(n11784) );
  NAND2_X1 U11231 ( .A1(n11305), .A2(n8760), .ZN(n11861) );
  NAND2_X1 U11232 ( .A1(n14280), .A2(n14259), .ZN(n11864) );
  NAND2_X1 U11233 ( .A1(n11861), .A2(n11864), .ZN(n14278) );
  NAND2_X1 U11234 ( .A1(n14267), .A2(n14274), .ZN(n11865) );
  NAND2_X1 U11235 ( .A1(n14266), .A2(n14264), .ZN(n8761) );
  NAND2_X1 U11236 ( .A1(n8761), .A2(n11871), .ZN(n11243) );
  NAND2_X1 U11237 ( .A1(n11243), .A2(n11872), .ZN(n8762) );
  NAND2_X1 U11238 ( .A1(n8762), .A2(n11873), .ZN(n11240) );
  INV_X1 U11239 ( .A(n11788), .ZN(n11875) );
  NAND2_X1 U11240 ( .A1(n11240), .A2(n11875), .ZN(n8764) );
  NAND2_X1 U11241 ( .A1(n12316), .A2(n12251), .ZN(n8763) );
  NAND2_X1 U11242 ( .A1(n8764), .A2(n8763), .ZN(n12246) );
  OR2_X1 U11243 ( .A1(n12313), .A2(n12239), .ZN(n11881) );
  NAND2_X1 U11244 ( .A1(n12313), .A2(n12239), .ZN(n11886) );
  NAND2_X1 U11245 ( .A1(n12236), .A2(n8765), .ZN(n12235) );
  INV_X1 U11246 ( .A(n12223), .ZN(n12253) );
  NAND2_X1 U11247 ( .A1(n12309), .A2(n12253), .ZN(n11887) );
  NAND2_X1 U11248 ( .A1(n12217), .A2(n12218), .ZN(n8766) );
  NAND2_X1 U11249 ( .A1(n12186), .A2(n11902), .ZN(n12173) );
  OR2_X1 U11250 ( .A1(n12293), .A2(n12166), .ZN(n11907) );
  NAND2_X1 U11251 ( .A1(n12289), .A2(n12179), .ZN(n8767) );
  NOR2_X1 U11252 ( .A1(n12285), .A2(n12165), .ZN(n11916) );
  NAND2_X1 U11253 ( .A1(n12285), .A2(n12165), .ZN(n11793) );
  INV_X1 U11254 ( .A(n11933), .ZN(n8768) );
  NAND2_X1 U11255 ( .A1(n8769), .A2(n11932), .ZN(n12101) );
  NOR2_X1 U11256 ( .A1(n12268), .A2(n12117), .ZN(n11937) );
  NAND2_X1 U11257 ( .A1(n12268), .A2(n12117), .ZN(n11791) );
  INV_X1 U11258 ( .A(n11943), .ZN(n8770) );
  AOI21_X1 U11259 ( .B1(n12090), .B2(n7092), .A(n8770), .ZN(n12075) );
  INV_X1 U11260 ( .A(n11946), .ZN(n8771) );
  XNOR2_X1 U11261 ( .A(n11768), .B(n11797), .ZN(n12073) );
  XNOR2_X1 U11262 ( .A(n8772), .B(n11966), .ZN(n8774) );
  OR2_X1 U11263 ( .A1(n12011), .A2(n11772), .ZN(n8773) );
  NAND2_X1 U11264 ( .A1(n8774), .A2(n8773), .ZN(n9430) );
  AND2_X1 U11265 ( .A1(n11960), .A2(n14988), .ZN(n8775) );
  NAND2_X1 U11266 ( .A1(n9430), .A2(n8775), .ZN(n8776) );
  NAND2_X1 U11267 ( .A1(n8776), .A2(n10578), .ZN(n12131) );
  NAND2_X1 U11268 ( .A1(n8777), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11269 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8935) );
  NOR2_X1 U11270 ( .A1(n8935), .A2(n9909), .ZN(n8934) );
  NAND2_X1 U11271 ( .A1(n8934), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8970) );
  INV_X1 U11272 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10121) );
  INV_X1 U11273 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9003) );
  AND2_X1 U11274 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n8780) );
  AND2_X1 U11275 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n8781) );
  INV_X1 U11276 ( .A(n9100), .ZN(n8782) );
  NAND2_X1 U11277 ( .A1(n8782), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9116) );
  INV_X1 U11278 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9115) );
  INV_X1 U11279 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8841) );
  INV_X1 U11280 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9159) );
  INV_X1 U11281 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9158) );
  INV_X1 U11282 ( .A(n9175), .ZN(n8785) );
  NAND2_X1 U11283 ( .A1(n8785), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9192) );
  INV_X1 U11284 ( .A(n9192), .ZN(n8786) );
  INV_X1 U11285 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12474) );
  INV_X1 U11286 ( .A(n9216), .ZN(n8788) );
  AND2_X1 U11287 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8787) );
  NAND2_X1 U11288 ( .A1(n8788), .A2(n8787), .ZN(n9234) );
  INV_X1 U11289 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8790) );
  INV_X1 U11290 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8789) );
  OAI21_X1 U11291 ( .B1(n9216), .B2(n8790), .A(n8789), .ZN(n8791) );
  NAND2_X1 U11292 ( .A1(n9234), .A2(n8791), .ZN(n12897) );
  NOR2_X2 U11293 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9048) );
  NOR3_X2 U11294 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .A3(
        P2_IR_REG_12__SCAN_IN), .ZN(n8795) );
  NOR2_X1 U11295 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8800) );
  NOR2_X1 U11296 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8799) );
  NOR2_X1 U11297 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8798) );
  NOR2_X1 U11298 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8801) );
  AND4_X2 U11299 ( .A1(n8801), .A2(n9277), .A3(n9244), .A4(n9249), .ZN(n8802)
         );
  INV_X1 U11300 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8803) );
  INV_X1 U11301 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8805) );
  OR2_X1 U11302 ( .A1(n12897), .A2(n11403), .ZN(n8817) );
  INV_X1 U11303 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U11304 ( .A1(n8811), .A2(n11334), .ZN(n8872) );
  INV_X2 U11305 ( .A(n9239), .ZN(n11429) );
  NAND2_X1 U11306 ( .A1(n11429), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11307 ( .A1(n11430), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8812) );
  OAI211_X1 U11308 ( .C1(n8814), .C2(n12668), .A(n8813), .B(n8812), .ZN(n8815)
         );
  INV_X1 U11309 ( .A(n8815), .ZN(n8816) );
  INV_X1 U11310 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8820) );
  NOR2_X1 U11311 ( .A1(n6619), .A2(n8805), .ZN(n8823) );
  XNOR2_X2 U11312 ( .A(n8823), .B(n9244), .ZN(n12778) );
  NAND2_X1 U11313 ( .A1(n8824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8825) );
  NOR2_X1 U11314 ( .A1(n12912), .A2(n12913), .ZN(n9229) );
  NAND2_X1 U11315 ( .A1(n12685), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8831) );
  NAND2_X2 U11316 ( .A1(n8832), .A2(n12767), .ZN(n12765) );
  OR2_X1 U11317 ( .A1(n8834), .A2(n15197), .ZN(n8835) );
  NAND2_X2 U11318 ( .A1(n8833), .A2(n8835), .ZN(n12762) );
  NAND2_X2 U11319 ( .A1(n9731), .A2(n12765), .ZN(n8901) );
  INV_X4 U11320 ( .A(n8849), .ZN(n12433) );
  XNOR2_X1 U11321 ( .A(n12900), .B(n12433), .ZN(n9227) );
  NAND2_X1 U11322 ( .A1(n8837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8838) );
  XNOR2_X1 U11323 ( .A(n8838), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14718) );
  AOI22_X1 U11324 ( .A1(n12685), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9135), 
        .B2(n14718), .ZN(n8839) );
  XNOR2_X1 U11325 ( .A(n13045), .B(n12433), .ZN(n9133) );
  NAND2_X1 U11326 ( .A1(n8852), .A2(n8841), .ZN(n8842) );
  NAND2_X1 U11327 ( .A1(n9139), .A2(n8842), .ZN(n13042) );
  AOI22_X1 U11328 ( .A1(n11429), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n11430), 
        .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n8844) );
  INV_X1 U11329 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14709) );
  OR2_X1 U11330 ( .A1(n12668), .A2(n14709), .ZN(n8843) );
  OAI211_X1 U11331 ( .C1(n13042), .C2(n11403), .A(n8844), .B(n8843), .ZN(
        n12788) );
  NAND2_X1 U11332 ( .A1(n12788), .A2(n9183), .ZN(n9134) );
  NAND2_X1 U11333 ( .A1(n10398), .A2(n12684), .ZN(n8848) );
  NAND2_X1 U11334 ( .A1(n9111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8845) );
  MUX2_X1 U11335 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8845), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8846) );
  AND2_X1 U11336 ( .A1(n8846), .A2(n8837), .ZN(n14703) );
  AOI22_X1 U11337 ( .A1(n12685), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9135), 
        .B2(n14703), .ZN(n8847) );
  XNOR2_X1 U11338 ( .A(n12618), .B(n8849), .ZN(n9132) );
  INV_X1 U11339 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U11340 ( .A1(n9118), .A2(n8850), .ZN(n8851) );
  NAND2_X1 U11341 ( .A1(n8852), .A2(n8851), .ZN(n11290) );
  OR2_X1 U11342 ( .A1(n11290), .A2(n11403), .ZN(n8857) );
  NAND2_X1 U11343 ( .A1(n11430), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8856) );
  INV_X1 U11344 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8853) );
  OR2_X1 U11345 ( .A1(n12668), .A2(n8853), .ZN(n8855) );
  INV_X1 U11346 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11291) );
  OR2_X1 U11347 ( .A1(n9239), .A2(n11291), .ZN(n8854) );
  NAND4_X1 U11348 ( .A1(n8857), .A2(n8856), .A3(n8855), .A4(n8854), .ZN(n13028) );
  NAND2_X1 U11349 ( .A1(n13028), .A2(n9183), .ZN(n9131) );
  NAND2_X1 U11350 ( .A1(n8896), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U11351 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8858) );
  XNOR2_X1 U11352 ( .A(n8858), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9550) );
  INV_X1 U11353 ( .A(n9550), .ZN(n8859) );
  NAND2_X1 U11354 ( .A1(n8917), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8864) );
  INV_X1 U11355 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9551) );
  NAND3_X1 U11356 ( .A1(n8864), .A2(n8863), .A3(n8862), .ZN(n8866) );
  INV_X1 U11357 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10052) );
  CLKBUF_X1 U11358 ( .A(n10013), .Z(n12513) );
  NOR2_X1 U11359 ( .A1(n12513), .A2(n12913), .ZN(n8879) );
  INV_X1 U11360 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U11361 ( .A1(n12680), .A2(SI_0_), .ZN(n8868) );
  NAND2_X1 U11362 ( .A1(n8868), .A2(n8867), .ZN(n8870) );
  NAND2_X1 U11363 ( .A1(n8870), .A2(n8869), .ZN(n13179) );
  MUX2_X1 U11364 ( .A(n8871), .B(n13179), .S(n9536), .Z(n10025) );
  INV_X1 U11365 ( .A(n10025), .ZN(n10024) );
  NOR2_X1 U11366 ( .A1(n8901), .A2(n10024), .ZN(n9856) );
  NAND2_X1 U11367 ( .A1(n8917), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8876) );
  INV_X1 U11368 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9849) );
  INV_X1 U11369 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9659) );
  OR2_X1 U11370 ( .A1(n8904), .A2(n9659), .ZN(n8874) );
  INV_X1 U11371 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U11372 ( .A1(n12805), .A2(n10024), .ZN(n10014) );
  AND2_X1 U11373 ( .A1(n10017), .A2(n8877), .ZN(n9901) );
  INV_X1 U11374 ( .A(n8878), .ZN(n8881) );
  INV_X1 U11375 ( .A(n8879), .ZN(n8880) );
  NAND2_X1 U11376 ( .A1(n8881), .A2(n8880), .ZN(n8882) );
  OR2_X1 U11377 ( .A1(n8883), .A2(n8805), .ZN(n8884) );
  XNOR2_X1 U11378 ( .A(n8884), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U11379 ( .A1(n9135), .A2(n9573), .ZN(n8885) );
  XNOR2_X1 U11380 ( .A(n8901), .B(n6589), .ZN(n8892) );
  NAND2_X1 U11381 ( .A1(n8917), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8891) );
  INV_X1 U11382 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10105) );
  OR2_X1 U11383 ( .A1(n8902), .A2(n10105), .ZN(n8890) );
  INV_X1 U11384 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8887) );
  OR2_X1 U11385 ( .A1(n8904), .A2(n8887), .ZN(n8889) );
  INV_X1 U11386 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9564) );
  OR2_X1 U11387 ( .A1(n9239), .A2(n9564), .ZN(n8888) );
  NAND4_X2 U11388 ( .A1(n8891), .A2(n8890), .A3(n8889), .A4(n8888), .ZN(n12802) );
  NAND2_X1 U11389 ( .A1(n12802), .A2(n8877), .ZN(n8893) );
  XNOR2_X1 U11390 ( .A(n8892), .B(n8893), .ZN(n9974) );
  INV_X1 U11391 ( .A(n8892), .ZN(n8894) );
  NAND2_X1 U11392 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  AND2_X1 U11393 ( .A1(n9982), .A2(n8895), .ZN(n9833) );
  NAND2_X1 U11394 ( .A1(n12685), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11395 ( .A1(n8883), .A2(n8897), .ZN(n9047) );
  NAND2_X1 U11396 ( .A1(n9047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8898) );
  XNOR2_X1 U11397 ( .A(n8898), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U11398 ( .A1(n9135), .A2(n9576), .ZN(n8899) );
  XNOR2_X1 U11399 ( .A(n8901), .B(n12511), .ZN(n8909) );
  NAND2_X1 U11400 ( .A1(n11430), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8908) );
  OR2_X1 U11401 ( .A1(n8902), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8907) );
  INV_X1 U11402 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8903) );
  OR2_X1 U11403 ( .A1(n8904), .A2(n8903), .ZN(n8906) );
  INV_X1 U11404 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9565) );
  OR2_X1 U11405 ( .A1(n9239), .A2(n9565), .ZN(n8905) );
  AND2_X1 U11406 ( .A1(n12801), .A2(n8877), .ZN(n8910) );
  NAND2_X1 U11407 ( .A1(n8909), .A2(n8910), .ZN(n8923) );
  INV_X1 U11408 ( .A(n8909), .ZN(n10003) );
  INV_X1 U11409 ( .A(n8910), .ZN(n8911) );
  NAND2_X1 U11410 ( .A1(n10003), .A2(n8911), .ZN(n8912) );
  AND2_X1 U11411 ( .A1(n8923), .A2(n8912), .ZN(n9832) );
  NAND2_X1 U11412 ( .A1(n8928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8914) );
  XNOR2_X1 U11413 ( .A(n8913), .B(n8914), .ZN(n14620) );
  NAND2_X1 U11414 ( .A1(n12685), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8915) );
  OAI211_X1 U11415 ( .C1(n9536), .C2(n14620), .A(n8916), .B(n8915), .ZN(n12536) );
  XNOR2_X1 U11416 ( .A(n12433), .B(n12536), .ZN(n8925) );
  NAND2_X1 U11417 ( .A1(n11429), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8922) );
  INV_X1 U11418 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8918) );
  OR2_X1 U11419 ( .A1(n12670), .A2(n8918), .ZN(n8921) );
  OAI21_X1 U11420 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8935), .ZN(n10426) );
  OR2_X1 U11421 ( .A1(n11403), .A2(n10426), .ZN(n8920) );
  INV_X1 U11422 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9578) );
  OR2_X1 U11423 ( .A1(n12668), .A2(n9578), .ZN(n8919) );
  NAND2_X1 U11424 ( .A1(n12800), .A2(n8877), .ZN(n8926) );
  XNOR2_X1 U11425 ( .A(n8925), .B(n8926), .ZN(n10004) );
  AND2_X1 U11426 ( .A1(n10004), .A2(n8923), .ZN(n8924) );
  NAND2_X1 U11427 ( .A1(n10002), .A2(n8924), .ZN(n10001) );
  INV_X1 U11428 ( .A(n8925), .ZN(n9914) );
  NAND2_X1 U11429 ( .A1(n9914), .A2(n8926), .ZN(n8927) );
  NAND2_X1 U11430 ( .A1(n10001), .A2(n8927), .ZN(n8941) );
  NAND2_X1 U11431 ( .A1(n9488), .A2(n12684), .ZN(n8932) );
  INV_X1 U11432 ( .A(n8928), .ZN(n8929) );
  NAND2_X1 U11433 ( .A1(n8929), .A2(n8913), .ZN(n8946) );
  NAND2_X1 U11434 ( .A1(n8946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8930) );
  XNOR2_X1 U11435 ( .A(n8930), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U11436 ( .A1(n12685), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9135), 
        .B2(n9590), .ZN(n8931) );
  NAND2_X1 U11437 ( .A1(n8932), .A2(n8931), .ZN(n12545) );
  XNOR2_X1 U11438 ( .A(n12433), .B(n12545), .ZN(n8942) );
  NAND2_X1 U11439 ( .A1(n11429), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8940) );
  INV_X1 U11440 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8933) );
  OR2_X1 U11441 ( .A1(n12670), .A2(n8933), .ZN(n8939) );
  INV_X1 U11442 ( .A(n8934), .ZN(n8953) );
  NAND2_X1 U11443 ( .A1(n8935), .A2(n9909), .ZN(n8936) );
  NAND2_X1 U11444 ( .A1(n8953), .A2(n8936), .ZN(n10440) );
  OR2_X1 U11445 ( .A1(n11403), .A2(n10440), .ZN(n8938) );
  OR2_X1 U11446 ( .A1(n12668), .A2(n14833), .ZN(n8937) );
  NAND4_X1 U11447 ( .A1(n8940), .A2(n8939), .A3(n8938), .A4(n8937), .ZN(n12799) );
  NAND2_X1 U11448 ( .A1(n12799), .A2(n9183), .ZN(n8943) );
  XNOR2_X1 U11449 ( .A(n8942), .B(n8943), .ZN(n9913) );
  INV_X1 U11450 ( .A(n8942), .ZN(n8944) );
  NAND2_X1 U11451 ( .A1(n8944), .A2(n8943), .ZN(n8945) );
  NAND2_X1 U11452 ( .A1(n9494), .A2(n12684), .ZN(n8949) );
  NAND2_X1 U11453 ( .A1(n8962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8947) );
  XNOR2_X1 U11454 ( .A(n8947), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14635) );
  AOI22_X1 U11455 ( .A1(n12685), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9135), 
        .B2(n14635), .ZN(n8948) );
  NAND2_X1 U11456 ( .A1(n8949), .A2(n8948), .ZN(n12549) );
  XNOR2_X1 U11457 ( .A(n12433), .B(n12549), .ZN(n10114) );
  NAND2_X1 U11458 ( .A1(n11430), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8958) );
  INV_X1 U11459 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8950) );
  OR2_X1 U11460 ( .A1(n12668), .A2(n8950), .ZN(n8957) );
  INV_X1 U11461 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8951) );
  OR2_X1 U11462 ( .A1(n9239), .A2(n8951), .ZN(n8956) );
  INV_X1 U11463 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U11464 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  NAND2_X1 U11465 ( .A1(n8970), .A2(n8954), .ZN(n10038) );
  OR2_X1 U11466 ( .A1(n11403), .A2(n10038), .ZN(n8955) );
  NAND4_X1 U11467 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(n12798) );
  AND2_X1 U11468 ( .A1(n12798), .A2(n8877), .ZN(n8959) );
  NAND2_X1 U11469 ( .A1(n10114), .A2(n8959), .ZN(n8961) );
  OR2_X1 U11470 ( .A1(n10114), .A2(n8959), .ZN(n8960) );
  NAND2_X1 U11471 ( .A1(n8961), .A2(n8960), .ZN(n10034) );
  NAND2_X1 U11472 ( .A1(n10036), .A2(n8961), .ZN(n8980) );
  NAND2_X1 U11473 ( .A1(n9516), .A2(n12684), .ZN(n8967) );
  INV_X1 U11474 ( .A(n8962), .ZN(n8964) );
  INV_X1 U11475 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11476 ( .A1(n8964), .A2(n8963), .ZN(n8981) );
  NAND2_X1 U11477 ( .A1(n8981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8965) );
  XNOR2_X1 U11478 ( .A(n8965), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9723) );
  AOI22_X1 U11479 ( .A1(n12685), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9135), 
        .B2(n9723), .ZN(n8966) );
  NAND2_X1 U11480 ( .A1(n8967), .A2(n8966), .ZN(n12558) );
  XNOR2_X1 U11481 ( .A(n12558), .B(n12433), .ZN(n8976) );
  NAND2_X1 U11482 ( .A1(n11430), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8975) );
  INV_X1 U11483 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8968) );
  OR2_X1 U11484 ( .A1(n12668), .A2(n8968), .ZN(n8974) );
  INV_X1 U11485 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8969) );
  OR2_X1 U11486 ( .A1(n9239), .A2(n8969), .ZN(n8973) );
  NAND2_X1 U11487 ( .A1(n8970), .A2(n10121), .ZN(n8971) );
  NAND2_X1 U11488 ( .A1(n8987), .A2(n8971), .ZN(n10118) );
  OR2_X1 U11489 ( .A1(n11403), .A2(n10118), .ZN(n8972) );
  NAND4_X1 U11490 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(n12797) );
  AND2_X1 U11491 ( .A1(n12797), .A2(n8877), .ZN(n8977) );
  NAND2_X1 U11492 ( .A1(n8976), .A2(n8977), .ZN(n8994) );
  INV_X1 U11493 ( .A(n8976), .ZN(n12451) );
  INV_X1 U11494 ( .A(n8977), .ZN(n8978) );
  NAND2_X1 U11495 ( .A1(n12451), .A2(n8978), .ZN(n8979) );
  AND2_X1 U11496 ( .A1(n8994), .A2(n8979), .ZN(n10113) );
  NAND2_X1 U11497 ( .A1(n9528), .A2(n12684), .ZN(n8984) );
  NAND2_X1 U11498 ( .A1(n8998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8982) );
  XNOR2_X1 U11499 ( .A(n8982), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U11500 ( .A1(n12685), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9135), 
        .B2(n9797), .ZN(n8983) );
  XNOR2_X1 U11501 ( .A(n12561), .B(n12433), .ZN(n8996) );
  NAND2_X1 U11502 ( .A1(n11429), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8993) );
  INV_X1 U11503 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8985) );
  OR2_X1 U11504 ( .A1(n12670), .A2(n8985), .ZN(n8992) );
  NAND2_X1 U11505 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  NAND2_X1 U11506 ( .A1(n9004), .A2(n8988), .ZN(n12449) );
  OR2_X1 U11507 ( .A1(n11403), .A2(n12449), .ZN(n8991) );
  INV_X1 U11508 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8989) );
  OR2_X1 U11509 ( .A1(n12668), .A2(n8989), .ZN(n8990) );
  NAND4_X1 U11510 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n12796) );
  NAND2_X1 U11511 ( .A1(n12796), .A2(n8877), .ZN(n8997) );
  XNOR2_X1 U11512 ( .A(n8996), .B(n8997), .ZN(n12452) );
  AND2_X1 U11513 ( .A1(n12452), .A2(n8994), .ZN(n8995) );
  INV_X1 U11514 ( .A(n8996), .ZN(n10382) );
  NAND2_X1 U11515 ( .A1(n9557), .A2(n12684), .ZN(n9001) );
  NAND2_X1 U11516 ( .A1(n9014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8999) );
  XNOR2_X1 U11517 ( .A(n8999), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U11518 ( .A1(n12685), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9135), 
        .B2(n9932), .ZN(n9000) );
  XNOR2_X1 U11519 ( .A(n14803), .B(n12433), .ZN(n9010) );
  NAND2_X1 U11520 ( .A1(n11430), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9009) );
  OR2_X1 U11521 ( .A1(n9239), .A2(n9798), .ZN(n9008) );
  INV_X1 U11522 ( .A(n9002), .ZN(n9036) );
  NAND2_X1 U11523 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  NAND2_X1 U11524 ( .A1(n9036), .A2(n9005), .ZN(n10701) );
  OR2_X1 U11525 ( .A1(n11403), .A2(n10701), .ZN(n9007) );
  INV_X1 U11526 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9936) );
  OR2_X1 U11527 ( .A1(n12668), .A2(n9936), .ZN(n9006) );
  NAND4_X1 U11528 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n12794) );
  NAND2_X1 U11529 ( .A1(n12794), .A2(n9183), .ZN(n9011) );
  INV_X1 U11530 ( .A(n9010), .ZN(n9012) );
  NAND2_X1 U11531 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  NAND2_X1 U11532 ( .A1(n10386), .A2(n9013), .ZN(n10882) );
  NAND2_X1 U11533 ( .A1(n9654), .A2(n12684), .ZN(n9019) );
  INV_X1 U11534 ( .A(n9014), .ZN(n9016) );
  INV_X1 U11535 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11536 ( .A1(n9016), .A2(n9015), .ZN(n9030) );
  NAND2_X1 U11537 ( .A1(n9030), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9017) );
  XNOR2_X1 U11538 ( .A(n9017), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U11539 ( .A1(n9135), .A2(n10929), .B1(n12685), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9018) );
  XNOR2_X1 U11540 ( .A(n14811), .B(n12433), .ZN(n9025) );
  NAND2_X1 U11541 ( .A1(n11429), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9024) );
  INV_X1 U11542 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9020) );
  OR2_X1 U11543 ( .A1(n12670), .A2(n9020), .ZN(n9023) );
  INV_X1 U11544 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9035) );
  XNOR2_X1 U11545 ( .A(n9036), .B(n9035), .ZN(n10876) );
  OR2_X1 U11546 ( .A1(n11403), .A2(n10876), .ZN(n9022) );
  INV_X1 U11547 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9935) );
  OR2_X1 U11548 ( .A1(n12668), .A2(n9935), .ZN(n9021) );
  NAND4_X1 U11549 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n12793) );
  AND2_X1 U11550 ( .A1(n12793), .A2(n9183), .ZN(n9026) );
  NAND2_X1 U11551 ( .A1(n9025), .A2(n9026), .ZN(n9044) );
  INV_X1 U11552 ( .A(n9025), .ZN(n10819) );
  INV_X1 U11553 ( .A(n9026), .ZN(n9027) );
  NAND2_X1 U11554 ( .A1(n10819), .A2(n9027), .ZN(n9028) );
  NAND2_X1 U11555 ( .A1(n9044), .A2(n9028), .ZN(n10883) );
  INV_X1 U11556 ( .A(n10883), .ZN(n9029) );
  NAND2_X1 U11557 ( .A1(n9696), .A2(n12684), .ZN(n9033) );
  OAI21_X1 U11558 ( .B1(n9030), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9031) );
  AOI22_X1 U11559 ( .A1(n12812), .A2(n9135), .B1(n12685), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U11560 ( .A1(n11430), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9043) );
  INV_X1 U11561 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10851) );
  OR2_X1 U11562 ( .A1(n9239), .A2(n10851), .ZN(n9042) );
  INV_X1 U11563 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9034) );
  OAI21_X1 U11564 ( .B1(n9036), .B2(n9035), .A(n9034), .ZN(n9038) );
  INV_X1 U11565 ( .A(n9037), .ZN(n9056) );
  NAND2_X1 U11566 ( .A1(n9038), .A2(n9056), .ZN(n10850) );
  OR2_X1 U11567 ( .A1(n11403), .A2(n10850), .ZN(n9041) );
  INV_X1 U11568 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9039) );
  OR2_X1 U11569 ( .A1(n12668), .A2(n9039), .ZN(n9040) );
  NAND4_X1 U11570 ( .A1(n9043), .A2(n9042), .A3(n9041), .A4(n9040), .ZN(n12792) );
  NAND2_X1 U11571 ( .A1(n12792), .A2(n9183), .ZN(n9045) );
  INV_X1 U11572 ( .A(n10888), .ZN(n9046) );
  NAND2_X1 U11573 ( .A1(n9786), .A2(n12684), .ZN(n9054) );
  INV_X1 U11574 ( .A(n9047), .ZN(n9051) );
  NAND4_X1 U11575 ( .A1(n9051), .A2(n9050), .A3(n9049), .A4(n9048), .ZN(n9068)
         );
  NAND2_X1 U11576 ( .A1(n9068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9052) );
  XNOR2_X1 U11577 ( .A(n9052), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U11578 ( .A1(n12685), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9135), 
        .B2(n10933), .ZN(n9053) );
  XNOR2_X1 U11579 ( .A(n12589), .B(n12433), .ZN(n9064) );
  NAND2_X1 U11580 ( .A1(n11430), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9062) );
  INV_X1 U11581 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10931) );
  OR2_X1 U11582 ( .A1(n9239), .A2(n10931), .ZN(n9061) );
  INV_X1 U11583 ( .A(n9055), .ZN(n9089) );
  INV_X1 U11584 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n15262) );
  NAND2_X1 U11585 ( .A1(n9056), .A2(n15262), .ZN(n9057) );
  NAND2_X1 U11586 ( .A1(n9089), .A2(n9057), .ZN(n11083) );
  OR2_X1 U11587 ( .A1(n11403), .A2(n11083), .ZN(n9060) );
  INV_X1 U11588 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9058) );
  OR2_X1 U11589 ( .A1(n12668), .A2(n9058), .ZN(n9059) );
  NAND4_X1 U11590 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n12791) );
  NAND2_X1 U11591 ( .A1(n12791), .A2(n9183), .ZN(n9065) );
  XNOR2_X1 U11592 ( .A(n9064), .B(n9065), .ZN(n10889) );
  NAND2_X1 U11593 ( .A1(n9063), .A2(n10889), .ZN(n10894) );
  INV_X1 U11594 ( .A(n9064), .ZN(n9066) );
  NAND2_X1 U11595 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  INV_X1 U11596 ( .A(n10986), .ZN(n9082) );
  NAND2_X1 U11597 ( .A1(n9826), .A2(n12684), .ZN(n9071) );
  OAI21_X1 U11598 ( .B1(n9068), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9069) );
  XNOR2_X1 U11599 ( .A(n9069), .B(P2_IR_REG_13__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U11600 ( .A1(n12685), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9135), 
        .B2(n14665), .ZN(n9070) );
  XNOR2_X1 U11601 ( .A(n12594), .B(n12433), .ZN(n9076) );
  NAND2_X1 U11602 ( .A1(n11430), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9075) );
  INV_X1 U11603 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10991) );
  XNOR2_X1 U11604 ( .A(n9089), .B(n10991), .ZN(n11032) );
  OR2_X1 U11605 ( .A1(n11403), .A2(n11032), .ZN(n9074) );
  INV_X1 U11606 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10919) );
  OR2_X1 U11607 ( .A1(n12668), .A2(n10919), .ZN(n9073) );
  INV_X1 U11608 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11033) );
  OR2_X1 U11609 ( .A1(n9239), .A2(n11033), .ZN(n9072) );
  NAND4_X1 U11610 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n14305) );
  AND2_X1 U11611 ( .A1(n14305), .A2(n9183), .ZN(n9077) );
  NAND2_X1 U11612 ( .A1(n9076), .A2(n9077), .ZN(n9083) );
  INV_X1 U11613 ( .A(n9076), .ZN(n9079) );
  INV_X1 U11614 ( .A(n9077), .ZN(n9078) );
  NAND2_X1 U11615 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  NAND2_X1 U11616 ( .A1(n9083), .A2(n9080), .ZN(n10985) );
  NAND2_X1 U11617 ( .A1(n9927), .A2(n12684), .ZN(n9087) );
  NAND2_X1 U11618 ( .A1(n9084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9085) );
  XNOR2_X1 U11619 ( .A(n9085), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U11620 ( .A1(n12685), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9135), 
        .B2(n12820), .ZN(n9086) );
  XNOR2_X1 U11621 ( .A(n12599), .B(n8849), .ZN(n9108) );
  NAND2_X1 U11622 ( .A1(n11430), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9094) );
  INV_X1 U11623 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9088) );
  OAI21_X1 U11624 ( .B1(n9089), .B2(n10991), .A(n9088), .ZN(n9090) );
  NAND2_X1 U11625 ( .A1(n9100), .A2(n9090), .ZN(n14315) );
  OR2_X1 U11626 ( .A1(n11403), .A2(n14315), .ZN(n9093) );
  INV_X1 U11627 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10923) );
  OR2_X1 U11628 ( .A1(n12668), .A2(n10923), .ZN(n9092) );
  INV_X1 U11629 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11156) );
  OR2_X1 U11630 ( .A1(n9239), .A2(n11156), .ZN(n9091) );
  NAND4_X1 U11631 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n12790) );
  NAND2_X1 U11632 ( .A1(n12790), .A2(n9183), .ZN(n9107) );
  XNOR2_X1 U11633 ( .A(n9108), .B(n9107), .ZN(n14300) );
  NAND2_X1 U11634 ( .A1(n10044), .A2(n12684), .ZN(n9098) );
  NAND2_X1 U11635 ( .A1(n9095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9096) );
  XNOR2_X1 U11636 ( .A(n9096), .B(n7417), .ZN(n12830) );
  INV_X1 U11637 ( .A(n12830), .ZN(n14676) );
  AOI22_X1 U11638 ( .A1(n12685), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9135), 
        .B2(n14676), .ZN(n9097) );
  XNOR2_X1 U11639 ( .A(n13137), .B(n8849), .ZN(n14317) );
  NAND2_X1 U11640 ( .A1(n11430), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9106) );
  INV_X1 U11641 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14672) );
  OR2_X1 U11642 ( .A1(n12668), .A2(n14672), .ZN(n9105) );
  INV_X1 U11643 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9099) );
  NAND2_X1 U11644 ( .A1(n9100), .A2(n9099), .ZN(n9101) );
  NAND2_X1 U11645 ( .A1(n9116), .A2(n9101), .ZN(n11259) );
  OR2_X1 U11646 ( .A1(n11403), .A2(n11259), .ZN(n9104) );
  INV_X1 U11647 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9102) );
  OR2_X1 U11648 ( .A1(n9239), .A2(n9102), .ZN(n9103) );
  NAND4_X1 U11649 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(n14307) );
  NAND2_X1 U11650 ( .A1(n14307), .A2(n9183), .ZN(n11207) );
  AND2_X1 U11651 ( .A1(n9108), .A2(n9107), .ZN(n11204) );
  AOI21_X1 U11652 ( .B1(n14317), .B2(n11207), .A(n11204), .ZN(n9109) );
  NAND2_X1 U11653 ( .A1(n10152), .A2(n12684), .ZN(n9114) );
  NAND2_X1 U11654 ( .A1(n6710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9110) );
  MUX2_X1 U11655 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9110), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9112) );
  AOI22_X1 U11656 ( .A1(n12685), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9135), 
        .B2(n14689), .ZN(n9113) );
  XNOR2_X1 U11657 ( .A(n14327), .B(n12433), .ZN(n9128) );
  NAND2_X1 U11658 ( .A1(n11429), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U11659 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  NAND2_X1 U11660 ( .A1(n9118), .A2(n9117), .ZN(n14330) );
  OR2_X1 U11661 ( .A1(n11403), .A2(n14330), .ZN(n9123) );
  INV_X1 U11662 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9119) );
  OR2_X1 U11663 ( .A1(n12668), .A2(n9119), .ZN(n9122) );
  INV_X1 U11664 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9120) );
  OR2_X1 U11665 ( .A1(n12670), .A2(n9120), .ZN(n9121) );
  NAND4_X1 U11666 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n12789) );
  NAND2_X1 U11667 ( .A1(n12789), .A2(n9183), .ZN(n9129) );
  XNOR2_X1 U11668 ( .A(n9128), .B(n9129), .ZN(n14322) );
  NAND2_X1 U11669 ( .A1(n9127), .A2(n9126), .ZN(n14321) );
  INV_X1 U11670 ( .A(n9128), .ZN(n11165) );
  NAND2_X1 U11671 ( .A1(n11165), .A2(n9129), .ZN(n9130) );
  XNOR2_X1 U11672 ( .A(n9132), .B(n9131), .ZN(n11167) );
  AOI21_X2 U11673 ( .B1(n14321), .B2(n9130), .A(n11167), .ZN(n11161) );
  NAND2_X1 U11674 ( .A1(n10831), .A2(n12684), .ZN(n9137) );
  AOI22_X1 U11675 ( .A1(n12685), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12842), 
        .B2(n9135), .ZN(n9136) );
  XNOR2_X1 U11676 ( .A(n13114), .B(n8849), .ZN(n9145) );
  INV_X1 U11677 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9143) );
  INV_X1 U11678 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11679 ( .A1(n9139), .A2(n9138), .ZN(n9140) );
  NAND2_X1 U11680 ( .A1(n9160), .A2(n9140), .ZN(n13014) );
  OR2_X1 U11681 ( .A1(n13014), .A2(n11403), .ZN(n9142) );
  AOI22_X1 U11682 ( .A1(n8861), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n11430), 
        .B2(P2_REG0_REG_19__SCAN_IN), .ZN(n9141) );
  OAI211_X1 U11683 ( .C1(n9239), .C2(n9143), .A(n9142), .B(n9141), .ZN(n13031)
         );
  NAND2_X1 U11684 ( .A1(n13031), .A2(n9183), .ZN(n9144) );
  NAND2_X1 U11685 ( .A1(n9145), .A2(n9144), .ZN(n12420) );
  NOR2_X1 U11686 ( .A1(n9145), .A2(n9144), .ZN(n12422) );
  OR2_X1 U11687 ( .A1(n11592), .A2(n12661), .ZN(n9147) );
  NAND2_X1 U11688 ( .A1(n12685), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9146) );
  XNOR2_X1 U11689 ( .A(n13109), .B(n12433), .ZN(n9155) );
  XNOR2_X1 U11690 ( .A(n9160), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U11691 ( .A1(n12991), .A2(n9236), .ZN(n9153) );
  INV_X1 U11692 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11693 ( .A1(n11429), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11694 ( .A1(n11430), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9148) );
  OAI211_X1 U11695 ( .C1(n9150), .C2(n12668), .A(n9149), .B(n9148), .ZN(n9151)
         );
  INV_X1 U11696 ( .A(n9151), .ZN(n9152) );
  NAND2_X1 U11697 ( .A1(n9153), .A2(n9152), .ZN(n12787) );
  AND2_X1 U11698 ( .A1(n12787), .A2(n9183), .ZN(n9154) );
  NOR2_X1 U11699 ( .A1(n9155), .A2(n9154), .ZN(n12484) );
  NAND2_X1 U11700 ( .A1(n9155), .A2(n9154), .ZN(n12485) );
  OR2_X1 U11701 ( .A1(n10970), .A2(n12661), .ZN(n9157) );
  NAND2_X1 U11702 ( .A1(n12685), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9156) );
  XNOR2_X1 U11703 ( .A(n13105), .B(n12433), .ZN(n9167) );
  OAI21_X1 U11704 ( .B1(n9160), .B2(n9159), .A(n9158), .ZN(n9161) );
  AND2_X1 U11705 ( .A1(n9161), .A2(n9175), .ZN(n12982) );
  NAND2_X1 U11706 ( .A1(n12982), .A2(n9236), .ZN(n9166) );
  INV_X1 U11707 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15361) );
  NAND2_X1 U11708 ( .A1(n11429), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11709 ( .A1(n8861), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9162) );
  OAI211_X1 U11710 ( .C1(n12670), .C2(n15361), .A(n9163), .B(n9162), .ZN(n9164) );
  INV_X1 U11711 ( .A(n9164), .ZN(n9165) );
  NAND2_X1 U11712 ( .A1(n9166), .A2(n9165), .ZN(n12997) );
  NAND2_X1 U11713 ( .A1(n12997), .A2(n9183), .ZN(n9168) );
  XNOR2_X1 U11714 ( .A(n9167), .B(n9168), .ZN(n12458) );
  XNOR2_X1 U11715 ( .A(n9172), .B(n9171), .ZN(n11106) );
  NAND2_X1 U11716 ( .A1(n11106), .A2(n12684), .ZN(n9174) );
  NAND2_X1 U11717 ( .A1(n12685), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9173) );
  XNOR2_X1 U11718 ( .A(n13099), .B(n12433), .ZN(n9185) );
  INV_X1 U11719 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U11720 ( .A1(n9175), .A2(n11578), .ZN(n9176) );
  AND2_X1 U11721 ( .A1(n9192), .A2(n9176), .ZN(n12967) );
  NAND2_X1 U11722 ( .A1(n12967), .A2(n9236), .ZN(n9182) );
  INV_X1 U11723 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11724 ( .A1(n11430), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11725 ( .A1(n11429), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9177) );
  OAI211_X1 U11726 ( .C1(n12668), .C2(n9179), .A(n9178), .B(n9177), .ZN(n9180)
         );
  INV_X1 U11727 ( .A(n9180), .ZN(n9181) );
  NAND2_X1 U11728 ( .A1(n9182), .A2(n9181), .ZN(n12945) );
  NAND2_X1 U11729 ( .A1(n12945), .A2(n9183), .ZN(n9184) );
  INV_X1 U11730 ( .A(n9190), .ZN(n9201) );
  NAND2_X1 U11731 ( .A1(n11171), .A2(n12684), .ZN(n9188) );
  NAND2_X1 U11732 ( .A1(n12685), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9187) );
  XNOR2_X1 U11733 ( .A(n13094), .B(n12433), .ZN(n9200) );
  INV_X1 U11734 ( .A(n9200), .ZN(n9189) );
  INV_X1 U11735 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U11736 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  NAND2_X1 U11737 ( .A1(n9204), .A2(n9193), .ZN(n12948) );
  OR2_X1 U11738 ( .A1(n12948), .A2(n11403), .ZN(n9199) );
  INV_X1 U11739 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U11740 ( .A1(n11430), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11741 ( .A1(n11429), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9194) );
  OAI211_X1 U11742 ( .C1(n9196), .C2(n12668), .A(n9195), .B(n9194), .ZN(n9197)
         );
  INV_X1 U11743 ( .A(n9197), .ZN(n9198) );
  NAND2_X1 U11744 ( .A1(n9199), .A2(n9198), .ZN(n12786) );
  INV_X1 U11745 ( .A(n12786), .ZN(n12927) );
  OR2_X1 U11746 ( .A1(n11202), .A2(n12661), .ZN(n9203) );
  NAND2_X1 U11747 ( .A1(n12685), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U11748 ( .A(n13089), .B(n12433), .ZN(n12466) );
  NAND2_X1 U11749 ( .A1(n9204), .A2(n12474), .ZN(n9205) );
  AND2_X1 U11750 ( .A1(n9216), .A2(n9205), .ZN(n12932) );
  NAND2_X1 U11751 ( .A1(n12932), .A2(n9236), .ZN(n9211) );
  INV_X1 U11752 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11753 ( .A1(n11430), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11754 ( .A1(n11429), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9206) );
  OAI211_X1 U11755 ( .C1(n12668), .C2(n9208), .A(n9207), .B(n9206), .ZN(n9209)
         );
  INV_X1 U11756 ( .A(n9209), .ZN(n9210) );
  AND2_X1 U11757 ( .A1(n12944), .A2(n9183), .ZN(n9212) );
  NAND2_X1 U11758 ( .A1(n12466), .A2(n9212), .ZN(n9213) );
  OAI21_X1 U11759 ( .B1(n12466), .B2(n9212), .A(n9213), .ZN(n12479) );
  NAND2_X1 U11760 ( .A1(n13176), .A2(n12684), .ZN(n9215) );
  NAND2_X1 U11761 ( .A1(n12685), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U11762 ( .A(n12915), .B(n8849), .ZN(n9223) );
  XNOR2_X1 U11763 ( .A(n9216), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n12918) );
  NAND2_X1 U11764 ( .A1(n12918), .A2(n9236), .ZN(n9222) );
  INV_X1 U11765 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11766 ( .A1(n11429), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11767 ( .A1(n11430), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9217) );
  OAI211_X1 U11768 ( .C1(n9219), .C2(n12668), .A(n9218), .B(n9217), .ZN(n9220)
         );
  INV_X1 U11769 ( .A(n9220), .ZN(n9221) );
  NOR2_X1 U11770 ( .A1(n12928), .A2(n12913), .ZN(n9224) );
  NAND2_X1 U11771 ( .A1(n9223), .A2(n9224), .ZN(n9228) );
  INV_X1 U11772 ( .A(n9223), .ZN(n12503) );
  INV_X1 U11773 ( .A(n9224), .ZN(n9225) );
  NAND2_X1 U11774 ( .A1(n12503), .A2(n9225), .ZN(n9226) );
  AND2_X1 U11775 ( .A1(n9228), .A2(n9226), .ZN(n12464) );
  XNOR2_X1 U11776 ( .A(n9227), .B(n9229), .ZN(n12504) );
  NAND2_X1 U11777 ( .A1(n13169), .A2(n12684), .ZN(n9231) );
  NAND2_X1 U11778 ( .A1(n12685), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9230) );
  XNOR2_X1 U11779 ( .A(n13072), .B(n8849), .ZN(n12430) );
  INV_X1 U11780 ( .A(n9234), .ZN(n9232) );
  INV_X1 U11781 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11782 ( .A1(n9234), .A2(n9233), .ZN(n9235) );
  NAND2_X1 U11783 ( .A1(n12884), .A2(n9236), .ZN(n9242) );
  INV_X1 U11784 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U11785 ( .A1(n8861), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11786 ( .A1(n11430), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9237) );
  OAI211_X1 U11787 ( .C1(n9239), .C2(n12886), .A(n9238), .B(n9237), .ZN(n9240)
         );
  INV_X1 U11788 ( .A(n9240), .ZN(n9241) );
  NOR2_X1 U11789 ( .A1(n12695), .A2(n12913), .ZN(n9243) );
  NAND2_X1 U11790 ( .A1(n12430), .A2(n9243), .ZN(n12441) );
  OAI21_X1 U11791 ( .B1(n12430), .B2(n9243), .A(n12441), .ZN(n9284) );
  NAND2_X1 U11792 ( .A1(n9251), .A2(n9245), .ZN(n9254) );
  NAND2_X1 U11793 ( .A1(n9254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9246) );
  MUX2_X1 U11794 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9246), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9247) );
  NAND2_X1 U11795 ( .A1(n9248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9250) );
  XNOR2_X1 U11796 ( .A(n11175), .B(P2_B_REG_SCAN_IN), .ZN(n9256) );
  INV_X1 U11797 ( .A(n9251), .ZN(n9252) );
  NAND2_X1 U11798 ( .A1(n9252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9253) );
  MUX2_X1 U11799 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9253), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9255) );
  NAND2_X1 U11800 ( .A1(n9255), .A2(n9254), .ZN(n13177) );
  NAND2_X1 U11801 ( .A1(n9256), .A2(n13177), .ZN(n9257) );
  NAND2_X1 U11802 ( .A1(n14724), .A2(n15260), .ZN(n9260) );
  INV_X1 U11803 ( .A(n11175), .ZN(n9258) );
  NAND2_X1 U11804 ( .A1(n9260), .A2(n9259), .ZN(n14750) );
  INV_X1 U11805 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15273) );
  NAND2_X1 U11806 ( .A1(n14724), .A2(n15273), .ZN(n9263) );
  INV_X1 U11807 ( .A(n13177), .ZN(n9261) );
  OR2_X1 U11808 ( .A1(n9261), .A2(n13174), .ZN(n9262) );
  NAND2_X1 U11809 ( .A1(n9263), .A2(n9262), .ZN(n9736) );
  INV_X1 U11810 ( .A(n9736), .ZN(n9842) );
  NOR2_X1 U11811 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .ZN(
        n9267) );
  NOR4_X1 U11812 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n9266) );
  NOR4_X1 U11813 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9265) );
  NOR4_X1 U11814 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9264) );
  NAND4_X1 U11815 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n9273)
         );
  NOR4_X1 U11816 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9271) );
  NOR4_X1 U11817 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n9270) );
  NOR4_X1 U11818 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n9269) );
  NOR4_X1 U11819 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9268) );
  NAND4_X1 U11820 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9272)
         );
  OAI21_X1 U11821 ( .B1(n9273), .B2(n9272), .A(n14724), .ZN(n9844) );
  NAND3_X1 U11822 ( .A1(n9739), .A2(n9842), .A3(n9844), .ZN(n9302) );
  NOR2_X1 U11823 ( .A1(n13177), .A2(n11175), .ZN(n9274) );
  NAND2_X1 U11824 ( .A1(n13174), .A2(n9274), .ZN(n9444) );
  INV_X1 U11825 ( .A(n9275), .ZN(n9276) );
  NAND2_X1 U11826 ( .A1(n9276), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9278) );
  AND2_X1 U11827 ( .A1(n9444), .A2(n11172), .ZN(n9289) );
  INV_X1 U11828 ( .A(n9534), .ZN(n9280) );
  NAND2_X1 U11829 ( .A1(n6559), .A2(n12762), .ZN(n12764) );
  NAND3_X1 U11830 ( .A1(n14751), .A2(n9280), .A3(n14797), .ZN(n9281) );
  NOR2_X1 U11831 ( .A1(n6559), .A2(n9730), .ZN(n10051) );
  NAND2_X1 U11832 ( .A1(n14751), .A2(n10051), .ZN(n9286) );
  OR2_X1 U11833 ( .A1(n9302), .A2(n9286), .ZN(n9288) );
  OR2_X1 U11834 ( .A1(n12725), .A2(n9730), .ZN(n9737) );
  INV_X1 U11835 ( .A(n9737), .ZN(n9287) );
  NAND2_X1 U11836 ( .A1(n9302), .A2(n9737), .ZN(n9291) );
  NAND2_X1 U11837 ( .A1(n12764), .A2(n9534), .ZN(n9843) );
  AND2_X1 U11838 ( .A1(n9289), .A2(n9843), .ZN(n9290) );
  NAND2_X1 U11839 ( .A1(n9291), .A2(n9290), .ZN(n9858) );
  INV_X1 U11840 ( .A(n14331), .ZN(n12489) );
  AOI22_X1 U11841 ( .A1(n12884), .A2(n12489), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9304) );
  NAND2_X1 U11842 ( .A1(n9292), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11442) );
  INV_X1 U11843 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11844 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NAND2_X1 U11845 ( .A1(n11442), .A2(n9295), .ZN(n12870) );
  INV_X1 U11846 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15195) );
  NAND2_X1 U11847 ( .A1(n11429), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11848 ( .A1(n11430), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9296) );
  OAI211_X1 U11849 ( .C1(n15195), .C2(n12668), .A(n9297), .B(n9296), .ZN(n9298) );
  INV_X1 U11850 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U11851 ( .A1(n9534), .A2(n9539), .ZN(n13006) );
  INV_X1 U11852 ( .A(n9539), .ZN(n9541) );
  OAI22_X1 U11853 ( .A1(n12692), .A2(n13006), .B1(n12912), .B2(n13004), .ZN(
        n12879) );
  INV_X1 U11854 ( .A(n12764), .ZN(n9301) );
  NAND2_X1 U11855 ( .A1(n14751), .A2(n9301), .ZN(n12777) );
  INV_X1 U11856 ( .A(n12438), .ZN(n14325) );
  NAND2_X1 U11857 ( .A1(n12879), .A2(n14325), .ZN(n9303) );
  OAI211_X1 U11858 ( .C1(n13072), .C2(n14310), .A(n9304), .B(n9303), .ZN(n9305) );
  INV_X1 U11859 ( .A(n9305), .ZN(n9306) );
  XNOR2_X1 U11860 ( .A(n12266), .B(n9316), .ZN(n11599) );
  NOR2_X1 U11861 ( .A1(n11599), .A2(n12079), .ZN(n11595) );
  AOI21_X1 U11862 ( .B1(n11599), .B2(n12079), .A(n11595), .ZN(n9402) );
  INV_X4 U11863 ( .A(n9316), .ZN(n11593) );
  XNOR2_X1 U11864 ( .A(n11593), .B(n9314), .ZN(n9336) );
  XNOR2_X1 U11865 ( .A(n9394), .B(n9315), .ZN(n9328) );
  XNOR2_X1 U11866 ( .A(n9328), .B(n12329), .ZN(n10400) );
  NAND2_X1 U11867 ( .A1(n9389), .A2(n8254), .ZN(n9318) );
  NOR2_X1 U11868 ( .A1(n6586), .A2(n9317), .ZN(n9320) );
  AND2_X1 U11869 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  NOR2_X1 U11870 ( .A1(n9324), .A2(n9321), .ZN(n10391) );
  INV_X1 U11871 ( .A(n9326), .ZN(n9389) );
  INV_X1 U11872 ( .A(n9324), .ZN(n9325) );
  XNOR2_X1 U11873 ( .A(n6586), .B(n12333), .ZN(n9327) );
  XNOR2_X1 U11874 ( .A(n9327), .B(n14979), .ZN(n10217) );
  XNOR2_X1 U11875 ( .A(n11593), .B(n9330), .ZN(n9332) );
  XNOR2_X1 U11876 ( .A(n9332), .B(n9331), .ZN(n10519) );
  XNOR2_X1 U11877 ( .A(n11593), .B(n11679), .ZN(n9335) );
  XNOR2_X1 U11878 ( .A(n9335), .B(n9334), .ZN(n11675) );
  XNOR2_X1 U11879 ( .A(n9336), .B(n11980), .ZN(n11719) );
  XNOR2_X1 U11880 ( .A(n9316), .B(n10779), .ZN(n11607) );
  XNOR2_X1 U11881 ( .A(n11593), .B(n9340), .ZN(n9341) );
  XNOR2_X1 U11882 ( .A(n9341), .B(n11126), .ZN(n11641) );
  INV_X1 U11883 ( .A(n9341), .ZN(n9342) );
  XNOR2_X1 U11884 ( .A(n11593), .B(n11125), .ZN(n9344) );
  XNOR2_X1 U11885 ( .A(n9344), .B(n14951), .ZN(n11124) );
  INV_X1 U11886 ( .A(n11124), .ZN(n9343) );
  INV_X1 U11887 ( .A(n9344), .ZN(n9346) );
  INV_X1 U11888 ( .A(n11624), .ZN(n9350) );
  XNOR2_X1 U11889 ( .A(n11593), .B(n11627), .ZN(n9351) );
  XNOR2_X1 U11890 ( .A(n9351), .B(n9348), .ZN(n11623) );
  INV_X1 U11891 ( .A(n11623), .ZN(n9349) );
  NAND2_X1 U11892 ( .A1(n9350), .A2(n9349), .ZN(n11625) );
  INV_X1 U11893 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U11894 ( .A1(n9352), .A2(n14275), .ZN(n9353) );
  XNOR2_X1 U11895 ( .A(n11593), .B(n14280), .ZN(n11313) );
  INV_X1 U11896 ( .A(n11313), .ZN(n9354) );
  XNOR2_X1 U11897 ( .A(n11593), .B(n14267), .ZN(n11315) );
  NAND2_X1 U11898 ( .A1(n11315), .A2(n14274), .ZN(n9356) );
  OAI21_X1 U11899 ( .B1(n9354), .B2(n11305), .A(n9356), .ZN(n9359) );
  NOR2_X1 U11900 ( .A1(n11313), .A2(n14259), .ZN(n9357) );
  INV_X1 U11901 ( .A(n11315), .ZN(n9355) );
  AOI22_X1 U11902 ( .A1(n9357), .A2(n9356), .B1(n11307), .B2(n9355), .ZN(n9358) );
  XNOR2_X1 U11903 ( .A(n11246), .B(n11593), .ZN(n9360) );
  NOR2_X1 U11904 ( .A1(n9360), .A2(n14258), .ZN(n11267) );
  NAND2_X1 U11905 ( .A1(n9360), .A2(n14258), .ZN(n11268) );
  XNOR2_X1 U11906 ( .A(n12316), .B(n11593), .ZN(n9361) );
  XNOR2_X1 U11907 ( .A(n9361), .B(n12251), .ZN(n11374) );
  INV_X1 U11908 ( .A(n9361), .ZN(n9362) );
  OAI22_X1 U11909 ( .A1(n11375), .A2(n11374), .B1(n9362), .B2(n11978), .ZN(
        n11739) );
  XNOR2_X1 U11910 ( .A(n12313), .B(n11593), .ZN(n9363) );
  XNOR2_X1 U11911 ( .A(n9363), .B(n11977), .ZN(n11738) );
  NAND2_X1 U11912 ( .A1(n11739), .A2(n11738), .ZN(n9365) );
  NAND2_X1 U11913 ( .A1(n9363), .A2(n12239), .ZN(n9364) );
  XOR2_X1 U11914 ( .A(n11593), .B(n12309), .Z(n11667) );
  NOR2_X1 U11915 ( .A1(n11667), .A2(n12223), .ZN(n11362) );
  XNOR2_X1 U11916 ( .A(n12303), .B(n11593), .ZN(n9366) );
  OR2_X1 U11917 ( .A1(n11362), .A2(n7547), .ZN(n9369) );
  NAND2_X1 U11918 ( .A1(n11667), .A2(n12223), .ZN(n11363) );
  NOR2_X1 U11919 ( .A1(n9366), .A2(n12240), .ZN(n11365) );
  INV_X1 U11920 ( .A(n11365), .ZN(n9367) );
  AND2_X1 U11921 ( .A1(n11363), .A2(n9367), .ZN(n9368) );
  XNOR2_X1 U11922 ( .A(n12300), .B(n9316), .ZN(n11712) );
  NAND2_X1 U11923 ( .A1(n11712), .A2(n12224), .ZN(n9371) );
  XNOR2_X1 U11924 ( .A(n12196), .B(n11593), .ZN(n9372) );
  XNOR2_X1 U11925 ( .A(n9372), .B(n12210), .ZN(n11633) );
  NAND2_X1 U11926 ( .A1(n11634), .A2(n11633), .ZN(n9374) );
  NAND2_X1 U11927 ( .A1(n9372), .A2(n11975), .ZN(n9373) );
  XNOR2_X1 U11928 ( .A(n12293), .B(n11593), .ZN(n9375) );
  XNOR2_X1 U11929 ( .A(n9375), .B(n12192), .ZN(n11695) );
  INV_X1 U11930 ( .A(n9375), .ZN(n9376) );
  NAND2_X1 U11931 ( .A1(n9376), .A2(n12192), .ZN(n9377) );
  XNOR2_X1 U11932 ( .A(n12289), .B(n11593), .ZN(n9378) );
  NAND2_X1 U11933 ( .A1(n9378), .A2(n12179), .ZN(n9379) );
  OAI21_X1 U11934 ( .B1(n9378), .B2(n12179), .A(n9379), .ZN(n11649) );
  INV_X1 U11935 ( .A(n9383), .ZN(n9381) );
  XNOR2_X1 U11936 ( .A(n12285), .B(n11593), .ZN(n9382) );
  INV_X1 U11937 ( .A(n9382), .ZN(n9380) );
  XNOR2_X1 U11938 ( .A(n12281), .B(n11593), .ZN(n9387) );
  INV_X1 U11939 ( .A(n9387), .ZN(n9386) );
  NAND2_X1 U11940 ( .A1(n6583), .A2(n9386), .ZN(n9388) );
  XNOR2_X1 U11941 ( .A(n9316), .B(n12279), .ZN(n9390) );
  NAND2_X1 U11942 ( .A1(n9390), .A2(n12139), .ZN(n11656) );
  INV_X1 U11943 ( .A(n9390), .ZN(n9391) );
  NAND2_X1 U11944 ( .A1(n9391), .A2(n11971), .ZN(n9392) );
  XNOR2_X1 U11945 ( .A(n12273), .B(n11593), .ZN(n9395) );
  NAND2_X1 U11946 ( .A1(n9395), .A2(n12125), .ZN(n9398) );
  INV_X1 U11947 ( .A(n9395), .ZN(n9396) );
  NAND2_X1 U11948 ( .A1(n9396), .A2(n11970), .ZN(n9397) );
  XNOR2_X1 U11949 ( .A(n12110), .B(n11593), .ZN(n9399) );
  NOR2_X1 U11950 ( .A1(n9399), .A2(n10445), .ZN(n9400) );
  AOI21_X1 U11951 ( .B1(n9399), .B2(n10445), .A(n9400), .ZN(n11729) );
  INV_X1 U11952 ( .A(n9400), .ZN(n9401) );
  NAND3_X1 U11953 ( .A1(n6564), .A2(n10581), .A3(n9403), .ZN(n9436) );
  NAND2_X1 U11954 ( .A1(n9430), .A2(n14988), .ZN(n9921) );
  NAND2_X1 U11955 ( .A1(n9308), .A2(n9403), .ZN(n9404) );
  INV_X1 U11956 ( .A(n9405), .ZN(n9406) );
  NAND2_X1 U11957 ( .A1(n9406), .A2(n11962), .ZN(n9407) );
  OR2_X1 U11958 ( .A1(n9407), .A2(n11772), .ZN(n9433) );
  OAI22_X1 U11959 ( .A1(n9436), .A2(n9921), .B1(n9432), .B2(n9433), .ZN(n9408)
         );
  INV_X1 U11960 ( .A(n14999), .ZN(n15008) );
  NAND2_X1 U11961 ( .A1(n9436), .A2(n15008), .ZN(n9409) );
  NAND2_X1 U11962 ( .A1(n9436), .A2(n9430), .ZN(n9414) );
  OAI211_X1 U11963 ( .C1(n11960), .C2(n11911), .A(n9446), .B(n10240), .ZN(
        n9410) );
  INV_X1 U11964 ( .A(n9410), .ZN(n9413) );
  INV_X1 U11965 ( .A(n9433), .ZN(n9411) );
  NAND2_X1 U11966 ( .A1(n9432), .A2(n9411), .ZN(n9412) );
  NAND3_X1 U11967 ( .A1(n9414), .A2(n9413), .A3(n9412), .ZN(n9415) );
  NAND2_X1 U11968 ( .A1(n9415), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9418) );
  AND2_X1 U11969 ( .A1(n10238), .A2(n11960), .ZN(n11964) );
  NAND2_X1 U11970 ( .A1(n11964), .A2(n11948), .ZN(n9435) );
  INV_X1 U11971 ( .A(n9435), .ZN(n9416) );
  NAND2_X1 U11972 ( .A1(n9432), .A2(n9416), .ZN(n9417) );
  NAND2_X2 U11973 ( .A1(n9418), .A2(n9417), .ZN(n11741) );
  INV_X1 U11974 ( .A(n9432), .ZN(n9420) );
  AND2_X1 U11975 ( .A1(n11964), .A2(n14977), .ZN(n9419) );
  NAND2_X1 U11976 ( .A1(n11964), .A2(n14980), .ZN(n9421) );
  NOR2_X2 U11977 ( .A1(n9432), .A2(n9421), .ZN(n11731) );
  AOI22_X1 U11978 ( .A1(n10445), .A2(n11731), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9422) );
  OAI21_X1 U11979 ( .B1(n12093), .B2(n11733), .A(n9422), .ZN(n9423) );
  AOI21_X1 U11980 ( .B1(n12094), .B2(n11741), .A(n9423), .ZN(n9424) );
  OAI21_X1 U11981 ( .B1(n9425), .B2(n11737), .A(n9424), .ZN(n9426) );
  NAND2_X1 U11982 ( .A1(n9428), .A2(n9427), .ZN(P3_U3154) );
  INV_X1 U11983 ( .A(n9430), .ZN(n9431) );
  OAI22_X1 U11984 ( .A1(n9436), .A2(n9433), .B1(n9432), .B2(n9431), .ZN(n9434)
         );
  NAND2_X1 U11985 ( .A1(n9434), .A2(n10238), .ZN(n9438) );
  NAND2_X1 U11986 ( .A1(n15056), .A2(n9439), .ZN(n9440) );
  NAND2_X1 U11987 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  INV_X1 U11988 ( .A(n15054), .ZN(n14288) );
  NAND2_X1 U11989 ( .A1(n9442), .A2(n7559), .ZN(P3_U3456) );
  INV_X1 U11990 ( .A(n11172), .ZN(n9443) );
  NOR2_X1 U11991 ( .A1(n9444), .A2(n9443), .ZN(n9538) );
  INV_X1 U11992 ( .A(n9486), .ZN(n9445) );
  NOR2_X1 U11993 ( .A1(n8042), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14162) );
  INV_X2 U11994 ( .A(n14162), .ZN(n14154) );
  INV_X1 U11995 ( .A(n9447), .ZN(n9449) );
  AND2_X1 U11996 ( .A1(n12680), .A2(P3_U3151), .ZN(n14161) );
  INV_X2 U11997 ( .A(n14161), .ZN(n12417) );
  OAI222_X1 U11998 ( .A1(n14154), .A2(n9449), .B1(n12417), .B2(n9448), .C1(
        n10675), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U11999 ( .A(n9450), .ZN(n9451) );
  OAI222_X1 U12000 ( .A1(P3_U3151), .A2(n10255), .B1(n12417), .B2(n9452), .C1(
        n14154), .C2(n9451), .ZN(P3_U3294) );
  INV_X1 U12001 ( .A(SI_5_), .ZN(n9453) );
  OAI222_X1 U12002 ( .A1(n14154), .A2(n9454), .B1(n12417), .B2(n9453), .C1(
        n10564), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12003 ( .A(SI_4_), .ZN(n9456) );
  OAI222_X1 U12004 ( .A1(P3_U3151), .A2(n10314), .B1(n12417), .B2(n9456), .C1(
        n14154), .C2(n9455), .ZN(P3_U3291) );
  INV_X1 U12005 ( .A(SI_7_), .ZN(n9457) );
  OAI222_X1 U12006 ( .A1(n10352), .A2(P3_U3151), .B1(n14154), .B2(n9458), .C1(
        n9457), .C2(n12417), .ZN(P3_U3288) );
  INV_X1 U12007 ( .A(n9459), .ZN(n9461) );
  OAI222_X1 U12008 ( .A1(n10550), .A2(P3_U3151), .B1(n14154), .B2(n9461), .C1(
        n9460), .C2(n12417), .ZN(P3_U3289) );
  INV_X1 U12009 ( .A(n9462), .ZN(n9464) );
  OAI222_X1 U12010 ( .A1(n15154), .A2(P3_U3151), .B1(n14154), .B2(n9464), .C1(
        n9463), .C2(n12417), .ZN(P3_U3295) );
  INV_X1 U12011 ( .A(n10374), .ZN(n10285) );
  INV_X1 U12012 ( .A(SI_3_), .ZN(n9465) );
  OAI222_X1 U12013 ( .A1(n10285), .A2(P3_U3151), .B1(n14154), .B2(n9466), .C1(
        n9465), .C2(n12417), .ZN(P3_U3292) );
  OAI222_X1 U12014 ( .A1(n7132), .A2(P3_U3151), .B1(n14154), .B2(n9468), .C1(
        n9467), .C2(n12417), .ZN(P3_U3293) );
  AND2_X1 U12015 ( .A1(n12680), .A2(P2_U3088), .ZN(n13164) );
  INV_X2 U12016 ( .A(n13164), .ZN(n13178) );
  INV_X1 U12017 ( .A(n9573), .ZN(n9563) );
  OAI222_X1 U12018 ( .A1(n13160), .A2(n9470), .B1(n13178), .B2(n9501), .C1(
        P2_U3088), .C2(n9563), .ZN(P2_U3325) );
  INV_X1 U12019 ( .A(n9576), .ZN(n9653) );
  OAI222_X1 U12020 ( .A1(n13160), .A2(n9471), .B1(n13178), .B2(n9475), .C1(
        P2_U3088), .C2(n9653), .ZN(P2_U3324) );
  INV_X1 U12021 ( .A(SI_9_), .ZN(n9472) );
  OAI222_X1 U12022 ( .A1(n14154), .A2(n9473), .B1(n12417), .B2(n9472), .C1(
        n12020), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12023 ( .A1(n14047), .A2(n9476), .B1(n14043), .B2(n9475), .C1(
        P1_U3086), .C2(n13606), .ZN(P1_U3352) );
  INV_X1 U12024 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9478) );
  INV_X1 U12025 ( .A(n9477), .ZN(n9491) );
  OAI222_X1 U12026 ( .A1(n13160), .A2(n9478), .B1(n13178), .B2(n9491), .C1(
        P2_U3088), .C2(n14620), .ZN(P2_U3323) );
  INV_X1 U12027 ( .A(SI_10_), .ZN(n9479) );
  OAI222_X1 U12028 ( .A1(n14154), .A2(n9480), .B1(n12417), .B2(n9479), .C1(
        n12018), .C2(P3_U3151), .ZN(P3_U3285) );
  NAND2_X1 U12029 ( .A1(n9481), .A2(n9691), .ZN(n14537) );
  AND2_X1 U12030 ( .A1(n9486), .A2(n14044), .ZN(n9483) );
  INV_X1 U12031 ( .A(n9482), .ZN(n11201) );
  AOI22_X1 U12032 ( .A1(n14537), .A2(n9484), .B1(n9483), .B2(n11201), .ZN(
        P1_U3445) );
  AOI22_X1 U12033 ( .A1(n14537), .A2(n9487), .B1(n9486), .B2(n9485), .ZN(
        P1_U3446) );
  INV_X1 U12034 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9489) );
  INV_X1 U12035 ( .A(n9488), .ZN(n9493) );
  OAI222_X1 U12036 ( .A1(n13160), .A2(n9489), .B1(n13178), .B2(n9493), .C1(
        P2_U3088), .C2(n6905), .ZN(P2_U3322) );
  INV_X1 U12037 ( .A(n14047), .ZN(n14035) );
  AOI22_X1 U12038 ( .A1(n13626), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n14035), .ZN(n9490) );
  OAI21_X1 U12039 ( .B1(n9491), .B2(n14043), .A(n9490), .ZN(P1_U3351) );
  AOI22_X1 U12040 ( .A1(n9633), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n14035), .ZN(n9492) );
  OAI21_X1 U12041 ( .B1(n9493), .B2(n14043), .A(n9492), .ZN(P1_U3350) );
  INV_X1 U12042 ( .A(n9494), .ZN(n9498) );
  INV_X1 U12043 ( .A(n14635), .ZN(n9495) );
  OAI222_X1 U12044 ( .A1(n13160), .A2(n9496), .B1(n13178), .B2(n9498), .C1(
        P2_U3088), .C2(n9495), .ZN(P2_U3321) );
  INV_X1 U12045 ( .A(n9622), .ZN(n9497) );
  OAI222_X1 U12046 ( .A1(n14047), .A2(n9499), .B1(n14043), .B2(n9498), .C1(
        P1_U3086), .C2(n9497), .ZN(P1_U3349) );
  INV_X1 U12047 ( .A(n13596), .ZN(n9500) );
  OAI222_X1 U12048 ( .A1(n14047), .A2(n9502), .B1(n14043), .B2(n9501), .C1(
        P1_U3086), .C2(n9500), .ZN(P1_U3353) );
  INV_X1 U12049 ( .A(n9691), .ZN(n9686) );
  INV_X1 U12050 ( .A(n9504), .ZN(n9503) );
  NAND2_X1 U12051 ( .A1(n9503), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13546) );
  NAND2_X1 U12052 ( .A1(n9686), .A2(n13546), .ZN(n9510) );
  INV_X1 U12053 ( .A(n13480), .ZN(n9505) );
  NAND2_X1 U12054 ( .A1(n9505), .A2(n9504), .ZN(n9507) );
  NAND2_X1 U12055 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  INV_X1 U12056 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9515) );
  INV_X1 U12057 ( .A(n9508), .ZN(n9509) );
  NAND2_X1 U12058 ( .A1(n9510), .A2(n9509), .ZN(n9612) );
  INV_X1 U12059 ( .A(n9612), .ZN(n9609) );
  INV_X1 U12060 ( .A(n14041), .ZN(n13586) );
  NOR2_X1 U12061 ( .A1(n14041), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9511) );
  NOR2_X1 U12062 ( .A1(n8115), .A2(n9511), .ZN(n13593) );
  OAI21_X1 U12063 ( .B1(n13586), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13593), .ZN(
        n9512) );
  XNOR2_X1 U12064 ( .A(n9512), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9513) );
  AOI22_X1 U12065 ( .A1(n9609), .A2(n9513), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9514) );
  OAI21_X1 U12066 ( .B1(n14499), .B2(n9515), .A(n9514), .ZN(P1_U3243) );
  INV_X1 U12067 ( .A(n9516), .ZN(n9523) );
  AOI22_X1 U12068 ( .A1(n9672), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14035), .ZN(n9517) );
  OAI21_X1 U12069 ( .B1(n9523), .B2(n14043), .A(n9517), .ZN(P1_U3348) );
  INV_X1 U12070 ( .A(n9518), .ZN(n9519) );
  OAI222_X1 U12071 ( .A1(n14154), .A2(n9519), .B1(n12417), .B2(n15182), .C1(
        n14880), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12072 ( .A(n13577), .ZN(n9521) );
  OAI222_X1 U12073 ( .A1(n9521), .A2(P1_U3086), .B1(n14043), .B2(n9525), .C1(
        n9520), .C2(n14047), .ZN(P1_U3354) );
  INV_X1 U12074 ( .A(n9723), .ZN(n9522) );
  OAI222_X1 U12075 ( .A1(n13160), .A2(n9524), .B1(n13178), .B2(n9523), .C1(
        P2_U3088), .C2(n9522), .ZN(P2_U3320) );
  OAI222_X1 U12076 ( .A1(n13160), .A2(n9526), .B1(n13178), .B2(n9525), .C1(
        P2_U3088), .C2(n8859), .ZN(P2_U3326) );
  OAI222_X1 U12077 ( .A1(n14154), .A2(n9527), .B1(n12417), .B2(n15245), .C1(
        n14899), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12078 ( .A(n9528), .ZN(n9532) );
  INV_X1 U12079 ( .A(n9814), .ZN(n9529) );
  OAI222_X1 U12080 ( .A1(n14047), .A2(n9530), .B1(n14043), .B2(n9532), .C1(
        P1_U3086), .C2(n9529), .ZN(P1_U3347) );
  INV_X1 U12081 ( .A(n9797), .ZN(n9531) );
  OAI222_X1 U12082 ( .A1(n13160), .A2(n9533), .B1(n13178), .B2(n9532), .C1(
        P2_U3088), .C2(n9531), .ZN(P2_U3319) );
  INV_X1 U12083 ( .A(n14499), .ZN(n13639) );
  CLKBUF_X2 U12084 ( .A(P1_U4016), .Z(n13591) );
  NOR2_X1 U12085 ( .A1(n13639), .A2(n13591), .ZN(P1_U3085) );
  NAND2_X1 U12086 ( .A1(n9534), .A2(n11172), .ZN(n9535) );
  AND2_X1 U12087 ( .A1(n9536), .A2(n9535), .ZN(n9537) );
  OR2_X1 U12088 ( .A1(n9538), .A2(n9537), .ZN(n9546) );
  AND2_X1 U12089 ( .A1(n9546), .A2(n9539), .ZN(n14639) );
  MUX2_X1 U12090 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8887), .S(n9573), .Z(n9545)
         );
  INV_X1 U12091 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10029) );
  MUX2_X1 U12092 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10029), .S(n9550), .Z(
        n14607) );
  AND2_X1 U12093 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n14606) );
  NAND2_X1 U12094 ( .A1(n14607), .A2(n14606), .ZN(n14605) );
  NAND2_X1 U12095 ( .A1(n9550), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U12096 ( .A1(n14605), .A2(n9540), .ZN(n9544) );
  NAND2_X1 U12097 ( .A1(n9541), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13166) );
  INV_X1 U12098 ( .A(n13166), .ZN(n9542) );
  NAND2_X1 U12099 ( .A1(n9546), .A2(n9542), .ZN(n9552) );
  INV_X1 U12100 ( .A(n9552), .ZN(n9543) );
  NAND2_X1 U12101 ( .A1(n9545), .A2(n9544), .ZN(n9575) );
  OAI211_X1 U12102 ( .C1(n9545), .C2(n9544), .A(n14655), .B(n9575), .ZN(n9548)
         );
  INV_X1 U12103 ( .A(n14722), .ZN(n14601) );
  NAND2_X1 U12104 ( .A1(n14601), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n9547) );
  OAI211_X1 U12105 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10105), .A(n9548), .B(
        n9547), .ZN(n9549) );
  INV_X1 U12106 ( .A(n9549), .ZN(n9556) );
  MUX2_X1 U12107 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9564), .S(n9573), .Z(n9554)
         );
  MUX2_X1 U12108 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9551), .S(n9550), .Z(n14604) );
  AND2_X1 U12109 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14603) );
  NAND2_X1 U12110 ( .A1(n14604), .A2(n14603), .ZN(n14602) );
  OAI21_X1 U12111 ( .B1(n8859), .B2(n9551), .A(n14602), .ZN(n9553) );
  NAND2_X1 U12112 ( .A1(n9554), .A2(n9553), .ZN(n9562) );
  OAI211_X1 U12113 ( .C1(n9554), .C2(n9553), .A(n14715), .B(n9562), .ZN(n9555)
         );
  OAI211_X1 U12114 ( .C1(n14621), .C2(n9563), .A(n9556), .B(n9555), .ZN(
        P2_U3216) );
  INV_X1 U12115 ( .A(n9557), .ZN(n9560) );
  INV_X1 U12116 ( .A(n9932), .ZN(n9937) );
  OAI222_X1 U12117 ( .A1(n13160), .A2(n9558), .B1(n13178), .B2(n9560), .C1(
        P2_U3088), .C2(n9937), .ZN(P2_U3318) );
  INV_X1 U12118 ( .A(n9894), .ZN(n9559) );
  OAI222_X1 U12119 ( .A1(n14047), .A2(n9561), .B1(n14043), .B2(n9560), .C1(
        P1_U3086), .C2(n9559), .ZN(P1_U3346) );
  AND2_X1 U12120 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n9572) );
  INV_X1 U12121 ( .A(n14620), .ZN(n9567) );
  OAI21_X1 U12122 ( .B1(n9564), .B2(n9563), .A(n9562), .ZN(n9643) );
  MUX2_X1 U12123 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9565), .S(n9576), .Z(n9644)
         );
  NAND2_X1 U12124 ( .A1(n9643), .A2(n9644), .ZN(n9642) );
  OAI21_X1 U12125 ( .B1(n9565), .B2(n9653), .A(n9642), .ZN(n14613) );
  INV_X1 U12126 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U12127 ( .A(n9566), .B(P2_REG2_REG_4__SCAN_IN), .S(n14620), .Z(
        n14614) );
  MUX2_X1 U12128 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6904), .S(n9590), .Z(n9568)
         );
  INV_X1 U12129 ( .A(n9568), .ZN(n9569) );
  AOI211_X1 U12130 ( .C1(n9570), .C2(n9569), .A(n9585), .B(n14695), .ZN(n9571)
         );
  AOI211_X1 U12131 ( .C1(n14601), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9572), .B(
        n9571), .ZN(n9583) );
  INV_X1 U12132 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14833) );
  MUX2_X1 U12133 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n14833), .S(n9590), .Z(n9581) );
  NAND2_X1 U12134 ( .A1(n9573), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U12135 ( .A1(n9575), .A2(n9574), .ZN(n9649) );
  MUX2_X1 U12136 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8903), .S(n9576), .Z(n9650)
         );
  NAND2_X1 U12137 ( .A1(n9649), .A2(n9650), .ZN(n9648) );
  NAND2_X1 U12138 ( .A1(n9576), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12139 ( .A1(n9648), .A2(n9577), .ZN(n14616) );
  MUX2_X1 U12140 ( .A(n9578), .B(P2_REG1_REG_4__SCAN_IN), .S(n14620), .Z(
        n14617) );
  NAND2_X1 U12141 ( .A1(n14616), .A2(n14617), .ZN(n14615) );
  OR2_X1 U12142 ( .A1(n14620), .A2(n9578), .ZN(n9579) );
  NAND2_X1 U12143 ( .A1(n14615), .A2(n9579), .ZN(n9580) );
  NAND2_X1 U12144 ( .A1(n9580), .A2(n9581), .ZN(n9592) );
  OAI211_X1 U12145 ( .C1(n9581), .C2(n9580), .A(n14655), .B(n9592), .ZN(n9582)
         );
  OAI211_X1 U12146 ( .C1(n14621), .C2(n6905), .A(n9583), .B(n9582), .ZN(
        P2_U3219) );
  INV_X1 U12147 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U12148 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n9584) );
  OAI21_X1 U12149 ( .B1(n14722), .B2(n14124), .A(n9584), .ZN(n9589) );
  XNOR2_X1 U12150 ( .A(n14635), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n14631) );
  NOR2_X1 U12151 ( .A1(n14632), .A2(n14631), .ZN(n14630) );
  AOI21_X1 U12152 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n14635), .A(n14630), .ZN(
        n9587) );
  XNOR2_X1 U12153 ( .A(n9723), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9586) );
  NOR2_X1 U12154 ( .A1(n9587), .A2(n9586), .ZN(n9718) );
  AOI211_X1 U12155 ( .C1(n9587), .C2(n9586), .A(n14695), .B(n9718), .ZN(n9588)
         );
  AOI211_X1 U12156 ( .C1(n14719), .C2(n9723), .A(n9589), .B(n9588), .ZN(n9597)
         );
  MUX2_X1 U12157 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8968), .S(n9723), .Z(n9595)
         );
  NAND2_X1 U12158 ( .A1(n9590), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U12159 ( .A1(n9592), .A2(n9591), .ZN(n14627) );
  MUX2_X1 U12160 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n8950), .S(n14635), .Z(
        n14628) );
  NAND2_X1 U12161 ( .A1(n14627), .A2(n14628), .ZN(n14626) );
  NAND2_X1 U12162 ( .A1(n14635), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U12163 ( .A1(n14626), .A2(n9593), .ZN(n9594) );
  NAND2_X1 U12164 ( .A1(n9594), .A2(n9595), .ZN(n9725) );
  OAI211_X1 U12165 ( .C1(n9595), .C2(n9594), .A(n14655), .B(n9725), .ZN(n9596)
         );
  NAND2_X1 U12166 ( .A1(n9597), .A2(n9596), .ZN(P2_U3221) );
  INV_X1 U12167 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10479) );
  MUX2_X1 U12168 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10479), .S(n13596), .Z(
        n13599) );
  INV_X1 U12169 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10468) );
  MUX2_X1 U12170 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10468), .S(n13577), .Z(
        n13582) );
  AND2_X1 U12171 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13587) );
  NAND2_X1 U12172 ( .A1(n13582), .A2(n13587), .ZN(n13581) );
  NAND2_X1 U12173 ( .A1(n13577), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9598) );
  NAND2_X1 U12174 ( .A1(n13581), .A2(n9598), .ZN(n13598) );
  NAND2_X1 U12175 ( .A1(n13599), .A2(n13598), .ZN(n13597) );
  NAND2_X1 U12176 ( .A1(n13596), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U12177 ( .A1(n13597), .A2(n9599), .ZN(n13611) );
  MUX2_X1 U12178 ( .A(n14509), .B(P1_REG2_REG_3__SCAN_IN), .S(n13606), .Z(
        n13612) );
  NAND2_X1 U12179 ( .A1(n13611), .A2(n13612), .ZN(n13610) );
  OR2_X1 U12180 ( .A1(n13606), .A2(n14509), .ZN(n9600) );
  NAND2_X1 U12181 ( .A1(n13610), .A2(n9600), .ZN(n13627) );
  MUX2_X1 U12182 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7630), .S(n13626), .Z(
        n13628) );
  XNOR2_X1 U12183 ( .A(n9633), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9636) );
  XNOR2_X1 U12184 ( .A(n9622), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U12185 ( .A1(n13589), .A2(n13586), .ZN(n9601) );
  NOR2_X1 U12186 ( .A1(n6627), .A2(n9602), .ZN(n9617) );
  AOI211_X1 U12187 ( .C1(n6627), .C2(n9602), .A(n14488), .B(n9617), .ZN(n9616)
         );
  INV_X1 U12188 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9603) );
  MUX2_X1 U12189 ( .A(n9603), .B(P1_REG1_REG_6__SCAN_IN), .S(n9622), .Z(n9611)
         );
  MUX2_X1 U12190 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7598), .S(n13596), .Z(
        n13602) );
  MUX2_X1 U12191 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7586), .S(n13577), .Z(
        n13580) );
  AND2_X1 U12192 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13579) );
  NAND2_X1 U12193 ( .A1(n13580), .A2(n13579), .ZN(n13578) );
  NAND2_X1 U12194 ( .A1(n13577), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U12195 ( .A1(n13578), .A2(n9604), .ZN(n13601) );
  NAND2_X1 U12196 ( .A1(n13602), .A2(n13601), .ZN(n13600) );
  NAND2_X1 U12197 ( .A1(n13596), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U12198 ( .A1(n13600), .A2(n9605), .ZN(n13614) );
  MUX2_X1 U12199 ( .A(n9606), .B(P1_REG1_REG_3__SCAN_IN), .S(n13606), .Z(
        n13615) );
  NAND2_X1 U12200 ( .A1(n13614), .A2(n13615), .ZN(n13613) );
  INV_X1 U12201 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9606) );
  OR2_X1 U12202 ( .A1(n13606), .A2(n9606), .ZN(n9607) );
  NAND2_X1 U12203 ( .A1(n13613), .A2(n9607), .ZN(n13622) );
  MUX2_X1 U12204 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7635), .S(n13626), .Z(
        n13621) );
  AND2_X1 U12205 ( .A1(n13622), .A2(n13621), .ZN(n13624) );
  XNOR2_X1 U12206 ( .A(n9633), .B(n9608), .ZN(n9632) );
  OAI21_X1 U12207 ( .B1(n9633), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9630), .ZN(
        n9610) );
  NOR2_X1 U12208 ( .A1(n9610), .A2(n9611), .ZN(n9621) );
  INV_X1 U12209 ( .A(n14483), .ZN(n14452) );
  AOI211_X1 U12210 ( .C1(n9611), .C2(n9610), .A(n9621), .B(n14452), .ZN(n9615)
         );
  INV_X1 U12211 ( .A(n14475), .ZN(n14493) );
  NAND2_X1 U12212 ( .A1(n14493), .A2(n9622), .ZN(n9613) );
  NAND2_X1 U12213 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10449) );
  OAI211_X1 U12214 ( .C1(n14116), .C2(n14499), .A(n9613), .B(n10449), .ZN(
        n9614) );
  OR3_X1 U12215 ( .A1(n9616), .A2(n9615), .A3(n9614), .ZN(P1_U3249) );
  AOI21_X1 U12216 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9622), .A(n9617), .ZN(
        n9620) );
  INV_X1 U12217 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9618) );
  MUX2_X1 U12218 ( .A(n9618), .B(P1_REG2_REG_7__SCAN_IN), .S(n9672), .Z(n9619)
         );
  AOI211_X1 U12219 ( .C1(n9620), .C2(n9619), .A(n14488), .B(n9671), .ZN(n9629)
         );
  INV_X1 U12220 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9623) );
  MUX2_X1 U12221 ( .A(n9623), .B(P1_REG1_REG_7__SCAN_IN), .S(n9672), .Z(n9624)
         );
  NOR2_X1 U12222 ( .A1(n9625), .A2(n9624), .ZN(n9666) );
  AOI211_X1 U12223 ( .C1(n9625), .C2(n9624), .A(n14452), .B(n9666), .ZN(n9628)
         );
  NAND2_X1 U12224 ( .A1(n14493), .A2(n9672), .ZN(n9626) );
  NAND2_X1 U12225 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10210) );
  OAI211_X1 U12226 ( .C1(n14122), .C2(n14499), .A(n9626), .B(n10210), .ZN(
        n9627) );
  OR3_X1 U12227 ( .A1(n9629), .A2(n9628), .A3(n9627), .ZN(P1_U3250) );
  OAI21_X1 U12228 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9640) );
  INV_X1 U12229 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15321) );
  NAND2_X1 U12230 ( .A1(n14493), .A2(n9633), .ZN(n9634) );
  NAND2_X1 U12231 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9965) );
  OAI211_X1 U12232 ( .C1(n15321), .C2(n14499), .A(n9634), .B(n9965), .ZN(n9639) );
  AOI211_X1 U12233 ( .C1(n9637), .C2(n9636), .A(n9635), .B(n14488), .ZN(n9638)
         );
  AOI211_X1 U12234 ( .C1(n14483), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9641)
         );
  INV_X1 U12235 ( .A(n9641), .ZN(P1_U3248) );
  INV_X1 U12236 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15398) );
  OAI211_X1 U12237 ( .C1(n9644), .C2(n9643), .A(n14715), .B(n9642), .ZN(n9646)
         );
  NAND2_X1 U12238 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n9645) );
  OAI211_X1 U12239 ( .C1(n15398), .C2(n14722), .A(n9646), .B(n9645), .ZN(n9647) );
  INV_X1 U12240 ( .A(n9647), .ZN(n9652) );
  OAI211_X1 U12241 ( .C1(n9650), .C2(n9649), .A(n14655), .B(n9648), .ZN(n9651)
         );
  OAI211_X1 U12242 ( .C1(n14621), .C2(n9653), .A(n9652), .B(n9651), .ZN(
        P2_U3217) );
  INV_X1 U12243 ( .A(n9654), .ZN(n9657) );
  INV_X1 U12244 ( .A(n10929), .ZN(n9944) );
  OAI222_X1 U12245 ( .A1(n13160), .A2(n9655), .B1(n13178), .B2(n9657), .C1(
        P2_U3088), .C2(n9944), .ZN(P2_U3317) );
  INV_X1 U12246 ( .A(n10067), .ZN(n9656) );
  OAI222_X1 U12247 ( .A1(n14047), .A2(n9658), .B1(n14043), .B2(n9657), .C1(
        P1_U3086), .C2(n9656), .ZN(P1_U3345) );
  AOI22_X1 U12248 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14715), .B1(n14655), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12249 ( .A1(n14655), .A2(n9659), .ZN(n9660) );
  OAI211_X1 U12250 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14695), .A(n14621), .B(
        n9660), .ZN(n9661) );
  INV_X1 U12251 ( .A(n9661), .ZN(n9662) );
  MUX2_X1 U12252 ( .A(n9663), .B(n9662), .S(P2_IR_REG_0__SCAN_IN), .Z(n9665)
         );
  AOI22_X1 U12253 ( .A1(n14601), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9664) );
  NAND2_X1 U12254 ( .A1(n9665), .A2(n9664), .ZN(P2_U3214) );
  AOI21_X1 U12255 ( .B1(n9672), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9666), .ZN(
        n9669) );
  MUX2_X1 U12256 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9667), .S(n9814), .Z(n9668)
         );
  NAND2_X1 U12257 ( .A1(n9669), .A2(n9668), .ZN(n9808) );
  OAI21_X1 U12258 ( .B1(n9669), .B2(n9668), .A(n9808), .ZN(n9678) );
  NAND2_X1 U12259 ( .A1(n14493), .A2(n9814), .ZN(n9670) );
  NAND2_X1 U12260 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10787) );
  OAI211_X1 U12261 ( .C1(n15151), .C2(n14499), .A(n9670), .B(n10787), .ZN(
        n9677) );
  INV_X1 U12262 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9673) );
  MUX2_X1 U12263 ( .A(n9673), .B(P1_REG2_REG_8__SCAN_IN), .S(n9814), .Z(n9674)
         );
  AOI211_X1 U12264 ( .C1(n9675), .C2(n9674), .A(n14488), .B(n9813), .ZN(n9676)
         );
  AOI211_X1 U12265 ( .C1(n14483), .C2(n9678), .A(n9677), .B(n9676), .ZN(n9679)
         );
  INV_X1 U12266 ( .A(n9679), .ZN(P1_U3251) );
  INV_X4 U12267 ( .A(n11564), .ZN(n11554) );
  INV_X1 U12268 ( .A(n9680), .ZN(n9681) );
  OAI21_X1 U12269 ( .B1(n10462), .B2(n11563), .A(n9682), .ZN(n9707) );
  INV_X1 U12270 ( .A(n9958), .ZN(n9685) );
  OAI22_X1 U12271 ( .A1(n11563), .A2(n14526), .B1(n9680), .B2(n9683), .ZN(
        n9684) );
  XOR2_X1 U12272 ( .A(n9707), .B(n9706), .Z(n13588) );
  NAND3_X1 U12273 ( .A1(n10079), .A2(n10078), .A3(n10076), .ZN(n9688) );
  OR2_X1 U12274 ( .A1(n9688), .A2(n9686), .ZN(n9692) );
  NAND2_X1 U12275 ( .A1(n14582), .A2(n13480), .ZN(n9687) );
  NOR2_X1 U12276 ( .A1(n9750), .A2(n13686), .ZN(n9984) );
  NAND2_X1 U12277 ( .A1(n9688), .A2(n9689), .ZN(n9869) );
  NAND2_X1 U12278 ( .A1(n9869), .A2(n10077), .ZN(n9753) );
  AOI22_X1 U12279 ( .A1(n14353), .A2(n9984), .B1(n9753), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U12280 ( .A1(n9693), .A2(n9986), .ZN(n9694) );
  OAI211_X1 U12281 ( .C1(n13588), .C2(n13286), .A(n9695), .B(n9694), .ZN(
        P1_U3232) );
  INV_X1 U12282 ( .A(n9696), .ZN(n9700) );
  INV_X1 U12283 ( .A(n12812), .ZN(n9697) );
  OAI222_X1 U12284 ( .A1(n13160), .A2(n9698), .B1(n13178), .B2(n9700), .C1(
        P2_U3088), .C2(n9697), .ZN(P2_U3316) );
  INV_X1 U12285 ( .A(n13642), .ZN(n9699) );
  OAI222_X1 U12286 ( .A1(n14047), .A2(n9701), .B1(n14043), .B2(n9700), .C1(
        P1_U3086), .C2(n9699), .ZN(P1_U3344) );
  INV_X1 U12287 ( .A(n9693), .ZN(n14362) );
  NAND2_X1 U12288 ( .A1(n14353), .A2(n13864), .ZN(n13274) );
  INV_X1 U12289 ( .A(n13274), .ZN(n9704) );
  INV_X1 U12290 ( .A(n9753), .ZN(n9702) );
  OR2_X1 U12291 ( .A1(n7611), .A2(n13686), .ZN(n10466) );
  OAI22_X1 U12292 ( .A1(n9702), .A2(n13575), .B1(n14360), .B2(n10466), .ZN(
        n9703) );
  AOI21_X1 U12293 ( .B1(n9704), .B2(n13574), .A(n9703), .ZN(n9715) );
  OAI22_X1 U12294 ( .A1(n9750), .A2(n11563), .B1(n14543), .B2(n11564), .ZN(
        n9705) );
  OAI22_X1 U12295 ( .A1(n9958), .A2(n9750), .B1(n14543), .B2(n11563), .ZN(
        n9742) );
  XNOR2_X1 U12296 ( .A(n9744), .B(n9742), .ZN(n9712) );
  NAND2_X1 U12297 ( .A1(n9706), .A2(n9707), .ZN(n9710) );
  INV_X1 U12298 ( .A(n9707), .ZN(n9708) );
  NAND2_X1 U12299 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  OAI21_X1 U12300 ( .B1(n9712), .B2(n9711), .A(n9746), .ZN(n9713) );
  NAND2_X1 U12301 ( .A1(n9713), .A2(n14365), .ZN(n9714) );
  OAI211_X1 U12302 ( .C1(n14543), .C2(n14362), .A(n9715), .B(n9714), .ZN(
        P1_U3222) );
  INV_X1 U12303 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12304 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n9716) );
  OAI21_X1 U12305 ( .B1(n14722), .B2(n9717), .A(n9716), .ZN(n9722) );
  INV_X1 U12306 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10613) );
  MUX2_X1 U12307 ( .A(n10613), .B(P2_REG2_REG_8__SCAN_IN), .S(n9797), .Z(n9719) );
  AOI211_X1 U12308 ( .C1(n9720), .C2(n9719), .A(n14695), .B(n9796), .ZN(n9721)
         );
  AOI211_X1 U12309 ( .C1(n14719), .C2(n9797), .A(n9722), .B(n9721), .ZN(n9729)
         );
  MUX2_X1 U12310 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n8989), .S(n9797), .Z(n9727)
         );
  NAND2_X1 U12311 ( .A1(n9723), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12312 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  NAND2_X1 U12313 ( .A1(n9726), .A2(n9727), .ZN(n9792) );
  OAI211_X1 U12314 ( .C1(n9727), .C2(n9726), .A(n14655), .B(n9792), .ZN(n9728)
         );
  NAND2_X1 U12315 ( .A1(n9729), .A2(n9728), .ZN(P2_U3222) );
  INV_X1 U12316 ( .A(n14822), .ZN(n14802) );
  AND2_X1 U12317 ( .A1(n12515), .A2(n12520), .ZN(n12729) );
  INV_X1 U12318 ( .A(n12729), .ZN(n9852) );
  NOR2_X1 U12319 ( .A1(n10025), .A2(n9730), .ZN(n9841) );
  INV_X1 U12320 ( .A(n9731), .ZN(n9734) );
  INV_X1 U12321 ( .A(n12767), .ZN(n10969) );
  OR2_X1 U12322 ( .A1(n6559), .A2(n10969), .ZN(n9733) );
  INV_X1 U12323 ( .A(n12778), .ZN(n12674) );
  OR2_X1 U12324 ( .A1(n12762), .A2(n12674), .ZN(n9732) );
  NOR2_X1 U12325 ( .A1(n9734), .A2(n13026), .ZN(n9735) );
  OR2_X1 U12326 ( .A1(n12513), .A2(n13006), .ZN(n9906) );
  OAI21_X1 U12327 ( .B1(n12729), .B2(n9735), .A(n9906), .ZN(n9840) );
  AOI211_X1 U12328 ( .C1(n14802), .C2(n9852), .A(n9841), .B(n9840), .ZN(n14755) );
  AND2_X1 U12329 ( .A1(n14751), .A2(n9736), .ZN(n14752) );
  AND3_X1 U12330 ( .A1(n9844), .A2(n9737), .A3(n9843), .ZN(n9738) );
  INV_X1 U12331 ( .A(n14842), .ZN(n14840) );
  NAND2_X1 U12332 ( .A1(n14840), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9740) );
  OAI21_X1 U12333 ( .B1(n14755), .B2(n14840), .A(n9740), .ZN(P2_U3499) );
  OAI22_X1 U12334 ( .A1(n7611), .A2(n11563), .B1(n10480), .B2(n11564), .ZN(
        n9741) );
  XNOR2_X1 U12335 ( .A(n9741), .B(n11476), .ZN(n9879) );
  OAI22_X1 U12336 ( .A1(n9958), .A2(n7611), .B1(n10480), .B2(n11563), .ZN(
        n9878) );
  XNOR2_X1 U12337 ( .A(n9879), .B(n9878), .ZN(n9748) );
  INV_X1 U12338 ( .A(n9742), .ZN(n9743) );
  NAND2_X1 U12339 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  NAND2_X1 U12340 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  OAI21_X1 U12341 ( .B1(n9748), .B2(n9747), .A(n9881), .ZN(n9749) );
  NAND2_X1 U12342 ( .A1(n9749), .A2(n14365), .ZN(n9755) );
  NOR2_X1 U12343 ( .A1(n9750), .A2(n13542), .ZN(n9752) );
  NOR2_X1 U12344 ( .A1(n9877), .A2(n13686), .ZN(n9751) );
  OR2_X1 U12345 ( .A1(n9752), .A2(n9751), .ZN(n10474) );
  AOI22_X1 U12346 ( .A1(n14353), .A2(n10474), .B1(n9753), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9754) );
  OAI211_X1 U12347 ( .C1(n10480), .C2(n14362), .A(n9755), .B(n9754), .ZN(
        P1_U3237) );
  INV_X1 U12348 ( .A(n8723), .ZN(n9757) );
  CLKBUF_X1 U12349 ( .A(n9759), .Z(n9775) );
  INV_X1 U12350 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15228) );
  NOR2_X1 U12351 ( .A1(n9775), .A2(n15228), .ZN(P3_U3254) );
  INV_X1 U12352 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9758) );
  NOR2_X1 U12353 ( .A1(n9775), .A2(n9758), .ZN(P3_U3263) );
  INV_X1 U12354 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9760) );
  NOR2_X1 U12355 ( .A1(n9775), .A2(n9760), .ZN(P3_U3262) );
  INV_X1 U12356 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9761) );
  NOR2_X1 U12357 ( .A1(n9759), .A2(n9761), .ZN(P3_U3260) );
  INV_X1 U12358 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9762) );
  NOR2_X1 U12359 ( .A1(n9775), .A2(n9762), .ZN(P3_U3259) );
  INV_X1 U12360 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9763) );
  NOR2_X1 U12361 ( .A1(n9759), .A2(n9763), .ZN(P3_U3258) );
  INV_X1 U12362 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9764) );
  NOR2_X1 U12363 ( .A1(n9775), .A2(n9764), .ZN(P3_U3257) );
  INV_X1 U12364 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9765) );
  NOR2_X1 U12365 ( .A1(n9775), .A2(n9765), .ZN(P3_U3256) );
  INV_X1 U12366 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9766) );
  NOR2_X1 U12367 ( .A1(n9775), .A2(n9766), .ZN(P3_U3255) );
  INV_X1 U12368 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9767) );
  NOR2_X1 U12369 ( .A1(n9775), .A2(n9767), .ZN(P3_U3261) );
  INV_X1 U12370 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9768) );
  NOR2_X1 U12371 ( .A1(n9775), .A2(n9768), .ZN(P3_U3253) );
  INV_X1 U12372 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9769) );
  NOR2_X1 U12373 ( .A1(n9759), .A2(n9769), .ZN(P3_U3237) );
  NOR2_X1 U12374 ( .A1(n9775), .A2(n15178), .ZN(P3_U3252) );
  NOR2_X1 U12375 ( .A1(n9775), .A2(n15303), .ZN(P3_U3251) );
  INV_X1 U12376 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9770) );
  NOR2_X1 U12377 ( .A1(n9775), .A2(n9770), .ZN(P3_U3250) );
  INV_X1 U12378 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9771) );
  NOR2_X1 U12379 ( .A1(n9775), .A2(n9771), .ZN(P3_U3249) );
  INV_X1 U12380 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9772) );
  NOR2_X1 U12381 ( .A1(n9775), .A2(n9772), .ZN(P3_U3248) );
  INV_X1 U12382 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9773) );
  NOR2_X1 U12383 ( .A1(n9775), .A2(n9773), .ZN(P3_U3247) );
  INV_X1 U12384 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9774) );
  NOR2_X1 U12385 ( .A1(n9775), .A2(n9774), .ZN(P3_U3246) );
  INV_X1 U12386 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9776) );
  NOR2_X1 U12387 ( .A1(n9759), .A2(n9776), .ZN(P3_U3245) );
  NOR2_X1 U12388 ( .A1(n9759), .A2(n15219), .ZN(P3_U3244) );
  INV_X1 U12389 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U12390 ( .A1(n9759), .A2(n9777), .ZN(P3_U3243) );
  INV_X1 U12391 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9778) );
  NOR2_X1 U12392 ( .A1(n9759), .A2(n9778), .ZN(P3_U3242) );
  INV_X1 U12393 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9779) );
  NOR2_X1 U12394 ( .A1(n9759), .A2(n9779), .ZN(P3_U3241) );
  NOR2_X1 U12395 ( .A1(n9759), .A2(n15336), .ZN(P3_U3238) );
  INV_X1 U12396 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9780) );
  NOR2_X1 U12397 ( .A1(n9759), .A2(n9780), .ZN(P3_U3235) );
  INV_X1 U12398 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n15243) );
  NOR2_X1 U12399 ( .A1(n9759), .A2(n15243), .ZN(P3_U3240) );
  INV_X1 U12400 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15225) );
  NOR2_X1 U12401 ( .A1(n9775), .A2(n15225), .ZN(P3_U3234) );
  INV_X1 U12402 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9781) );
  NOR2_X1 U12403 ( .A1(n9775), .A2(n9781), .ZN(P3_U3239) );
  INV_X1 U12404 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9782) );
  NOR2_X1 U12405 ( .A1(n9775), .A2(n9782), .ZN(P3_U3236) );
  INV_X1 U12406 ( .A(n9783), .ZN(n9785) );
  OAI222_X1 U12407 ( .A1(n14938), .A2(P3_U3151), .B1(n14154), .B2(n9785), .C1(
        n9784), .C2(n12417), .ZN(P3_U3281) );
  INV_X1 U12408 ( .A(n9786), .ZN(n9789) );
  INV_X1 U12409 ( .A(n13666), .ZN(n9787) );
  OAI222_X1 U12410 ( .A1(n14047), .A2(n9788), .B1(n14043), .B2(n9789), .C1(
        n9787), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12411 ( .A(n10933), .ZN(n14640) );
  OAI222_X1 U12412 ( .A1(n13160), .A2(n9790), .B1(n14640), .B2(P2_U3088), .C1(
        n13178), .C2(n9789), .ZN(P2_U3315) );
  MUX2_X1 U12413 ( .A(n9936), .B(P2_REG1_REG_9__SCAN_IN), .S(n9932), .Z(n9795)
         );
  NAND2_X1 U12414 ( .A1(n9797), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U12415 ( .A1(n9792), .A2(n9791), .ZN(n9794) );
  OR2_X1 U12416 ( .A1(n9794), .A2(n9795), .ZN(n9939) );
  INV_X1 U12417 ( .A(n9939), .ZN(n9793) );
  AOI21_X1 U12418 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n9806) );
  INV_X1 U12419 ( .A(n14655), .ZN(n14707) );
  INV_X1 U12420 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9798) );
  MUX2_X1 U12421 ( .A(n9798), .B(P2_REG2_REG_9__SCAN_IN), .S(n9932), .Z(n9799)
         );
  INV_X1 U12422 ( .A(n9799), .ZN(n9800) );
  OAI21_X1 U12423 ( .B1(n9801), .B2(n9800), .A(n9931), .ZN(n9804) );
  NAND2_X1 U12424 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U12425 ( .A1(n14601), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9802) );
  OAI211_X1 U12426 ( .C1(n14621), .C2(n9937), .A(n10379), .B(n9802), .ZN(n9803) );
  AOI21_X1 U12427 ( .B1(n9804), .B2(n14715), .A(n9803), .ZN(n9805) );
  OAI21_X1 U12428 ( .B1(n9806), .B2(n14707), .A(n9805), .ZN(P2_U3223) );
  MUX2_X1 U12429 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9807), .S(n9894), .Z(n9810)
         );
  OAI21_X1 U12430 ( .B1(n9814), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9808), .ZN(
        n9809) );
  NAND2_X1 U12431 ( .A1(n9809), .A2(n9810), .ZN(n9893) );
  OAI21_X1 U12432 ( .B1(n9810), .B2(n9809), .A(n9893), .ZN(n9821) );
  INV_X1 U12433 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9812) );
  NAND2_X1 U12434 ( .A1(n14493), .A2(n9894), .ZN(n9811) );
  NAND2_X1 U12435 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11041) );
  OAI211_X1 U12436 ( .C1(n9812), .C2(n14499), .A(n9811), .B(n11041), .ZN(n9820) );
  INV_X1 U12437 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U12438 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9815), .S(n9894), .Z(n9816)
         );
  INV_X1 U12439 ( .A(n9816), .ZN(n9817) );
  NOR2_X1 U12440 ( .A1(n9818), .A2(n9817), .ZN(n9889) );
  AOI211_X1 U12441 ( .C1(n9818), .C2(n9817), .A(n14488), .B(n9889), .ZN(n9819)
         );
  AOI211_X1 U12442 ( .C1(n14483), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9822)
         );
  INV_X1 U12443 ( .A(n9822), .ZN(P1_U3252) );
  INV_X1 U12444 ( .A(n9823), .ZN(n9825) );
  OAI222_X1 U12445 ( .A1(n12039), .A2(P3_U3151), .B1(n14154), .B2(n9825), .C1(
        n9824), .C2(n12417), .ZN(P3_U3280) );
  INV_X1 U12446 ( .A(n9826), .ZN(n9829) );
  INV_X1 U12447 ( .A(n14425), .ZN(n9827) );
  OAI222_X1 U12448 ( .A1(n14047), .A2(n9828), .B1(n14043), .B2(n9829), .C1(
        n9827), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12449 ( .A(n14665), .ZN(n9830) );
  OAI222_X1 U12450 ( .A1(n13160), .A2(n9831), .B1(n9830), .B2(P2_U3088), .C1(
        n13178), .C2(n9829), .ZN(P2_U3314) );
  OAI211_X1 U12451 ( .C1(n9833), .C2(n9832), .A(n10002), .B(n9282), .ZN(n9839)
         );
  INV_X1 U12452 ( .A(n12511), .ZN(n14763) );
  NOR2_X1 U12453 ( .A1(n12438), .A2(n13006), .ZN(n14308) );
  NAND2_X1 U12454 ( .A1(n14308), .A2(n12800), .ZN(n9835) );
  NOR2_X1 U12455 ( .A1(n12438), .A2(n13004), .ZN(n14306) );
  NAND2_X1 U12456 ( .A1(n14306), .A2(n12802), .ZN(n9834) );
  OAI211_X1 U12457 ( .C1(n14763), .C2(n14310), .A(n9835), .B(n9834), .ZN(n9837) );
  INV_X1 U12458 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U12459 ( .A1(n14331), .A2(n10535), .B1(P2_STATE_REG_SCAN_IN), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n9836) );
  NOR2_X1 U12460 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  NAND2_X1 U12461 ( .A1(n9839), .A2(n9838), .ZN(P2_U3190) );
  AOI21_X1 U12462 ( .B1(n9841), .B2(n12725), .A(n9840), .ZN(n9855) );
  NAND2_X1 U12463 ( .A1(n9842), .A2(n14750), .ZN(n9846) );
  NAND3_X1 U12464 ( .A1(n14751), .A2(n9844), .A3(n9843), .ZN(n9845) );
  OR2_X1 U12465 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  OR2_X1 U12466 ( .A1(n12725), .A2(n10969), .ZN(n10424) );
  INV_X1 U12467 ( .A(n10424), .ZN(n9848) );
  NAND2_X1 U12468 ( .A1(n12979), .A2(n9848), .ZN(n13020) );
  INV_X1 U12469 ( .A(n13020), .ZN(n9853) );
  OAI22_X1 U12470 ( .A1(n12979), .A2(n9850), .B1(n9849), .B2(n13041), .ZN(
        n9851) );
  AOI21_X1 U12471 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9854) );
  OAI21_X1 U12472 ( .B1(n9855), .B2(n13051), .A(n9854), .ZN(P2_U3265) );
  NAND2_X1 U12473 ( .A1(n9282), .A2(n9183), .ZN(n12502) );
  INV_X1 U12474 ( .A(n9856), .ZN(n9857) );
  OAI22_X1 U12475 ( .A1(n12502), .A2(n10014), .B1(n14302), .B2(n9857), .ZN(
        n9862) );
  NOR2_X1 U12476 ( .A1(n9858), .A2(P2_U3088), .ZN(n9976) );
  AOI22_X1 U12477 ( .A1(n14308), .A2(n12802), .B1(n6560), .B2(n14328), .ZN(
        n9860) );
  NAND2_X1 U12478 ( .A1(n14306), .A2(n12805), .ZN(n9859) );
  OAI211_X1 U12479 ( .C1(n9976), .C2(n10052), .A(n9860), .B(n9859), .ZN(n9861)
         );
  AOI21_X1 U12480 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9864) );
  OAI21_X1 U12481 ( .B1(n14302), .B2(n9979), .A(n9864), .ZN(P2_U3194) );
  INV_X1 U12482 ( .A(n9865), .ZN(n9867) );
  OAI222_X1 U12483 ( .A1(n14154), .A2(n9867), .B1(n12417), .B2(n9866), .C1(
        n14229), .C2(P3_U3151), .ZN(P3_U3278) );
  NAND3_X1 U12484 ( .A1(n9869), .A2(n9680), .A3(n9868), .ZN(n9870) );
  NAND2_X1 U12485 ( .A1(n9870), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9871) );
  NAND2_X1 U12486 ( .A1(n13573), .A2(n13864), .ZN(n9873) );
  NAND2_X1 U12487 ( .A1(n13571), .A2(n13262), .ZN(n9872) );
  AND2_X1 U12488 ( .A1(n9873), .A2(n9872), .ZN(n14504) );
  NAND2_X1 U12489 ( .A1(n9693), .A2(n14511), .ZN(n9874) );
  NAND2_X1 U12490 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13607) );
  OAI211_X1 U12491 ( .C1(n14504), .C2(n14360), .A(n9874), .B(n13607), .ZN(
        n9887) );
  NAND2_X1 U12492 ( .A1(n11554), .A2(n14511), .ZN(n9875) );
  OAI21_X1 U12493 ( .B1(n9877), .B2(n11563), .A(n9875), .ZN(n9876) );
  XNOR2_X1 U12494 ( .A(n9876), .B(n9952), .ZN(n9955) );
  OAI22_X1 U12495 ( .A1(n9958), .A2(n9877), .B1(n14559), .B2(n11563), .ZN(
        n9954) );
  XNOR2_X1 U12496 ( .A(n9955), .B(n9954), .ZN(n9885) );
  INV_X1 U12497 ( .A(n9957), .ZN(n9883) );
  AOI211_X1 U12498 ( .C1(n9885), .C2(n9884), .A(n13286), .B(n9883), .ZN(n9886)
         );
  AOI211_X1 U12499 ( .C1(n7632), .C2(n13293), .A(n9887), .B(n9886), .ZN(n9888)
         );
  INV_X1 U12500 ( .A(n9888), .ZN(P1_U3218) );
  MUX2_X1 U12501 ( .A(n15337), .B(P1_REG2_REG_10__SCAN_IN), .S(n10067), .Z(
        n9890) );
  AOI211_X1 U12502 ( .C1(n9891), .C2(n9890), .A(n14488), .B(n10066), .ZN(n9900) );
  INV_X1 U12503 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9892) );
  MUX2_X1 U12504 ( .A(n9892), .B(P1_REG1_REG_10__SCAN_IN), .S(n10067), .Z(
        n9896) );
  OAI21_X1 U12505 ( .B1(n9894), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9893), .ZN(
        n9895) );
  NOR2_X1 U12506 ( .A1(n9895), .A2(n9896), .ZN(n10060) );
  AOI211_X1 U12507 ( .C1(n9896), .C2(n9895), .A(n14452), .B(n10060), .ZN(n9899) );
  INV_X1 U12508 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14073) );
  NAND2_X1 U12509 ( .A1(n14493), .A2(n10067), .ZN(n9897) );
  NAND2_X1 U12510 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10958)
         );
  OAI211_X1 U12511 ( .C1(n14073), .C2(n14499), .A(n9897), .B(n10958), .ZN(
        n9898) );
  OR3_X1 U12512 ( .A1(n9900), .A2(n9899), .A3(n9898), .ZN(P1_U3253) );
  INV_X1 U12513 ( .A(n9976), .ZN(n9903) );
  OAI21_X1 U12514 ( .B1(n9901), .B2(n14302), .A(n14310), .ZN(n9902) );
  AOI22_X1 U12515 ( .A1(n9903), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n10024), .B2(
        n9902), .ZN(n9905) );
  INV_X1 U12516 ( .A(n12502), .ZN(n12465) );
  NAND3_X1 U12517 ( .A1(n12465), .A2(n12805), .A3(n10014), .ZN(n9904) );
  OAI211_X1 U12518 ( .C1(n9906), .C2(n12438), .A(n9905), .B(n9904), .ZN(
        P2_U3204) );
  NAND2_X1 U12519 ( .A1(n12798), .A2(n13030), .ZN(n9908) );
  NAND2_X1 U12520 ( .A1(n12800), .A2(n13029), .ZN(n9907) );
  NAND2_X1 U12521 ( .A1(n9908), .A2(n9907), .ZN(n10436) );
  INV_X1 U12522 ( .A(n10436), .ZN(n9910) );
  OAI22_X1 U12523 ( .A1(n12438), .A2(n9910), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9909), .ZN(n9912) );
  NOR2_X1 U12524 ( .A1(n14331), .A2(n10440), .ZN(n9911) );
  AOI211_X1 U12525 ( .C1(n12545), .C2(n14328), .A(n9912), .B(n9911), .ZN(n9918) );
  INV_X1 U12526 ( .A(n9913), .ZN(n9916) );
  INV_X1 U12527 ( .A(n12800), .ZN(n10433) );
  OAI22_X1 U12528 ( .A1(n12502), .A2(n10433), .B1(n9914), .B2(n14302), .ZN(
        n9915) );
  NAND3_X1 U12529 ( .A1(n10001), .A2(n9916), .A3(n9915), .ZN(n9917) );
  OAI211_X1 U12530 ( .C1(n9919), .C2(n14302), .A(n9918), .B(n9917), .ZN(
        P2_U3199) );
  INV_X1 U12531 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U12532 ( .A1(n12337), .A2(n10740), .ZN(n11806) );
  INV_X1 U12533 ( .A(n11806), .ZN(n9920) );
  NOR2_X1 U12534 ( .A1(n12342), .A2(n9920), .ZN(n11780) );
  AND2_X1 U12535 ( .A1(n9921), .A2(n12249), .ZN(n9922) );
  OR2_X1 U12536 ( .A1(n11780), .A2(n9922), .ZN(n9924) );
  NAND2_X1 U12537 ( .A1(n9319), .A2(n14977), .ZN(n9923) );
  NAND2_X1 U12538 ( .A1(n9924), .A2(n9923), .ZN(n10738) );
  INV_X1 U12539 ( .A(n10738), .ZN(n9925) );
  OAI21_X1 U12540 ( .B1(n10740), .B2(n14988), .A(n9925), .ZN(n9948) );
  NAND2_X1 U12541 ( .A1(n9948), .A2(n15072), .ZN(n9926) );
  OAI21_X1 U12542 ( .B1(n15072), .B2(n15347), .A(n9926), .ZN(P3_U3459) );
  INV_X1 U12543 ( .A(n9927), .ZN(n9929) );
  INV_X1 U12544 ( .A(n12820), .ZN(n10935) );
  OAI222_X1 U12545 ( .A1(n13178), .A2(n9929), .B1(n10935), .B2(P2_U3088), .C1(
        n9928), .C2(n13160), .ZN(P2_U3313) );
  INV_X1 U12546 ( .A(n13667), .ZN(n14432) );
  OAI222_X1 U12547 ( .A1(n14047), .A2(n9930), .B1(n14043), .B2(n9929), .C1(
        n14432), .C2(P1_U3086), .ZN(P1_U3341) );
  XNOR2_X1 U12548 ( .A(n10929), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n9934) );
  OAI21_X1 U12549 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n9932), .A(n9931), .ZN(
        n9933) );
  NOR2_X1 U12550 ( .A1(n9933), .A2(n9934), .ZN(n10928) );
  AOI211_X1 U12551 ( .C1(n9934), .C2(n9933), .A(n14695), .B(n10928), .ZN(n9947) );
  MUX2_X1 U12552 ( .A(n9935), .B(P2_REG1_REG_10__SCAN_IN), .S(n10929), .Z(
        n9942) );
  NAND2_X1 U12553 ( .A1(n9937), .A2(n9936), .ZN(n9938) );
  NAND2_X1 U12554 ( .A1(n9939), .A2(n9938), .ZN(n9941) );
  OR2_X1 U12555 ( .A1(n9941), .A2(n9942), .ZN(n10915) );
  INV_X1 U12556 ( .A(n10915), .ZN(n9940) );
  AOI211_X1 U12557 ( .C1(n9942), .C2(n9941), .A(n14707), .B(n9940), .ZN(n9946)
         );
  NAND2_X1 U12558 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10878)
         );
  NAND2_X1 U12559 ( .A1(n14601), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n9943) );
  OAI211_X1 U12560 ( .C1(n14621), .C2(n9944), .A(n10878), .B(n9943), .ZN(n9945) );
  OR3_X1 U12561 ( .A1(n9947), .A2(n9946), .A3(n9945), .ZN(P2_U3224) );
  NAND2_X1 U12562 ( .A1(n9948), .A2(n15055), .ZN(n9949) );
  OAI21_X1 U12563 ( .B1(n8248), .B2(n15055), .A(n9949), .ZN(P3_U3390) );
  INV_X1 U12564 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15226) );
  NAND2_X1 U12565 ( .A1(n14951), .A2(P3_U3897), .ZN(n9950) );
  OAI21_X1 U12566 ( .B1(n11973), .B2(n15226), .A(n9950), .ZN(P3_U3500) );
  INV_X1 U12567 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15277) );
  NAND2_X1 U12568 ( .A1(n14274), .A2(P3_U3897), .ZN(n9951) );
  OAI21_X1 U12569 ( .B1(P3_U3897), .B2(n15277), .A(n9951), .ZN(P3_U3503) );
  OAI22_X1 U12570 ( .A1(n14565), .A2(n11564), .B1(n13321), .B2(n11563), .ZN(
        n9953) );
  XOR2_X1 U12571 ( .A(n9952), .B(n9953), .Z(n9993) );
  NAND2_X1 U12572 ( .A1(n9955), .A2(n9954), .ZN(n9956) );
  NAND2_X1 U12573 ( .A1(n9957), .A2(n9956), .ZN(n9961) );
  OR2_X1 U12574 ( .A1(n14565), .A2(n11563), .ZN(n9959) );
  OAI21_X1 U12575 ( .B1(n9958), .B2(n13321), .A(n9959), .ZN(n9960) );
  NAND2_X1 U12576 ( .A1(n9961), .A2(n9960), .ZN(n9991) );
  AOI21_X1 U12577 ( .B1(n9993), .B2(n9991), .A(n9990), .ZN(n10191) );
  AOI22_X1 U12578 ( .A1(n14571), .A2(n11554), .B1(n9963), .B2(n13570), .ZN(
        n9962) );
  XOR2_X1 U12579 ( .A(n9952), .B(n9962), .Z(n10188) );
  AOI22_X1 U12580 ( .A1(n14571), .A2(n11559), .B1(n11558), .B2(n13570), .ZN(
        n10187) );
  XNOR2_X1 U12581 ( .A(n10188), .B(n10187), .ZN(n9964) );
  XNOR2_X1 U12582 ( .A(n10191), .B(n9964), .ZN(n9970) );
  INV_X1 U12583 ( .A(n10131), .ZN(n9967) );
  AOI22_X1 U12584 ( .A1(n13571), .A2(n13864), .B1(n13262), .B2(n13569), .ZN(
        n10130) );
  OAI21_X1 U12585 ( .B1(n14360), .B2(n10130), .A(n9965), .ZN(n9966) );
  AOI21_X1 U12586 ( .B1(n13293), .B2(n9967), .A(n9966), .ZN(n9969) );
  NAND2_X1 U12587 ( .A1(n9693), .A2(n14571), .ZN(n9968) );
  OAI211_X1 U12588 ( .C1(n9970), .C2(n13286), .A(n9969), .B(n9968), .ZN(
        P1_U3227) );
  INV_X1 U12589 ( .A(n9971), .ZN(n9973) );
  OAI222_X1 U12590 ( .A1(n14239), .A2(P3_U3151), .B1(n14154), .B2(n9973), .C1(
        n9972), .C2(n12417), .ZN(P3_U3277) );
  AOI22_X1 U12591 ( .A1(n12465), .A2(n12803), .B1(n9282), .B2(n8878), .ZN(
        n9975) );
  NOR2_X1 U12592 ( .A1(n9975), .A2(n9974), .ZN(n9980) );
  INV_X1 U12593 ( .A(n14308), .ZN(n12493) );
  INV_X1 U12594 ( .A(n12801), .ZN(n12510) );
  INV_X1 U12595 ( .A(n6589), .ZN(n14757) );
  OAI22_X1 U12596 ( .A1(n12493), .A2(n12510), .B1(n14757), .B2(n14310), .ZN(
        n9978) );
  INV_X1 U12597 ( .A(n14306), .ZN(n12475) );
  OAI22_X1 U12598 ( .A1(n12475), .A2(n12513), .B1(n9976), .B2(n10105), .ZN(
        n9977) );
  AOI211_X1 U12599 ( .C1(n9980), .C2(n9979), .A(n9978), .B(n9977), .ZN(n9981)
         );
  OAI21_X1 U12600 ( .B1(n14302), .B2(n9982), .A(n9981), .ZN(P2_U3209) );
  NAND2_X1 U12601 ( .A1(n13574), .A2(n14526), .ZN(n13308) );
  AND2_X1 U12602 ( .A1(n13310), .A2(n13308), .ZN(n14530) );
  AND2_X1 U12603 ( .A1(n13991), .A2(n14505), .ZN(n9983) );
  OR2_X1 U12604 ( .A1(n14530), .A2(n9983), .ZN(n9988) );
  INV_X1 U12605 ( .A(n9984), .ZN(n14525) );
  INV_X1 U12606 ( .A(n9985), .ZN(n14524) );
  NAND2_X1 U12607 ( .A1(n9986), .A2(n14524), .ZN(n9987) );
  AND3_X1 U12608 ( .A1(n9988), .A2(n14525), .A3(n9987), .ZN(n14540) );
  NAND2_X1 U12609 ( .A1(n14598), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9989) );
  OAI21_X1 U12610 ( .B1(n14598), .B2(n14540), .A(n9989), .ZN(P1_U3528) );
  INV_X1 U12611 ( .A(n9991), .ZN(n9992) );
  NOR2_X1 U12612 ( .A1(n9990), .A2(n9992), .ZN(n9994) );
  XNOR2_X1 U12613 ( .A(n9994), .B(n9993), .ZN(n9995) );
  NAND2_X1 U12614 ( .A1(n9995), .A2(n14365), .ZN(n9999) );
  AND2_X1 U12615 ( .A1(n13570), .A2(n13262), .ZN(n9996) );
  AOI21_X1 U12616 ( .B1(n13572), .B2(n13864), .A(n9996), .ZN(n10086) );
  NAND2_X1 U12617 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13619) );
  OAI21_X1 U12618 ( .B1(n14360), .B2(n10086), .A(n13619), .ZN(n9997) );
  AOI21_X1 U12619 ( .B1(n9693), .B2(n13322), .A(n9997), .ZN(n9998) );
  OAI211_X1 U12620 ( .C1(n14369), .C2(n10090), .A(n9999), .B(n9998), .ZN(
        P1_U3230) );
  INV_X1 U12621 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15152) );
  NAND2_X1 U12622 ( .A1(n11617), .A2(n11973), .ZN(n10000) );
  OAI21_X1 U12623 ( .B1(P3_U3897), .B2(n15152), .A(n10000), .ZN(P3_U3514) );
  OAI21_X1 U12624 ( .B1(n10004), .B2(n10002), .A(n10001), .ZN(n10010) );
  NOR3_X1 U12625 ( .A1(n10004), .A2(n12502), .A3(n10003), .ZN(n10005) );
  OAI21_X1 U12626 ( .B1(n10005), .B2(n14306), .A(n12801), .ZN(n10008) );
  NAND2_X1 U12627 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14623) );
  OAI21_X1 U12628 ( .B1(n14310), .B2(n14769), .A(n14623), .ZN(n10006) );
  AOI21_X1 U12629 ( .B1(n14308), .B2(n12799), .A(n10006), .ZN(n10007) );
  OAI211_X1 U12630 ( .C1(n14331), .C2(n10426), .A(n10008), .B(n10007), .ZN(
        n10009) );
  AOI21_X1 U12631 ( .B1(n10010), .B2(n9282), .A(n10009), .ZN(n10011) );
  INV_X1 U12632 ( .A(n10011), .ZN(P2_U3202) );
  OAI222_X1 U12633 ( .A1(n14154), .A2(n10012), .B1(n12057), .B2(P3_U3151), 
        .C1(n12417), .C2(n15339), .ZN(P3_U3276) );
  NAND2_X1 U12634 ( .A1(n12512), .A2(n12803), .ZN(n12521) );
  NAND2_X1 U12635 ( .A1(n10013), .A2(n12514), .ZN(n12517) );
  NAND2_X1 U12636 ( .A1(n10015), .A2(n10014), .ZN(n10097) );
  INV_X1 U12637 ( .A(n10097), .ZN(n10016) );
  AOI21_X1 U12638 ( .B1(n10017), .B2(n12728), .A(n10016), .ZN(n10055) );
  INV_X1 U12639 ( .A(n12515), .ZN(n10019) );
  OAI21_X1 U12640 ( .B1(n10019), .B2(n12728), .A(n10100), .ZN(n10023) );
  INV_X1 U12641 ( .A(n12802), .ZN(n10419) );
  OAI22_X1 U12642 ( .A1(n10020), .A2(n13004), .B1(n10419), .B2(n13006), .ZN(
        n10022) );
  NOR2_X1 U12643 ( .A1(n10055), .A2(n9731), .ZN(n10021) );
  AOI211_X1 U12644 ( .C1(n13026), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10059) );
  AOI21_X1 U12645 ( .B1(n10024), .B2(n6560), .A(n9183), .ZN(n10026) );
  NAND2_X1 U12646 ( .A1(n12512), .A2(n10025), .ZN(n10106) );
  AND2_X1 U12647 ( .A1(n10026), .A2(n10106), .ZN(n10053) );
  AOI21_X1 U12648 ( .B1(n14818), .B2(n6560), .A(n10053), .ZN(n10027) );
  OAI211_X1 U12649 ( .C1(n10055), .C2(n14822), .A(n10059), .B(n10027), .ZN(
        n10031) );
  NAND2_X1 U12650 ( .A1(n10031), .A2(n14842), .ZN(n10028) );
  OAI21_X1 U12651 ( .B1(n14842), .B2(n10029), .A(n10028), .ZN(P2_U3500) );
  INV_X1 U12652 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U12653 ( .A1(n10031), .A2(n14829), .ZN(n10032) );
  OAI21_X1 U12654 ( .B1(n14829), .B2(n10033), .A(n10032), .ZN(P2_U3433) );
  INV_X1 U12655 ( .A(n12549), .ZN(n14781) );
  AOI21_X1 U12656 ( .B1(n10035), .B2(n10034), .A(n14302), .ZN(n10037) );
  NAND2_X1 U12657 ( .A1(n10037), .A2(n10036), .ZN(n10043) );
  INV_X1 U12658 ( .A(n10038), .ZN(n10510) );
  NAND2_X1 U12659 ( .A1(n12797), .A2(n13030), .ZN(n10040) );
  NAND2_X1 U12660 ( .A1(n12799), .A2(n13029), .ZN(n10039) );
  AND2_X1 U12661 ( .A1(n10040), .A2(n10039), .ZN(n10507) );
  NAND2_X1 U12662 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14636) );
  OAI21_X1 U12663 ( .B1(n12438), .B2(n10507), .A(n14636), .ZN(n10041) );
  AOI21_X1 U12664 ( .B1(n12489), .B2(n10510), .A(n10041), .ZN(n10042) );
  OAI211_X1 U12665 ( .C1(n14781), .C2(n14310), .A(n10043), .B(n10042), .ZN(
        P2_U3211) );
  INV_X1 U12666 ( .A(n10044), .ZN(n10046) );
  OAI222_X1 U12667 ( .A1(n14047), .A2(n10045), .B1(n14043), .B2(n10046), .C1(
        P1_U3086), .C2(n14445), .ZN(P1_U3340) );
  OAI222_X1 U12668 ( .A1(n13160), .A2(n10047), .B1(n13178), .B2(n10046), .C1(
        P2_U3088), .C2(n12830), .ZN(P2_U3312) );
  INV_X1 U12669 ( .A(n11741), .ZN(n10407) );
  NAND2_X1 U12670 ( .A1(n10407), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10387) );
  NAND2_X1 U12671 ( .A1(n10387), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U12672 ( .A1(n11746), .A2(n10048), .B1(n11740), .B2(n9319), .ZN(
        n10049) );
  OAI211_X1 U12673 ( .C1(n11780), .C2(n11748), .A(n10050), .B(n10049), .ZN(
        P3_U3172) );
  OAI22_X1 U12674 ( .A1(n12979), .A2(n9551), .B1(n10052), .B2(n13041), .ZN(
        n10057) );
  INV_X1 U12675 ( .A(n10053), .ZN(n10054) );
  OAI22_X1 U12676 ( .A1(n10055), .A2(n13020), .B1(n13047), .B2(n10054), .ZN(
        n10056) );
  AOI211_X1 U12677 ( .C1(n13044), .C2(n6560), .A(n10057), .B(n10056), .ZN(
        n10058) );
  OAI21_X1 U12678 ( .B1(n10059), .B2(n13051), .A(n10058), .ZN(P2_U3264) );
  MUX2_X1 U12679 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10061), .S(n13642), .Z(
        n10062) );
  NAND2_X1 U12680 ( .A1(n10063), .A2(n10062), .ZN(n13641) );
  OAI21_X1 U12681 ( .B1(n10063), .B2(n10062), .A(n13641), .ZN(n10074) );
  INV_X1 U12682 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U12683 ( .A1(n14493), .A2(n13642), .ZN(n10065) );
  NAND2_X1 U12684 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10064)
         );
  OAI211_X1 U12685 ( .C1(n14076), .C2(n14499), .A(n10065), .B(n10064), .ZN(
        n10073) );
  INV_X1 U12686 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10068) );
  MUX2_X1 U12687 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10068), .S(n13642), .Z(
        n10069) );
  INV_X1 U12688 ( .A(n10069), .ZN(n10070) );
  AOI211_X1 U12689 ( .C1(n10071), .C2(n10070), .A(n14488), .B(n13633), .ZN(
        n10072) );
  AOI211_X1 U12690 ( .C1(n14483), .C2(n10074), .A(n10073), .B(n10072), .ZN(
        n10075) );
  INV_X1 U12691 ( .A(n10075), .ZN(P1_U3254) );
  NAND3_X1 U12692 ( .A1(n10078), .A2(n10077), .A3(n10076), .ZN(n10080) );
  AND2_X1 U12693 ( .A1(n10083), .A2(n10082), .ZN(n13496) );
  XNOR2_X1 U12694 ( .A(n10084), .B(n13496), .ZN(n14568) );
  INV_X1 U12695 ( .A(n14568), .ZN(n10095) );
  XNOR2_X1 U12696 ( .A(n10085), .B(n13496), .ZN(n10087) );
  OAI21_X1 U12697 ( .B1(n10087), .B2(n14505), .A(n10086), .ZN(n14566) );
  NAND2_X1 U12698 ( .A1(n14536), .A2(n14523), .ZN(n13888) );
  AOI21_X1 U12699 ( .B1(n14514), .B2(n13322), .A(n13884), .ZN(n10088) );
  NAND2_X1 U12700 ( .A1(n10088), .A2(n10133), .ZN(n14564) );
  INV_X1 U12701 ( .A(n10089), .ZN(n14522) );
  OAI22_X1 U12702 ( .A1(n14536), .A2(n7630), .B1(n10090), .B2(n14508), .ZN(
        n10091) );
  AOI21_X1 U12703 ( .B1(n14512), .B2(n13322), .A(n10091), .ZN(n10092) );
  OAI21_X1 U12704 ( .B1(n13888), .B2(n14564), .A(n10092), .ZN(n10093) );
  AOI21_X1 U12705 ( .B1(n14536), .B2(n14566), .A(n10093), .ZN(n10094) );
  OAI21_X1 U12706 ( .B1(n13895), .B2(n10095), .A(n10094), .ZN(P1_U3289) );
  NAND2_X1 U12707 ( .A1(n12513), .A2(n12512), .ZN(n10096) );
  NAND2_X1 U12708 ( .A1(n10097), .A2(n10096), .ZN(n10099) );
  OAI21_X1 U12709 ( .B1(n10099), .B2(n10098), .A(n10421), .ZN(n14760) );
  INV_X1 U12710 ( .A(n14760), .ZN(n10112) );
  NAND2_X1 U12711 ( .A1(n10100), .A2(n12517), .ZN(n10101) );
  NAND2_X1 U12712 ( .A1(n10101), .A2(n12727), .ZN(n10414) );
  OAI21_X1 U12713 ( .B1(n10101), .B2(n12727), .A(n10414), .ZN(n10103) );
  OAI22_X1 U12714 ( .A1(n12510), .A2(n13006), .B1(n12513), .B2(n13004), .ZN(
        n10102) );
  AOI21_X1 U12715 ( .B1(n10103), .B2(n13026), .A(n10102), .ZN(n10104) );
  OAI21_X1 U12716 ( .B1(n10112), .B2(n9731), .A(n10104), .ZN(n14758) );
  NAND2_X1 U12717 ( .A1(n14758), .A2(n12979), .ZN(n10111) );
  OAI22_X1 U12718 ( .A1(n12979), .A2(n9564), .B1(n10105), .B2(n13041), .ZN(
        n10109) );
  INV_X1 U12719 ( .A(n10106), .ZN(n10107) );
  OAI211_X1 U12720 ( .C1(n10107), .C2(n14757), .A(n12913), .B(n10531), .ZN(
        n14756) );
  NOR2_X1 U12721 ( .A1(n13047), .A2(n14756), .ZN(n10108) );
  AOI211_X1 U12722 ( .C1(n13044), .C2(n6589), .A(n10109), .B(n10108), .ZN(
        n10110) );
  OAI211_X1 U12723 ( .C1(n10112), .C2(n13020), .A(n10111), .B(n10110), .ZN(
        P2_U3263) );
  INV_X1 U12724 ( .A(n12558), .ZN(n14790) );
  AOI21_X1 U12725 ( .B1(n10036), .B2(n7414), .A(n14302), .ZN(n10117) );
  INV_X1 U12726 ( .A(n12798), .ZN(n10605) );
  INV_X1 U12727 ( .A(n10114), .ZN(n10115) );
  NOR3_X1 U12728 ( .A1(n12502), .A2(n10605), .A3(n10115), .ZN(n10116) );
  OAI21_X1 U12729 ( .B1(n10117), .B2(n10116), .A(n12446), .ZN(n10124) );
  INV_X1 U12730 ( .A(n10118), .ZN(n10638) );
  NAND2_X1 U12731 ( .A1(n12796), .A2(n13030), .ZN(n10120) );
  NAND2_X1 U12732 ( .A1(n12798), .A2(n13029), .ZN(n10119) );
  AND2_X1 U12733 ( .A1(n10120), .A2(n10119), .ZN(n10631) );
  OAI22_X1 U12734 ( .A1(n12438), .A2(n10631), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10121), .ZN(n10122) );
  AOI21_X1 U12735 ( .B1(n12489), .B2(n10638), .A(n10122), .ZN(n10123) );
  OAI211_X1 U12736 ( .C1(n14790), .C2(n14310), .A(n10124), .B(n10123), .ZN(
        P2_U3185) );
  AOI21_X1 U12737 ( .B1(n13497), .B2(n10125), .A(n6718), .ZN(n14570) );
  NAND2_X1 U12738 ( .A1(n10126), .A2(n13525), .ZN(n13481) );
  XOR2_X1 U12739 ( .A(n13497), .B(n10127), .Z(n10128) );
  NAND2_X1 U12740 ( .A1(n10128), .A2(n14585), .ZN(n10129) );
  OAI211_X1 U12741 ( .C1(n14570), .C2(n11340), .A(n10130), .B(n10129), .ZN(
        n14573) );
  NAND2_X1 U12742 ( .A1(n14573), .A2(n14536), .ZN(n10138) );
  INV_X1 U12743 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10132) );
  OAI22_X1 U12744 ( .A1(n14536), .A2(n10132), .B1(n10131), .B2(n14508), .ZN(
        n10136) );
  AOI21_X1 U12745 ( .B1(n10133), .B2(n14571), .A(n13884), .ZN(n10134) );
  NAND2_X1 U12746 ( .A1(n10134), .A2(n10226), .ZN(n14572) );
  NOR2_X1 U12747 ( .A1(n13888), .A2(n14572), .ZN(n10135) );
  AOI211_X1 U12748 ( .C1(n14512), .C2(n14571), .A(n10136), .B(n10135), .ZN(
        n10137) );
  OAI211_X1 U12749 ( .C1(n14570), .C2(n13877), .A(n10138), .B(n10137), .ZN(
        P1_U3288) );
  OAI21_X1 U12750 ( .B1(n10140), .B2(n13502), .A(n10139), .ZN(n14589) );
  INV_X1 U12751 ( .A(n14589), .ZN(n10151) );
  NAND2_X1 U12752 ( .A1(n13568), .A2(n13864), .ZN(n10142) );
  NAND2_X1 U12753 ( .A1(n13566), .A2(n13262), .ZN(n10141) );
  NAND2_X1 U12754 ( .A1(n10142), .A2(n10141), .ZN(n14579) );
  INV_X1 U12755 ( .A(n10788), .ZN(n10143) );
  INV_X1 U12756 ( .A(n14508), .ZN(n14528) );
  AOI22_X1 U12757 ( .A1(n14536), .A2(n14579), .B1(n10143), .B2(n14528), .ZN(
        n10144) );
  OAI21_X1 U12758 ( .B1(n9673), .B2(n14536), .A(n10144), .ZN(n10147) );
  AOI21_X1 U12759 ( .B1(n10163), .B2(n14578), .A(n13884), .ZN(n10145) );
  NAND2_X1 U12760 ( .A1(n10145), .A2(n6608), .ZN(n14581) );
  NOR2_X1 U12761 ( .A1(n14581), .A2(n13888), .ZN(n10146) );
  AOI211_X1 U12762 ( .C1(n14512), .C2(n14578), .A(n10147), .B(n10146), .ZN(
        n10150) );
  NAND2_X1 U12763 ( .A1(n10148), .A2(n13502), .ZN(n14584) );
  NAND3_X1 U12764 ( .A1(n14586), .A2(n14584), .A3(n14532), .ZN(n10149) );
  OAI211_X1 U12765 ( .C1(n10151), .C2(n13895), .A(n10150), .B(n10149), .ZN(
        P1_U3285) );
  INV_X1 U12766 ( .A(n10152), .ZN(n10183) );
  INV_X1 U12767 ( .A(n14461), .ZN(n10153) );
  OAI222_X1 U12768 ( .A1(n14047), .A2(n10154), .B1(n14043), .B2(n10183), .C1(
        n10153), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI21_X1 U12769 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(n10158) );
  INV_X1 U12770 ( .A(n10158), .ZN(n10171) );
  NAND2_X1 U12771 ( .A1(n13569), .A2(n13864), .ZN(n10160) );
  NAND2_X1 U12772 ( .A1(n13567), .A2(n13262), .ZN(n10159) );
  NAND2_X1 U12773 ( .A1(n10160), .A2(n10159), .ZN(n10208) );
  INV_X1 U12774 ( .A(n10211), .ZN(n10161) );
  AOI22_X1 U12775 ( .A1(n14536), .A2(n10208), .B1(n10161), .B2(n14528), .ZN(
        n10162) );
  OAI21_X1 U12776 ( .B1(n9618), .B2(n14536), .A(n10162), .ZN(n10165) );
  OAI211_X1 U12777 ( .C1(n10225), .C2(n10215), .A(n14513), .B(n10163), .ZN(
        n10169) );
  NOR2_X1 U12778 ( .A1(n10169), .A2(n13888), .ZN(n10164) );
  AOI211_X1 U12779 ( .C1(n14512), .C2(n13333), .A(n10165), .B(n10164), .ZN(
        n10168) );
  XNOR2_X1 U12780 ( .A(n10166), .B(n13500), .ZN(n10173) );
  NAND2_X1 U12781 ( .A1(n10173), .A2(n14532), .ZN(n10167) );
  OAI211_X1 U12782 ( .C1(n10171), .C2(n13895), .A(n10168), .B(n10167), .ZN(
        P1_U3286) );
  INV_X1 U12783 ( .A(n10208), .ZN(n10170) );
  OAI211_X1 U12784 ( .C1(n10171), .C2(n13991), .A(n10170), .B(n10169), .ZN(
        n10172) );
  AOI21_X1 U12785 ( .B1(n14585), .B2(n10173), .A(n10172), .ZN(n10179) );
  OAI22_X1 U12786 ( .A1(n13976), .A2(n10215), .B1(n14600), .B2(n9623), .ZN(
        n10174) );
  INV_X1 U12787 ( .A(n10174), .ZN(n10175) );
  OAI21_X1 U12788 ( .B1(n10179), .B2(n14598), .A(n10175), .ZN(P1_U3535) );
  INV_X1 U12789 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10176) );
  OAI22_X1 U12790 ( .A1(n14028), .A2(n10215), .B1(n8150), .B2(n10176), .ZN(
        n10177) );
  INV_X1 U12791 ( .A(n10177), .ZN(n10178) );
  OAI21_X1 U12792 ( .B1(n10179), .B2(n14577), .A(n10178), .ZN(P1_U3480) );
  INV_X1 U12793 ( .A(n10180), .ZN(n10181) );
  OAI222_X1 U12794 ( .A1(P3_U3151), .A2(n10182), .B1(n12417), .B2(n15138), 
        .C1(n14154), .C2(n10181), .ZN(P3_U3275) );
  INV_X1 U12795 ( .A(n14689), .ZN(n10184) );
  OAI222_X1 U12796 ( .A1(n13160), .A2(n10185), .B1(n10184), .B2(P2_U3088), 
        .C1(n13178), .C2(n10183), .ZN(P2_U3311) );
  INV_X1 U12797 ( .A(n10188), .ZN(n10186) );
  NAND2_X1 U12798 ( .A1(n10186), .A2(n10187), .ZN(n10190) );
  NAND2_X1 U12799 ( .A1(n13330), .A2(n11554), .ZN(n10193) );
  NAND2_X1 U12800 ( .A1(n13569), .A2(n11559), .ZN(n10192) );
  NAND2_X1 U12801 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  XNOR2_X1 U12802 ( .A(n10194), .B(n11476), .ZN(n10200) );
  INV_X1 U12803 ( .A(n10200), .ZN(n10198) );
  NOR2_X1 U12804 ( .A1(n9958), .A2(n10195), .ZN(n10196) );
  AOI21_X1 U12805 ( .B1(n13330), .B2(n11559), .A(n10196), .ZN(n10199) );
  INV_X1 U12806 ( .A(n10199), .ZN(n10197) );
  NAND2_X1 U12807 ( .A1(n10198), .A2(n10197), .ZN(n10451) );
  AND2_X1 U12808 ( .A1(n10200), .A2(n10199), .ZN(n10450) );
  NAND2_X1 U12809 ( .A1(n13333), .A2(n11554), .ZN(n10202) );
  NAND2_X1 U12810 ( .A1(n13568), .A2(n11559), .ZN(n10201) );
  NAND2_X1 U12811 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  XNOR2_X1 U12812 ( .A(n10203), .B(n9952), .ZN(n10792) );
  NOR2_X1 U12813 ( .A1(n9958), .A2(n10204), .ZN(n10205) );
  AOI21_X1 U12814 ( .B1(n13333), .B2(n11559), .A(n10205), .ZN(n10794) );
  XNOR2_X1 U12815 ( .A(n10792), .B(n10794), .ZN(n10206) );
  OAI211_X1 U12816 ( .C1(n10207), .C2(n10206), .A(n10793), .B(n14365), .ZN(
        n10214) );
  NAND2_X1 U12817 ( .A1(n14353), .A2(n10208), .ZN(n10209) );
  OAI211_X1 U12818 ( .C1(n14369), .C2(n10211), .A(n10210), .B(n10209), .ZN(
        n10212) );
  INV_X1 U12819 ( .A(n10212), .ZN(n10213) );
  OAI211_X1 U12820 ( .C1(n10215), .C2(n14362), .A(n10214), .B(n10213), .ZN(
        P1_U3213) );
  XOR2_X1 U12821 ( .A(n10216), .B(n10217), .Z(n10222) );
  AOI22_X1 U12822 ( .A1(n11740), .A2(n12329), .B1(n11731), .B2(n9319), .ZN(
        n10218) );
  OAI21_X1 U12823 ( .B1(n10219), .B2(n11737), .A(n10218), .ZN(n10220) );
  AOI21_X1 U12824 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10387), .A(n10220), .ZN(
        n10221) );
  OAI21_X1 U12825 ( .B1(n10222), .B2(n11748), .A(n10221), .ZN(P3_U3177) );
  INV_X1 U12826 ( .A(n14553), .ZN(n14576) );
  OAI21_X1 U12827 ( .B1(n10224), .B2(n10228), .A(n10223), .ZN(n10487) );
  AOI211_X1 U12828 ( .C1(n13330), .C2(n10226), .A(n13884), .B(n10225), .ZN(
        n10494) );
  XNOR2_X1 U12829 ( .A(n10227), .B(n10228), .ZN(n10232) );
  INV_X1 U12830 ( .A(n11340), .ZN(n14557) );
  NAND2_X1 U12831 ( .A1(n13568), .A2(n13262), .ZN(n10230) );
  NAND2_X1 U12832 ( .A1(n13570), .A2(n13864), .ZN(n10229) );
  NAND2_X1 U12833 ( .A1(n10230), .A2(n10229), .ZN(n10447) );
  AOI21_X1 U12834 ( .B1(n10487), .B2(n14557), .A(n10447), .ZN(n10231) );
  OAI21_X1 U12835 ( .B1(n14505), .B2(n10232), .A(n10231), .ZN(n10488) );
  AOI211_X1 U12836 ( .C1(n14576), .C2(n10487), .A(n10494), .B(n10488), .ZN(
        n10237) );
  INV_X1 U12837 ( .A(n13330), .ZN(n10489) );
  INV_X1 U12838 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U12839 ( .A1(n14028), .A2(n10489), .B1(n8150), .B2(n15233), .ZN(
        n10233) );
  INV_X1 U12840 ( .A(n10233), .ZN(n10234) );
  OAI21_X1 U12841 ( .B1(n10237), .B2(n14577), .A(n10234), .ZN(P1_U3477) );
  OAI22_X1 U12842 ( .A1(n13976), .A2(n10489), .B1(n14600), .B2(n9603), .ZN(
        n10235) );
  INV_X1 U12843 ( .A(n10235), .ZN(n10236) );
  OAI21_X1 U12844 ( .B1(n10237), .B2(n14598), .A(n10236), .ZN(P1_U3534) );
  NAND2_X1 U12845 ( .A1(P3_U3897), .A2(n11329), .ZN(n14933) );
  INV_X1 U12846 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10253) );
  MUX2_X1 U12847 ( .A(n10253), .B(n15347), .S(n6590), .Z(n14843) );
  AND2_X1 U12848 ( .A1(n14843), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14847) );
  MUX2_X1 U12849 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6590), .Z(n10265) );
  XOR2_X1 U12850 ( .A(n10255), .B(n10265), .Z(n10268) );
  XOR2_X1 U12851 ( .A(n14847), .B(n10268), .Z(n10264) );
  INV_X2 U12852 ( .A(n11973), .ZN(n11981) );
  INV_X1 U12853 ( .A(n10238), .ZN(n10239) );
  OR2_X1 U12854 ( .A1(n10240), .A2(P3_U3151), .ZN(n11968) );
  NAND2_X1 U12855 ( .A1(n10239), .A2(n11968), .ZN(n10250) );
  INV_X1 U12856 ( .A(n10240), .ZN(n10241) );
  OR2_X1 U12857 ( .A1(n11911), .A2(n10241), .ZN(n10242) );
  INV_X1 U12858 ( .A(n10259), .ZN(n10243) );
  MUX2_X1 U12859 ( .A(n11981), .B(n10243), .S(n11329), .Z(n14939) );
  INV_X1 U12860 ( .A(n14939), .ZN(n14866) );
  INV_X1 U12861 ( .A(n10255), .ZN(n10267) );
  INV_X1 U12862 ( .A(n14929), .ZN(n14844) );
  INV_X1 U12863 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10247) );
  AND2_X1 U12864 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n15154), .ZN(n10244) );
  OR3_X1 U12865 ( .A1(n15347), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n10280) );
  OAI21_X1 U12866 ( .B1(n10255), .B2(n10244), .A(n10280), .ZN(n10246) );
  OR2_X1 U12867 ( .A1(n10246), .A2(n10247), .ZN(n10281) );
  INV_X1 U12868 ( .A(n10281), .ZN(n10245) );
  AOI21_X1 U12869 ( .B1(n10247), .B2(n10246), .A(n10245), .ZN(n10252) );
  INV_X1 U12870 ( .A(n10248), .ZN(n10249) );
  AOI22_X1 U12871 ( .A1(n14860), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10251) );
  OAI21_X1 U12872 ( .B1(n14844), .B2(n10252), .A(n10251), .ZN(n10262) );
  NOR2_X1 U12873 ( .A1(n10253), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10254) );
  OAI21_X1 U12874 ( .B1(n10255), .B2(n10254), .A(n6613), .ZN(n10256) );
  INV_X1 U12875 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15016) );
  OR2_X1 U12876 ( .A1(n10256), .A2(n15016), .ZN(n10272) );
  NAND2_X1 U12877 ( .A1(n10256), .A2(n15016), .ZN(n10260) );
  INV_X1 U12878 ( .A(n10257), .ZN(n10258) );
  AND2_X1 U12879 ( .A1(n10259), .A2(n10258), .ZN(n14192) );
  AOI21_X1 U12880 ( .B1(n10272), .B2(n10260), .A(n14945), .ZN(n10261) );
  AOI211_X1 U12881 ( .C1(n14866), .C2(n10267), .A(n10262), .B(n10261), .ZN(
        n10263) );
  OAI21_X1 U12882 ( .B1(n14933), .B2(n10264), .A(n10263), .ZN(P3_U3183) );
  MUX2_X1 U12883 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n6590), .Z(n10300) );
  XOR2_X1 U12884 ( .A(n10297), .B(n10300), .Z(n10301) );
  INV_X1 U12885 ( .A(n10265), .ZN(n10266) );
  AOI22_X1 U12886 ( .A1(n10268), .A2(n14847), .B1(n10267), .B2(n10266), .ZN(
        n10331) );
  MUX2_X1 U12887 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n6590), .Z(n10269) );
  XOR2_X1 U12888 ( .A(n10343), .B(n10269), .Z(n10332) );
  OAI22_X1 U12889 ( .A1(n10331), .A2(n10332), .B1(n10269), .B2(n7132), .ZN(
        n10365) );
  MUX2_X1 U12890 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n6590), .Z(n10270) );
  XNOR2_X1 U12891 ( .A(n10270), .B(n10374), .ZN(n10366) );
  INV_X1 U12892 ( .A(n10270), .ZN(n10271) );
  AOI22_X1 U12893 ( .A1(n10365), .A2(n10366), .B1(n10374), .B2(n10271), .ZN(
        n10302) );
  XOR2_X1 U12894 ( .A(n10301), .B(n10302), .Z(n10299) );
  INV_X1 U12895 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10592) );
  MUX2_X1 U12896 ( .A(n10592), .B(P3_REG2_REG_4__SCAN_IN), .S(n10297), .Z(
        n10277) );
  INV_X1 U12897 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U12898 ( .A1(n10272), .A2(n6613), .ZN(n10336) );
  OR2_X1 U12899 ( .A1(n10343), .A2(n15005), .ZN(n10273) );
  INV_X1 U12900 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14994) );
  NAND2_X1 U12901 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  OAI21_X1 U12902 ( .B1(n10277), .B2(n10276), .A(n10316), .ZN(n10278) );
  NAND2_X1 U12903 ( .A1(n14192), .A2(n10278), .ZN(n10295) );
  INV_X1 U12904 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10279) );
  MUX2_X1 U12905 ( .A(n10279), .B(P3_REG1_REG_4__SCAN_IN), .S(n10297), .Z(
        n10290) );
  NAND2_X1 U12906 ( .A1(n10281), .A2(n10280), .ZN(n10334) );
  NAND2_X1 U12907 ( .A1(n10333), .A2(n10334), .ZN(n10284) );
  INV_X1 U12908 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10282) );
  OR2_X1 U12909 ( .A1(n10343), .A2(n10282), .ZN(n10283) );
  XNOR2_X1 U12910 ( .A(n10286), .B(n10374), .ZN(n10368) );
  NAND2_X1 U12911 ( .A1(n10368), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U12912 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  NAND2_X1 U12913 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  NAND2_X1 U12914 ( .A1(n10289), .A2(n10290), .ZN(n10307) );
  OAI21_X1 U12915 ( .B1(n10290), .B2(n10289), .A(n10307), .ZN(n10291) );
  NAND2_X1 U12916 ( .A1(n14929), .A2(n10291), .ZN(n10294) );
  INV_X1 U12917 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10292) );
  NOR2_X1 U12918 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10292), .ZN(n10522) );
  AOI21_X1 U12919 ( .B1(n14860), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10522), .ZN(
        n10293) );
  NAND3_X1 U12920 ( .A1(n10295), .A2(n10294), .A3(n10293), .ZN(n10296) );
  AOI21_X1 U12921 ( .B1(n14866), .B2(n10297), .A(n10296), .ZN(n10298) );
  OAI21_X1 U12922 ( .B1(n10299), .B2(n14933), .A(n10298), .ZN(P3_U3186) );
  MUX2_X1 U12923 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6590), .Z(n10346) );
  XNOR2_X1 U12924 ( .A(n10346), .B(n10348), .ZN(n10349) );
  OAI22_X1 U12925 ( .A1(n10302), .A2(n10301), .B1(n10300), .B2(n10314), .ZN(
        n10565) );
  MUX2_X1 U12926 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n6590), .Z(n10303) );
  XNOR2_X1 U12927 ( .A(n10303), .B(n10308), .ZN(n10566) );
  INV_X1 U12928 ( .A(n10303), .ZN(n10304) );
  MUX2_X1 U12929 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6590), .Z(n10305) );
  XNOR2_X1 U12930 ( .A(n10305), .B(n10550), .ZN(n10552) );
  OAI22_X1 U12931 ( .A1(n10551), .A2(n10552), .B1(n10305), .B2(n10550), .ZN(
        n10350) );
  XOR2_X1 U12932 ( .A(n10349), .B(n10350), .Z(n10330) );
  INV_X1 U12933 ( .A(n10550), .ZN(n10312) );
  INV_X1 U12934 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15062) );
  NAND2_X1 U12935 ( .A1(n10314), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12936 ( .A1(n10558), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U12937 ( .A1(n10309), .A2(n10564), .ZN(n10310) );
  NAND2_X1 U12938 ( .A1(n10311), .A2(n10310), .ZN(n10542) );
  MUX2_X1 U12939 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15062), .S(n10550), .Z(
        n10543) );
  NAND2_X1 U12940 ( .A1(n10542), .A2(n10543), .ZN(n10541) );
  XNOR2_X1 U12941 ( .A(n10353), .B(n10348), .ZN(n10313) );
  NAND2_X1 U12942 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10313), .ZN(n10354) );
  OAI21_X1 U12943 ( .B1(n10313), .B2(P3_REG1_REG_7__SCAN_IN), .A(n10354), .ZN(
        n10328) );
  NAND2_X1 U12944 ( .A1(n10314), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10315) );
  INV_X1 U12945 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U12946 ( .A1(n10319), .A2(n10318), .ZN(n10545) );
  INV_X1 U12947 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n14974) );
  MUX2_X1 U12948 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n14974), .S(n10550), .Z(
        n10546) );
  NAND2_X1 U12949 ( .A1(n10545), .A2(n10546), .ZN(n10544) );
  NAND2_X1 U12950 ( .A1(n10550), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U12951 ( .A1(n10544), .A2(n10320), .ZN(n10321) );
  OR2_X1 U12952 ( .A1(n10321), .A2(n10352), .ZN(n10322) );
  INV_X1 U12953 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10783) );
  XNOR2_X1 U12954 ( .A(n10351), .B(n10783), .ZN(n10323) );
  NAND2_X1 U12955 ( .A1(n10323), .A2(n14192), .ZN(n10326) );
  INV_X1 U12956 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10324) );
  NOR2_X1 U12957 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10324), .ZN(n11609) );
  AOI21_X1 U12958 ( .B1(n14860), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11609), .ZN(
        n10325) );
  OAI211_X1 U12959 ( .C1(n14939), .C2(n10352), .A(n10326), .B(n10325), .ZN(
        n10327) );
  AOI21_X1 U12960 ( .B1(n14929), .B2(n10328), .A(n10327), .ZN(n10329) );
  OAI21_X1 U12961 ( .B1(n10330), .B2(n14933), .A(n10329), .ZN(P3_U3189) );
  XOR2_X1 U12962 ( .A(n10332), .B(n10331), .Z(n10345) );
  XOR2_X1 U12963 ( .A(n10334), .B(n10333), .Z(n10341) );
  AOI22_X1 U12964 ( .A1(n14860), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10340) );
  OAI21_X1 U12965 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10338) );
  NAND2_X1 U12966 ( .A1(n14192), .A2(n10338), .ZN(n10339) );
  OAI211_X1 U12967 ( .C1(n14844), .C2(n10341), .A(n10340), .B(n10339), .ZN(
        n10342) );
  AOI21_X1 U12968 ( .B1(n10343), .B2(n14866), .A(n10342), .ZN(n10344) );
  OAI21_X1 U12969 ( .B1(n10345), .B2(n14933), .A(n10344), .ZN(P3_U3184) );
  MUX2_X1 U12970 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n6590), .Z(n10667) );
  XNOR2_X1 U12971 ( .A(n10667), .B(n10675), .ZN(n10668) );
  INV_X1 U12972 ( .A(n10346), .ZN(n10347) );
  AOI22_X1 U12973 ( .A1(n10350), .A2(n10349), .B1(n10348), .B2(n10347), .ZN(
        n10669) );
  XOR2_X1 U12974 ( .A(n10668), .B(n10669), .Z(n10364) );
  INV_X1 U12975 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U12976 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10677), .B1(n10675), 
        .B2(n14958), .ZN(n10673) );
  XNOR2_X1 U12977 ( .A(n10674), .B(n10673), .ZN(n10362) );
  INV_X1 U12978 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U12979 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10675), .B1(n10677), 
        .B2(n15066), .ZN(n10357) );
  NAND2_X1 U12980 ( .A1(n10353), .A2(n10352), .ZN(n10355) );
  NAND2_X1 U12981 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NAND2_X1 U12982 ( .A1(n10357), .A2(n10356), .ZN(n10676) );
  OAI21_X1 U12983 ( .B1(n10357), .B2(n10356), .A(n10676), .ZN(n10358) );
  NAND2_X1 U12984 ( .A1(n10358), .A2(n14929), .ZN(n10360) );
  AND2_X1 U12985 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11643) );
  AOI21_X1 U12986 ( .B1(n14860), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11643), .ZN(
        n10359) );
  OAI211_X1 U12987 ( .C1(n14939), .C2(n10675), .A(n10360), .B(n10359), .ZN(
        n10361) );
  AOI21_X1 U12988 ( .B1(n14192), .B2(n10362), .A(n10361), .ZN(n10363) );
  OAI21_X1 U12989 ( .B1(n10364), .B2(n14933), .A(n10363), .ZN(P3_U3190) );
  XOR2_X1 U12990 ( .A(n10366), .B(n10365), .Z(n10376) );
  XNOR2_X1 U12991 ( .A(n10367), .B(P3_REG2_REG_3__SCAN_IN), .ZN(n10372) );
  NOR2_X1 U12992 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14990), .ZN(n10404) );
  AOI21_X1 U12993 ( .B1(n14860), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10404), .ZN(
        n10371) );
  XNOR2_X1 U12994 ( .A(n10368), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U12995 ( .A1(n14929), .A2(n10369), .ZN(n10370) );
  OAI211_X1 U12996 ( .C1(n14945), .C2(n10372), .A(n10371), .B(n10370), .ZN(
        n10373) );
  AOI21_X1 U12997 ( .B1(n10374), .B2(n14866), .A(n10373), .ZN(n10375) );
  OAI21_X1 U12998 ( .B1(n10376), .B2(n14933), .A(n10375), .ZN(P3_U3185) );
  NAND2_X1 U12999 ( .A1(n12793), .A2(n13030), .ZN(n10378) );
  NAND2_X1 U13000 ( .A1(n12796), .A2(n13029), .ZN(n10377) );
  AND2_X1 U13001 ( .A1(n10378), .A2(n10377), .ZN(n10693) );
  OAI21_X1 U13002 ( .B1(n12438), .B2(n10693), .A(n10379), .ZN(n10381) );
  NOR2_X1 U13003 ( .A1(n14331), .A2(n10701), .ZN(n10380) );
  AOI211_X1 U13004 ( .C1(n14803), .C2(n14328), .A(n10381), .B(n10380), .ZN(
        n10385) );
  OAI22_X1 U13005 ( .A1(n10382), .A2(n14302), .B1(n10686), .B2(n12502), .ZN(
        n10383) );
  NAND3_X1 U13006 ( .A1(n12445), .A2(n6724), .A3(n10383), .ZN(n10384) );
  OAI211_X1 U13007 ( .C1(n10386), .C2(n14302), .A(n10385), .B(n10384), .ZN(
        P2_U3203) );
  INV_X1 U13008 ( .A(n10387), .ZN(n10397) );
  INV_X1 U13009 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15011) );
  INV_X1 U13010 ( .A(n12342), .ZN(n10389) );
  NAND3_X1 U13011 ( .A1(n10389), .A2(n10388), .A3(n11593), .ZN(n10390) );
  NAND2_X1 U13012 ( .A1(n10392), .A2(n11730), .ZN(n10396) );
  OAI22_X1 U13013 ( .A1(n11744), .A2(n7267), .B1(n10402), .B2(n11733), .ZN(
        n10394) );
  AOI21_X1 U13014 ( .B1(n11746), .B2(n10393), .A(n10394), .ZN(n10395) );
  OAI211_X1 U13015 ( .C1(n10397), .C2(n15011), .A(n10396), .B(n10395), .ZN(
        P3_U3162) );
  INV_X1 U13016 ( .A(n10398), .ZN(n10411) );
  INV_X1 U13017 ( .A(n13671), .ZN(n14474) );
  OAI222_X1 U13018 ( .A1(n14047), .A2(n15334), .B1(n14043), .B2(n10411), .C1(
        n14474), .C2(P1_U3086), .ZN(P1_U3338) );
  OAI211_X1 U13019 ( .C1(n10401), .C2(n10400), .A(n10399), .B(n11730), .ZN(
        n10406) );
  OAI22_X1 U13020 ( .A1(n11744), .A2(n10402), .B1(n11737), .B2(n14989), .ZN(
        n10403) );
  AOI211_X1 U13021 ( .C1(n11740), .C2(n14978), .A(n10404), .B(n10403), .ZN(
        n10405) );
  OAI211_X1 U13022 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n10407), .A(n10406), .B(
        n10405), .ZN(P3_U3158) );
  INV_X1 U13023 ( .A(n10408), .ZN(n10409) );
  OAI222_X1 U13024 ( .A1(P3_U3151), .A2(n11801), .B1(n12417), .B2(n10410), 
        .C1(n14154), .C2(n10409), .ZN(P3_U3274) );
  OAI222_X1 U13025 ( .A1(n13160), .A2(n10412), .B1(n6894), .B2(P2_U3088), .C1(
        n13178), .C2(n10411), .ZN(P2_U3310) );
  NAND2_X1 U13026 ( .A1(n10419), .A2(n6589), .ZN(n10413) );
  NAND2_X1 U13027 ( .A1(n10527), .A2(n12529), .ZN(n10526) );
  NAND2_X1 U13028 ( .A1(n12510), .A2(n12511), .ZN(n10415) );
  INV_X1 U13029 ( .A(n12730), .ZN(n10416) );
  NAND2_X1 U13030 ( .A1(n10417), .A2(n10416), .ZN(n10435) );
  OAI21_X1 U13031 ( .B1(n10417), .B2(n10416), .A(n10435), .ZN(n10418) );
  AOI222_X1 U13032 ( .A1(n13026), .A2(n10418), .B1(n12799), .B2(n13030), .C1(
        n12801), .C2(n13029), .ZN(n14770) );
  MUX2_X1 U13033 ( .A(n9566), .B(n14770), .S(n12979), .Z(n10430) );
  NAND2_X1 U13034 ( .A1(n10419), .A2(n14757), .ZN(n10420) );
  NAND2_X1 U13035 ( .A1(n10421), .A2(n10420), .ZN(n10530) );
  INV_X1 U13036 ( .A(n12529), .ZN(n12731) );
  NAND2_X1 U13037 ( .A1(n12510), .A2(n14763), .ZN(n10422) );
  OAI21_X1 U13038 ( .B1(n10423), .B2(n12730), .A(n10432), .ZN(n14773) );
  NAND2_X1 U13039 ( .A1(n9731), .A2(n10424), .ZN(n10425) );
  NAND2_X1 U13040 ( .A1(n10533), .A2(n14769), .ZN(n10438) );
  OAI211_X1 U13041 ( .C1(n10533), .C2(n14769), .A(n10438), .B(n12913), .ZN(
        n14768) );
  NOR2_X1 U13042 ( .A1(n14768), .A2(n13047), .ZN(n10428) );
  OAI22_X1 U13043 ( .A1(n13018), .A2(n14769), .B1(n13041), .B2(n10426), .ZN(
        n10427) );
  AOI211_X1 U13044 ( .C1(n14773), .C2(n13049), .A(n10428), .B(n10427), .ZN(
        n10429) );
  NAND2_X1 U13045 ( .A1(n10430), .A2(n10429), .ZN(P2_U3261) );
  NAND2_X1 U13046 ( .A1(n10433), .A2(n14769), .ZN(n10431) );
  XNOR2_X1 U13047 ( .A(n12799), .B(n12545), .ZN(n12733) );
  XNOR2_X1 U13048 ( .A(n10499), .B(n12733), .ZN(n14777) );
  NAND2_X1 U13049 ( .A1(n10433), .A2(n12536), .ZN(n10434) );
  NAND2_X1 U13050 ( .A1(n10435), .A2(n10434), .ZN(n10503) );
  XNOR2_X1 U13051 ( .A(n10503), .B(n12733), .ZN(n10437) );
  AOI21_X1 U13052 ( .B1(n10437), .B2(n13026), .A(n10436), .ZN(n14775) );
  MUX2_X1 U13053 ( .A(n6904), .B(n14775), .S(n12979), .Z(n10444) );
  INV_X1 U13054 ( .A(n10438), .ZN(n10439) );
  INV_X1 U13055 ( .A(n12545), .ZN(n14776) );
  OAI211_X1 U13056 ( .C1(n10439), .C2(n14776), .A(n12913), .B(n10509), .ZN(
        n14774) );
  INV_X1 U13057 ( .A(n14774), .ZN(n10442) );
  OAI22_X1 U13058 ( .A1(n13018), .A2(n14776), .B1(n10440), .B2(n13041), .ZN(
        n10441) );
  AOI21_X1 U13059 ( .B1(n13023), .B2(n10442), .A(n10441), .ZN(n10443) );
  OAI211_X1 U13060 ( .C1(n13002), .C2(n14777), .A(n10444), .B(n10443), .ZN(
        P2_U3260) );
  INV_X1 U13061 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n15203) );
  NAND2_X1 U13062 ( .A1(n10445), .A2(P3_U3897), .ZN(n10446) );
  OAI21_X1 U13063 ( .B1(P3_U3897), .B2(n15203), .A(n10446), .ZN(P3_U3517) );
  NAND2_X1 U13064 ( .A1(n14353), .A2(n10447), .ZN(n10448) );
  OAI211_X1 U13065 ( .C1(n14369), .C2(n10490), .A(n10449), .B(n10448), .ZN(
        n10457) );
  INV_X1 U13066 ( .A(n10450), .ZN(n10452) );
  NAND2_X1 U13067 ( .A1(n10452), .A2(n10451), .ZN(n10453) );
  XNOR2_X1 U13068 ( .A(n10454), .B(n10453), .ZN(n10455) );
  NOR2_X1 U13069 ( .A1(n10455), .A2(n13286), .ZN(n10456) );
  AOI211_X1 U13070 ( .C1(n13330), .C2(n9693), .A(n10457), .B(n10456), .ZN(
        n10458) );
  INV_X1 U13071 ( .A(n10458), .ZN(P1_U3239) );
  XNOR2_X1 U13072 ( .A(n10459), .B(n13493), .ZN(n14547) );
  NAND2_X1 U13073 ( .A1(n13493), .A2(n13542), .ZN(n10461) );
  OAI21_X1 U13074 ( .B1(n14543), .B2(n14526), .A(n10476), .ZN(n10465) );
  MUX2_X1 U13075 ( .A(n10461), .B(n10460), .S(n10462), .Z(n10464) );
  OAI21_X1 U13076 ( .B1(n10462), .B2(n13542), .A(n14505), .ZN(n10463) );
  AOI22_X1 U13077 ( .A1(n14557), .A2(n14547), .B1(n10464), .B2(n10463), .ZN(
        n14544) );
  OR2_X1 U13078 ( .A1(n10465), .A2(n13884), .ZN(n10467) );
  NAND2_X1 U13079 ( .A1(n10467), .A2(n10466), .ZN(n14541) );
  OAI22_X1 U13080 ( .A1(n14536), .A2(n10468), .B1(n13575), .B2(n14508), .ZN(
        n10470) );
  NOR2_X1 U13081 ( .A1(n14376), .A2(n14543), .ZN(n10469) );
  AOI211_X1 U13082 ( .C1(n14517), .C2(n14541), .A(n10470), .B(n10469), .ZN(
        n10472) );
  INV_X1 U13083 ( .A(n13877), .ZN(n14518) );
  NAND2_X1 U13084 ( .A1(n14518), .A2(n14547), .ZN(n10471) );
  OAI211_X1 U13085 ( .C1(n14521), .C2(n14544), .A(n10472), .B(n10471), .ZN(
        P1_U3292) );
  XNOR2_X1 U13086 ( .A(n10473), .B(n10484), .ZN(n10475) );
  AOI21_X1 U13087 ( .B1(n10475), .B2(n14585), .A(n10474), .ZN(n14552) );
  NAND2_X1 U13088 ( .A1(n10476), .A2(n14550), .ZN(n10477) );
  NAND2_X1 U13089 ( .A1(n10477), .A2(n14513), .ZN(n10478) );
  NOR2_X1 U13090 ( .A1(n14515), .A2(n10478), .ZN(n14548) );
  OAI22_X1 U13091 ( .A1(n14536), .A2(n10479), .B1(n13594), .B2(n14508), .ZN(
        n10482) );
  NOR2_X1 U13092 ( .A1(n14376), .A2(n10480), .ZN(n10481) );
  AOI211_X1 U13093 ( .C1(n14548), .C2(n14517), .A(n10482), .B(n10481), .ZN(
        n10486) );
  OAI21_X1 U13094 ( .B1(n14521), .B2(n11340), .A(n13877), .ZN(n13775) );
  XNOR2_X1 U13095 ( .A(n10484), .B(n10483), .ZN(n14554) );
  INV_X1 U13096 ( .A(n14554), .ZN(n14556) );
  NAND2_X1 U13097 ( .A1(n13775), .A2(n14556), .ZN(n10485) );
  OAI211_X1 U13098 ( .C1(n14521), .C2(n14552), .A(n10486), .B(n10485), .ZN(
        P1_U3291) );
  INV_X1 U13099 ( .A(n10487), .ZN(n10497) );
  NAND2_X1 U13100 ( .A1(n10488), .A2(n14536), .ZN(n10496) );
  NOR2_X1 U13101 ( .A1(n14376), .A2(n10489), .ZN(n10493) );
  INV_X1 U13102 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10491) );
  OAI22_X1 U13103 ( .A1(n14536), .A2(n10491), .B1(n10490), .B2(n14508), .ZN(
        n10492) );
  AOI211_X1 U13104 ( .C1(n10494), .C2(n14517), .A(n10493), .B(n10492), .ZN(
        n10495) );
  OAI211_X1 U13105 ( .C1(n10497), .C2(n13877), .A(n10496), .B(n10495), .ZN(
        P1_U3287) );
  NAND2_X1 U13106 ( .A1(n12799), .A2(n12545), .ZN(n10498) );
  INV_X1 U13107 ( .A(n12799), .ZN(n10504) );
  NAND2_X1 U13108 ( .A1(n10504), .A2(n14776), .ZN(n10500) );
  NAND2_X1 U13109 ( .A1(n10501), .A2(n10500), .ZN(n10597) );
  XNOR2_X1 U13110 ( .A(n12549), .B(n12798), .ZN(n12734) );
  XNOR2_X1 U13111 ( .A(n10597), .B(n12734), .ZN(n14780) );
  NAND2_X1 U13112 ( .A1(n14776), .A2(n12799), .ZN(n10502) );
  NAND2_X1 U13113 ( .A1(n10503), .A2(n10502), .ZN(n10506) );
  NAND2_X1 U13114 ( .A1(n10504), .A2(n12545), .ZN(n10505) );
  INV_X1 U13115 ( .A(n12734), .ZN(n10596) );
  XNOR2_X1 U13116 ( .A(n10604), .B(n10596), .ZN(n10508) );
  INV_X1 U13117 ( .A(n13026), .ZN(n12977) );
  OAI21_X1 U13118 ( .B1(n10508), .B2(n12977), .A(n10507), .ZN(n14784) );
  NAND2_X1 U13119 ( .A1(n14784), .A2(n12979), .ZN(n10514) );
  AOI211_X1 U13120 ( .C1(n12549), .C2(n10509), .A(n8877), .B(n10635), .ZN(
        n14783) );
  INV_X1 U13121 ( .A(n13041), .ZN(n13015) );
  AOI22_X1 U13122 ( .A1(n13051), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n10510), 
        .B2(n13015), .ZN(n10511) );
  OAI21_X1 U13123 ( .B1(n13018), .B2(n14781), .A(n10511), .ZN(n10512) );
  AOI21_X1 U13124 ( .B1(n14783), .B2(n13023), .A(n10512), .ZN(n10513) );
  OAI211_X1 U13125 ( .C1(n13002), .C2(n14780), .A(n10514), .B(n10513), .ZN(
        P2_U3259) );
  INV_X1 U13126 ( .A(n10515), .ZN(n10517) );
  OAI22_X1 U13127 ( .A1(n11966), .A2(P3_U3151), .B1(SI_22_), .B2(n12417), .ZN(
        n10516) );
  AOI21_X1 U13128 ( .B1(n10517), .B2(n14162), .A(n10516), .ZN(P3_U3273) );
  AOI21_X1 U13129 ( .B1(n10519), .B2(n6584), .A(n10518), .ZN(n10525) );
  OAI22_X1 U13130 ( .A1(n11744), .A2(n10520), .B1(n11737), .B2(n10589), .ZN(
        n10521) );
  AOI211_X1 U13131 ( .C1(n11740), .C2(n14965), .A(n10522), .B(n10521), .ZN(
        n10524) );
  NAND2_X1 U13132 ( .A1(n11741), .A2(n10590), .ZN(n10523) );
  OAI211_X1 U13133 ( .C1(n10525), .C2(n11748), .A(n10524), .B(n10523), .ZN(
        P3_U3170) );
  OAI21_X1 U13134 ( .B1(n10527), .B2(n12529), .A(n10526), .ZN(n10528) );
  AOI222_X1 U13135 ( .A1(n13026), .A2(n10528), .B1(n12800), .B2(n13030), .C1(
        n12802), .C2(n13029), .ZN(n14764) );
  OAI21_X1 U13136 ( .B1(n10530), .B2(n12731), .A(n10529), .ZN(n14767) );
  NAND2_X1 U13137 ( .A1(n10531), .A2(n12511), .ZN(n10532) );
  NAND2_X1 U13138 ( .A1(n10532), .A2(n12913), .ZN(n10534) );
  OR2_X1 U13139 ( .A1(n10534), .A2(n10533), .ZN(n14762) );
  AOI22_X1 U13140 ( .A1(n13051), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n13015), 
        .B2(n10535), .ZN(n10537) );
  NAND2_X1 U13141 ( .A1(n13044), .A2(n12511), .ZN(n10536) );
  OAI211_X1 U13142 ( .C1(n14762), .C2(n13047), .A(n10537), .B(n10536), .ZN(
        n10538) );
  AOI21_X1 U13143 ( .B1(n14767), .B2(n13049), .A(n10538), .ZN(n10539) );
  OAI21_X1 U13144 ( .B1(n14764), .B2(n13051), .A(n10539), .ZN(P2_U3262) );
  NAND2_X1 U13145 ( .A1(n11981), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10540) );
  OAI21_X1 U13146 ( .B1(n12093), .B2(n11981), .A(n10540), .ZN(P3_U3519) );
  OAI21_X1 U13147 ( .B1(n10543), .B2(n10542), .A(n10541), .ZN(n10556) );
  AND2_X1 U13148 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11723) );
  AOI21_X1 U13149 ( .B1(n14860), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11723), .ZN(
        n10549) );
  OAI21_X1 U13150 ( .B1(n10546), .B2(n10545), .A(n10544), .ZN(n10547) );
  NAND2_X1 U13151 ( .A1(n14192), .A2(n10547), .ZN(n10548) );
  OAI211_X1 U13152 ( .C1(n14939), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10555) );
  XOR2_X1 U13153 ( .A(n10552), .B(n10551), .Z(n10553) );
  NOR2_X1 U13154 ( .A1(n10553), .A2(n14933), .ZN(n10554) );
  AOI211_X1 U13155 ( .C1(n14929), .C2(n10556), .A(n10555), .B(n10554), .ZN(
        n10557) );
  INV_X1 U13156 ( .A(n10557), .ZN(P3_U3188) );
  XNOR2_X1 U13157 ( .A(n10558), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U13158 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10559), .ZN(n11678) );
  AOI21_X1 U13159 ( .B1(n14860), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11678), .ZN(
        n10563) );
  XNOR2_X1 U13160 ( .A(n10560), .B(n10317), .ZN(n10561) );
  NAND2_X1 U13161 ( .A1(n14192), .A2(n10561), .ZN(n10562) );
  OAI211_X1 U13162 ( .C1(n14939), .C2(n10564), .A(n10563), .B(n10562), .ZN(
        n10569) );
  XOR2_X1 U13163 ( .A(n10566), .B(n10565), .Z(n10567) );
  NOR2_X1 U13164 ( .A1(n10567), .A2(n14933), .ZN(n10568) );
  AOI211_X1 U13165 ( .C1(n14929), .C2(n10570), .A(n10569), .B(n10568), .ZN(
        n10571) );
  INV_X1 U13166 ( .A(n10571), .ZN(P3_U3187) );
  XNOR2_X1 U13167 ( .A(n11779), .B(n10572), .ZN(n10587) );
  AOI22_X1 U13168 ( .A1(n14977), .A2(n14965), .B1(n12329), .B2(n14980), .ZN(
        n10576) );
  OAI211_X1 U13169 ( .C1(n10574), .C2(n11779), .A(n10573), .B(n14982), .ZN(
        n10575) );
  OAI211_X1 U13170 ( .C1(n10587), .C2(n15038), .A(n10576), .B(n10575), .ZN(
        n15025) );
  INV_X1 U13171 ( .A(n15025), .ZN(n10595) );
  INV_X1 U13172 ( .A(n10577), .ZN(n10582) );
  NAND2_X1 U13173 ( .A1(n11911), .A2(n10578), .ZN(n10579) );
  NAND2_X1 U13174 ( .A1(n10581), .A2(n10579), .ZN(n10580) );
  OAI21_X1 U13175 ( .B1(n10582), .B2(n10581), .A(n10580), .ZN(n10583) );
  INV_X1 U13176 ( .A(n10583), .ZN(n10584) );
  INV_X1 U13177 ( .A(n10587), .ZN(n15027) );
  AND2_X1 U13178 ( .A1(n14999), .A2(n11772), .ZN(n15003) );
  NAND2_X1 U13179 ( .A1(n14995), .A2(n15003), .ZN(n15013) );
  INV_X1 U13180 ( .A(n15013), .ZN(n14971) );
  INV_X1 U13181 ( .A(n14268), .ZN(n14992) );
  NOR2_X1 U13182 ( .A1(n10589), .A2(n14988), .ZN(n15026) );
  AOI22_X1 U13183 ( .A1(n14992), .A2(n15026), .B1(n14991), .B2(n10590), .ZN(
        n10591) );
  OAI21_X1 U13184 ( .B1(n10592), .B2(n14995), .A(n10591), .ZN(n10593) );
  AOI21_X1 U13185 ( .B1(n15027), .B2(n14971), .A(n10593), .ZN(n10594) );
  OAI21_X1 U13186 ( .B1(n10595), .B2(n15018), .A(n10594), .ZN(P3_U3229) );
  NAND2_X1 U13187 ( .A1(n10597), .A2(n10596), .ZN(n10599) );
  OR2_X1 U13188 ( .A1(n12798), .A2(n12549), .ZN(n10598) );
  NAND2_X1 U13189 ( .A1(n10599), .A2(n10598), .ZN(n10634) );
  XNOR2_X1 U13190 ( .A(n12558), .B(n12797), .ZN(n12735) );
  INV_X1 U13191 ( .A(n12735), .ZN(n10633) );
  OR2_X1 U13192 ( .A1(n12558), .A2(n12797), .ZN(n10600) );
  XNOR2_X1 U13193 ( .A(n12561), .B(n10686), .ZN(n12737) );
  INV_X1 U13194 ( .A(n12737), .ZN(n10601) );
  NAND2_X1 U13195 ( .A1(n10602), .A2(n10601), .ZN(n10603) );
  NAND2_X1 U13196 ( .A1(n10696), .A2(n10603), .ZN(n14795) );
  AOI22_X1 U13197 ( .A1(n13029), .A2(n12797), .B1(n12794), .B2(n13030), .ZN(
        n10612) );
  NAND2_X1 U13198 ( .A1(n12549), .A2(n10605), .ZN(n10606) );
  INV_X1 U13199 ( .A(n12797), .ZN(n10608) );
  AND2_X1 U13200 ( .A1(n12558), .A2(n10608), .ZN(n10609) );
  XNOR2_X1 U13201 ( .A(n10688), .B(n12737), .ZN(n10610) );
  NAND2_X1 U13202 ( .A1(n10610), .A2(n13026), .ZN(n10611) );
  OAI211_X1 U13203 ( .C1(n14795), .C2(n9731), .A(n10612), .B(n10611), .ZN(
        n14799) );
  NAND2_X1 U13204 ( .A1(n14799), .A2(n12979), .ZN(n10617) );
  OAI22_X1 U13205 ( .A1(n12979), .A2(n10613), .B1(n12449), .B2(n13041), .ZN(
        n10615) );
  AND2_X1 U13206 ( .A1(n10635), .A2(n14790), .ZN(n10636) );
  INV_X1 U13207 ( .A(n12561), .ZN(n14798) );
  NAND2_X1 U13208 ( .A1(n10636), .A2(n14798), .ZN(n10699) );
  OAI211_X1 U13209 ( .C1(n10636), .C2(n14798), .A(n12913), .B(n10699), .ZN(
        n14796) );
  NOR2_X1 U13210 ( .A1(n14796), .A2(n13047), .ZN(n10614) );
  AOI211_X1 U13211 ( .C1(n13044), .C2(n12561), .A(n10615), .B(n10614), .ZN(
        n10616) );
  OAI211_X1 U13212 ( .C1(n14795), .C2(n13020), .A(n10617), .B(n10616), .ZN(
        P2_U3257) );
  XNOR2_X1 U13213 ( .A(n10618), .B(n8313), .ZN(n15028) );
  NAND2_X1 U13214 ( .A1(n10620), .A2(n11825), .ZN(n10621) );
  NAND2_X1 U13215 ( .A1(n10619), .A2(n10621), .ZN(n10622) );
  NAND2_X1 U13216 ( .A1(n10622), .A2(n14982), .ZN(n10624) );
  AOI22_X1 U13217 ( .A1(n14980), .A2(n14978), .B1(n11980), .B2(n14977), .ZN(
        n10623) );
  OAI211_X1 U13218 ( .C1(n15028), .C2(n15038), .A(n10624), .B(n10623), .ZN(
        n15029) );
  MUX2_X1 U13219 ( .A(n15029), .B(P3_REG2_REG_5__SCAN_IN), .S(n15018), .Z(
        n10625) );
  INV_X1 U13220 ( .A(n10625), .ZN(n10628) );
  NOR2_X1 U13221 ( .A1(n10626), .A2(n14988), .ZN(n15030) );
  AOI22_X1 U13222 ( .A1(n14992), .A2(n15030), .B1(n14991), .B2(n11680), .ZN(
        n10627) );
  OAI211_X1 U13223 ( .C1(n15028), .C2(n15013), .A(n10628), .B(n10627), .ZN(
        P3_U3228) );
  XNOR2_X1 U13224 ( .A(n10629), .B(n12735), .ZN(n10630) );
  NAND2_X1 U13225 ( .A1(n10630), .A2(n13026), .ZN(n10632) );
  NAND2_X1 U13226 ( .A1(n10632), .A2(n10631), .ZN(n14792) );
  INV_X1 U13227 ( .A(n14792), .ZN(n10643) );
  INV_X2 U13228 ( .A(n12979), .ZN(n13051) );
  XNOR2_X1 U13229 ( .A(n10634), .B(n10633), .ZN(n14788) );
  OAI21_X1 U13230 ( .B1(n10635), .B2(n14790), .A(n12913), .ZN(n10637) );
  OR2_X1 U13231 ( .A1(n10637), .A2(n10636), .ZN(n14789) );
  AOI22_X1 U13232 ( .A1(n13051), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n10638), 
        .B2(n13015), .ZN(n10640) );
  NAND2_X1 U13233 ( .A1(n13044), .A2(n12558), .ZN(n10639) );
  OAI211_X1 U13234 ( .C1(n14789), .C2(n13047), .A(n10640), .B(n10639), .ZN(
        n10641) );
  AOI21_X1 U13235 ( .B1(n14788), .B2(n13049), .A(n10641), .ZN(n10642) );
  OAI21_X1 U13236 ( .B1(n10643), .B2(n13051), .A(n10642), .ZN(P2_U3258) );
  INV_X1 U13237 ( .A(n13775), .ZN(n10657) );
  OAI21_X1 U13238 ( .B1(n10645), .B2(n13503), .A(n10644), .ZN(n10717) );
  INV_X1 U13239 ( .A(n10717), .ZN(n10656) );
  OAI21_X1 U13240 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(n10651) );
  NAND2_X1 U13241 ( .A1(n13565), .A2(n13262), .ZN(n10650) );
  NAND2_X1 U13242 ( .A1(n13567), .A2(n13864), .ZN(n10649) );
  NAND2_X1 U13243 ( .A1(n10650), .A2(n10649), .ZN(n11039) );
  AOI21_X1 U13244 ( .B1(n10651), .B2(n14585), .A(n11039), .ZN(n10714) );
  MUX2_X1 U13245 ( .A(n10714), .B(n9815), .S(n14521), .Z(n10655) );
  AOI211_X1 U13246 ( .C1(n13345), .C2(n6608), .A(n13884), .B(n10727), .ZN(
        n10716) );
  INV_X1 U13247 ( .A(n13345), .ZN(n10652) );
  OAI22_X1 U13248 ( .A1(n10652), .A2(n14376), .B1(n14508), .B2(n11042), .ZN(
        n10653) );
  AOI21_X1 U13249 ( .B1(n10716), .B2(n14517), .A(n10653), .ZN(n10654) );
  OAI211_X1 U13250 ( .C1(n10657), .C2(n10656), .A(n10655), .B(n10654), .ZN(
        P1_U3284) );
  INV_X1 U13251 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15302) );
  INV_X1 U13252 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U13253 ( .A1(n10658), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10660) );
  NAND2_X1 U13254 ( .A1(n8264), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10659) );
  OAI211_X1 U13255 ( .C1(n10662), .C2(n10661), .A(n10660), .B(n10659), .ZN(
        n10663) );
  INV_X1 U13256 ( .A(n10663), .ZN(n10664) );
  NAND2_X1 U13257 ( .A1(n10665), .A2(n10664), .ZN(n12065) );
  NAND2_X1 U13258 ( .A1(n12065), .A2(P3_U3897), .ZN(n10666) );
  OAI21_X1 U13259 ( .B1(P3_U3897), .B2(n15302), .A(n10666), .ZN(P3_U3522) );
  OAI22_X1 U13260 ( .A1(n10669), .A2(n10668), .B1(n10667), .B2(n10675), .ZN(
        n10671) );
  MUX2_X1 U13261 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n6590), .Z(n12021) );
  XNOR2_X1 U13262 ( .A(n12021), .B(n11983), .ZN(n10670) );
  NAND2_X1 U13263 ( .A1(n10671), .A2(n10670), .ZN(n12022) );
  OAI21_X1 U13264 ( .B1(n10671), .B2(n10670), .A(n12022), .ZN(n10672) );
  INV_X1 U13265 ( .A(n14933), .ZN(n14893) );
  NAND2_X1 U13266 ( .A1(n10672), .A2(n14893), .ZN(n10685) );
  XOR2_X1 U13267 ( .A(n12020), .B(n11982), .Z(n11984) );
  XOR2_X1 U13268 ( .A(P3_REG2_REG_9__SCAN_IN), .B(n11984), .Z(n10683) );
  XNOR2_X1 U13269 ( .A(n11983), .B(n11998), .ZN(n10678) );
  NAND2_X1 U13270 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n10678), .ZN(n11999) );
  OAI21_X1 U13271 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n10678), .A(n11999), .ZN(
        n10679) );
  NAND2_X1 U13272 ( .A1(n10679), .A2(n14929), .ZN(n10681) );
  NOR2_X1 U13273 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15364), .ZN(n11128) );
  AOI21_X1 U13274 ( .B1(n14860), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11128), .ZN(
        n10680) );
  OAI211_X1 U13275 ( .C1(n14939), .C2(n12020), .A(n10681), .B(n10680), .ZN(
        n10682) );
  AOI21_X1 U13276 ( .B1(n14192), .B2(n10683), .A(n10682), .ZN(n10684) );
  NAND2_X1 U13277 ( .A1(n10685), .A2(n10684), .ZN(P3_U3191) );
  NOR2_X1 U13278 ( .A1(n12561), .A2(n10686), .ZN(n10687) );
  INV_X1 U13279 ( .A(n12794), .ZN(n10755) );
  XNOR2_X1 U13280 ( .A(n14803), .B(n10755), .ZN(n12738) );
  INV_X1 U13281 ( .A(n12738), .ZN(n10689) );
  NAND2_X1 U13282 ( .A1(n10691), .A2(n12738), .ZN(n10692) );
  NAND3_X1 U13283 ( .A1(n10757), .A2(n13026), .A3(n10692), .ZN(n10694) );
  NAND2_X1 U13284 ( .A1(n10694), .A2(n10693), .ZN(n14807) );
  INV_X1 U13285 ( .A(n14807), .ZN(n10707) );
  NAND2_X1 U13286 ( .A1(n12561), .A2(n12796), .ZN(n10695) );
  NAND2_X1 U13287 ( .A1(n10696), .A2(n10695), .ZN(n10697) );
  NAND2_X1 U13288 ( .A1(n10697), .A2(n12738), .ZN(n10764) );
  OR2_X1 U13289 ( .A1(n10697), .A2(n12738), .ZN(n10698) );
  NAND2_X1 U13290 ( .A1(n10764), .A2(n10698), .ZN(n14806) );
  INV_X1 U13291 ( .A(n14806), .ZN(n10705) );
  AOI21_X1 U13292 ( .B1(n10699), .B2(n14803), .A(n9183), .ZN(n10700) );
  NAND2_X1 U13293 ( .A1(n10700), .A2(n10767), .ZN(n14804) );
  OAI22_X1 U13294 ( .A1(n12979), .A2(n9798), .B1(n10701), .B2(n13041), .ZN(
        n10702) );
  AOI21_X1 U13295 ( .B1(n14803), .B2(n13044), .A(n10702), .ZN(n10703) );
  OAI21_X1 U13296 ( .B1(n14804), .B2(n13047), .A(n10703), .ZN(n10704) );
  AOI21_X1 U13297 ( .B1(n10705), .B2(n13049), .A(n10704), .ZN(n10706) );
  OAI21_X1 U13298 ( .B1(n10707), .B2(n13051), .A(n10706), .ZN(P2_U3256) );
  NAND2_X1 U13299 ( .A1(n10708), .A2(n14162), .ZN(n10709) );
  OAI211_X1 U13300 ( .C1(n15288), .C2(n12417), .A(n10709), .B(n11968), .ZN(
        P3_U3272) );
  INV_X1 U13301 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15212) );
  INV_X1 U13302 ( .A(n11766), .ZN(n11770) );
  NAND2_X1 U13303 ( .A1(n11770), .A2(P3_U3897), .ZN(n10710) );
  OAI21_X1 U13304 ( .B1(P3_U3897), .B2(n15212), .A(n10710), .ZN(P3_U3521) );
  INV_X1 U13305 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n15179) );
  INV_X1 U13306 ( .A(n12082), .ZN(n10711) );
  NAND2_X1 U13307 ( .A1(n10711), .A2(n11973), .ZN(n10712) );
  OAI21_X1 U13308 ( .B1(P3_U3897), .B2(n15179), .A(n10712), .ZN(P3_U3520) );
  INV_X1 U13309 ( .A(n14718), .ZN(n12835) );
  OAI222_X1 U13310 ( .A1(n13178), .A2(n10723), .B1(n12835), .B2(P2_U3088), 
        .C1(n10713), .C2(n13160), .ZN(P2_U3309) );
  INV_X1 U13311 ( .A(n10714), .ZN(n10715) );
  AOI211_X1 U13312 ( .C1(n14590), .C2(n10717), .A(n10716), .B(n10715), .ZN(
        n10722) );
  AOI22_X1 U13313 ( .A1(n13345), .A2(n13969), .B1(n14598), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n10718) );
  OAI21_X1 U13314 ( .B1(n10722), .B2(n14598), .A(n10718), .ZN(P1_U3537) );
  INV_X1 U13315 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10719) );
  NOR2_X1 U13316 ( .A1(n8150), .A2(n10719), .ZN(n10720) );
  AOI21_X1 U13317 ( .B1(n14023), .B2(n13345), .A(n10720), .ZN(n10721) );
  OAI21_X1 U13318 ( .B1(n10722), .B2(n14577), .A(n10721), .ZN(P1_U3486) );
  OAI222_X1 U13319 ( .A1(n14047), .A2(n10724), .B1(n14043), .B2(n10723), .C1(
        n14491), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13320 ( .A(n13895), .ZN(n14533) );
  OAI21_X1 U13321 ( .B1(n10726), .B2(n13504), .A(n10725), .ZN(n10749) );
  OAI21_X1 U13322 ( .B1(n10727), .B2(n10967), .A(n14513), .ZN(n10728) );
  OR2_X1 U13323 ( .A1(n10728), .A2(n10807), .ZN(n10730) );
  AND2_X1 U13324 ( .A1(n13564), .A2(n13262), .ZN(n10960) );
  INV_X1 U13325 ( .A(n10960), .ZN(n10729) );
  AND2_X1 U13326 ( .A1(n10730), .A2(n10729), .ZN(n10746) );
  NAND2_X1 U13327 ( .A1(n10731), .A2(n13504), .ZN(n10743) );
  NAND3_X1 U13328 ( .A1(n10744), .A2(n14532), .A3(n10743), .ZN(n10735) );
  NAND2_X1 U13329 ( .A1(n13566), .A2(n13864), .ZN(n10745) );
  OAI22_X1 U13330 ( .A1(n14521), .A2(n10745), .B1(n10957), .B2(n14508), .ZN(
        n10733) );
  NOR2_X1 U13331 ( .A1(n10967), .A2(n14376), .ZN(n10732) );
  AOI211_X1 U13332 ( .C1(n14521), .C2(P1_REG2_REG_10__SCAN_IN), .A(n10733), 
        .B(n10732), .ZN(n10734) );
  OAI211_X1 U13333 ( .C1(n10746), .C2(n13888), .A(n10735), .B(n10734), .ZN(
        n10736) );
  AOI21_X1 U13334 ( .B1(n14533), .B2(n10749), .A(n10736), .ZN(n10737) );
  INV_X1 U13335 ( .A(n10737), .ZN(P1_U3283) );
  MUX2_X1 U13336 ( .A(P3_REG2_REG_0__SCAN_IN), .B(n10738), .S(n14995), .Z(
        n10742) );
  INV_X1 U13337 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10739) );
  OAI22_X1 U13338 ( .A1(n12134), .A2(n10740), .B1(n15010), .B2(n10739), .ZN(
        n10741) );
  OR2_X1 U13339 ( .A1(n10742), .A2(n10741), .ZN(P3_U3233) );
  NAND3_X1 U13340 ( .A1(n10744), .A2(n14585), .A3(n10743), .ZN(n10747) );
  NAND3_X1 U13341 ( .A1(n10747), .A2(n10746), .A3(n10745), .ZN(n10748) );
  AOI21_X1 U13342 ( .B1(n14590), .B2(n10749), .A(n10748), .ZN(n10754) );
  AOI22_X1 U13343 ( .A1(n13352), .A2(n13969), .B1(n14598), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n10750) );
  OAI21_X1 U13344 ( .B1(n10754), .B2(n14598), .A(n10750), .ZN(P1_U3538) );
  INV_X1 U13345 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10751) );
  OAI22_X1 U13346 ( .A1(n10967), .A2(n14028), .B1(n8150), .B2(n10751), .ZN(
        n10752) );
  INV_X1 U13347 ( .A(n10752), .ZN(n10753) );
  OAI21_X1 U13348 ( .B1(n10754), .B2(n14577), .A(n10753), .ZN(P1_U3489) );
  OR2_X1 U13349 ( .A1(n14803), .A2(n10755), .ZN(n10756) );
  NAND2_X1 U13350 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  INV_X1 U13351 ( .A(n12793), .ZN(n10842) );
  XNOR2_X1 U13352 ( .A(n14811), .B(n10842), .ZN(n12740) );
  INV_X1 U13353 ( .A(n12740), .ZN(n10758) );
  NAND2_X1 U13354 ( .A1(n10759), .A2(n10758), .ZN(n10844) );
  OAI211_X1 U13355 ( .C1(n10759), .C2(n10758), .A(n10844), .B(n13026), .ZN(
        n10762) );
  NAND2_X1 U13356 ( .A1(n12792), .A2(n13030), .ZN(n10761) );
  NAND2_X1 U13357 ( .A1(n12794), .A2(n13029), .ZN(n10760) );
  AND2_X1 U13358 ( .A1(n10761), .A2(n10760), .ZN(n10880) );
  NAND2_X1 U13359 ( .A1(n10762), .A2(n10880), .ZN(n14815) );
  INV_X1 U13360 ( .A(n14815), .ZN(n10775) );
  NAND2_X1 U13361 ( .A1(n14803), .A2(n12794), .ZN(n10763) );
  NAND2_X1 U13362 ( .A1(n10764), .A2(n10763), .ZN(n10765) );
  NAND2_X1 U13363 ( .A1(n10765), .A2(n12740), .ZN(n10839) );
  OR2_X1 U13364 ( .A1(n10765), .A2(n12740), .ZN(n10766) );
  NAND2_X1 U13365 ( .A1(n10839), .A2(n10766), .ZN(n14814) );
  INV_X1 U13366 ( .A(n14814), .ZN(n10773) );
  AOI21_X1 U13367 ( .B1(n10767), .B2(n14811), .A(n9183), .ZN(n10768) );
  NAND2_X1 U13368 ( .A1(n10768), .A2(n10852), .ZN(n14812) );
  INV_X1 U13369 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10769) );
  OAI22_X1 U13370 ( .A1(n12979), .A2(n10769), .B1(n10876), .B2(n13041), .ZN(
        n10770) );
  AOI21_X1 U13371 ( .B1(n14811), .B2(n13044), .A(n10770), .ZN(n10771) );
  OAI21_X1 U13372 ( .B1(n14812), .B2(n13047), .A(n10771), .ZN(n10772) );
  AOI21_X1 U13373 ( .B1(n10773), .B2(n13049), .A(n10772), .ZN(n10774) );
  OAI21_X1 U13374 ( .B1(n10775), .B2(n13051), .A(n10774), .ZN(P2_U3255) );
  NAND2_X1 U13375 ( .A1(n14995), .A2(n12131), .ZN(n10776) );
  XNOR2_X1 U13376 ( .A(n10777), .B(n10779), .ZN(n15036) );
  OAI211_X1 U13377 ( .C1(n10780), .C2(n10779), .A(n10778), .B(n14982), .ZN(
        n10782) );
  AOI22_X1 U13378 ( .A1(n14980), .A2(n11980), .B1(n11979), .B2(n14977), .ZN(
        n10781) );
  AND2_X1 U13379 ( .A1(n10782), .A2(n10781), .ZN(n15039) );
  MUX2_X1 U13380 ( .A(n15039), .B(n10783), .S(n15018), .Z(n10785) );
  AOI22_X1 U13381 ( .A1(n14253), .A2(n15042), .B1(n14991), .B2(n11610), .ZN(
        n10784) );
  OAI211_X1 U13382 ( .C1(n14269), .C2(n15036), .A(n10785), .B(n10784), .ZN(
        P3_U3226) );
  NAND2_X1 U13383 ( .A1(n14353), .A2(n14579), .ZN(n10786) );
  OAI211_X1 U13384 ( .C1(n14369), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        n10799) );
  AOI22_X1 U13385 ( .A1(n14578), .A2(n11559), .B1(n11558), .B2(n13567), .ZN(
        n10943) );
  NAND2_X1 U13386 ( .A1(n14578), .A2(n11554), .ZN(n10790) );
  NAND2_X1 U13387 ( .A1(n11559), .A2(n13567), .ZN(n10789) );
  NAND2_X1 U13388 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  XNOR2_X1 U13389 ( .A(n10791), .B(n9952), .ZN(n10942) );
  XOR2_X1 U13390 ( .A(n10943), .B(n10942), .Z(n10796) );
  AOI21_X1 U13391 ( .B1(n10796), .B2(n10795), .A(n6701), .ZN(n10797) );
  NOR2_X1 U13392 ( .A1(n10797), .A2(n13286), .ZN(n10798) );
  AOI211_X1 U13393 ( .C1(n14578), .C2(n9693), .A(n10799), .B(n10798), .ZN(
        n10800) );
  INV_X1 U13394 ( .A(n10800), .ZN(P1_U3221) );
  OAI211_X1 U13395 ( .C1(n10802), .C2(n13505), .A(n10801), .B(n14585), .ZN(
        n10806) );
  NAND2_X1 U13396 ( .A1(n13565), .A2(n13864), .ZN(n10804) );
  NAND2_X1 U13397 ( .A1(n13563), .A2(n13262), .ZN(n10803) );
  NAND2_X1 U13398 ( .A1(n10804), .A2(n10803), .ZN(n11062) );
  INV_X1 U13399 ( .A(n11062), .ZN(n10805) );
  NAND2_X1 U13400 ( .A1(n10806), .A2(n10805), .ZN(n10905) );
  INV_X1 U13401 ( .A(n10905), .ZN(n10817) );
  INV_X1 U13402 ( .A(n10807), .ZN(n10809) );
  INV_X1 U13403 ( .A(n10866), .ZN(n10808) );
  AOI211_X1 U13404 ( .C1(n13355), .C2(n10809), .A(n13884), .B(n10808), .ZN(
        n10906) );
  NOR2_X1 U13405 ( .A1(n10909), .A2(n14376), .ZN(n10811) );
  OAI22_X1 U13406 ( .A1(n14536), .A2(n10068), .B1(n11064), .B2(n14508), .ZN(
        n10810) );
  AOI211_X1 U13407 ( .C1(n10906), .C2(n14517), .A(n10811), .B(n10810), .ZN(
        n10816) );
  OAI21_X1 U13408 ( .B1(n10814), .B2(n10813), .A(n10812), .ZN(n10907) );
  NAND2_X1 U13409 ( .A1(n10907), .A2(n14533), .ZN(n10815) );
  OAI211_X1 U13410 ( .C1(n10817), .C2(n14521), .A(n10816), .B(n10815), .ZN(
        P1_U3282) );
  INV_X1 U13411 ( .A(n10818), .ZN(n10881) );
  NOR3_X1 U13412 ( .A1(n10819), .A2(n10842), .A3(n12502), .ZN(n10820) );
  AOI21_X1 U13413 ( .B1(n10881), .B2(n9282), .A(n10820), .ZN(n10829) );
  NAND2_X1 U13414 ( .A1(n14819), .A2(n14328), .ZN(n10825) );
  NAND2_X1 U13415 ( .A1(n12791), .A2(n13030), .ZN(n10822) );
  NAND2_X1 U13416 ( .A1(n12793), .A2(n13029), .ZN(n10821) );
  AND2_X1 U13417 ( .A1(n10822), .A2(n10821), .ZN(n10848) );
  INV_X1 U13418 ( .A(n10848), .ZN(n10823) );
  AOI22_X1 U13419 ( .A1(n14325), .A2(n10823), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10824) );
  OAI211_X1 U13420 ( .C1(n14331), .C2(n10850), .A(n10825), .B(n10824), .ZN(
        n10826) );
  AOI21_X1 U13421 ( .B1(n6715), .B2(n9282), .A(n10826), .ZN(n10827) );
  OAI21_X1 U13422 ( .B1(n10829), .B2(n10828), .A(n10827), .ZN(P2_U3208) );
  OAI222_X1 U13423 ( .A1(n14047), .A2(n10830), .B1(n14043), .B2(n11592), .C1(
        n13477), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13424 ( .A(n10831), .ZN(n10833) );
  OAI222_X1 U13425 ( .A1(n13160), .A2(n10832), .B1(n13178), .B2(n10833), .C1(
        P2_U3088), .C2(n12762), .ZN(P2_U3308) );
  OAI222_X1 U13426 ( .A1(n14047), .A2(n15176), .B1(n14043), .B2(n10833), .C1(
        P1_U3086), .C2(n14523), .ZN(P1_U3336) );
  INV_X1 U13427 ( .A(n10834), .ZN(n10837) );
  OAI222_X1 U13428 ( .A1(n14154), .A2(n10837), .B1(P3_U3151), .B2(n10836), 
        .C1(n10835), .C2(n12417), .ZN(P3_U3270) );
  NAND2_X1 U13429 ( .A1(n14811), .A2(n12793), .ZN(n10838) );
  NAND2_X1 U13430 ( .A1(n10839), .A2(n10838), .ZN(n10840) );
  INV_X1 U13431 ( .A(n12792), .ZN(n10998) );
  XNOR2_X1 U13432 ( .A(n14819), .B(n10998), .ZN(n12742) );
  NAND2_X1 U13433 ( .A1(n10840), .A2(n12742), .ZN(n10997) );
  OR2_X1 U13434 ( .A1(n10840), .A2(n12742), .ZN(n10841) );
  NAND2_X1 U13435 ( .A1(n10997), .A2(n10841), .ZN(n14823) );
  OR2_X1 U13436 ( .A1(n14811), .A2(n10842), .ZN(n10843) );
  NAND2_X1 U13437 ( .A1(n10845), .A2(n12742), .ZN(n10846) );
  NAND2_X1 U13438 ( .A1(n11000), .A2(n10846), .ZN(n10847) );
  NAND2_X1 U13439 ( .A1(n10847), .A2(n13026), .ZN(n10849) );
  NAND2_X1 U13440 ( .A1(n10849), .A2(n10848), .ZN(n14824) );
  NAND2_X1 U13441 ( .A1(n14824), .A2(n12979), .ZN(n10858) );
  OAI22_X1 U13442 ( .A1(n12979), .A2(n10851), .B1(n10850), .B2(n13041), .ZN(
        n10856) );
  INV_X1 U13443 ( .A(n11004), .ZN(n10854) );
  AOI21_X1 U13444 ( .B1(n10852), .B2(n14819), .A(n9183), .ZN(n10853) );
  NAND2_X1 U13445 ( .A1(n10854), .A2(n10853), .ZN(n14820) );
  NOR2_X1 U13446 ( .A1(n14820), .A2(n13047), .ZN(n10855) );
  AOI211_X1 U13447 ( .C1(n13044), .C2(n14819), .A(n10856), .B(n10855), .ZN(
        n10857) );
  OAI211_X1 U13448 ( .C1(n13002), .C2(n14823), .A(n10858), .B(n10857), .ZN(
        P2_U3254) );
  OAI211_X1 U13449 ( .C1(n10860), .C2(n13506), .A(n10859), .B(n14585), .ZN(
        n10864) );
  NAND2_X1 U13450 ( .A1(n13562), .A2(n13262), .ZN(n10862) );
  NAND2_X1 U13451 ( .A1(n13564), .A2(n13864), .ZN(n10861) );
  NAND2_X1 U13452 ( .A1(n10862), .A2(n10861), .ZN(n11143) );
  INV_X1 U13453 ( .A(n11143), .ZN(n10863) );
  NAND2_X1 U13454 ( .A1(n10864), .A2(n10863), .ZN(n11011) );
  INV_X1 U13455 ( .A(n11011), .ZN(n10875) );
  INV_X1 U13456 ( .A(n11074), .ZN(n10865) );
  AOI211_X1 U13457 ( .C1(n13363), .C2(n10866), .A(n13884), .B(n10865), .ZN(
        n11012) );
  NOR2_X1 U13458 ( .A1(n6876), .A2(n14376), .ZN(n10869) );
  OAI22_X1 U13459 ( .A1(n14536), .A2(n10867), .B1(n11141), .B2(n14508), .ZN(
        n10868) );
  AOI211_X1 U13460 ( .C1(n11012), .C2(n14517), .A(n10869), .B(n10868), .ZN(
        n10874) );
  OAI21_X1 U13461 ( .B1(n10872), .B2(n10871), .A(n10870), .ZN(n11013) );
  NAND2_X1 U13462 ( .A1(n11013), .A2(n13775), .ZN(n10873) );
  OAI211_X1 U13463 ( .C1(n10875), .C2(n14521), .A(n10874), .B(n10873), .ZN(
        P1_U3281) );
  INV_X1 U13464 ( .A(n10876), .ZN(n10877) );
  NAND2_X1 U13465 ( .A1(n12489), .A2(n10877), .ZN(n10879) );
  OAI211_X1 U13466 ( .C1(n10880), .C2(n12438), .A(n10879), .B(n10878), .ZN(
        n10885) );
  AOI211_X1 U13467 ( .C1(n10883), .C2(n10882), .A(n14302), .B(n10881), .ZN(
        n10884) );
  AOI211_X1 U13468 ( .C1(n14811), .C2(n14328), .A(n10885), .B(n10884), .ZN(
        n10886) );
  INV_X1 U13469 ( .A(n10886), .ZN(P2_U3189) );
  INV_X1 U13470 ( .A(n14305), .ZN(n11150) );
  OAI22_X1 U13471 ( .A1(n10998), .A2(n13004), .B1(n11150), .B2(n13006), .ZN(
        n11002) );
  AOI22_X1 U13472 ( .A1(n14325), .A2(n11002), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10887) );
  OAI21_X1 U13473 ( .B1(n11083), .B2(n14331), .A(n10887), .ZN(n10892) );
  AOI22_X1 U13474 ( .A1(n10888), .A2(n9282), .B1(n12465), .B2(n12792), .ZN(
        n10890) );
  NOR3_X1 U13475 ( .A1(n6715), .A2(n10890), .A3(n10889), .ZN(n10891) );
  AOI211_X1 U13476 ( .C1(n12589), .C2(n14328), .A(n10892), .B(n10891), .ZN(
        n10893) );
  OAI21_X1 U13477 ( .B1(n14302), .B2(n10894), .A(n10893), .ZN(P2_U3196) );
  XOR2_X1 U13478 ( .A(n10895), .B(n11847), .Z(n10899) );
  OAI211_X1 U13479 ( .C1(n6721), .C2(n8385), .A(n14982), .B(n10896), .ZN(
        n10898) );
  AOI22_X1 U13480 ( .A1(n14980), .A2(n11979), .B1(n14275), .B2(n14977), .ZN(
        n10897) );
  OAI211_X1 U13481 ( .C1(n10899), .C2(n15038), .A(n10898), .B(n10897), .ZN(
        n15047) );
  INV_X1 U13482 ( .A(n15047), .ZN(n10904) );
  INV_X1 U13483 ( .A(n10899), .ZN(n15050) );
  INV_X1 U13484 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10901) );
  NOR2_X1 U13485 ( .A1(n11125), .A2(n14988), .ZN(n15048) );
  AOI22_X1 U13486 ( .A1(n14992), .A2(n15048), .B1(n14991), .B2(n11129), .ZN(
        n10900) );
  OAI21_X1 U13487 ( .B1(n10901), .B2(n14995), .A(n10900), .ZN(n10902) );
  AOI21_X1 U13488 ( .B1(n15050), .B2(n14971), .A(n10902), .ZN(n10903) );
  OAI21_X1 U13489 ( .B1(n10904), .B2(n15018), .A(n10903), .ZN(P3_U3224) );
  AOI211_X1 U13490 ( .C1(n14590), .C2(n10907), .A(n10906), .B(n10905), .ZN(
        n10913) );
  INV_X1 U13491 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10908) );
  OAI22_X1 U13492 ( .A1(n10909), .A2(n14028), .B1(n8150), .B2(n10908), .ZN(
        n10910) );
  INV_X1 U13493 ( .A(n10910), .ZN(n10911) );
  OAI21_X1 U13494 ( .B1(n10913), .B2(n14577), .A(n10911), .ZN(P1_U3492) );
  AOI22_X1 U13495 ( .A1(n13355), .A2(n13969), .B1(n14598), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n10912) );
  OAI21_X1 U13496 ( .B1(n10913), .B2(n14598), .A(n10912), .ZN(P1_U3539) );
  NAND2_X1 U13497 ( .A1(n10929), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U13498 ( .A1(n10915), .A2(n10914), .ZN(n12815) );
  MUX2_X1 U13499 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9039), .S(n12812), .Z(
        n12814) );
  NAND2_X1 U13500 ( .A1(n12815), .A2(n12814), .ZN(n12813) );
  NAND2_X1 U13501 ( .A1(n12812), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10916) );
  NAND2_X1 U13502 ( .A1(n12813), .A2(n10916), .ZN(n14647) );
  OR2_X1 U13503 ( .A1(n10933), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U13504 ( .A1(n10933), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U13505 ( .A1(n10918), .A2(n10917), .ZN(n14646) );
  OR2_X1 U13506 ( .A1(n14665), .A2(n10919), .ZN(n10921) );
  NAND2_X1 U13507 ( .A1(n14665), .A2(n10919), .ZN(n10920) );
  NAND2_X1 U13508 ( .A1(n10921), .A2(n10920), .ZN(n14657) );
  NAND2_X1 U13509 ( .A1(n14658), .A2(n14657), .ZN(n14656) );
  NAND2_X1 U13510 ( .A1(n14665), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10922) );
  NAND2_X1 U13511 ( .A1(n14656), .A2(n10922), .ZN(n10927) );
  OR2_X1 U13512 ( .A1(n12820), .A2(n10923), .ZN(n10925) );
  NAND2_X1 U13513 ( .A1(n12820), .A2(n10923), .ZN(n10924) );
  NAND2_X1 U13514 ( .A1(n10925), .A2(n10924), .ZN(n10926) );
  OAI21_X1 U13515 ( .B1(n10927), .B2(n10926), .A(n14655), .ZN(n10941) );
  MUX2_X1 U13516 ( .A(n10851), .B(P2_REG2_REG_11__SCAN_IN), .S(n12812), .Z(
        n10930) );
  INV_X1 U13517 ( .A(n10930), .ZN(n12807) );
  NOR2_X1 U13518 ( .A1(n14640), .A2(n10931), .ZN(n10932) );
  AOI21_X1 U13519 ( .B1(n10931), .B2(n14640), .A(n10932), .ZN(n14645) );
  OAI21_X1 U13520 ( .B1(n10933), .B2(P2_REG2_REG_12__SCAN_IN), .A(n14643), 
        .ZN(n14661) );
  NOR2_X1 U13521 ( .A1(n14665), .A2(n11033), .ZN(n10934) );
  AOI21_X1 U13522 ( .B1(n14665), .B2(n11033), .A(n10934), .ZN(n14662) );
  NOR2_X1 U13523 ( .A1(n6611), .A2(n11156), .ZN(n12827) );
  AOI211_X1 U13524 ( .C1(n11156), .C2(n6611), .A(n14695), .B(n12827), .ZN(
        n10936) );
  INV_X1 U13525 ( .A(n10936), .ZN(n10940) );
  INV_X1 U13526 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U13527 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14313)
         );
  OAI21_X1 U13528 ( .B1(n14722), .B2(n10937), .A(n14313), .ZN(n10938) );
  AOI21_X1 U13529 ( .B1(n12820), .B2(n14719), .A(n10938), .ZN(n10939) );
  OAI211_X1 U13530 ( .C1(n12819), .C2(n10941), .A(n10940), .B(n10939), .ZN(
        P2_U3228) );
  INV_X1 U13531 ( .A(n10942), .ZN(n10944) );
  NOR2_X1 U13532 ( .A1(n9958), .A2(n10962), .ZN(n10945) );
  AOI21_X1 U13533 ( .B1(n13345), .B2(n11559), .A(n10945), .ZN(n10948) );
  XNOR2_X1 U13534 ( .A(n10947), .B(n10948), .ZN(n11044) );
  AOI22_X1 U13535 ( .A1(n13345), .A2(n11554), .B1(n11559), .B2(n13566), .ZN(
        n10946) );
  XNOR2_X1 U13536 ( .A(n10946), .B(n9952), .ZN(n11043) );
  INV_X1 U13537 ( .A(n10947), .ZN(n10949) );
  NAND2_X1 U13538 ( .A1(n13352), .A2(n11554), .ZN(n10951) );
  NAND2_X1 U13539 ( .A1(n13565), .A2(n11559), .ZN(n10950) );
  NAND2_X1 U13540 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  XNOR2_X1 U13541 ( .A(n10952), .B(n9952), .ZN(n11055) );
  NOR2_X1 U13542 ( .A1(n9958), .A2(n10953), .ZN(n10954) );
  AOI21_X1 U13543 ( .B1(n13352), .B2(n11559), .A(n10954), .ZN(n11056) );
  XNOR2_X1 U13544 ( .A(n11055), .B(n11056), .ZN(n10955) );
  NAND2_X1 U13545 ( .A1(n10956), .A2(n10955), .ZN(n11059) );
  OAI211_X1 U13546 ( .C1(n10956), .C2(n10955), .A(n11059), .B(n14365), .ZN(
        n10966) );
  INV_X1 U13547 ( .A(n10957), .ZN(n10964) );
  INV_X1 U13548 ( .A(n10958), .ZN(n10959) );
  AOI21_X1 U13549 ( .B1(n14353), .B2(n10960), .A(n10959), .ZN(n10961) );
  OAI21_X1 U13550 ( .B1(n13274), .B2(n10962), .A(n10961), .ZN(n10963) );
  AOI21_X1 U13551 ( .B1(n13293), .B2(n10964), .A(n10963), .ZN(n10965) );
  OAI211_X1 U13552 ( .C1(n10967), .C2(n14362), .A(n10966), .B(n10965), .ZN(
        P1_U3217) );
  OAI222_X1 U13553 ( .A1(n13178), .A2(n10970), .B1(n10969), .B2(P2_U3088), 
        .C1(n10968), .C2(n13160), .ZN(P2_U3306) );
  INV_X1 U13554 ( .A(n13450), .ZN(n13484) );
  OAI222_X1 U13555 ( .A1(n14047), .A2(n15292), .B1(n14043), .B2(n10970), .C1(
        n13484), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI211_X1 U13556 ( .C1(n10972), .C2(n11854), .A(n10971), .B(n14982), .ZN(
        n10974) );
  AOI22_X1 U13557 ( .A1(n14977), .A2(n14259), .B1(n14951), .B2(n14980), .ZN(
        n10973) );
  NAND2_X1 U13558 ( .A1(n10974), .A2(n10973), .ZN(n15051) );
  INV_X1 U13559 ( .A(n15051), .ZN(n10980) );
  XNOR2_X1 U13560 ( .A(n10975), .B(n11854), .ZN(n15053) );
  INV_X1 U13561 ( .A(n14269), .ZN(n14281) );
  INV_X1 U13562 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12017) );
  NOR2_X1 U13563 ( .A1(n10976), .A2(n14988), .ZN(n15052) );
  AOI22_X1 U13564 ( .A1(n14992), .A2(n15052), .B1(n14991), .B2(n11628), .ZN(
        n10977) );
  OAI21_X1 U13565 ( .B1(n12017), .B2(n14995), .A(n10977), .ZN(n10978) );
  AOI21_X1 U13566 ( .B1(n15053), .B2(n14281), .A(n10978), .ZN(n10979) );
  OAI21_X1 U13567 ( .B1(n10980), .B2(n15018), .A(n10979), .ZN(P3_U3223) );
  INV_X1 U13568 ( .A(n10981), .ZN(n10982) );
  OAI222_X1 U13569 ( .A1(n10984), .A2(P3_U3151), .B1(n12417), .B2(n10983), 
        .C1(n14154), .C2(n10982), .ZN(P3_U3269) );
  AOI21_X1 U13570 ( .B1(n10986), .B2(n10985), .A(n14302), .ZN(n10988) );
  NAND2_X1 U13571 ( .A1(n10988), .A2(n10987), .ZN(n10995) );
  INV_X1 U13572 ( .A(n11032), .ZN(n10993) );
  NAND2_X1 U13573 ( .A1(n12790), .A2(n13030), .ZN(n10990) );
  NAND2_X1 U13574 ( .A1(n12791), .A2(n13029), .ZN(n10989) );
  AND2_X1 U13575 ( .A1(n10990), .A2(n10989), .ZN(n11024) );
  OAI22_X1 U13576 ( .A1(n12438), .A2(n11024), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10991), .ZN(n10992) );
  AOI21_X1 U13577 ( .B1(n12489), .B2(n10993), .A(n10992), .ZN(n10994) );
  OAI211_X1 U13578 ( .C1(n14340), .C2(n14310), .A(n10995), .B(n10994), .ZN(
        P2_U3206) );
  NAND2_X1 U13579 ( .A1(n14819), .A2(n12792), .ZN(n10996) );
  XNOR2_X1 U13580 ( .A(n12589), .B(n12791), .ZN(n12743) );
  XNOR2_X1 U13581 ( .A(n11027), .B(n7467), .ZN(n11092) );
  NAND2_X1 U13582 ( .A1(n14819), .A2(n10998), .ZN(n10999) );
  AOI21_X1 U13583 ( .B1(n11001), .B2(n7467), .A(n12977), .ZN(n11003) );
  AOI21_X1 U13584 ( .B1(n11003), .B2(n11021), .A(n11002), .ZN(n11087) );
  INV_X1 U13585 ( .A(n12589), .ZN(n11086) );
  OAI21_X1 U13586 ( .B1(n11004), .B2(n11086), .A(n12913), .ZN(n11005) );
  NOR2_X1 U13587 ( .A1(n11005), .A2(n11030), .ZN(n11090) );
  AOI21_X1 U13588 ( .B1(n14818), .B2(n12589), .A(n11090), .ZN(n11006) );
  OAI211_X1 U13589 ( .C1(n13140), .C2(n11092), .A(n11087), .B(n11006), .ZN(
        n11008) );
  NAND2_X1 U13590 ( .A1(n11008), .A2(n14842), .ZN(n11007) );
  OAI21_X1 U13591 ( .B1(n14842), .B2(n9058), .A(n11007), .ZN(P2_U3511) );
  INV_X1 U13592 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13593 ( .A1(n11008), .A2(n14829), .ZN(n11009) );
  OAI21_X1 U13594 ( .B1(n14829), .B2(n11010), .A(n11009), .ZN(P2_U3466) );
  AOI211_X1 U13595 ( .C1(n14590), .C2(n11013), .A(n11012), .B(n11011), .ZN(
        n11018) );
  AOI22_X1 U13596 ( .A1(n13363), .A2(n13969), .B1(n14598), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11014) );
  OAI21_X1 U13597 ( .B1(n11018), .B2(n14598), .A(n11014), .ZN(P1_U3540) );
  INV_X1 U13598 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11015) );
  OAI22_X1 U13599 ( .A1(n6876), .A2(n14028), .B1(n8150), .B2(n11015), .ZN(
        n11016) );
  INV_X1 U13600 ( .A(n11016), .ZN(n11017) );
  OAI21_X1 U13601 ( .B1(n11018), .B2(n14577), .A(n11017), .ZN(P1_U3495) );
  INV_X1 U13602 ( .A(n12791), .ZN(n11019) );
  OR2_X1 U13603 ( .A1(n12589), .A2(n11019), .ZN(n11020) );
  XNOR2_X1 U13604 ( .A(n12594), .B(n14305), .ZN(n12744) );
  INV_X1 U13605 ( .A(n12744), .ZN(n11022) );
  XNOR2_X1 U13606 ( .A(n11149), .B(n11022), .ZN(n11023) );
  NAND2_X1 U13607 ( .A1(n11023), .A2(n13026), .ZN(n11025) );
  NAND2_X1 U13608 ( .A1(n11025), .A2(n11024), .ZN(n14343) );
  INV_X1 U13609 ( .A(n14343), .ZN(n11038) );
  OR2_X1 U13610 ( .A1(n12589), .A2(n12791), .ZN(n11026) );
  NAND2_X1 U13611 ( .A1(n11027), .A2(n11026), .ZN(n11029) );
  NAND2_X1 U13612 ( .A1(n12589), .A2(n12791), .ZN(n11028) );
  NAND2_X1 U13613 ( .A1(n11029), .A2(n11028), .ZN(n11154) );
  XNOR2_X1 U13614 ( .A(n11154), .B(n12744), .ZN(n14338) );
  OAI21_X1 U13615 ( .B1(n11030), .B2(n14340), .A(n12913), .ZN(n11031) );
  OR2_X1 U13616 ( .A1(n11155), .A2(n11031), .ZN(n14339) );
  OAI22_X1 U13617 ( .A1(n12979), .A2(n11033), .B1(n11032), .B2(n13041), .ZN(
        n11034) );
  AOI21_X1 U13618 ( .B1(n12594), .B2(n13044), .A(n11034), .ZN(n11035) );
  OAI21_X1 U13619 ( .B1(n14339), .B2(n13047), .A(n11035), .ZN(n11036) );
  AOI21_X1 U13620 ( .B1(n14338), .B2(n13049), .A(n11036), .ZN(n11037) );
  OAI21_X1 U13621 ( .B1(n11038), .B2(n13051), .A(n11037), .ZN(P2_U3252) );
  NAND2_X1 U13622 ( .A1(n14353), .A2(n11039), .ZN(n11040) );
  OAI211_X1 U13623 ( .C1(n14369), .C2(n11042), .A(n11041), .B(n11040), .ZN(
        n11047) );
  XOR2_X1 U13624 ( .A(n11044), .B(n11043), .Z(n11045) );
  NOR2_X1 U13625 ( .A1(n11045), .A2(n13286), .ZN(n11046) );
  AOI211_X1 U13626 ( .C1(n13345), .C2(n9693), .A(n11047), .B(n11046), .ZN(
        n11048) );
  INV_X1 U13627 ( .A(n11048), .ZN(P1_U3231) );
  INV_X1 U13628 ( .A(n11049), .ZN(n11050) );
  OAI222_X1 U13629 ( .A1(P3_U3151), .A2(n6590), .B1(n12417), .B2(n11051), .C1(
        n14154), .C2(n11050), .ZN(P3_U3268) );
  AOI22_X1 U13630 ( .A1(n13355), .A2(n11559), .B1(n11558), .B2(n13564), .ZN(
        n11134) );
  NAND2_X1 U13631 ( .A1(n13355), .A2(n11554), .ZN(n11053) );
  NAND2_X1 U13632 ( .A1(n11559), .A2(n13564), .ZN(n11052) );
  NAND2_X1 U13633 ( .A1(n11053), .A2(n11052), .ZN(n11054) );
  XNOR2_X1 U13634 ( .A(n11054), .B(n9952), .ZN(n11133) );
  XOR2_X1 U13635 ( .A(n11134), .B(n11133), .Z(n11061) );
  AOI21_X1 U13636 ( .B1(n11061), .B2(n11060), .A(n11136), .ZN(n11067) );
  AOI22_X1 U13637 ( .A1(n14353), .A2(n11062), .B1(P1_REG3_REG_11__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11063) );
  OAI21_X1 U13638 ( .B1(n14369), .B2(n11064), .A(n11063), .ZN(n11065) );
  AOI21_X1 U13639 ( .B1(n13355), .B2(n9693), .A(n11065), .ZN(n11066) );
  OAI21_X1 U13640 ( .B1(n11067), .B2(n13286), .A(n11066), .ZN(P1_U3236) );
  INV_X1 U13641 ( .A(n13252), .ZN(n11072) );
  OAI211_X1 U13642 ( .C1(n13508), .C2(n11068), .A(n11191), .B(n14585), .ZN(
        n11071) );
  NAND2_X1 U13643 ( .A1(n13563), .A2(n13864), .ZN(n11069) );
  OAI21_X1 U13644 ( .B1(n11464), .B2(n13686), .A(n11069), .ZN(n13255) );
  INV_X1 U13645 ( .A(n13255), .ZN(n11070) );
  NAND2_X1 U13646 ( .A1(n11071), .A2(n11070), .ZN(n11109) );
  AOI21_X1 U13647 ( .B1(n11072), .B2(n14528), .A(n11109), .ZN(n11082) );
  INV_X1 U13648 ( .A(n11189), .ZN(n11073) );
  AOI211_X1 U13649 ( .C1(n13366), .C2(n11074), .A(n13884), .B(n11073), .ZN(
        n11110) );
  INV_X1 U13650 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11075) );
  OAI22_X1 U13651 ( .A1(n6875), .A2(n14376), .B1(n11075), .B2(n14536), .ZN(
        n11076) );
  AOI21_X1 U13652 ( .B1(n11110), .B2(n14517), .A(n11076), .ZN(n11081) );
  OAI21_X1 U13653 ( .B1(n11079), .B2(n11078), .A(n11077), .ZN(n11111) );
  NAND2_X1 U13654 ( .A1(n11111), .A2(n14533), .ZN(n11080) );
  OAI211_X1 U13655 ( .C1(n11082), .C2(n14521), .A(n11081), .B(n11080), .ZN(
        P1_U3280) );
  INV_X1 U13656 ( .A(n11083), .ZN(n11084) );
  AOI22_X1 U13657 ( .A1(n13051), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11084), 
        .B2(n13015), .ZN(n11085) );
  OAI21_X1 U13658 ( .B1(n11086), .B2(n13018), .A(n11085), .ZN(n11089) );
  NOR2_X1 U13659 ( .A1(n11087), .A2(n13051), .ZN(n11088) );
  AOI211_X1 U13660 ( .C1(n11090), .C2(n13023), .A(n11089), .B(n11088), .ZN(
        n11091) );
  OAI21_X1 U13661 ( .B1(n13002), .B2(n11092), .A(n11091), .ZN(P2_U3253) );
  OAI21_X1 U13662 ( .B1(n6704), .B2(n13510), .A(n11093), .ZN(n14390) );
  INV_X1 U13663 ( .A(n14390), .ZN(n11105) );
  NAND2_X1 U13664 ( .A1(n13559), .A2(n13262), .ZN(n11095) );
  NAND2_X1 U13665 ( .A1(n13561), .A2(n13864), .ZN(n11094) );
  AND2_X1 U13666 ( .A1(n11095), .A2(n11094), .ZN(n14387) );
  INV_X1 U13667 ( .A(n14387), .ZN(n11097) );
  INV_X1 U13668 ( .A(n11096), .ZN(n13292) );
  AOI22_X1 U13669 ( .A1(n14536), .A2(n11097), .B1(n13292), .B2(n14528), .ZN(
        n11098) );
  OAI21_X1 U13670 ( .B1(n7840), .B2(n14536), .A(n11098), .ZN(n11100) );
  OAI211_X1 U13671 ( .C1(n13296), .C2(n11188), .A(n14513), .B(n11179), .ZN(
        n14386) );
  NOR2_X1 U13672 ( .A1(n14386), .A2(n13888), .ZN(n11099) );
  AOI211_X1 U13673 ( .C1(n14512), .C2(n14384), .A(n11100), .B(n11099), .ZN(
        n11104) );
  OR2_X1 U13674 ( .A1(n11102), .A2(n11101), .ZN(n14383) );
  NAND3_X1 U13675 ( .A1(n14383), .A2(n14382), .A3(n14532), .ZN(n11103) );
  OAI211_X1 U13676 ( .C1(n11105), .C2(n13895), .A(n11104), .B(n11103), .ZN(
        P1_U3278) );
  INV_X1 U13677 ( .A(n11106), .ZN(n11107) );
  OAI222_X1 U13678 ( .A1(n13160), .A2(n11108), .B1(n13178), .B2(n11107), .C1(
        P2_U3088), .C2(n12674), .ZN(P2_U3305) );
  AOI211_X1 U13679 ( .C1(n14590), .C2(n11111), .A(n11110), .B(n11109), .ZN(
        n11116) );
  INV_X1 U13680 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11112) );
  OAI22_X1 U13681 ( .A1(n6875), .A2(n14028), .B1(n8150), .B2(n11112), .ZN(
        n11113) );
  INV_X1 U13682 ( .A(n11113), .ZN(n11114) );
  OAI21_X1 U13683 ( .B1(n11116), .B2(n14577), .A(n11114), .ZN(P1_U3498) );
  INV_X1 U13684 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U13685 ( .A1(n13366), .A2(n13969), .B1(n14598), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11115) );
  OAI21_X1 U13686 ( .B1(n11116), .B2(n14598), .A(n11115), .ZN(P1_U3541) );
  INV_X1 U13687 ( .A(n11117), .ZN(n11119) );
  OAI222_X1 U13688 ( .A1(n12417), .A2(n11120), .B1(n14154), .B2(n11119), .C1(
        P3_U3151), .C2(n11118), .ZN(P3_U3266) );
  INV_X1 U13689 ( .A(n11121), .ZN(n11122) );
  AOI21_X1 U13690 ( .B1(n11124), .B2(n11123), .A(n11122), .ZN(n11132) );
  OAI22_X1 U13691 ( .A1(n11744), .A2(n11126), .B1(n11737), .B2(n11125), .ZN(
        n11127) );
  AOI211_X1 U13692 ( .C1(n11740), .C2(n14275), .A(n11128), .B(n11127), .ZN(
        n11131) );
  NAND2_X1 U13693 ( .A1(n11741), .A2(n11129), .ZN(n11130) );
  OAI211_X1 U13694 ( .C1(n11132), .C2(n11748), .A(n11131), .B(n11130), .ZN(
        P3_U3171) );
  INV_X1 U13695 ( .A(n11133), .ZN(n11135) );
  NOR2_X1 U13696 ( .A1(n9958), .A2(n11137), .ZN(n11138) );
  AOI21_X1 U13697 ( .B1(n13363), .B2(n11559), .A(n11138), .ZN(n11453) );
  AOI22_X1 U13698 ( .A1(n13363), .A2(n11554), .B1(n11559), .B2(n13563), .ZN(
        n11139) );
  XNOR2_X1 U13699 ( .A(n11139), .B(n9952), .ZN(n11452) );
  XOR2_X1 U13700 ( .A(n11453), .B(n11452), .Z(n11140) );
  OAI211_X1 U13701 ( .C1(n6705), .C2(n11140), .A(n11457), .B(n14365), .ZN(
        n11145) );
  AND2_X1 U13702 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13638) );
  NOR2_X1 U13703 ( .A1(n14369), .A2(n11141), .ZN(n11142) );
  AOI211_X1 U13704 ( .C1(n14353), .C2(n11143), .A(n13638), .B(n11142), .ZN(
        n11144) );
  OAI211_X1 U13705 ( .C1(n6876), .C2(n14362), .A(n11145), .B(n11144), .ZN(
        P1_U3224) );
  INV_X1 U13706 ( .A(n11171), .ZN(n11147) );
  NAND2_X1 U13707 ( .A1(n14035), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11146) );
  OAI211_X1 U13708 ( .C1(n11147), .C2(n14043), .A(n13546), .B(n11146), .ZN(
        P1_U3332) );
  NAND2_X1 U13709 ( .A1(n12594), .A2(n11150), .ZN(n11148) );
  OR2_X1 U13710 ( .A1(n12594), .A2(n11150), .ZN(n11151) );
  INV_X1 U13711 ( .A(n12790), .ZN(n11215) );
  XNOR2_X1 U13712 ( .A(n12599), .B(n11215), .ZN(n12747) );
  XNOR2_X1 U13713 ( .A(n11218), .B(n12747), .ZN(n11153) );
  AOI222_X1 U13714 ( .A1(n14305), .A2(n13029), .B1(n14307), .B2(n13030), .C1(
        n13026), .C2(n11153), .ZN(n14334) );
  XNOR2_X1 U13715 ( .A(n11225), .B(n12747), .ZN(n14337) );
  OAI211_X1 U13716 ( .C1(n14333), .C2(n11155), .A(n12913), .B(n11258), .ZN(
        n14332) );
  OAI22_X1 U13717 ( .A1(n12979), .A2(n11156), .B1(n14315), .B2(n13041), .ZN(
        n11157) );
  AOI21_X1 U13718 ( .B1(n12599), .B2(n13044), .A(n11157), .ZN(n11158) );
  OAI21_X1 U13719 ( .B1(n14332), .B2(n13047), .A(n11158), .ZN(n11159) );
  AOI21_X1 U13720 ( .B1(n14337), .B2(n13049), .A(n11159), .ZN(n11160) );
  OAI21_X1 U13721 ( .B1(n14334), .B2(n13051), .A(n11160), .ZN(P2_U3251) );
  INV_X1 U13722 ( .A(n11161), .ZN(n11170) );
  INV_X1 U13723 ( .A(n12788), .ZN(n13005) );
  NAND2_X1 U13724 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14704)
         );
  OAI21_X1 U13725 ( .B1(n12493), .B2(n13005), .A(n14704), .ZN(n11162) );
  AOI21_X1 U13726 ( .B1(n14306), .B2(n12789), .A(n11162), .ZN(n11163) );
  OAI21_X1 U13727 ( .B1(n11290), .B2(n14331), .A(n11163), .ZN(n11164) );
  AOI21_X1 U13728 ( .B1(n12618), .B2(n14328), .A(n11164), .ZN(n11169) );
  INV_X1 U13729 ( .A(n12789), .ZN(n11281) );
  OAI22_X1 U13730 ( .A1(n11165), .A2(n14302), .B1(n11281), .B2(n12502), .ZN(
        n11166) );
  NAND3_X1 U13731 ( .A1(n14321), .A2(n11167), .A3(n11166), .ZN(n11168) );
  OAI211_X1 U13732 ( .C1(n11170), .C2(n14302), .A(n11169), .B(n11168), .ZN(
        P2_U3200) );
  NAND2_X1 U13733 ( .A1(n11171), .A2(n13164), .ZN(n11173) );
  OR2_X1 U13734 ( .A1(n11172), .A2(P2_U3088), .ZN(n12781) );
  OAI211_X1 U13735 ( .C1(n15285), .C2(n13160), .A(n11173), .B(n12781), .ZN(
        P2_U3304) );
  OAI222_X1 U13736 ( .A1(n13178), .A2(n11202), .B1(n11175), .B2(P2_U3088), 
        .C1(n11174), .C2(n13160), .ZN(P2_U3303) );
  XNOR2_X1 U13737 ( .A(n11176), .B(n13511), .ZN(n13990) );
  XNOR2_X1 U13738 ( .A(n11177), .B(n13511), .ZN(n11178) );
  AOI22_X1 U13739 ( .A1(n13865), .A2(n13262), .B1(n13560), .B2(n13864), .ZN(
        n14361) );
  OAI21_X1 U13740 ( .B1(n11178), .B2(n14505), .A(n14361), .ZN(n13986) );
  NAND2_X1 U13741 ( .A1(n13986), .A2(n14536), .ZN(n11184) );
  AOI211_X1 U13742 ( .C1(n13988), .C2(n11179), .A(n13884), .B(n6881), .ZN(
        n13987) );
  INV_X1 U13743 ( .A(n13988), .ZN(n14363) );
  NOR2_X1 U13744 ( .A1(n14363), .A2(n14376), .ZN(n11182) );
  INV_X1 U13745 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11180) );
  OAI22_X1 U13746 ( .A1(n14536), .A2(n11180), .B1(n14368), .B2(n14508), .ZN(
        n11181) );
  AOI211_X1 U13747 ( .C1(n13987), .C2(n14517), .A(n11182), .B(n11181), .ZN(
        n11183) );
  OAI211_X1 U13748 ( .C1(n13990), .C2(n13895), .A(n11184), .B(n11183), .ZN(
        P1_U3277) );
  NAND2_X1 U13749 ( .A1(n11185), .A2(n13377), .ZN(n11186) );
  AND2_X1 U13750 ( .A1(n11187), .A2(n11186), .ZN(n14379) );
  AOI211_X1 U13751 ( .C1(n14370), .C2(n11189), .A(n13884), .B(n11188), .ZN(
        n14371) );
  NAND3_X1 U13752 ( .A1(n11191), .A2(n6984), .A3(n11190), .ZN(n11192) );
  AND3_X1 U13753 ( .A1(n11193), .A2(n14585), .A3(n11192), .ZN(n11194) );
  OAI22_X1 U13754 ( .A1(n11478), .A2(n13686), .B1(n11458), .B2(n13542), .ZN(
        n14354) );
  NOR2_X1 U13755 ( .A1(n11194), .A2(n14354), .ZN(n14381) );
  INV_X1 U13756 ( .A(n14381), .ZN(n11195) );
  AOI211_X1 U13757 ( .C1(n14379), .C2(n14590), .A(n14371), .B(n11195), .ZN(
        n11200) );
  AOI22_X1 U13758 ( .A1(n14370), .A2(n13969), .B1(n14598), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n11196) );
  OAI21_X1 U13759 ( .B1(n11200), .B2(n14598), .A(n11196), .ZN(P1_U3542) );
  INV_X1 U13760 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11197) );
  NOR2_X1 U13761 ( .A1(n8150), .A2(n11197), .ZN(n11198) );
  AOI21_X1 U13762 ( .B1(n14370), .B2(n14023), .A(n11198), .ZN(n11199) );
  OAI21_X1 U13763 ( .B1(n11200), .B2(n14577), .A(n11199), .ZN(P1_U3501) );
  OAI222_X1 U13764 ( .A1(n14047), .A2(n11203), .B1(n14043), .B2(n11202), .C1(
        n11201), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U13765 ( .A(n11204), .ZN(n11205) );
  NAND2_X1 U13766 ( .A1(n14304), .A2(n11205), .ZN(n14316) );
  XNOR2_X1 U13767 ( .A(n14316), .B(n14317), .ZN(n11208) );
  INV_X1 U13768 ( .A(n11208), .ZN(n11206) );
  AOI22_X1 U13769 ( .A1(n11206), .A2(n9282), .B1(n12465), .B2(n14307), .ZN(
        n11214) );
  NOR2_X1 U13770 ( .A1(n11208), .A2(n11207), .ZN(n14318) );
  NAND2_X1 U13771 ( .A1(n12789), .A2(n13030), .ZN(n11210) );
  NAND2_X1 U13772 ( .A1(n12790), .A2(n13029), .ZN(n11209) );
  NAND2_X1 U13773 ( .A1(n11210), .A2(n11209), .ZN(n11254) );
  AOI22_X1 U13774 ( .A1(n14325), .A2(n11254), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11211) );
  OAI21_X1 U13775 ( .B1(n11259), .B2(n14331), .A(n11211), .ZN(n11212) );
  AOI21_X1 U13776 ( .B1(n13137), .B2(n14328), .A(n11212), .ZN(n11213) );
  OAI21_X1 U13777 ( .B1(n11214), .B2(n14318), .A(n11213), .ZN(P2_U3213) );
  NOR2_X1 U13778 ( .A1(n12599), .A2(n11215), .ZN(n11217) );
  NAND2_X1 U13779 ( .A1(n12599), .A2(n11215), .ZN(n11216) );
  XNOR2_X1 U13780 ( .A(n13137), .B(n14307), .ZN(n12746) );
  INV_X1 U13781 ( .A(n12746), .ZN(n11252) );
  INV_X1 U13782 ( .A(n14307), .ZN(n11219) );
  OR2_X1 U13783 ( .A1(n13137), .A2(n11219), .ZN(n11280) );
  NAND2_X1 U13784 ( .A1(n11283), .A2(n11280), .ZN(n11220) );
  XNOR2_X1 U13785 ( .A(n14327), .B(n11281), .ZN(n12748) );
  XNOR2_X1 U13786 ( .A(n11220), .B(n12748), .ZN(n11223) );
  NAND2_X1 U13787 ( .A1(n13028), .A2(n13030), .ZN(n11222) );
  NAND2_X1 U13788 ( .A1(n14307), .A2(n13029), .ZN(n11221) );
  NAND2_X1 U13789 ( .A1(n11222), .A2(n11221), .ZN(n14326) );
  AOI21_X1 U13790 ( .B1(n11223), .B2(n13026), .A(n14326), .ZN(n13135) );
  NOR2_X1 U13791 ( .A1(n12599), .A2(n12790), .ZN(n11224) );
  XNOR2_X1 U13792 ( .A(n11289), .B(n12748), .ZN(n13133) );
  NAND2_X1 U13793 ( .A1(n14327), .A2(n11256), .ZN(n11226) );
  NAND2_X1 U13794 ( .A1(n11226), .A2(n12913), .ZN(n11227) );
  OR2_X1 U13795 ( .A1(n6700), .A2(n11227), .ZN(n13130) );
  INV_X1 U13796 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11228) );
  OAI22_X1 U13797 ( .A1(n12979), .A2(n11228), .B1(n14330), .B2(n13041), .ZN(
        n11229) );
  AOI21_X1 U13798 ( .B1(n14327), .B2(n13044), .A(n11229), .ZN(n11230) );
  OAI21_X1 U13799 ( .B1(n13130), .B2(n13047), .A(n11230), .ZN(n11231) );
  AOI21_X1 U13800 ( .B1(n13133), .B2(n13049), .A(n11231), .ZN(n11232) );
  OAI21_X1 U13801 ( .B1(n13135), .B2(n13051), .A(n11232), .ZN(P2_U3249) );
  OAI211_X1 U13802 ( .C1(n11234), .C2(n11788), .A(n11233), .B(n14982), .ZN(
        n11236) );
  AOI22_X1 U13803 ( .A1(n14977), .A2(n11977), .B1(n14258), .B2(n14980), .ZN(
        n11235) );
  AND2_X1 U13804 ( .A1(n11236), .A2(n11235), .ZN(n12318) );
  INV_X1 U13805 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11238) );
  INV_X1 U13806 ( .A(n11376), .ZN(n11237) );
  OAI22_X1 U13807 ( .A1(n14995), .A2(n11238), .B1(n11237), .B2(n15010), .ZN(
        n11239) );
  AOI21_X1 U13808 ( .B1(n12316), .B2(n14253), .A(n11239), .ZN(n11242) );
  XNOR2_X1 U13809 ( .A(n11240), .B(n11788), .ZN(n12401) );
  OR2_X1 U13810 ( .A1(n12401), .A2(n14269), .ZN(n11241) );
  OAI211_X1 U13811 ( .C1(n12318), .C2(n15018), .A(n11242), .B(n11241), .ZN(
        P3_U3219) );
  XNOR2_X1 U13812 ( .A(n11243), .B(n11787), .ZN(n12406) );
  INV_X1 U13813 ( .A(n11787), .ZN(n11869) );
  XNOR2_X1 U13814 ( .A(n11244), .B(n11869), .ZN(n11245) );
  OAI222_X1 U13815 ( .A1(n12254), .A2(n12251), .B1(n12252), .B2(n11307), .C1(
        n12249), .C2(n11245), .ZN(n12321) );
  NAND2_X1 U13816 ( .A1(n12321), .A2(n14995), .ZN(n11251) );
  INV_X1 U13817 ( .A(n11246), .ZN(n12322) );
  INV_X1 U13818 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11248) );
  INV_X1 U13819 ( .A(n11272), .ZN(n11247) );
  OAI22_X1 U13820 ( .A1(n14995), .A2(n11248), .B1(n11247), .B2(n15010), .ZN(
        n11249) );
  AOI21_X1 U13821 ( .B1(n12322), .B2(n14253), .A(n11249), .ZN(n11250) );
  OAI211_X1 U13822 ( .C1(n14269), .C2(n12406), .A(n11251), .B(n11250), .ZN(
        P3_U3220) );
  AOI21_X1 U13823 ( .B1(n11253), .B2(n11252), .A(n12977), .ZN(n11255) );
  AOI21_X1 U13824 ( .B1(n11255), .B2(n11283), .A(n11254), .ZN(n13139) );
  INV_X1 U13825 ( .A(n11256), .ZN(n11257) );
  AOI211_X1 U13826 ( .C1(n13137), .C2(n11258), .A(n9183), .B(n11257), .ZN(
        n13136) );
  INV_X1 U13827 ( .A(n13137), .ZN(n11262) );
  INV_X1 U13828 ( .A(n11259), .ZN(n11260) );
  AOI22_X1 U13829 ( .A1(n13051), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11260), 
        .B2(n13015), .ZN(n11261) );
  OAI21_X1 U13830 ( .B1(n11262), .B2(n13018), .A(n11261), .ZN(n11265) );
  AOI21_X1 U13831 ( .B1(n12746), .B2(n11263), .A(n6707), .ZN(n13141) );
  NOR2_X1 U13832 ( .A1(n13141), .A2(n13002), .ZN(n11264) );
  AOI211_X1 U13833 ( .C1(n13136), .C2(n13023), .A(n11265), .B(n11264), .ZN(
        n11266) );
  OAI21_X1 U13834 ( .B1(n13051), .B2(n13139), .A(n11266), .ZN(P2_U3250) );
  INV_X1 U13835 ( .A(n11267), .ZN(n11269) );
  NAND2_X1 U13836 ( .A1(n11269), .A2(n11268), .ZN(n11270) );
  XNOR2_X1 U13837 ( .A(n11271), .B(n11270), .ZN(n11278) );
  NAND2_X1 U13838 ( .A1(n11741), .A2(n11272), .ZN(n11275) );
  NOR2_X1 U13839 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11273), .ZN(n14920) );
  AOI21_X1 U13840 ( .B1(n11740), .B2(n11978), .A(n14920), .ZN(n11274) );
  OAI211_X1 U13841 ( .C1(n11307), .C2(n11744), .A(n11275), .B(n11274), .ZN(
        n11276) );
  AOI21_X1 U13842 ( .B1(n12322), .B2(n11746), .A(n11276), .ZN(n11277) );
  OAI21_X1 U13843 ( .B1(n11278), .B2(n11748), .A(n11277), .ZN(P3_U3174) );
  OR2_X1 U13844 ( .A1(n14327), .A2(n11281), .ZN(n11279) );
  AND2_X1 U13845 ( .A1(n11280), .A2(n11279), .ZN(n11282) );
  INV_X1 U13846 ( .A(n13028), .ZN(n11410) );
  XNOR2_X1 U13847 ( .A(n12618), .B(n11410), .ZN(n12750) );
  XNOR2_X1 U13848 ( .A(n11413), .B(n12750), .ZN(n11284) );
  NAND2_X1 U13849 ( .A1(n11284), .A2(n13026), .ZN(n11286) );
  AOI22_X1 U13850 ( .A1(n12788), .A2(n13030), .B1(n13029), .B2(n12789), .ZN(
        n11285) );
  NAND2_X1 U13851 ( .A1(n11286), .A2(n11285), .ZN(n13129) );
  INV_X1 U13852 ( .A(n13129), .ZN(n11296) );
  INV_X1 U13853 ( .A(n12748), .ZN(n11288) );
  NAND2_X1 U13854 ( .A1(n14327), .A2(n12789), .ZN(n11287) );
  INV_X1 U13855 ( .A(n12750), .ZN(n11412) );
  XNOR2_X1 U13856 ( .A(n11383), .B(n11412), .ZN(n13124) );
  INV_X1 U13857 ( .A(n12618), .ZN(n13126) );
  OAI211_X1 U13858 ( .C1(n13126), .C2(n6700), .A(n12913), .B(n13038), .ZN(
        n13125) );
  OAI22_X1 U13859 ( .A1(n12979), .A2(n11291), .B1(n11290), .B2(n13041), .ZN(
        n11292) );
  AOI21_X1 U13860 ( .B1(n12618), .B2(n13044), .A(n11292), .ZN(n11293) );
  OAI21_X1 U13861 ( .B1(n13125), .B2(n13047), .A(n11293), .ZN(n11294) );
  AOI21_X1 U13862 ( .B1(n13124), .B2(n13049), .A(n11294), .ZN(n11295) );
  OAI21_X1 U13863 ( .B1(n11296), .B2(n13051), .A(n11295), .ZN(P2_U3248) );
  INV_X1 U13864 ( .A(n13045), .ZN(n13120) );
  OAI211_X1 U13865 ( .C1(n11299), .C2(n11298), .A(n11297), .B(n9282), .ZN(
        n11303) );
  NOR2_X1 U13866 ( .A1(n14331), .A2(n13042), .ZN(n11301) );
  INV_X1 U13867 ( .A(n13031), .ZN(n11415) );
  NAND2_X1 U13868 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14720)
         );
  OAI21_X1 U13869 ( .B1(n12493), .B2(n11415), .A(n14720), .ZN(n11300) );
  AOI211_X1 U13870 ( .C1(n14306), .C2(n13028), .A(n11301), .B(n11300), .ZN(
        n11302) );
  OAI211_X1 U13871 ( .C1(n13120), .C2(n14310), .A(n11303), .B(n11302), .ZN(
        P2_U3210) );
  XNOR2_X1 U13872 ( .A(n11304), .B(n11313), .ZN(n11314) );
  XNOR2_X1 U13873 ( .A(n11314), .B(n11305), .ZN(n11312) );
  INV_X1 U13874 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11306) );
  NOR2_X1 U13875 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11306), .ZN(n14884) );
  NOR2_X1 U13876 ( .A1(n11733), .A2(n11307), .ZN(n11308) );
  AOI211_X1 U13877 ( .C1(n11731), .C2(n14275), .A(n14884), .B(n11308), .ZN(
        n11309) );
  OAI21_X1 U13878 ( .B1(n14280), .B2(n11737), .A(n11309), .ZN(n11310) );
  AOI21_X1 U13879 ( .B1(n14277), .B2(n11741), .A(n11310), .ZN(n11311) );
  OAI21_X1 U13880 ( .B1(n11312), .B2(n11748), .A(n11311), .ZN(P3_U3176) );
  OAI22_X1 U13881 ( .A1(n11314), .A2(n14259), .B1(n11313), .B2(n11304), .ZN(
        n11317) );
  XNOR2_X1 U13882 ( .A(n11315), .B(n14274), .ZN(n11316) );
  XNOR2_X1 U13883 ( .A(n11317), .B(n11316), .ZN(n11323) );
  AND2_X1 U13884 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n14903) );
  NOR2_X1 U13885 ( .A1(n11733), .A2(n11379), .ZN(n11318) );
  AOI211_X1 U13886 ( .C1(n11731), .C2(n14259), .A(n14903), .B(n11318), .ZN(
        n11319) );
  OAI21_X1 U13887 ( .B1(n14267), .B2(n11737), .A(n11319), .ZN(n11320) );
  AOI21_X1 U13888 ( .B1(n11321), .B2(n11741), .A(n11320), .ZN(n11322) );
  OAI21_X1 U13889 ( .B1(n11323), .B2(n11748), .A(n11322), .ZN(P3_U3164) );
  INV_X1 U13890 ( .A(n13165), .ZN(n11324) );
  OAI222_X1 U13891 ( .A1(n14047), .A2(n11325), .B1(n14043), .B2(n11324), .C1(
        P1_U3086), .C2(n8115), .ZN(P1_U3327) );
  INV_X1 U13892 ( .A(n11326), .ZN(n11328) );
  OAI222_X1 U13893 ( .A1(n11329), .A2(P3_U3151), .B1(n14154), .B2(n11328), 
        .C1(n11327), .C2(n12417), .ZN(P3_U3267) );
  INV_X1 U13894 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14038) );
  INV_X1 U13895 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11333) );
  MUX2_X1 U13896 ( .A(n14038), .B(n11333), .S(n8042), .Z(n11349) );
  XNOR2_X1 U13897 ( .A(n11349), .B(SI_29_), .ZN(n11352) );
  INV_X1 U13898 ( .A(n13454), .ZN(n14039) );
  OAI222_X1 U13899 ( .A1(n13178), .A2(n14039), .B1(n11334), .B2(P2_U3088), 
        .C1(n11333), .C2(n13160), .ZN(P2_U3298) );
  XNOR2_X1 U13900 ( .A(n11335), .B(n13518), .ZN(n11341) );
  OAI22_X1 U13901 ( .A1(n11336), .A2(n13542), .B1(n13430), .B2(n13686), .ZN(
        n13183) );
  AOI211_X1 U13902 ( .C1(n13915), .C2(n13727), .A(n13884), .B(n11342), .ZN(
        n13914) );
  INV_X1 U13903 ( .A(n13185), .ZN(n11343) );
  AOI22_X1 U13904 ( .A1(n14521), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n11343), 
        .B2(n14528), .ZN(n11344) );
  OAI21_X1 U13905 ( .B1(n11345), .B2(n14376), .A(n11344), .ZN(n11347) );
  NOR2_X1 U13906 ( .A1(n13918), .A2(n13877), .ZN(n11346) );
  AOI211_X1 U13907 ( .C1(n13914), .C2(n14517), .A(n11347), .B(n11346), .ZN(
        n11348) );
  OAI21_X1 U13908 ( .B1(n13917), .B2(n14521), .A(n11348), .ZN(P1_U3266) );
  INV_X1 U13909 ( .A(n11349), .ZN(n11350) );
  NOR2_X1 U13910 ( .A1(n11350), .A2(SI_29_), .ZN(n11351) );
  INV_X1 U13911 ( .A(n11358), .ZN(n11355) );
  MUX2_X1 U13912 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8042), .Z(n11354) );
  NAND2_X1 U13913 ( .A1(n11354), .A2(SI_30_), .ZN(n12678) );
  OAI21_X1 U13914 ( .B1(n11354), .B2(SI_30_), .A(n12678), .ZN(n11356) );
  NAND2_X1 U13915 ( .A1(n11355), .A2(n11356), .ZN(n11359) );
  INV_X1 U13916 ( .A(n11356), .ZN(n11357) );
  NAND2_X1 U13917 ( .A1(n11358), .A2(n11357), .ZN(n12679) );
  INV_X1 U13918 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11759) );
  OAI222_X1 U13919 ( .A1(n11360), .A2(P1_U3086), .B1(n14043), .B2(n13445), 
        .C1(n11759), .C2(n14047), .ZN(P1_U3325) );
  OR2_X1 U13920 ( .A1(n11361), .A2(n11362), .ZN(n11364) );
  NAND2_X1 U13921 ( .A1(n11364), .A2(n11363), .ZN(n11367) );
  NOR2_X1 U13922 ( .A1(n11365), .A2(n7547), .ZN(n11366) );
  XNOR2_X1 U13923 ( .A(n11367), .B(n11366), .ZN(n11373) );
  NAND2_X1 U13924 ( .A1(n11741), .A2(n12227), .ZN(n11370) );
  NOR2_X1 U13925 ( .A1(n11368), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14233) );
  AOI21_X1 U13926 ( .B1(n11740), .B2(n12224), .A(n14233), .ZN(n11369) );
  OAI211_X1 U13927 ( .C1(n12253), .C2(n11744), .A(n11370), .B(n11369), .ZN(
        n11371) );
  AOI21_X1 U13928 ( .B1(n12303), .B2(n11746), .A(n11371), .ZN(n11372) );
  OAI21_X1 U13929 ( .B1(n11373), .B2(n11748), .A(n11372), .ZN(P3_U3168) );
  XOR2_X1 U13930 ( .A(n11375), .B(n11374), .Z(n11382) );
  AOI22_X1 U13931 ( .A1(n11740), .A2(n11977), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11378) );
  NAND2_X1 U13932 ( .A1(n11741), .A2(n11376), .ZN(n11377) );
  OAI211_X1 U13933 ( .C1(n11379), .C2(n11744), .A(n11378), .B(n11377), .ZN(
        n11380) );
  AOI21_X1 U13934 ( .B1(n12316), .B2(n11746), .A(n11380), .ZN(n11381) );
  OAI21_X1 U13935 ( .B1(n11382), .B2(n11748), .A(n11381), .ZN(P3_U3155) );
  NAND2_X1 U13936 ( .A1(n11383), .A2(n12750), .ZN(n11385) );
  NAND2_X1 U13937 ( .A1(n12618), .A2(n13028), .ZN(n11384) );
  NAND2_X1 U13938 ( .A1(n11385), .A2(n11384), .ZN(n13035) );
  INV_X1 U13939 ( .A(n13035), .ZN(n11386) );
  XNOR2_X1 U13940 ( .A(n13045), .B(n13005), .ZN(n12752) );
  OR2_X1 U13941 ( .A1(n13045), .A2(n12788), .ZN(n11387) );
  NAND2_X1 U13942 ( .A1(n13037), .A2(n11387), .ZN(n13009) );
  NAND2_X1 U13943 ( .A1(n13114), .A2(n13031), .ZN(n11388) );
  OR2_X1 U13944 ( .A1(n13114), .A2(n13031), .ZN(n11389) );
  NAND2_X1 U13945 ( .A1(n13109), .A2(n12787), .ZN(n11390) );
  INV_X1 U13946 ( .A(n12997), .ZN(n12492) );
  XNOR2_X1 U13947 ( .A(n13105), .B(n12492), .ZN(n12974) );
  INV_X1 U13948 ( .A(n12974), .ZN(n11393) );
  OR2_X1 U13949 ( .A1(n13105), .A2(n12997), .ZN(n11392) );
  NAND2_X1 U13950 ( .A1(n13099), .A2(n12978), .ZN(n11394) );
  NAND2_X1 U13951 ( .A1(n13094), .A2(n12786), .ZN(n12755) );
  OR2_X1 U13952 ( .A1(n13094), .A2(n12786), .ZN(n12756) );
  XNOR2_X1 U13953 ( .A(n13089), .B(n12944), .ZN(n12937) );
  NOR2_X1 U13954 ( .A1(n13084), .A2(n12893), .ZN(n11395) );
  INV_X1 U13955 ( .A(n12877), .ZN(n12883) );
  NAND2_X1 U13956 ( .A1(n13165), .A2(n12684), .ZN(n11398) );
  NAND2_X1 U13957 ( .A1(n12685), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U13958 ( .A1(n12872), .A2(n11425), .ZN(n11400) );
  INV_X1 U13959 ( .A(n12861), .ZN(n12866) );
  NAND2_X1 U13960 ( .A1(n12867), .A2(n12866), .ZN(n12865) );
  NAND2_X1 U13961 ( .A1(n13454), .A2(n12684), .ZN(n11402) );
  NAND2_X1 U13962 ( .A1(n12685), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11401) );
  NAND2_X2 U13963 ( .A1(n11402), .A2(n11401), .ZN(n13059) );
  OR2_X1 U13964 ( .A1(n11442), .A2(n11403), .ZN(n11408) );
  INV_X1 U13965 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n15240) );
  NAND2_X1 U13966 ( .A1(n11429), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U13967 ( .A1(n8861), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11404) );
  OAI211_X1 U13968 ( .C1(n12670), .C2(n15240), .A(n11405), .B(n11404), .ZN(
        n11406) );
  INV_X1 U13969 ( .A(n11406), .ZN(n11407) );
  NAND2_X1 U13970 ( .A1(n11408), .A2(n11407), .ZN(n12784) );
  INV_X1 U13971 ( .A(n12784), .ZN(n11409) );
  INV_X1 U13972 ( .A(n12944), .ZN(n12911) );
  INV_X1 U13973 ( .A(n13114), .ZN(n13019) );
  NOR2_X1 U13974 ( .A1(n12618), .A2(n11410), .ZN(n11411) );
  INV_X1 U13975 ( .A(n12787), .ZN(n13007) );
  NAND2_X1 U13976 ( .A1(n13109), .A2(n13007), .ZN(n11418) );
  OR2_X1 U13977 ( .A1(n13109), .A2(n13007), .ZN(n11417) );
  NAND2_X1 U13978 ( .A1(n12995), .A2(n12996), .ZN(n12994) );
  INV_X1 U13979 ( .A(n13105), .ZN(n12984) );
  NAND2_X1 U13980 ( .A1(n12984), .A2(n12997), .ZN(n11419) );
  INV_X1 U13981 ( .A(n13094), .ZN(n12951) );
  OAI21_X1 U13982 ( .B1(n12927), .B2(n13094), .A(n11422), .ZN(n12924) );
  INV_X1 U13983 ( .A(n12937), .ZN(n12925) );
  AOI21_X1 U13984 ( .B1(n12911), .B2(n13089), .A(n12923), .ZN(n12909) );
  XNOR2_X1 U13985 ( .A(n13084), .B(n12928), .ZN(n12908) );
  NOR2_X1 U13986 ( .A1(n13078), .A2(n12912), .ZN(n11424) );
  NAND2_X1 U13987 ( .A1(n12860), .A2(n11426), .ZN(n11427) );
  XNOR2_X1 U13988 ( .A(n11427), .B(n12760), .ZN(n11428) );
  NAND2_X1 U13989 ( .A1(n11428), .A2(n13026), .ZN(n11439) );
  INV_X1 U13990 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n11433) );
  NAND2_X1 U13991 ( .A1(n11429), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U13992 ( .A1(n11430), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11431) );
  OAI211_X1 U13993 ( .C1(n12668), .C2(n11433), .A(n11432), .B(n11431), .ZN(
        n12783) );
  INV_X1 U13994 ( .A(P2_B_REG_SCAN_IN), .ZN(n11434) );
  NOR2_X1 U13995 ( .A1(n6777), .A2(n11434), .ZN(n11435) );
  NOR2_X1 U13996 ( .A1(n13006), .A2(n11435), .ZN(n12848) );
  NAND2_X1 U13997 ( .A1(n12783), .A2(n12848), .ZN(n11436) );
  INV_X1 U13998 ( .A(n11437), .ZN(n11438) );
  NAND2_X1 U13999 ( .A1(n13058), .A2(n12979), .ZN(n11447) );
  INV_X1 U14000 ( .A(n13109), .ZN(n12993) );
  NAND2_X1 U14001 ( .A1(n13013), .A2(n12993), .ZN(n12990) );
  AND2_X2 U14002 ( .A1(n13072), .A2(n12895), .ZN(n12882) );
  AOI21_X1 U14003 ( .B1(n13059), .B2(n12868), .A(n9183), .ZN(n11440) );
  NAND2_X1 U14004 ( .A1(n11440), .A2(n12854), .ZN(n13060) );
  INV_X1 U14005 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11441) );
  OAI22_X1 U14006 ( .A1(n11442), .A2(n13041), .B1(n11441), .B2(n12979), .ZN(
        n11443) );
  AOI21_X1 U14007 ( .B1(n13059), .B2(n13044), .A(n11443), .ZN(n11444) );
  OAI21_X1 U14008 ( .B1(n13060), .B2(n13047), .A(n11444), .ZN(n11445) );
  INV_X1 U14009 ( .A(n11445), .ZN(n11446) );
  OAI211_X1 U14010 ( .C1(n13063), .C2(n13002), .A(n11447), .B(n11446), .ZN(
        P2_U3236) );
  NOR2_X1 U14011 ( .A1(n13271), .A2(n9958), .ZN(n11448) );
  AOI21_X1 U14012 ( .B1(n14022), .B2(n11559), .A(n11448), .ZN(n11505) );
  NAND2_X1 U14013 ( .A1(n14022), .A2(n11554), .ZN(n11450) );
  OR2_X1 U14014 ( .A1(n13271), .A2(n11563), .ZN(n11449) );
  NAND2_X1 U14015 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  XNOR2_X1 U14016 ( .A(n11451), .B(n9952), .ZN(n11503) );
  INV_X1 U14017 ( .A(n11503), .ZN(n11504) );
  INV_X1 U14018 ( .A(n11452), .ZN(n11455) );
  INV_X1 U14019 ( .A(n11453), .ZN(n11454) );
  NAND2_X1 U14020 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  NOR2_X1 U14021 ( .A1(n9958), .A2(n11458), .ZN(n11459) );
  AOI21_X1 U14022 ( .B1(n13366), .B2(n11559), .A(n11459), .ZN(n11467) );
  AOI22_X1 U14023 ( .A1(n13366), .A2(n11554), .B1(n11559), .B2(n13562), .ZN(
        n11460) );
  XNOR2_X1 U14024 ( .A(n11460), .B(n9952), .ZN(n11466) );
  XOR2_X1 U14025 ( .A(n11467), .B(n11466), .Z(n13250) );
  NAND2_X1 U14026 ( .A1(n14370), .A2(n11554), .ZN(n11462) );
  NAND2_X1 U14027 ( .A1(n13561), .A2(n11559), .ZN(n11461) );
  NAND2_X1 U14028 ( .A1(n11462), .A2(n11461), .ZN(n11463) );
  XNOR2_X1 U14029 ( .A(n11463), .B(n9952), .ZN(n11471) );
  NOR2_X1 U14030 ( .A1(n9958), .A2(n11464), .ZN(n11465) );
  AOI21_X1 U14031 ( .B1(n14370), .B2(n11559), .A(n11465), .ZN(n11472) );
  XNOR2_X1 U14032 ( .A(n11471), .B(n11472), .ZN(n14348) );
  INV_X1 U14033 ( .A(n11466), .ZN(n11469) );
  INV_X1 U14034 ( .A(n11467), .ZN(n11468) );
  NAND2_X1 U14035 ( .A1(n11469), .A2(n11468), .ZN(n14349) );
  INV_X1 U14036 ( .A(n11471), .ZN(n11473) );
  NAND2_X1 U14037 ( .A1(n14384), .A2(n11554), .ZN(n11475) );
  OR2_X1 U14038 ( .A1(n11478), .A2(n11563), .ZN(n11474) );
  NAND2_X1 U14039 ( .A1(n11475), .A2(n11474), .ZN(n11477) );
  XNOR2_X1 U14040 ( .A(n11477), .B(n11476), .ZN(n11483) );
  OAI22_X1 U14041 ( .A1(n13296), .A2(n11563), .B1(n11478), .B2(n9958), .ZN(
        n13289) );
  NAND2_X1 U14042 ( .A1(n13290), .A2(n13289), .ZN(n13288) );
  NAND2_X1 U14043 ( .A1(n13988), .A2(n11554), .ZN(n11480) );
  NAND2_X1 U14044 ( .A1(n13559), .A2(n11559), .ZN(n11479) );
  NAND2_X1 U14045 ( .A1(n11480), .A2(n11479), .ZN(n11481) );
  XNOR2_X1 U14046 ( .A(n11481), .B(n9952), .ZN(n11488) );
  AND2_X1 U14047 ( .A1(n13559), .A2(n11558), .ZN(n11482) );
  AOI21_X1 U14048 ( .B1(n13988), .B2(n11559), .A(n11482), .ZN(n11486) );
  XNOR2_X1 U14049 ( .A(n11488), .B(n11486), .ZN(n14358) );
  INV_X1 U14050 ( .A(n11483), .ZN(n11484) );
  NAND2_X1 U14051 ( .A1(n11485), .A2(n11484), .ZN(n14356) );
  INV_X1 U14052 ( .A(n11486), .ZN(n11487) );
  OR2_X1 U14053 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  NAND2_X1 U14054 ( .A1(n13979), .A2(n11554), .ZN(n11491) );
  NAND2_X1 U14055 ( .A1(n13865), .A2(n11559), .ZN(n11490) );
  NAND2_X1 U14056 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  XNOR2_X1 U14057 ( .A(n11492), .B(n9952), .ZN(n11495) );
  AOI22_X1 U14058 ( .A1(n13979), .A2(n11559), .B1(n11558), .B2(n13865), .ZN(
        n11493) );
  XNOR2_X1 U14059 ( .A(n11495), .B(n11493), .ZN(n13226) );
  INV_X1 U14060 ( .A(n11493), .ZN(n11494) );
  NAND2_X1 U14061 ( .A1(n13873), .A2(n11554), .ZN(n11498) );
  NAND2_X1 U14062 ( .A1(n13558), .A2(n11559), .ZN(n11497) );
  NAND2_X1 U14063 ( .A1(n11498), .A2(n11497), .ZN(n11499) );
  XNOR2_X1 U14064 ( .A(n11499), .B(n9952), .ZN(n11500) );
  AOI22_X1 U14065 ( .A1(n13873), .A2(n11559), .B1(n11558), .B2(n13558), .ZN(
        n11501) );
  XNOR2_X1 U14066 ( .A(n11500), .B(n11501), .ZN(n13270) );
  INV_X1 U14067 ( .A(n11500), .ZN(n11502) );
  XNOR2_X1 U14068 ( .A(n11503), .B(n11505), .ZN(n13198) );
  OR2_X1 U14069 ( .A1(n13831), .A2(n11563), .ZN(n11507) );
  OR2_X1 U14070 ( .A1(n13400), .A2(n9958), .ZN(n11506) );
  NAND2_X1 U14071 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  OAI22_X1 U14072 ( .A1(n13831), .A2(n11564), .B1(n13400), .B2(n11563), .ZN(
        n11508) );
  XNOR2_X1 U14073 ( .A(n11508), .B(n9952), .ZN(n11510) );
  XOR2_X1 U14074 ( .A(n11509), .B(n11510), .Z(n13242) );
  NAND2_X1 U14075 ( .A1(n13243), .A2(n13242), .ZN(n13241) );
  NAND2_X1 U14076 ( .A1(n11510), .A2(n11509), .ZN(n11511) );
  AOI22_X1 U14077 ( .A1(n13950), .A2(n11554), .B1(n9963), .B2(n13555), .ZN(
        n11512) );
  XNOR2_X1 U14078 ( .A(n11512), .B(n9952), .ZN(n11515) );
  AOI22_X1 U14079 ( .A1(n13950), .A2(n11559), .B1(n11558), .B2(n13555), .ZN(
        n11514) );
  XNOR2_X1 U14080 ( .A(n11515), .B(n11514), .ZN(n13209) );
  INV_X1 U14081 ( .A(n13209), .ZN(n11513) );
  NAND2_X1 U14082 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  NAND2_X1 U14083 ( .A1(n13946), .A2(n11554), .ZN(n11518) );
  NAND2_X1 U14084 ( .A1(n13554), .A2(n11559), .ZN(n11517) );
  NAND2_X1 U14085 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  XNOR2_X1 U14086 ( .A(n11519), .B(n9952), .ZN(n11520) );
  AOI22_X1 U14087 ( .A1(n13946), .A2(n11559), .B1(n11558), .B2(n13554), .ZN(
        n11521) );
  XNOR2_X1 U14088 ( .A(n11520), .B(n11521), .ZN(n13260) );
  INV_X1 U14089 ( .A(n11520), .ZN(n11522) );
  NAND2_X1 U14090 ( .A1(n11522), .A2(n11521), .ZN(n11523) );
  NAND2_X1 U14091 ( .A1(n13939), .A2(n11554), .ZN(n11525) );
  NAND2_X1 U14092 ( .A1(n11559), .A2(n13553), .ZN(n11524) );
  NAND2_X1 U14093 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  XNOR2_X1 U14094 ( .A(n11526), .B(n9952), .ZN(n11527) );
  AOI22_X1 U14095 ( .A1(n13939), .A2(n11559), .B1(n11558), .B2(n13553), .ZN(
        n11528) );
  XNOR2_X1 U14096 ( .A(n11527), .B(n11528), .ZN(n13190) );
  INV_X1 U14097 ( .A(n11527), .ZN(n11529) );
  NAND2_X1 U14098 ( .A1(n11529), .A2(n11528), .ZN(n11530) );
  NAND2_X1 U14099 ( .A1(n11531), .A2(n11530), .ZN(n13233) );
  NAND2_X1 U14100 ( .A1(n14011), .A2(n11554), .ZN(n11533) );
  NAND2_X1 U14101 ( .A1(n11559), .A2(n13552), .ZN(n11532) );
  NAND2_X1 U14102 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  XNOR2_X1 U14103 ( .A(n11534), .B(n9952), .ZN(n11535) );
  AOI22_X1 U14104 ( .A1(n14011), .A2(n11559), .B1(n11558), .B2(n13552), .ZN(
        n11536) );
  XNOR2_X1 U14105 ( .A(n11535), .B(n11536), .ZN(n13234) );
  INV_X1 U14106 ( .A(n11535), .ZN(n11537) );
  NAND2_X1 U14107 ( .A1(n11537), .A2(n11536), .ZN(n11538) );
  NAND2_X1 U14108 ( .A1(n14007), .A2(n11554), .ZN(n11540) );
  NAND2_X1 U14109 ( .A1(n13551), .A2(n11559), .ZN(n11539) );
  NAND2_X1 U14110 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  XNOR2_X1 U14111 ( .A(n11541), .B(n9952), .ZN(n11542) );
  AOI22_X1 U14112 ( .A1(n14007), .A2(n11559), .B1(n11558), .B2(n13551), .ZN(
        n11543) );
  XNOR2_X1 U14113 ( .A(n11542), .B(n11543), .ZN(n13217) );
  INV_X1 U14114 ( .A(n11542), .ZN(n11544) );
  NAND2_X1 U14115 ( .A1(n11544), .A2(n11543), .ZN(n11545) );
  NAND2_X1 U14116 ( .A1(n13729), .A2(n11554), .ZN(n11548) );
  NAND2_X1 U14117 ( .A1(n13550), .A2(n11559), .ZN(n11547) );
  NAND2_X1 U14118 ( .A1(n11548), .A2(n11547), .ZN(n11549) );
  XNOR2_X1 U14119 ( .A(n11549), .B(n9952), .ZN(n11550) );
  AOI22_X1 U14120 ( .A1(n13729), .A2(n11559), .B1(n11558), .B2(n13550), .ZN(
        n11551) );
  XNOR2_X1 U14121 ( .A(n11550), .B(n11551), .ZN(n13280) );
  INV_X1 U14122 ( .A(n11550), .ZN(n11552) );
  NAND2_X1 U14123 ( .A1(n11552), .A2(n11551), .ZN(n11553) );
  NAND2_X1 U14124 ( .A1(n13915), .A2(n11554), .ZN(n11556) );
  NAND2_X1 U14125 ( .A1(n11559), .A2(n13549), .ZN(n11555) );
  NAND2_X1 U14126 ( .A1(n11556), .A2(n11555), .ZN(n11557) );
  XNOR2_X1 U14127 ( .A(n11557), .B(n9952), .ZN(n11560) );
  AOI22_X1 U14128 ( .A1(n13915), .A2(n11559), .B1(n11558), .B2(n13549), .ZN(
        n11561) );
  XNOR2_X1 U14129 ( .A(n11560), .B(n11561), .ZN(n13182) );
  INV_X1 U14130 ( .A(n11560), .ZN(n11562) );
  OAI22_X1 U14131 ( .A1(n13429), .A2(n11563), .B1(n13430), .B2(n9958), .ZN(
        n11567) );
  OAI22_X1 U14132 ( .A1(n13429), .A2(n11564), .B1(n13430), .B2(n11563), .ZN(
        n11565) );
  XNOR2_X1 U14133 ( .A(n11565), .B(n9952), .ZN(n11566) );
  XOR2_X1 U14134 ( .A(n11567), .B(n11566), .Z(n11568) );
  XNOR2_X1 U14135 ( .A(n11569), .B(n11568), .ZN(n11574) );
  AOI22_X1 U14136 ( .A1(n14353), .A2(n11570), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11571) );
  OAI21_X1 U14137 ( .B1(n14369), .B2(n13716), .A(n11571), .ZN(n11572) );
  AOI21_X1 U14138 ( .B1(n13721), .B2(n9693), .A(n11572), .ZN(n11573) );
  OAI21_X1 U14139 ( .B1(n11574), .B2(n13286), .A(n11573), .ZN(P1_U3220) );
  INV_X1 U14140 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11575) );
  OAI222_X1 U14141 ( .A1(n13178), .A2(n13445), .B1(n11576), .B2(P2_U3088), 
        .C1(n11575), .C2(n13160), .ZN(P2_U3297) );
  AOI22_X1 U14142 ( .A1(n6703), .A2(n9282), .B1(n12465), .B2(n12945), .ZN(
        n11582) );
  AND2_X1 U14143 ( .A1(n12997), .A2(n13029), .ZN(n11577) );
  AOI21_X1 U14144 ( .B1(n12786), .B2(n13030), .A(n11577), .ZN(n12959) );
  OAI22_X1 U14145 ( .A1(n12959), .A2(n12438), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11578), .ZN(n11580) );
  NOR2_X1 U14146 ( .A1(n6885), .A2(n14310), .ZN(n11579) );
  AOI211_X1 U14147 ( .C1(n12489), .C2(n12967), .A(n11580), .B(n11579), .ZN(
        n11581) );
  OAI21_X1 U14148 ( .B1(n11583), .B2(n11582), .A(n11581), .ZN(P2_U3207) );
  INV_X1 U14149 ( .A(n11584), .ZN(n11585) );
  AOI22_X1 U14150 ( .A1(n11585), .A2(n9282), .B1(n12465), .B2(n12786), .ZN(
        n11590) );
  AOI22_X1 U14151 ( .A1(n12944), .A2(n14308), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11587) );
  NAND2_X1 U14152 ( .A1(n14306), .A2(n12945), .ZN(n11586) );
  OAI211_X1 U14153 ( .C1(n14331), .C2(n12948), .A(n11587), .B(n11586), .ZN(
        n11588) );
  AOI21_X1 U14154 ( .B1(n13094), .B2(n14328), .A(n11588), .ZN(n11589) );
  OAI21_X1 U14155 ( .B1(n11591), .B2(n11590), .A(n11589), .ZN(P2_U3188) );
  OAI222_X1 U14156 ( .A1(n13178), .A2(n11592), .B1(n6559), .B2(P2_U3088), .C1(
        n15175), .C2(n13160), .ZN(P2_U3307) );
  XNOR2_X1 U14157 ( .A(n12077), .B(n9394), .ZN(n11600) );
  INV_X1 U14158 ( .A(n11600), .ZN(n11594) );
  NAND2_X1 U14159 ( .A1(n11594), .A2(n11730), .ZN(n11605) );
  INV_X1 U14160 ( .A(n11595), .ZN(n11596) );
  AOI22_X1 U14161 ( .A1(n12079), .A2(n11731), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11598) );
  NAND2_X1 U14162 ( .A1(n12083), .A2(n11741), .ZN(n11597) );
  OAI211_X1 U14163 ( .C1(n12082), .C2(n11733), .A(n11598), .B(n11597), .ZN(
        n11602) );
  NOR4_X1 U14164 ( .A1(n11600), .A2(n11599), .A3(n12079), .A4(n11748), .ZN(
        n11601) );
  AOI211_X1 U14165 ( .C1(n11746), .C2(n12263), .A(n11602), .B(n11601), .ZN(
        n11603) );
  OAI211_X1 U14166 ( .C1(n11608), .C2(n11607), .A(n11606), .B(n11730), .ZN(
        n11614) );
  AOI21_X1 U14167 ( .B1(n11740), .B2(n11979), .A(n11609), .ZN(n11613) );
  AOI22_X1 U14168 ( .A1(n11746), .A2(n15042), .B1(n11731), .B2(n11980), .ZN(
        n11612) );
  NAND2_X1 U14169 ( .A1(n11741), .A2(n11610), .ZN(n11611) );
  NAND4_X1 U14170 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        P3_U3153) );
  INV_X1 U14171 ( .A(n11615), .ZN(n11688) );
  AOI21_X1 U14172 ( .B1(n11617), .B2(n11616), .A(n11688), .ZN(n11622) );
  AOI22_X1 U14173 ( .A1(n11971), .A2(n11740), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11619) );
  NAND2_X1 U14174 ( .A1(n11741), .A2(n12144), .ZN(n11618) );
  OAI211_X1 U14175 ( .C1(n12165), .C2(n11744), .A(n11619), .B(n11618), .ZN(
        n11620) );
  AOI21_X1 U14176 ( .B1(n12281), .B2(n11746), .A(n11620), .ZN(n11621) );
  OAI21_X1 U14177 ( .B1(n11622), .B2(n11748), .A(n11621), .ZN(P3_U3156) );
  AOI21_X1 U14178 ( .B1(n11624), .B2(n11623), .A(n11748), .ZN(n11626) );
  NAND2_X1 U14179 ( .A1(n11626), .A2(n11625), .ZN(n11632) );
  INV_X1 U14180 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15163) );
  NOR2_X1 U14181 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15163), .ZN(n14859) );
  AOI21_X1 U14182 ( .B1(n11740), .B2(n14259), .A(n14859), .ZN(n11631) );
  AOI22_X1 U14183 ( .A1(n11746), .A2(n11627), .B1(n11731), .B2(n14951), .ZN(
        n11630) );
  NAND2_X1 U14184 ( .A1(n11741), .A2(n11628), .ZN(n11629) );
  NAND4_X1 U14185 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        P3_U3157) );
  XNOR2_X1 U14186 ( .A(n11634), .B(n11633), .ZN(n11639) );
  NAND2_X1 U14187 ( .A1(n11731), .A2(n12224), .ZN(n11635) );
  NAND2_X1 U14188 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12056)
         );
  OAI211_X1 U14189 ( .C1(n12166), .C2(n11733), .A(n11635), .B(n12056), .ZN(
        n11637) );
  NOR2_X1 U14190 ( .A1(n12196), .A2(n11737), .ZN(n11636) );
  AOI211_X1 U14191 ( .C1(n12197), .C2(n11741), .A(n11637), .B(n11636), .ZN(
        n11638) );
  OAI21_X1 U14192 ( .B1(n11639), .B2(n11748), .A(n11638), .ZN(P3_U3159) );
  OAI211_X1 U14193 ( .C1(n11642), .C2(n11641), .A(n11640), .B(n11730), .ZN(
        n11647) );
  AOI21_X1 U14194 ( .B1(n11740), .B2(n14951), .A(n11643), .ZN(n11646) );
  AOI22_X1 U14195 ( .A1(n11746), .A2(n14955), .B1(n11731), .B2(n14964), .ZN(
        n11645) );
  NAND2_X1 U14196 ( .A1(n11741), .A2(n14956), .ZN(n11644) );
  NAND4_X1 U14197 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        P3_U3161) );
  AOI21_X1 U14198 ( .B1(n11649), .B2(n11648), .A(n6654), .ZN(n11654) );
  AOI22_X1 U14199 ( .A1(n12192), .A2(n11731), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11651) );
  NAND2_X1 U14200 ( .A1(n11741), .A2(n12167), .ZN(n11650) );
  OAI211_X1 U14201 ( .C1(n12165), .C2(n11733), .A(n11651), .B(n11650), .ZN(
        n11652) );
  AOI21_X1 U14202 ( .B1(n12289), .B2(n11746), .A(n11652), .ZN(n11653) );
  OAI21_X1 U14203 ( .B1(n11654), .B2(n11748), .A(n11653), .ZN(P3_U3163) );
  INV_X1 U14204 ( .A(n12273), .ZN(n11666) );
  INV_X1 U14205 ( .A(n11656), .ZN(n11658) );
  NOR3_X1 U14206 ( .A1(n11655), .A2(n11658), .A3(n11657), .ZN(n11661) );
  INV_X1 U14207 ( .A(n11659), .ZN(n11660) );
  OAI21_X1 U14208 ( .B1(n11661), .B2(n11660), .A(n11730), .ZN(n11665) );
  AOI22_X1 U14209 ( .A1(n11971), .A2(n11731), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11662) );
  OAI21_X1 U14210 ( .B1(n12117), .B2(n11733), .A(n11662), .ZN(n11663) );
  AOI21_X1 U14211 ( .B1(n12118), .B2(n11741), .A(n11663), .ZN(n11664) );
  OAI211_X1 U14212 ( .C1(n11666), .C2(n11737), .A(n11665), .B(n11664), .ZN(
        P3_U3165) );
  XNOR2_X1 U14213 ( .A(n11667), .B(n12223), .ZN(n11668) );
  XNOR2_X1 U14214 ( .A(n11361), .B(n11668), .ZN(n11674) );
  NAND2_X1 U14215 ( .A1(n11741), .A2(n12241), .ZN(n11671) );
  NOR2_X1 U14216 ( .A1(n11669), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14215) );
  AOI21_X1 U14217 ( .B1(n11740), .B2(n11976), .A(n14215), .ZN(n11670) );
  OAI211_X1 U14218 ( .C1(n12239), .C2(n11744), .A(n11671), .B(n11670), .ZN(
        n11672) );
  AOI21_X1 U14219 ( .B1(n12309), .B2(n11746), .A(n11672), .ZN(n11673) );
  OAI21_X1 U14220 ( .B1(n11674), .B2(n11748), .A(n11673), .ZN(P3_U3166) );
  XNOR2_X1 U14221 ( .A(n11676), .B(n11675), .ZN(n11677) );
  NAND2_X1 U14222 ( .A1(n11677), .A2(n11730), .ZN(n11684) );
  AOI21_X1 U14223 ( .B1(n11740), .B2(n11980), .A(n11678), .ZN(n11683) );
  AOI22_X1 U14224 ( .A1(n11746), .A2(n11679), .B1(n11731), .B2(n14978), .ZN(
        n11682) );
  NAND2_X1 U14225 ( .A1(n11741), .A2(n11680), .ZN(n11681) );
  NAND4_X1 U14226 ( .A1(n11684), .A2(n11683), .A3(n11682), .A4(n11681), .ZN(
        P3_U3167) );
  INV_X1 U14227 ( .A(n11685), .ZN(n11687) );
  NOR3_X1 U14228 ( .A1(n11688), .A2(n11687), .A3(n11686), .ZN(n11689) );
  OAI21_X1 U14229 ( .B1(n11689), .B2(n11655), .A(n11730), .ZN(n11694) );
  NOR2_X1 U14230 ( .A1(n12154), .A2(n11744), .ZN(n11692) );
  OAI22_X1 U14231 ( .A1(n12125), .A2(n11733), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11690), .ZN(n11691) );
  AOI211_X1 U14232 ( .C1(n12132), .C2(n11741), .A(n11692), .B(n11691), .ZN(
        n11693) );
  OAI211_X1 U14233 ( .C1(n11737), .C2(n12279), .A(n11694), .B(n11693), .ZN(
        P3_U3169) );
  XNOR2_X1 U14234 ( .A(n6585), .B(n11695), .ZN(n11701) );
  NAND2_X1 U14235 ( .A1(n11741), .A2(n12180), .ZN(n11698) );
  AOI22_X1 U14236 ( .A1(n11731), .A2(n11975), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11697) );
  OAI211_X1 U14237 ( .C1(n12179), .C2(n11733), .A(n11698), .B(n11697), .ZN(
        n11699) );
  AOI21_X1 U14238 ( .B1(n12293), .B2(n11746), .A(n11699), .ZN(n11700) );
  OAI21_X1 U14239 ( .B1(n11701), .B2(n11748), .A(n11700), .ZN(P3_U3173) );
  INV_X1 U14240 ( .A(n11702), .ZN(n11703) );
  AOI21_X1 U14241 ( .B1(n11972), .B2(n11704), .A(n11703), .ZN(n11709) );
  AOI22_X1 U14242 ( .A1(n11974), .A2(n11731), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11706) );
  NAND2_X1 U14243 ( .A1(n11741), .A2(n12155), .ZN(n11705) );
  OAI211_X1 U14244 ( .C1(n12154), .C2(n11733), .A(n11706), .B(n11705), .ZN(
        n11707) );
  AOI21_X1 U14245 ( .B1(n12285), .B2(n11746), .A(n11707), .ZN(n11708) );
  OAI21_X1 U14246 ( .B1(n11709), .B2(n11748), .A(n11708), .ZN(P3_U3175) );
  XNOR2_X1 U14247 ( .A(n11712), .B(n11711), .ZN(n11713) );
  XNOR2_X1 U14248 ( .A(n11710), .B(n11713), .ZN(n11718) );
  NAND2_X1 U14249 ( .A1(n11741), .A2(n12211), .ZN(n11715) );
  INV_X1 U14250 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15242) );
  NOR2_X1 U14251 ( .A1(n15242), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14241) );
  AOI21_X1 U14252 ( .B1(n11740), .B2(n11975), .A(n14241), .ZN(n11714) );
  OAI211_X1 U14253 ( .C1(n12240), .C2(n11744), .A(n11715), .B(n11714), .ZN(
        n11716) );
  AOI21_X1 U14254 ( .B1(n12300), .B2(n11746), .A(n11716), .ZN(n11717) );
  OAI21_X1 U14255 ( .B1(n11718), .B2(n11748), .A(n11717), .ZN(P3_U3178) );
  AOI21_X1 U14256 ( .B1(n11720), .B2(n11719), .A(n11748), .ZN(n11722) );
  NAND2_X1 U14257 ( .A1(n11722), .A2(n11721), .ZN(n11727) );
  AOI21_X1 U14258 ( .B1(n11740), .B2(n14964), .A(n11723), .ZN(n11726) );
  AOI22_X1 U14259 ( .A1(n11746), .A2(n14960), .B1(n11731), .B2(n14965), .ZN(
        n11725) );
  NAND2_X1 U14260 ( .A1(n11741), .A2(n14961), .ZN(n11724) );
  NAND4_X1 U14261 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        P3_U3179) );
  AOI22_X1 U14262 ( .A1(n11970), .A2(n11731), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11732) );
  OAI21_X1 U14263 ( .B1(n12102), .B2(n11733), .A(n11732), .ZN(n11734) );
  AOI21_X1 U14264 ( .B1(n12108), .B2(n11741), .A(n11734), .ZN(n11735) );
  OAI211_X1 U14265 ( .C1(n12110), .C2(n11737), .A(n11736), .B(n11735), .ZN(
        P3_U3180) );
  XOR2_X1 U14266 ( .A(n11739), .B(n11738), .Z(n11749) );
  AOI22_X1 U14267 ( .A1(n11740), .A2(n12223), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11743) );
  NAND2_X1 U14268 ( .A1(n11741), .A2(n12255), .ZN(n11742) );
  OAI211_X1 U14269 ( .C1(n12251), .C2(n11744), .A(n11743), .B(n11742), .ZN(
        n11745) );
  AOI21_X1 U14270 ( .B1(n12313), .B2(n11746), .A(n11745), .ZN(n11747) );
  OAI21_X1 U14271 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(P3_U3181) );
  INV_X1 U14272 ( .A(n11750), .ZN(n11751) );
  NAND2_X1 U14273 ( .A1(n14038), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11753) );
  XNOR2_X1 U14274 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n11757) );
  INV_X1 U14275 ( .A(n11757), .ZN(n11754) );
  XNOR2_X1 U14276 ( .A(n11758), .B(n11754), .ZN(n12414) );
  NAND2_X1 U14277 ( .A1(n12414), .A2(n8307), .ZN(n11756) );
  INV_X1 U14278 ( .A(SI_30_), .ZN(n12416) );
  OR2_X1 U14279 ( .A1(n11764), .A2(n12416), .ZN(n11755) );
  NAND2_X1 U14280 ( .A1(n11758), .A2(n11757), .ZN(n11761) );
  NAND2_X1 U14281 ( .A1(n11759), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14282 ( .A1(n11761), .A2(n11760), .ZN(n11763) );
  INV_X1 U14283 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n15354) );
  XNOR2_X1 U14284 ( .A(n15354), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n11762) );
  XNOR2_X1 U14285 ( .A(n11763), .B(n11762), .ZN(n12412) );
  INV_X1 U14286 ( .A(SI_31_), .ZN(n12408) );
  NOR2_X1 U14287 ( .A1(n11764), .A2(n12408), .ZN(n11765) );
  AOI22_X1 U14288 ( .A1(n12261), .A2(n12065), .B1(n11766), .B2(n14285), .ZN(
        n11957) );
  OAI211_X1 U14289 ( .C1(n11771), .C2(n12065), .A(n11957), .B(n11951), .ZN(
        n11767) );
  INV_X1 U14290 ( .A(n12261), .ZN(n11773) );
  INV_X1 U14291 ( .A(n12065), .ZN(n11769) );
  INV_X1 U14292 ( .A(n12218), .ZN(n12216) );
  NAND3_X1 U14293 ( .A1(n11836), .A2(n11843), .A3(n11825), .ZN(n11778) );
  INV_X1 U14294 ( .A(n10388), .ZN(n11776) );
  NAND2_X1 U14295 ( .A1(n11776), .A2(n8753), .ZN(n11777) );
  OR2_X1 U14296 ( .A1(n11778), .A2(n11777), .ZN(n11783) );
  NOR2_X1 U14297 ( .A1(n11779), .A2(n8749), .ZN(n11781) );
  NAND4_X1 U14298 ( .A1(n11781), .A2(n14966), .A3(n11847), .A4(n11780), .ZN(
        n11782) );
  NOR2_X1 U14299 ( .A1(n11783), .A2(n11782), .ZN(n11785) );
  NAND4_X1 U14300 ( .A1(n11785), .A2(n11784), .A3(n7257), .A4(n14264), .ZN(
        n11786) );
  NOR4_X1 U14301 ( .A1(n12216), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11789) );
  NAND4_X1 U14302 ( .A1(n12208), .A2(n12247), .A3(n11789), .A4(n12235), .ZN(
        n11790) );
  NOR4_X1 U14303 ( .A1(n12190), .A2(n12176), .A3(n12140), .A4(n11790), .ZN(
        n11796) );
  INV_X1 U14304 ( .A(n11791), .ZN(n11936) );
  INV_X1 U14305 ( .A(n12100), .ZN(n12103) );
  INV_X1 U14306 ( .A(n12162), .ZN(n11794) );
  INV_X1 U14307 ( .A(n11793), .ZN(n11917) );
  NOR3_X1 U14308 ( .A1(n12114), .A2(n11794), .A3(n12151), .ZN(n11795) );
  NAND4_X1 U14309 ( .A1(n11796), .A2(n12103), .A3(n11795), .A4(n12126), .ZN(
        n11798) );
  NOR4_X1 U14310 ( .A1(n11798), .A2(n11797), .A3(n12077), .A4(n12089), .ZN(
        n11800) );
  INV_X1 U14311 ( .A(n11799), .ZN(n11954) );
  AND4_X1 U14312 ( .A1(n11957), .A2(n11800), .A3(n11954), .A4(n11775), .ZN(
        n11802) );
  NAND2_X1 U14313 ( .A1(n8748), .A2(n11806), .ZN(n11807) );
  MUX2_X1 U14314 ( .A(n11807), .B(n11806), .S(n11805), .Z(n11808) );
  MUX2_X1 U14315 ( .A(n11808), .B(n12342), .S(n11801), .Z(n11810) );
  MUX2_X1 U14316 ( .A(n11911), .B(n11810), .S(n11809), .Z(n11817) );
  NOR2_X1 U14317 ( .A1(n8748), .A2(n11948), .ZN(n11811) );
  NOR2_X1 U14318 ( .A1(n8749), .A2(n11811), .ZN(n11816) );
  NAND2_X1 U14319 ( .A1(n11819), .A2(n8751), .ZN(n11814) );
  NAND2_X1 U14320 ( .A1(n11818), .A2(n11812), .ZN(n11813) );
  MUX2_X1 U14321 ( .A(n11814), .B(n11813), .S(n11948), .Z(n11815) );
  AOI21_X1 U14322 ( .B1(n11817), .B2(n11816), .A(n11815), .ZN(n11827) );
  MUX2_X1 U14323 ( .A(n11819), .B(n11818), .S(n11911), .Z(n11820) );
  NAND2_X1 U14324 ( .A1(n11821), .A2(n11820), .ZN(n11826) );
  MUX2_X1 U14325 ( .A(n11823), .B(n11822), .S(n11948), .Z(n11824) );
  OAI211_X1 U14326 ( .C1(n11827), .C2(n11826), .A(n11825), .B(n11824), .ZN(
        n11839) );
  NAND2_X1 U14327 ( .A1(n11833), .A2(n11828), .ZN(n11831) );
  NAND2_X1 U14328 ( .A1(n11834), .A2(n11829), .ZN(n11830) );
  MUX2_X1 U14329 ( .A(n11831), .B(n11830), .S(n11948), .Z(n11832) );
  INV_X1 U14330 ( .A(n11832), .ZN(n11838) );
  MUX2_X1 U14331 ( .A(n11834), .B(n11833), .S(n11948), .Z(n11835) );
  NAND2_X1 U14332 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  AOI21_X1 U14333 ( .B1(n11839), .B2(n11838), .A(n11837), .ZN(n11849) );
  MUX2_X1 U14334 ( .A(n11841), .B(n11840), .S(n11911), .Z(n11842) );
  NAND2_X1 U14335 ( .A1(n11843), .A2(n11842), .ZN(n11848) );
  MUX2_X1 U14336 ( .A(n11845), .B(n11844), .S(n11948), .Z(n11846) );
  OAI211_X1 U14337 ( .C1(n11849), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        n11856) );
  AND2_X1 U14338 ( .A1(n11850), .A2(n11948), .ZN(n11852) );
  NOR2_X1 U14339 ( .A1(n11850), .A2(n11948), .ZN(n11851) );
  MUX2_X1 U14340 ( .A(n11852), .B(n11851), .S(n14951), .Z(n11853) );
  NOR2_X1 U14341 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  NAND2_X1 U14342 ( .A1(n11856), .A2(n11855), .ZN(n11860) );
  MUX2_X1 U14343 ( .A(n11858), .B(n11857), .S(n11948), .Z(n11859) );
  AOI21_X1 U14344 ( .B1(n11860), .B2(n11859), .A(n14278), .ZN(n11863) );
  AOI21_X1 U14345 ( .B1(n11871), .B2(n11861), .A(n11948), .ZN(n11862) );
  OAI21_X1 U14346 ( .B1(n11863), .B2(n11862), .A(n11865), .ZN(n11868) );
  NAND2_X1 U14347 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  NAND2_X1 U14348 ( .A1(n11866), .A2(n11948), .ZN(n11867) );
  NAND2_X1 U14349 ( .A1(n11868), .A2(n11867), .ZN(n11870) );
  OAI211_X1 U14350 ( .C1(n11871), .C2(n11911), .A(n11870), .B(n11869), .ZN(
        n11876) );
  MUX2_X1 U14351 ( .A(n11873), .B(n11872), .S(n11948), .Z(n11874) );
  NAND3_X1 U14352 ( .A1(n11876), .A2(n11875), .A3(n11874), .ZN(n11878) );
  NAND3_X1 U14353 ( .A1(n12316), .A2(n12251), .A3(n11948), .ZN(n11877) );
  NAND2_X1 U14354 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  NAND2_X1 U14355 ( .A1(n11879), .A2(n12247), .ZN(n11885) );
  INV_X1 U14356 ( .A(n12316), .ZN(n11880) );
  NAND3_X1 U14357 ( .A1(n12247), .A2(n11880), .A3(n11978), .ZN(n11882) );
  OAI211_X1 U14358 ( .C1(n12253), .C2(n12309), .A(n11882), .B(n11881), .ZN(
        n11883) );
  NAND2_X1 U14359 ( .A1(n11883), .A2(n11911), .ZN(n11884) );
  AOI21_X1 U14360 ( .B1(n11885), .B2(n11884), .A(n7231), .ZN(n11890) );
  AOI21_X1 U14361 ( .B1(n11887), .B2(n11886), .A(n11911), .ZN(n11889) );
  NAND2_X1 U14362 ( .A1(n12223), .A2(n11948), .ZN(n11888) );
  OAI22_X1 U14363 ( .A1(n11890), .A2(n11889), .B1(n12309), .B2(n11888), .ZN(
        n11896) );
  INV_X1 U14364 ( .A(n11892), .ZN(n11893) );
  NAND2_X1 U14365 ( .A1(n11897), .A2(n11893), .ZN(n11894) );
  NAND4_X1 U14366 ( .A1(n11903), .A2(n11948), .A3(n11895), .A4(n11894), .ZN(
        n11899) );
  AOI22_X1 U14367 ( .A1(n11896), .A2(n12218), .B1(n7269), .B2(n11899), .ZN(
        n11901) );
  NAND3_X1 U14368 ( .A1(n11902), .A2(n11911), .A3(n11897), .ZN(n11898) );
  NAND2_X1 U14369 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  OAI21_X1 U14370 ( .B1(n11901), .B2(n12202), .A(n11900), .ZN(n11906) );
  INV_X1 U14371 ( .A(n12176), .ZN(n11905) );
  MUX2_X1 U14372 ( .A(n11903), .B(n11902), .S(n11948), .Z(n11904) );
  NAND3_X1 U14373 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n11910) );
  NAND2_X1 U14374 ( .A1(n12293), .A2(n12166), .ZN(n11908) );
  MUX2_X1 U14375 ( .A(n11908), .B(n11907), .S(n11948), .Z(n11909) );
  NAND3_X1 U14376 ( .A1(n11910), .A2(n12162), .A3(n11909), .ZN(n11915) );
  INV_X1 U14377 ( .A(n12151), .ZN(n12149) );
  NAND2_X1 U14378 ( .A1(n11974), .A2(n11911), .ZN(n11913) );
  OR2_X1 U14379 ( .A1(n11974), .A2(n11911), .ZN(n11912) );
  MUX2_X1 U14380 ( .A(n11913), .B(n11912), .S(n12289), .Z(n11914) );
  NAND3_X1 U14381 ( .A1(n11915), .A2(n12149), .A3(n11914), .ZN(n11920) );
  MUX2_X1 U14382 ( .A(n11917), .B(n11916), .S(n11948), .Z(n11918) );
  NOR2_X1 U14383 ( .A1(n12140), .A2(n11918), .ZN(n11919) );
  NAND2_X1 U14384 ( .A1(n11920), .A2(n11919), .ZN(n11922) );
  NAND3_X1 U14385 ( .A1(n12281), .A2(n12154), .A3(n11948), .ZN(n11921) );
  NAND2_X1 U14386 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  NAND2_X1 U14387 ( .A1(n11923), .A2(n12126), .ZN(n11931) );
  INV_X1 U14388 ( .A(n12114), .ZN(n11930) );
  NAND2_X1 U14389 ( .A1(n11925), .A2(n11924), .ZN(n11926) );
  NAND2_X1 U14390 ( .A1(n11926), .A2(n11927), .ZN(n11928) );
  MUX2_X1 U14391 ( .A(n11928), .B(n11927), .S(n11948), .Z(n11929) );
  NAND3_X1 U14392 ( .A1(n11931), .A2(n11930), .A3(n11929), .ZN(n11935) );
  MUX2_X1 U14393 ( .A(n11933), .B(n11932), .S(n11948), .Z(n11934) );
  NAND3_X1 U14394 ( .A1(n11935), .A2(n12103), .A3(n11934), .ZN(n11940) );
  MUX2_X1 U14395 ( .A(n11937), .B(n11936), .S(n11948), .Z(n11938) );
  INV_X1 U14396 ( .A(n11938), .ZN(n11939) );
  AOI21_X1 U14397 ( .B1(n11940), .B2(n11939), .A(n12089), .ZN(n11949) );
  INV_X1 U14398 ( .A(n11941), .ZN(n11942) );
  NOR2_X1 U14399 ( .A1(n11949), .A2(n11942), .ZN(n11947) );
  NAND3_X1 U14400 ( .A1(n11944), .A2(n11948), .A3(n11943), .ZN(n11945) );
  OAI211_X1 U14401 ( .C1(n11947), .C2(n12077), .A(n11946), .B(n11945), .ZN(
        n11952) );
  INV_X1 U14402 ( .A(n12077), .ZN(n12074) );
  NAND3_X1 U14403 ( .A1(n11949), .A2(n11948), .A3(n12074), .ZN(n11950) );
  NAND3_X1 U14404 ( .A1(n11952), .A2(n11951), .A3(n11950), .ZN(n11955) );
  NAND3_X1 U14405 ( .A1(n11955), .A2(n11954), .A3(n11953), .ZN(n11958) );
  AOI21_X1 U14406 ( .B1(n11958), .B2(n11957), .A(n11956), .ZN(n11959) );
  MUX2_X1 U14407 ( .A(n14999), .B(n11960), .S(n11959), .Z(n11961) );
  AOI21_X1 U14408 ( .B1(n11963), .B2(n11962), .A(n11961), .ZN(n11969) );
  NAND3_X1 U14409 ( .A1(n11964), .A2(n14980), .A3(n6590), .ZN(n11965) );
  OAI211_X1 U14410 ( .C1(n11966), .C2(n11968), .A(n11965), .B(P3_B_REG_SCAN_IN), .ZN(n11967) );
  OAI21_X1 U14411 ( .B1(n11969), .B2(n11968), .A(n11967), .ZN(P3_U3296) );
  MUX2_X1 U14412 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12079), .S(n11973), .Z(
        P3_U3518) );
  MUX2_X1 U14413 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n11970), .S(n11973), .Z(
        P3_U3516) );
  MUX2_X1 U14414 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n11971), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14415 ( .A(n11972), .B(P3_DATAO_REG_22__SCAN_IN), .S(n11981), .Z(
        P3_U3513) );
  MUX2_X1 U14416 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n11974), .S(n11973), .Z(
        P3_U3512) );
  MUX2_X1 U14417 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12192), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14418 ( .A(n11975), .B(P3_DATAO_REG_19__SCAN_IN), .S(n11981), .Z(
        P3_U3510) );
  MUX2_X1 U14419 ( .A(n12224), .B(P3_DATAO_REG_18__SCAN_IN), .S(n11981), .Z(
        P3_U3509) );
  MUX2_X1 U14420 ( .A(n11976), .B(P3_DATAO_REG_17__SCAN_IN), .S(n11981), .Z(
        P3_U3508) );
  MUX2_X1 U14421 ( .A(n12223), .B(P3_DATAO_REG_16__SCAN_IN), .S(n11981), .Z(
        P3_U3507) );
  MUX2_X1 U14422 ( .A(n11977), .B(P3_DATAO_REG_15__SCAN_IN), .S(n11981), .Z(
        P3_U3506) );
  MUX2_X1 U14423 ( .A(n11978), .B(P3_DATAO_REG_14__SCAN_IN), .S(n11981), .Z(
        P3_U3505) );
  MUX2_X1 U14424 ( .A(n14258), .B(P3_DATAO_REG_13__SCAN_IN), .S(n11981), .Z(
        P3_U3504) );
  MUX2_X1 U14425 ( .A(n14259), .B(P3_DATAO_REG_11__SCAN_IN), .S(n11981), .Z(
        P3_U3502) );
  MUX2_X1 U14426 ( .A(n14275), .B(P3_DATAO_REG_10__SCAN_IN), .S(n11981), .Z(
        P3_U3501) );
  MUX2_X1 U14427 ( .A(n11979), .B(P3_DATAO_REG_8__SCAN_IN), .S(n11981), .Z(
        P3_U3499) );
  MUX2_X1 U14428 ( .A(n14964), .B(P3_DATAO_REG_7__SCAN_IN), .S(n11981), .Z(
        P3_U3498) );
  MUX2_X1 U14429 ( .A(n11980), .B(P3_DATAO_REG_6__SCAN_IN), .S(n11981), .Z(
        P3_U3497) );
  MUX2_X1 U14430 ( .A(n14965), .B(P3_DATAO_REG_5__SCAN_IN), .S(n11981), .Z(
        P3_U3496) );
  MUX2_X1 U14431 ( .A(n14978), .B(P3_DATAO_REG_4__SCAN_IN), .S(n11981), .Z(
        P3_U3495) );
  MUX2_X1 U14432 ( .A(n12329), .B(P3_DATAO_REG_3__SCAN_IN), .S(n11981), .Z(
        P3_U3494) );
  MUX2_X1 U14433 ( .A(n14979), .B(P3_DATAO_REG_2__SCAN_IN), .S(n11981), .Z(
        P3_U3493) );
  MUX2_X1 U14434 ( .A(n9319), .B(P3_DATAO_REG_1__SCAN_IN), .S(n11981), .Z(
        P3_U3492) );
  MUX2_X1 U14435 ( .A(n12337), .B(P3_DATAO_REG_0__SCAN_IN), .S(n11981), .Z(
        P3_U3491) );
  INV_X1 U14436 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n15368) );
  MUX2_X1 U14437 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n15368), .S(n12011), .Z(
        n12015) );
  MUX2_X1 U14438 ( .A(n12017), .B(P3_REG2_REG_10__SCAN_IN), .S(n12018), .Z(
        n14852) );
  NOR2_X1 U14439 ( .A1(n12016), .A2(n11985), .ZN(n11986) );
  INV_X1 U14440 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14872) );
  XOR2_X1 U14441 ( .A(n14880), .B(n11985), .Z(n14871) );
  INV_X1 U14442 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14263) );
  AOI22_X1 U14443 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12027), .B1(n14899), 
        .B2(n14263), .ZN(n14888) );
  NOR2_X1 U14444 ( .A1(n12031), .A2(n11987), .ZN(n11988) );
  XOR2_X1 U14445 ( .A(n14916), .B(n11987), .Z(n14907) );
  NOR2_X1 U14446 ( .A1(n11248), .A2(n14907), .ZN(n14906) );
  XNOR2_X1 U14447 ( .A(n14938), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n14924) );
  NOR2_X1 U14448 ( .A1(n14925), .A2(n14924), .ZN(n14923) );
  AOI21_X1 U14449 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n14938), .A(n14923), 
        .ZN(n11989) );
  NOR2_X1 U14450 ( .A1(n14185), .A2(n11989), .ZN(n11990) );
  INV_X1 U14451 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14194) );
  INV_X1 U14452 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U14453 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12045), .B1(n14211), 
        .B2(n11991), .ZN(n14201) );
  INV_X1 U14454 ( .A(n14200), .ZN(n11992) );
  NAND2_X1 U14455 ( .A1(n11993), .A2(n14229), .ZN(n11994) );
  OAI21_X1 U14456 ( .B1(n11993), .B2(n14229), .A(n11994), .ZN(n14219) );
  INV_X1 U14457 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14220) );
  INV_X1 U14458 ( .A(n11994), .ZN(n11995) );
  INV_X1 U14459 ( .A(n14239), .ZN(n12050) );
  INV_X1 U14460 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n15210) );
  AOI22_X1 U14461 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n12050), .B1(n14239), 
        .B2(n15210), .ZN(n14237) );
  NOR2_X1 U14462 ( .A1(n14238), .A2(n14237), .ZN(n14236) );
  AOI21_X1 U14463 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n14239), .A(n14236), 
        .ZN(n11996) );
  XOR2_X1 U14464 ( .A(n12015), .B(n11996), .Z(n12062) );
  INV_X1 U14465 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U14466 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n14239), .B1(n12050), 
        .B2(n12301), .ZN(n14244) );
  INV_X1 U14467 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12310) );
  XNOR2_X1 U14468 ( .A(n12045), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14203) );
  AND2_X1 U14469 ( .A1(n14938), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12006) );
  NOR2_X1 U14470 ( .A1(n14938), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11997) );
  OR2_X1 U14471 ( .A1(n12006), .A2(n11997), .ZN(n12034) );
  INV_X1 U14472 ( .A(n12034), .ZN(n14927) );
  INV_X1 U14473 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15274) );
  MUX2_X1 U14474 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n15274), .S(n14899), .Z(
        n14890) );
  INV_X1 U14475 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U14476 ( .A1(n12020), .A2(n11998), .ZN(n12000) );
  MUX2_X1 U14477 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n15070), .S(n12018), .Z(
        n14855) );
  NAND2_X1 U14478 ( .A1(n14856), .A2(n14855), .ZN(n14854) );
  NAND2_X1 U14479 ( .A1(n14880), .A2(n12001), .ZN(n12002) );
  XNOR2_X1 U14480 ( .A(n12001), .B(n12016), .ZN(n14874) );
  NAND2_X1 U14481 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n14874), .ZN(n14873) );
  NAND2_X1 U14482 ( .A1(n12002), .A2(n14873), .ZN(n14891) );
  NAND2_X1 U14483 ( .A1(n14890), .A2(n14891), .ZN(n14889) );
  NAND2_X1 U14484 ( .A1(n14916), .A2(n12003), .ZN(n12004) );
  XNOR2_X1 U14485 ( .A(n12031), .B(n12003), .ZN(n14909) );
  NAND2_X1 U14486 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n14909), .ZN(n14908) );
  NAND2_X1 U14487 ( .A1(n12004), .A2(n14908), .ZN(n14928) );
  NAND2_X1 U14488 ( .A1(n14927), .A2(n14928), .ZN(n14926) );
  INV_X1 U14489 ( .A(n14926), .ZN(n12005) );
  OR2_X1 U14490 ( .A1(n14185), .A2(n12007), .ZN(n12008) );
  XOR2_X1 U14491 ( .A(n12007), .B(n14185), .Z(n14187) );
  NAND2_X1 U14492 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14187), .ZN(n14186) );
  NAND2_X1 U14493 ( .A1(n12008), .A2(n14186), .ZN(n14204) );
  NAND2_X1 U14494 ( .A1(n14203), .A2(n14204), .ZN(n14202) );
  NAND2_X1 U14495 ( .A1(n12009), .A2(n14229), .ZN(n12010) );
  INV_X1 U14496 ( .A(n14229), .ZN(n12047) );
  XNOR2_X1 U14497 ( .A(n12009), .B(n12047), .ZN(n14222) );
  NAND2_X1 U14498 ( .A1(n14222), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14221) );
  NAND2_X1 U14499 ( .A1(n12010), .A2(n14221), .ZN(n14243) );
  XNOR2_X1 U14500 ( .A(n12011), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12013) );
  XNOR2_X1 U14501 ( .A(n12012), .B(n12013), .ZN(n12060) );
  INV_X1 U14502 ( .A(n12013), .ZN(n12014) );
  MUX2_X1 U14503 ( .A(n12015), .B(n12014), .S(n6590), .Z(n12053) );
  MUX2_X1 U14504 ( .A(n15210), .B(n12301), .S(n6590), .Z(n14246) );
  INV_X1 U14505 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12306) );
  MUX2_X1 U14506 ( .A(n14220), .B(n12306), .S(n6590), .Z(n12046) );
  NOR2_X1 U14507 ( .A1(n12046), .A2(n12047), .ZN(n12048) );
  MUX2_X1 U14508 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n6590), .Z(n12043) );
  INV_X1 U14509 ( .A(n12043), .ZN(n12044) );
  MUX2_X1 U14510 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6590), .Z(n12025) );
  XNOR2_X1 U14511 ( .A(n12025), .B(n12016), .ZN(n14877) );
  MUX2_X1 U14512 ( .A(n12017), .B(n15070), .S(n6590), .Z(n12019) );
  NAND2_X1 U14513 ( .A1(n12019), .A2(n14865), .ZN(n12024) );
  XNOR2_X1 U14514 ( .A(n12019), .B(n12018), .ZN(n14863) );
  OR2_X1 U14515 ( .A1(n12021), .A2(n12020), .ZN(n12023) );
  NAND2_X1 U14516 ( .A1(n12023), .A2(n12022), .ZN(n14862) );
  NAND2_X1 U14517 ( .A1(n14863), .A2(n14862), .ZN(n14861) );
  NAND2_X1 U14518 ( .A1(n12024), .A2(n14861), .ZN(n14876) );
  NOR2_X1 U14519 ( .A1(n12025), .A2(n14880), .ZN(n12026) );
  AOI21_X1 U14520 ( .B1(n14877), .B2(n14876), .A(n12026), .ZN(n14896) );
  MUX2_X1 U14521 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6590), .Z(n12028) );
  XNOR2_X1 U14522 ( .A(n12028), .B(n12027), .ZN(n14895) );
  NAND2_X1 U14523 ( .A1(n14896), .A2(n14895), .ZN(n14894) );
  NAND2_X1 U14524 ( .A1(n12028), .A2(n14899), .ZN(n12029) );
  NAND2_X1 U14525 ( .A1(n14894), .A2(n12029), .ZN(n14912) );
  MUX2_X1 U14526 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6590), .Z(n12030) );
  XNOR2_X1 U14527 ( .A(n12030), .B(n14916), .ZN(n14911) );
  INV_X1 U14528 ( .A(n12030), .ZN(n12032) );
  NAND2_X1 U14529 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  NAND2_X1 U14530 ( .A1(n14914), .A2(n12033), .ZN(n14934) );
  MUX2_X1 U14531 ( .A(n14924), .B(n12034), .S(n6590), .Z(n14935) );
  MUX2_X1 U14532 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n6590), .Z(n12035) );
  NAND2_X1 U14533 ( .A1(n12035), .A2(n14938), .ZN(n12036) );
  NAND2_X1 U14534 ( .A1(n14931), .A2(n12036), .ZN(n12040) );
  XNOR2_X1 U14535 ( .A(n12040), .B(n14185), .ZN(n14189) );
  INV_X1 U14536 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12314) );
  MUX2_X1 U14537 ( .A(n14194), .B(n12314), .S(n6590), .Z(n14188) );
  INV_X1 U14538 ( .A(n14188), .ZN(n12038) );
  NAND2_X1 U14539 ( .A1(n14189), .A2(n12038), .ZN(n12042) );
  NAND2_X1 U14540 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  NAND2_X1 U14541 ( .A1(n12042), .A2(n12041), .ZN(n14208) );
  XNOR2_X1 U14542 ( .A(n12043), .B(n12045), .ZN(n14207) );
  NAND2_X1 U14543 ( .A1(n14208), .A2(n14207), .ZN(n14206) );
  OAI21_X1 U14544 ( .B1(n12045), .B2(n12044), .A(n14206), .ZN(n14225) );
  AOI21_X1 U14545 ( .B1(n12047), .B2(n12046), .A(n12048), .ZN(n14224) );
  AND2_X1 U14546 ( .A1(n14225), .A2(n14224), .ZN(n14226) );
  NOR2_X1 U14547 ( .A1(n12048), .A2(n14226), .ZN(n12049) );
  XNOR2_X1 U14548 ( .A(n14239), .B(n12049), .ZN(n14247) );
  NAND2_X1 U14549 ( .A1(n14246), .A2(n14247), .ZN(n14245) );
  NAND2_X1 U14550 ( .A1(n12050), .A2(n12049), .ZN(n12051) );
  NAND2_X1 U14551 ( .A1(n14245), .A2(n12051), .ZN(n12052) );
  XNOR2_X1 U14552 ( .A(n12053), .B(n12052), .ZN(n12054) );
  NOR2_X1 U14553 ( .A1(n12054), .A2(n14933), .ZN(n12059) );
  NAND2_X1 U14554 ( .A1(n14860), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12055) );
  OAI211_X1 U14555 ( .C1(n14939), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n12058) );
  OAI21_X1 U14556 ( .B1(n12062), .B2(n14945), .A(n12061), .ZN(P3_U3201) );
  INV_X1 U14557 ( .A(n12063), .ZN(n12064) );
  NAND2_X1 U14558 ( .A1(n12065), .A2(n12064), .ZN(n12260) );
  INV_X1 U14559 ( .A(n12260), .ZN(n14284) );
  NOR2_X1 U14560 ( .A1(n12066), .A2(n15010), .ZN(n12070) );
  AOI21_X1 U14561 ( .B1(n14284), .B2(n14995), .A(n12070), .ZN(n14255) );
  NAND2_X1 U14562 ( .A1(n15018), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12067) );
  OAI211_X1 U14563 ( .C1(n12261), .C2(n12134), .A(n14255), .B(n12067), .ZN(
        P3_U3202) );
  NAND2_X1 U14564 ( .A1(n12068), .A2(n14995), .ZN(n12072) );
  NOR2_X1 U14565 ( .A1(n6633), .A2(n14268), .ZN(n12069) );
  AOI211_X1 U14566 ( .C1(n15018), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12070), 
        .B(n12069), .ZN(n12071) );
  OAI211_X1 U14567 ( .C1(n12073), .C2(n14269), .A(n12072), .B(n12071), .ZN(
        P3_U3204) );
  XNOR2_X1 U14568 ( .A(n12075), .B(n12074), .ZN(n12352) );
  OAI211_X1 U14569 ( .C1(n12078), .C2(n12077), .A(n12076), .B(n14982), .ZN(
        n12081) );
  NAND2_X1 U14570 ( .A1(n12079), .A2(n14980), .ZN(n12080) );
  OAI211_X1 U14571 ( .C1(n12082), .C2(n12254), .A(n12081), .B(n12080), .ZN(
        n12262) );
  NAND2_X1 U14572 ( .A1(n12262), .A2(n14995), .ZN(n12088) );
  INV_X1 U14573 ( .A(n12083), .ZN(n12085) );
  INV_X1 U14574 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12084) );
  OAI22_X1 U14575 ( .A1(n12085), .A2(n15010), .B1(n14995), .B2(n12084), .ZN(
        n12086) );
  AOI21_X1 U14576 ( .B1(n12263), .B2(n14253), .A(n12086), .ZN(n12087) );
  OAI211_X1 U14577 ( .C1(n14269), .C2(n12352), .A(n12088), .B(n12087), .ZN(
        P3_U3205) );
  XNOR2_X1 U14578 ( .A(n12090), .B(n12089), .ZN(n12356) );
  XNOR2_X1 U14579 ( .A(n12091), .B(n7092), .ZN(n12092) );
  OAI222_X1 U14580 ( .A1(n12252), .A2(n12117), .B1(n12254), .B2(n12093), .C1(
        n12092), .C2(n12249), .ZN(n12265) );
  NAND2_X1 U14581 ( .A1(n12265), .A2(n14995), .ZN(n12099) );
  INV_X1 U14582 ( .A(n12094), .ZN(n12096) );
  INV_X1 U14583 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12095) );
  OAI22_X1 U14584 ( .A1(n12096), .A2(n15010), .B1(n14995), .B2(n12095), .ZN(
        n12097) );
  AOI21_X1 U14585 ( .B1(n12266), .B2(n14253), .A(n12097), .ZN(n12098) );
  OAI211_X1 U14586 ( .C1(n14269), .C2(n12356), .A(n12099), .B(n12098), .ZN(
        P3_U3206) );
  XNOR2_X1 U14587 ( .A(n12101), .B(n12100), .ZN(n12269) );
  OAI22_X1 U14588 ( .A1(n12102), .A2(n12254), .B1(n12125), .B2(n12252), .ZN(
        n12107) );
  XNOR2_X1 U14589 ( .A(n12104), .B(n12103), .ZN(n12105) );
  NOR2_X1 U14590 ( .A1(n12105), .A2(n12249), .ZN(n12106) );
  AOI211_X1 U14591 ( .C1(n12131), .C2(n12269), .A(n12107), .B(n12106), .ZN(
        n12271) );
  AOI22_X1 U14592 ( .A1(n12108), .A2(n14991), .B1(n15018), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12109) );
  OAI21_X1 U14593 ( .B1(n12110), .B2(n12134), .A(n12109), .ZN(n12111) );
  AOI21_X1 U14594 ( .B1(n12269), .B2(n14971), .A(n12111), .ZN(n12112) );
  OAI21_X1 U14595 ( .B1(n12271), .B2(n15018), .A(n12112), .ZN(P3_U3207) );
  XNOR2_X1 U14596 ( .A(n12113), .B(n12114), .ZN(n12361) );
  XNOR2_X1 U14597 ( .A(n12115), .B(n12114), .ZN(n12116) );
  OAI222_X1 U14598 ( .A1(n12254), .A2(n12117), .B1(n12252), .B2(n12139), .C1(
        n12116), .C2(n12249), .ZN(n12272) );
  NAND2_X1 U14599 ( .A1(n12272), .A2(n14995), .ZN(n12123) );
  INV_X1 U14600 ( .A(n12118), .ZN(n12120) );
  INV_X1 U14601 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12119) );
  OAI22_X1 U14602 ( .A1(n12120), .A2(n15010), .B1(n14995), .B2(n12119), .ZN(
        n12121) );
  AOI21_X1 U14603 ( .B1(n12273), .B2(n14253), .A(n12121), .ZN(n12122) );
  OAI211_X1 U14604 ( .C1(n14269), .C2(n12361), .A(n12123), .B(n12122), .ZN(
        P3_U3208) );
  OAI22_X1 U14605 ( .A1(n12125), .A2(n12254), .B1(n12154), .B2(n12252), .ZN(
        n12130) );
  XNOR2_X1 U14606 ( .A(n12127), .B(n12126), .ZN(n12128) );
  NOR2_X1 U14607 ( .A1(n12128), .A2(n12249), .ZN(n12129) );
  AOI211_X1 U14608 ( .C1(n12131), .C2(n12276), .A(n12130), .B(n12129), .ZN(
        n12278) );
  AOI22_X1 U14609 ( .A1(n15018), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12132), 
        .B2(n14991), .ZN(n12133) );
  OAI21_X1 U14610 ( .B1(n12279), .B2(n12134), .A(n12133), .ZN(n12135) );
  AOI21_X1 U14611 ( .B1(n12276), .B2(n14971), .A(n12135), .ZN(n12136) );
  OAI21_X1 U14612 ( .B1(n12278), .B2(n15018), .A(n12136), .ZN(P3_U3209) );
  XNOR2_X1 U14613 ( .A(n12137), .B(n12140), .ZN(n12138) );
  OAI222_X1 U14614 ( .A1(n12254), .A2(n12139), .B1(n12252), .B2(n12165), .C1(
        n12138), .C2(n12249), .ZN(n12280) );
  NAND2_X1 U14615 ( .A1(n12141), .A2(n12140), .ZN(n12142) );
  NAND2_X1 U14616 ( .A1(n12143), .A2(n12142), .ZN(n12366) );
  AOI22_X1 U14617 ( .A1(n15018), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n14991), 
        .B2(n12144), .ZN(n12146) );
  NAND2_X1 U14618 ( .A1(n12281), .A2(n14253), .ZN(n12145) );
  OAI211_X1 U14619 ( .C1(n12366), .C2(n14269), .A(n12146), .B(n12145), .ZN(
        n12147) );
  AOI21_X1 U14620 ( .B1(n12280), .B2(n14995), .A(n12147), .ZN(n12148) );
  INV_X1 U14621 ( .A(n12148), .ZN(P3_U3210) );
  XNOR2_X1 U14622 ( .A(n12150), .B(n12149), .ZN(n12370) );
  XNOR2_X1 U14623 ( .A(n12152), .B(n12151), .ZN(n12153) );
  OAI222_X1 U14624 ( .A1(n12252), .A2(n12179), .B1(n12254), .B2(n12154), .C1(
        n12249), .C2(n12153), .ZN(n12284) );
  NAND2_X1 U14625 ( .A1(n12284), .A2(n14995), .ZN(n12160) );
  INV_X1 U14626 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12157) );
  INV_X1 U14627 ( .A(n12155), .ZN(n12156) );
  OAI22_X1 U14628 ( .A1(n14995), .A2(n12157), .B1(n12156), .B2(n15010), .ZN(
        n12158) );
  AOI21_X1 U14629 ( .B1(n12285), .B2(n14253), .A(n12158), .ZN(n12159) );
  OAI211_X1 U14630 ( .C1(n14269), .C2(n12370), .A(n12160), .B(n12159), .ZN(
        P3_U3211) );
  XNOR2_X1 U14631 ( .A(n12161), .B(n12162), .ZN(n12374) );
  XNOR2_X1 U14632 ( .A(n12163), .B(n12162), .ZN(n12164) );
  OAI222_X1 U14633 ( .A1(n12252), .A2(n12166), .B1(n12254), .B2(n12165), .C1(
        n12249), .C2(n12164), .ZN(n12288) );
  NAND2_X1 U14634 ( .A1(n12288), .A2(n14995), .ZN(n12172) );
  INV_X1 U14635 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12169) );
  INV_X1 U14636 ( .A(n12167), .ZN(n12168) );
  OAI22_X1 U14637 ( .A1(n14995), .A2(n12169), .B1(n12168), .B2(n15010), .ZN(
        n12170) );
  AOI21_X1 U14638 ( .B1(n12289), .B2(n14253), .A(n12170), .ZN(n12171) );
  OAI211_X1 U14639 ( .C1(n14269), .C2(n12374), .A(n12172), .B(n12171), .ZN(
        P3_U3212) );
  NAND2_X1 U14640 ( .A1(n12173), .A2(n12176), .ZN(n12174) );
  NAND2_X1 U14641 ( .A1(n12175), .A2(n12174), .ZN(n12377) );
  XNOR2_X1 U14642 ( .A(n12177), .B(n12176), .ZN(n12178) );
  OAI222_X1 U14643 ( .A1(n12254), .A2(n12179), .B1(n12252), .B2(n12210), .C1(
        n12249), .C2(n12178), .ZN(n12292) );
  NAND2_X1 U14644 ( .A1(n12292), .A2(n14995), .ZN(n12185) );
  INV_X1 U14645 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12182) );
  INV_X1 U14646 ( .A(n12180), .ZN(n12181) );
  OAI22_X1 U14647 ( .A1(n14995), .A2(n12182), .B1(n12181), .B2(n15010), .ZN(
        n12183) );
  AOI21_X1 U14648 ( .B1(n12293), .B2(n14253), .A(n12183), .ZN(n12184) );
  OAI211_X1 U14649 ( .C1(n14269), .C2(n12377), .A(n12185), .B(n12184), .ZN(
        P3_U3213) );
  INV_X1 U14650 ( .A(n12186), .ZN(n12187) );
  AOI21_X1 U14651 ( .B1(n12190), .B2(n12188), .A(n12187), .ZN(n12381) );
  NAND2_X1 U14652 ( .A1(n12189), .A2(n14982), .ZN(n12195) );
  AOI21_X1 U14653 ( .B1(n12206), .B2(n12191), .A(n12190), .ZN(n12194) );
  AOI22_X1 U14654 ( .A1(n12192), .A2(n14977), .B1(n14980), .B2(n12224), .ZN(
        n12193) );
  OAI21_X1 U14655 ( .B1(n12195), .B2(n12194), .A(n12193), .ZN(n12296) );
  NAND2_X1 U14656 ( .A1(n12296), .A2(n14995), .ZN(n12201) );
  INV_X1 U14657 ( .A(n12197), .ZN(n12198) );
  OAI22_X1 U14658 ( .A1(n14995), .A2(n15368), .B1(n12198), .B2(n15010), .ZN(
        n12199) );
  AOI21_X1 U14659 ( .B1(n8535), .B2(n14253), .A(n12199), .ZN(n12200) );
  OAI211_X1 U14660 ( .C1(n14269), .C2(n12381), .A(n12201), .B(n12200), .ZN(
        P3_U3214) );
  NAND2_X1 U14661 ( .A1(n12203), .A2(n12202), .ZN(n12204) );
  NAND2_X1 U14662 ( .A1(n12205), .A2(n12204), .ZN(n12385) );
  INV_X1 U14663 ( .A(n12206), .ZN(n12207) );
  AOI21_X1 U14664 ( .B1(n12208), .B2(n6702), .A(n12207), .ZN(n12209) );
  OAI222_X1 U14665 ( .A1(n12252), .A2(n12240), .B1(n12254), .B2(n12210), .C1(
        n12249), .C2(n12209), .ZN(n12299) );
  NAND2_X1 U14666 ( .A1(n12299), .A2(n14995), .ZN(n12215) );
  INV_X1 U14667 ( .A(n12211), .ZN(n12212) );
  OAI22_X1 U14668 ( .A1(n14995), .A2(n15210), .B1(n12212), .B2(n15010), .ZN(
        n12213) );
  AOI21_X1 U14669 ( .B1(n12300), .B2(n14253), .A(n12213), .ZN(n12214) );
  OAI211_X1 U14670 ( .C1(n14269), .C2(n12385), .A(n12215), .B(n12214), .ZN(
        P3_U3215) );
  XNOR2_X1 U14671 ( .A(n12217), .B(n12216), .ZN(n12389) );
  NAND2_X1 U14672 ( .A1(n12219), .A2(n12218), .ZN(n12220) );
  NAND2_X1 U14673 ( .A1(n12220), .A2(n14982), .ZN(n12221) );
  OR2_X1 U14674 ( .A1(n12222), .A2(n12221), .ZN(n12226) );
  AOI22_X1 U14675 ( .A1(n14977), .A2(n12224), .B1(n12223), .B2(n14980), .ZN(
        n12225) );
  NAND2_X1 U14676 ( .A1(n12226), .A2(n12225), .ZN(n12305) );
  NAND2_X1 U14677 ( .A1(n12305), .A2(n14995), .ZN(n12231) );
  INV_X1 U14678 ( .A(n12227), .ZN(n12228) );
  OAI22_X1 U14679 ( .A1(n14995), .A2(n14220), .B1(n12228), .B2(n15010), .ZN(
        n12229) );
  AOI21_X1 U14680 ( .B1(n12303), .B2(n14253), .A(n12229), .ZN(n12230) );
  OAI211_X1 U14681 ( .C1(n14269), .C2(n12389), .A(n12231), .B(n12230), .ZN(
        P3_U3216) );
  XNOR2_X1 U14682 ( .A(n12232), .B(n7233), .ZN(n12393) );
  INV_X1 U14683 ( .A(n12233), .ZN(n12237) );
  AOI22_X1 U14684 ( .A1(n12237), .A2(n12236), .B1(n12235), .B2(n12234), .ZN(
        n12238) );
  OAI222_X1 U14685 ( .A1(n12254), .A2(n12240), .B1(n12252), .B2(n12239), .C1(
        n12249), .C2(n12238), .ZN(n12308) );
  NAND2_X1 U14686 ( .A1(n12308), .A2(n14995), .ZN(n12245) );
  INV_X1 U14687 ( .A(n12241), .ZN(n12242) );
  OAI22_X1 U14688 ( .A1(n14995), .A2(n11991), .B1(n12242), .B2(n15010), .ZN(
        n12243) );
  AOI21_X1 U14689 ( .B1(n12309), .B2(n14253), .A(n12243), .ZN(n12244) );
  OAI211_X1 U14690 ( .C1(n14269), .C2(n12393), .A(n12245), .B(n12244), .ZN(
        P3_U3217) );
  XNOR2_X1 U14691 ( .A(n12246), .B(n7229), .ZN(n12397) );
  XOR2_X1 U14692 ( .A(n12248), .B(n12247), .Z(n12250) );
  OAI222_X1 U14693 ( .A1(n12254), .A2(n12253), .B1(n12252), .B2(n12251), .C1(
        n12250), .C2(n12249), .ZN(n12312) );
  NAND2_X1 U14694 ( .A1(n12312), .A2(n14995), .ZN(n12259) );
  INV_X1 U14695 ( .A(n12255), .ZN(n12256) );
  OAI22_X1 U14696 ( .A1(n14995), .A2(n14194), .B1(n12256), .B2(n15010), .ZN(
        n12257) );
  AOI21_X1 U14697 ( .B1(n12313), .B2(n14253), .A(n12257), .ZN(n12258) );
  OAI211_X1 U14698 ( .C1(n14269), .C2(n12397), .A(n12259), .B(n12258), .ZN(
        P3_U3218) );
  OAI21_X1 U14699 ( .B1(n12261), .B2(n14988), .A(n12260), .ZN(n12348) );
  MUX2_X1 U14700 ( .A(P3_REG1_REG_31__SCAN_IN), .B(n12348), .S(n15072), .Z(
        P3_U3490) );
  AOI21_X1 U14701 ( .B1(n15043), .B2(n12263), .A(n12262), .ZN(n12349) );
  MUX2_X1 U14702 ( .A(n15276), .B(n12349), .S(n15072), .Z(n12264) );
  OAI21_X1 U14703 ( .B1(n12325), .B2(n12352), .A(n12264), .ZN(P3_U3487) );
  AOI21_X1 U14704 ( .B1(n15043), .B2(n12266), .A(n12265), .ZN(n12353) );
  MUX2_X1 U14705 ( .A(n15246), .B(n12353), .S(n15072), .Z(n12267) );
  OAI21_X1 U14706 ( .B1(n12325), .B2(n12356), .A(n12267), .ZN(P3_U3486) );
  AOI22_X1 U14707 ( .A1(n12269), .A2(n15049), .B1(n15043), .B2(n12268), .ZN(
        n12270) );
  NAND2_X1 U14708 ( .A1(n12271), .A2(n12270), .ZN(n12357) );
  MUX2_X1 U14709 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12357), .S(n15072), .Z(
        P3_U3485) );
  INV_X1 U14710 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12274) );
  AOI21_X1 U14711 ( .B1(n15043), .B2(n12273), .A(n12272), .ZN(n12358) );
  MUX2_X1 U14712 ( .A(n12274), .B(n12358), .S(n15072), .Z(n12275) );
  OAI21_X1 U14713 ( .B1(n12325), .B2(n12361), .A(n12275), .ZN(P3_U3484) );
  NAND2_X1 U14714 ( .A1(n12276), .A2(n15049), .ZN(n12277) );
  OAI211_X1 U14715 ( .C1(n12279), .C2(n14988), .A(n12278), .B(n12277), .ZN(
        n12362) );
  MUX2_X1 U14716 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12362), .S(n15072), .Z(
        P3_U3483) );
  INV_X1 U14717 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12282) );
  AOI21_X1 U14718 ( .B1(n15043), .B2(n12281), .A(n12280), .ZN(n12363) );
  MUX2_X1 U14719 ( .A(n12282), .B(n12363), .S(n15072), .Z(n12283) );
  OAI21_X1 U14720 ( .B1(n12325), .B2(n12366), .A(n12283), .ZN(P3_U3482) );
  INV_X1 U14721 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12286) );
  AOI21_X1 U14722 ( .B1(n15043), .B2(n12285), .A(n12284), .ZN(n12367) );
  MUX2_X1 U14723 ( .A(n12286), .B(n12367), .S(n15072), .Z(n12287) );
  OAI21_X1 U14724 ( .B1(n12370), .B2(n12325), .A(n12287), .ZN(P3_U3481) );
  INV_X1 U14725 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12290) );
  AOI21_X1 U14726 ( .B1(n15043), .B2(n12289), .A(n12288), .ZN(n12371) );
  MUX2_X1 U14727 ( .A(n12290), .B(n12371), .S(n15072), .Z(n12291) );
  OAI21_X1 U14728 ( .B1(n12325), .B2(n12374), .A(n12291), .ZN(P3_U3480) );
  INV_X1 U14729 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12294) );
  AOI21_X1 U14730 ( .B1(n15043), .B2(n12293), .A(n12292), .ZN(n12375) );
  MUX2_X1 U14731 ( .A(n12294), .B(n12375), .S(n15072), .Z(n12295) );
  OAI21_X1 U14732 ( .B1(n12325), .B2(n12377), .A(n12295), .ZN(P3_U3479) );
  INV_X1 U14733 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12297) );
  AOI21_X1 U14734 ( .B1(n15043), .B2(n8535), .A(n12296), .ZN(n12378) );
  MUX2_X1 U14735 ( .A(n12297), .B(n12378), .S(n15072), .Z(n12298) );
  OAI21_X1 U14736 ( .B1(n12381), .B2(n12325), .A(n12298), .ZN(P3_U3478) );
  AOI21_X1 U14737 ( .B1(n15043), .B2(n12300), .A(n12299), .ZN(n12382) );
  MUX2_X1 U14738 ( .A(n12301), .B(n12382), .S(n15072), .Z(n12302) );
  OAI21_X1 U14739 ( .B1(n12325), .B2(n12385), .A(n12302), .ZN(P3_U3477) );
  AND2_X1 U14740 ( .A1(n12303), .A2(n15043), .ZN(n12304) );
  NOR2_X1 U14741 ( .A1(n12305), .A2(n12304), .ZN(n12386) );
  MUX2_X1 U14742 ( .A(n12306), .B(n12386), .S(n15072), .Z(n12307) );
  OAI21_X1 U14743 ( .B1(n12325), .B2(n12389), .A(n12307), .ZN(P3_U3476) );
  AOI21_X1 U14744 ( .B1(n15043), .B2(n12309), .A(n12308), .ZN(n12390) );
  MUX2_X1 U14745 ( .A(n12310), .B(n12390), .S(n15072), .Z(n12311) );
  OAI21_X1 U14746 ( .B1(n12393), .B2(n12325), .A(n12311), .ZN(P3_U3475) );
  AOI21_X1 U14747 ( .B1(n15043), .B2(n12313), .A(n12312), .ZN(n12394) );
  MUX2_X1 U14748 ( .A(n12314), .B(n12394), .S(n15072), .Z(n12315) );
  OAI21_X1 U14749 ( .B1(n12325), .B2(n12397), .A(n12315), .ZN(P3_U3474) );
  INV_X1 U14750 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U14751 ( .A1(n12316), .A2(n15043), .ZN(n12317) );
  AND2_X1 U14752 ( .A1(n12318), .A2(n12317), .ZN(n12399) );
  MUX2_X1 U14753 ( .A(n12319), .B(n12399), .S(n15072), .Z(n12320) );
  OAI21_X1 U14754 ( .B1(n12401), .B2(n12325), .A(n12320), .ZN(P3_U3473) );
  INV_X1 U14755 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12323) );
  AOI21_X1 U14756 ( .B1(n15043), .B2(n12322), .A(n12321), .ZN(n12402) );
  MUX2_X1 U14757 ( .A(n12323), .B(n12402), .S(n15072), .Z(n12324) );
  OAI21_X1 U14758 ( .B1(n12325), .B2(n12406), .A(n12324), .ZN(P3_U3472) );
  XNOR2_X1 U14759 ( .A(n12326), .B(n8749), .ZN(n14997) );
  OR2_X1 U14760 ( .A1(n14997), .A2(n15038), .ZN(n12332) );
  XNOR2_X1 U14761 ( .A(n12327), .B(n8749), .ZN(n12328) );
  NAND2_X1 U14762 ( .A1(n12328), .A2(n14982), .ZN(n12331) );
  AOI22_X1 U14763 ( .A1(n14980), .A2(n9319), .B1(n12329), .B2(n14977), .ZN(
        n12330) );
  NAND3_X1 U14764 ( .A1(n12332), .A2(n12331), .A3(n12330), .ZN(n15000) );
  INV_X1 U14765 ( .A(n15049), .ZN(n15037) );
  NAND2_X1 U14766 ( .A1(n12333), .A2(n15043), .ZN(n14998) );
  OAI21_X1 U14767 ( .B1(n14997), .B2(n15037), .A(n14998), .ZN(n12334) );
  NOR2_X1 U14768 ( .A1(n15000), .A2(n12334), .ZN(n15021) );
  INV_X1 U14769 ( .A(n15021), .ZN(n12335) );
  MUX2_X1 U14770 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n12335), .S(n15072), .Z(
        P3_U3461) );
  XNOR2_X1 U14771 ( .A(n12336), .B(n10388), .ZN(n12341) );
  NAND2_X1 U14772 ( .A1(n12337), .A2(n14980), .ZN(n12339) );
  NAND2_X1 U14773 ( .A1(n14979), .A2(n14977), .ZN(n12338) );
  NAND2_X1 U14774 ( .A1(n12339), .A2(n12338), .ZN(n12340) );
  AOI21_X1 U14775 ( .B1(n12341), .B2(n14982), .A(n12340), .ZN(n12344) );
  XNOR2_X1 U14776 ( .A(n10388), .B(n12342), .ZN(n15012) );
  OR2_X1 U14777 ( .A1(n15012), .A2(n15038), .ZN(n12343) );
  AND2_X1 U14778 ( .A1(n12344), .A2(n12343), .ZN(n15006) );
  INV_X1 U14779 ( .A(n15012), .ZN(n12345) );
  AND2_X1 U14780 ( .A1(n10393), .A2(n15043), .ZN(n15009) );
  AOI21_X1 U14781 ( .B1(n12345), .B2(n15049), .A(n15009), .ZN(n12346) );
  AND2_X1 U14782 ( .A1(n15006), .A2(n12346), .ZN(n15019) );
  INV_X1 U14783 ( .A(n15019), .ZN(n12347) );
  MUX2_X1 U14784 ( .A(n12347), .B(P3_REG1_REG_1__SCAN_IN), .S(n8777), .Z(
        P3_U3460) );
  MUX2_X1 U14785 ( .A(P3_REG0_REG_31__SCAN_IN), .B(n12348), .S(n15055), .Z(
        P3_U3458) );
  INV_X1 U14786 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12350) );
  MUX2_X1 U14787 ( .A(n12350), .B(n12349), .S(n15055), .Z(n12351) );
  OAI21_X1 U14788 ( .B1(n12352), .B2(n12405), .A(n12351), .ZN(P3_U3455) );
  INV_X1 U14789 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12354) );
  MUX2_X1 U14790 ( .A(n12354), .B(n12353), .S(n15055), .Z(n12355) );
  OAI21_X1 U14791 ( .B1(n12356), .B2(n12405), .A(n12355), .ZN(P3_U3454) );
  MUX2_X1 U14792 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12357), .S(n15055), .Z(
        P3_U3453) );
  MUX2_X1 U14793 ( .A(n12359), .B(n12358), .S(n15055), .Z(n12360) );
  OAI21_X1 U14794 ( .B1(n12361), .B2(n12405), .A(n12360), .ZN(P3_U3452) );
  MUX2_X1 U14795 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12362), .S(n15055), .Z(
        P3_U3451) );
  MUX2_X1 U14796 ( .A(n12364), .B(n12363), .S(n15055), .Z(n12365) );
  OAI21_X1 U14797 ( .B1(n12366), .B2(n12405), .A(n12365), .ZN(P3_U3450) );
  MUX2_X1 U14798 ( .A(n12368), .B(n12367), .S(n15055), .Z(n12369) );
  OAI21_X1 U14799 ( .B1(n12370), .B2(n12405), .A(n12369), .ZN(P3_U3449) );
  MUX2_X1 U14800 ( .A(n12372), .B(n12371), .S(n15055), .Z(n12373) );
  OAI21_X1 U14801 ( .B1(n12374), .B2(n12405), .A(n12373), .ZN(P3_U3448) );
  MUX2_X1 U14802 ( .A(n15385), .B(n12375), .S(n15055), .Z(n12376) );
  OAI21_X1 U14803 ( .B1(n12377), .B2(n12405), .A(n12376), .ZN(P3_U3447) );
  MUX2_X1 U14804 ( .A(n12379), .B(n12378), .S(n15055), .Z(n12380) );
  OAI21_X1 U14805 ( .B1(n12381), .B2(n12405), .A(n12380), .ZN(P3_U3446) );
  MUX2_X1 U14806 ( .A(n12383), .B(n12382), .S(n15055), .Z(n12384) );
  OAI21_X1 U14807 ( .B1(n12385), .B2(n12405), .A(n12384), .ZN(P3_U3444) );
  MUX2_X1 U14808 ( .A(n12387), .B(n12386), .S(n15055), .Z(n12388) );
  OAI21_X1 U14809 ( .B1(n12389), .B2(n12405), .A(n12388), .ZN(P3_U3441) );
  MUX2_X1 U14810 ( .A(n12391), .B(n12390), .S(n15055), .Z(n12392) );
  OAI21_X1 U14811 ( .B1(n12393), .B2(n12405), .A(n12392), .ZN(P3_U3438) );
  MUX2_X1 U14812 ( .A(n12395), .B(n12394), .S(n15055), .Z(n12396) );
  OAI21_X1 U14813 ( .B1(n12397), .B2(n12405), .A(n12396), .ZN(P3_U3435) );
  MUX2_X1 U14814 ( .A(n12399), .B(n12398), .S(n15056), .Z(n12400) );
  OAI21_X1 U14815 ( .B1(n12401), .B2(n12405), .A(n12400), .ZN(P3_U3432) );
  MUX2_X1 U14816 ( .A(n12403), .B(n12402), .S(n15055), .Z(n12404) );
  OAI21_X1 U14817 ( .B1(n12406), .B2(n12405), .A(n12404), .ZN(P3_U3429) );
  MUX2_X1 U14818 ( .A(P3_D_REG_0__SCAN_IN), .B(n6564), .S(n15075), .Z(P3_U3376) );
  INV_X1 U14819 ( .A(n12407), .ZN(n12410) );
  NAND3_X1 U14820 ( .A1(n8172), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n12409) );
  OAI22_X1 U14821 ( .A1(n12410), .A2(n12409), .B1(n12408), .B2(n12417), .ZN(
        n12411) );
  AOI21_X1 U14822 ( .B1(n12412), .B2(n14162), .A(n12411), .ZN(n12413) );
  INV_X1 U14823 ( .A(n12413), .ZN(P3_U3264) );
  INV_X1 U14824 ( .A(n12414), .ZN(n12415) );
  OAI222_X1 U14825 ( .A1(P3_U3151), .A2(n8179), .B1(n12417), .B2(n12416), .C1(
        n14154), .C2(n12415), .ZN(P3_U3265) );
  MUX2_X1 U14826 ( .A(n12419), .B(n12418), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3271) );
  INV_X1 U14827 ( .A(n12420), .ZN(n12421) );
  NOR2_X1 U14828 ( .A1(n12422), .A2(n12421), .ZN(n12423) );
  XNOR2_X1 U14829 ( .A(n12424), .B(n12423), .ZN(n12429) );
  NAND2_X1 U14830 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12844)
         );
  OAI21_X1 U14831 ( .B1(n12475), .B2(n13005), .A(n12844), .ZN(n12425) );
  AOI21_X1 U14832 ( .B1(n14308), .B2(n12787), .A(n12425), .ZN(n12426) );
  OAI21_X1 U14833 ( .B1(n13014), .B2(n14331), .A(n12426), .ZN(n12427) );
  AOI21_X1 U14834 ( .B1(n13114), .B2(n14328), .A(n12427), .ZN(n12428) );
  OAI21_X1 U14835 ( .B1(n12429), .B2(n14302), .A(n12428), .ZN(P2_U3191) );
  INV_X1 U14836 ( .A(n12430), .ZN(n12431) );
  NOR3_X1 U14837 ( .A1(n12431), .A2(n12695), .A3(n12502), .ZN(n12432) );
  AOI21_X1 U14838 ( .B1(n12440), .B2(n9282), .A(n12432), .ZN(n12444) );
  NOR2_X1 U14839 ( .A1(n12692), .A2(n12913), .ZN(n12434) );
  XNOR2_X1 U14840 ( .A(n12434), .B(n12433), .ZN(n12435) );
  XNOR2_X1 U14841 ( .A(n13065), .B(n12435), .ZN(n12443) );
  AOI22_X1 U14842 ( .A1(n12894), .A2(n13029), .B1(n13030), .B2(n12784), .ZN(
        n12863) );
  INV_X1 U14843 ( .A(n12870), .ZN(n12436) );
  AOI22_X1 U14844 ( .A1(n12436), .A2(n12489), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12437) );
  OAI21_X1 U14845 ( .B1(n12863), .B2(n12438), .A(n12437), .ZN(n12439) );
  AOI21_X1 U14846 ( .B1(n12872), .B2(n14328), .A(n12439), .ZN(n12442) );
  OAI21_X1 U14847 ( .B1(n12452), .B2(n12446), .A(n12445), .ZN(n12447) );
  NAND2_X1 U14848 ( .A1(n12447), .A2(n9282), .ZN(n12456) );
  AOI22_X1 U14849 ( .A1(n14308), .A2(n12794), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12448) );
  OAI21_X1 U14850 ( .B1(n12449), .B2(n14331), .A(n12448), .ZN(n12450) );
  AOI21_X1 U14851 ( .B1(n12561), .B2(n14328), .A(n12450), .ZN(n12455) );
  NOR3_X1 U14852 ( .A1(n12452), .A2(n12451), .A3(n12502), .ZN(n12453) );
  OAI21_X1 U14853 ( .B1(n12453), .B2(n14306), .A(n12797), .ZN(n12454) );
  NAND3_X1 U14854 ( .A1(n12456), .A2(n12455), .A3(n12454), .ZN(P2_U3193) );
  OAI211_X1 U14855 ( .C1(n12459), .C2(n12458), .A(n12457), .B(n9282), .ZN(
        n12463) );
  AOI22_X1 U14856 ( .A1(n14308), .A2(n12945), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12460) );
  OAI21_X1 U14857 ( .B1(n13007), .B2(n12475), .A(n12460), .ZN(n12461) );
  AOI21_X1 U14858 ( .B1(n12982), .B2(n12489), .A(n12461), .ZN(n12462) );
  OAI211_X1 U14859 ( .C1(n12984), .C2(n14310), .A(n12463), .B(n12462), .ZN(
        P2_U3195) );
  OAI21_X1 U14860 ( .B1(n12478), .B2(n12464), .A(n9282), .ZN(n12468) );
  NAND3_X1 U14861 ( .A1(n12466), .A2(n12465), .A3(n12944), .ZN(n12467) );
  NAND2_X1 U14862 ( .A1(n12468), .A2(n12467), .ZN(n12469) );
  NAND2_X1 U14863 ( .A1(n12498), .A2(n12469), .ZN(n12473) );
  AOI22_X1 U14864 ( .A1(n12785), .A2(n14308), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12470) );
  OAI21_X1 U14865 ( .B1(n12911), .B2(n12475), .A(n12470), .ZN(n12471) );
  AOI21_X1 U14866 ( .B1(n12918), .B2(n12489), .A(n12471), .ZN(n12472) );
  OAI211_X1 U14867 ( .C1(n12915), .C2(n14310), .A(n12473), .B(n12472), .ZN(
        P2_U3197) );
  OAI22_X1 U14868 ( .A1(n12475), .A2(n12927), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12474), .ZN(n12476) );
  AOI21_X1 U14869 ( .B1(n12932), .B2(n12489), .A(n12476), .ZN(n12477) );
  OAI21_X1 U14870 ( .B1(n12928), .B2(n12493), .A(n12477), .ZN(n12482) );
  AOI211_X1 U14871 ( .C1(n12480), .C2(n12479), .A(n14302), .B(n12478), .ZN(
        n12481) );
  AOI211_X1 U14872 ( .C1(n13089), .C2(n14328), .A(n12482), .B(n12481), .ZN(
        n12483) );
  INV_X1 U14873 ( .A(n12483), .ZN(P2_U3201) );
  INV_X1 U14874 ( .A(n12484), .ZN(n12486) );
  NAND2_X1 U14875 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  XNOR2_X1 U14876 ( .A(n12488), .B(n12487), .ZN(n12496) );
  AOI22_X1 U14877 ( .A1(n14306), .A2(n13031), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12491) );
  NAND2_X1 U14878 ( .A1(n12489), .A2(n12991), .ZN(n12490) );
  OAI211_X1 U14879 ( .C1(n12493), .C2(n12492), .A(n12491), .B(n12490), .ZN(
        n12494) );
  AOI21_X1 U14880 ( .B1(n13109), .B2(n14328), .A(n12494), .ZN(n12495) );
  OAI21_X1 U14881 ( .B1(n12496), .B2(n14302), .A(n12495), .ZN(P2_U3205) );
  OAI21_X1 U14882 ( .B1(n12504), .B2(n12498), .A(n12497), .ZN(n12499) );
  NAND2_X1 U14883 ( .A1(n12499), .A2(n9282), .ZN(n12508) );
  AOI22_X1 U14884 ( .A1(n12894), .A2(n14308), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12500) );
  OAI21_X1 U14885 ( .B1(n12897), .B2(n14331), .A(n12500), .ZN(n12501) );
  AOI21_X1 U14886 ( .B1(n13078), .B2(n14328), .A(n12501), .ZN(n12507) );
  NOR3_X1 U14887 ( .A1(n12504), .A2(n12503), .A3(n12502), .ZN(n12505) );
  OAI21_X1 U14888 ( .B1(n12505), .B2(n14306), .A(n12893), .ZN(n12506) );
  NAND3_X1 U14889 ( .A1(n12508), .A2(n12507), .A3(n12506), .ZN(P2_U3212) );
  INV_X1 U14890 ( .A(n12765), .ZN(n12509) );
  NOR2_X1 U14891 ( .A1(n12762), .A2(n12778), .ZN(n12516) );
  AOI21_X1 U14892 ( .B1(n12510), .B2(n12664), .A(n14763), .ZN(n12535) );
  INV_X1 U14893 ( .A(n12528), .ZN(n12691) );
  INV_X2 U14894 ( .A(n12691), .ZN(n12719) );
  AOI21_X1 U14895 ( .B1(n12801), .B2(n12719), .A(n12511), .ZN(n12534) );
  AOI21_X1 U14896 ( .B1(n12513), .B2(n12691), .A(n12512), .ZN(n12527) );
  AOI21_X1 U14897 ( .B1(n12803), .B2(n12528), .A(n6560), .ZN(n12526) );
  NAND2_X1 U14898 ( .A1(n12515), .A2(n12765), .ZN(n12524) );
  NAND2_X1 U14899 ( .A1(n12517), .A2(n12516), .ZN(n12519) );
  NAND2_X1 U14900 ( .A1(n12519), .A2(n12518), .ZN(n12523) );
  NAND2_X1 U14901 ( .A1(n12520), .A2(n12528), .ZN(n12522) );
  NAND4_X1 U14902 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12525) );
  MUX2_X1 U14903 ( .A(n12802), .B(n6589), .S(n12691), .Z(n12530) );
  MUX2_X1 U14904 ( .A(n12802), .B(n6589), .S(n12719), .Z(n12532) );
  MUX2_X1 U14905 ( .A(n12536), .B(n12800), .S(n12606), .Z(n12540) );
  MUX2_X1 U14906 ( .A(n12800), .B(n12536), .S(n12606), .Z(n12537) );
  NAND2_X1 U14907 ( .A1(n12538), .A2(n12537), .ZN(n12544) );
  INV_X1 U14908 ( .A(n12539), .ZN(n12542) );
  INV_X1 U14909 ( .A(n12540), .ZN(n12541) );
  NAND2_X1 U14910 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  MUX2_X1 U14911 ( .A(n12799), .B(n12545), .S(n12606), .Z(n12547) );
  MUX2_X1 U14912 ( .A(n12545), .B(n12799), .S(n12606), .Z(n12546) );
  INV_X1 U14913 ( .A(n12547), .ZN(n12548) );
  MUX2_X1 U14914 ( .A(n12798), .B(n12549), .S(n12664), .Z(n12553) );
  NAND2_X1 U14915 ( .A1(n12552), .A2(n12553), .ZN(n12551) );
  MUX2_X1 U14916 ( .A(n12798), .B(n12549), .S(n12606), .Z(n12550) );
  NAND2_X1 U14917 ( .A1(n12551), .A2(n12550), .ZN(n12557) );
  INV_X1 U14918 ( .A(n12552), .ZN(n12555) );
  INV_X1 U14919 ( .A(n12553), .ZN(n12554) );
  NAND2_X1 U14920 ( .A1(n12555), .A2(n12554), .ZN(n12556) );
  MUX2_X1 U14921 ( .A(n12797), .B(n12558), .S(n12606), .Z(n12560) );
  MUX2_X1 U14922 ( .A(n12797), .B(n12558), .S(n12664), .Z(n12559) );
  MUX2_X1 U14923 ( .A(n12796), .B(n12561), .S(n12694), .Z(n12565) );
  NAND2_X1 U14924 ( .A1(n12564), .A2(n12565), .ZN(n12563) );
  MUX2_X1 U14925 ( .A(n12796), .B(n12561), .S(n12606), .Z(n12562) );
  NAND2_X1 U14926 ( .A1(n12563), .A2(n12562), .ZN(n12569) );
  INV_X1 U14927 ( .A(n12564), .ZN(n12567) );
  INV_X1 U14928 ( .A(n12565), .ZN(n12566) );
  NAND2_X1 U14929 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  MUX2_X1 U14930 ( .A(n12794), .B(n14803), .S(n12606), .Z(n12571) );
  MUX2_X1 U14931 ( .A(n12794), .B(n14803), .S(n12694), .Z(n12570) );
  MUX2_X1 U14932 ( .A(n12793), .B(n14811), .S(n12694), .Z(n12576) );
  MUX2_X1 U14933 ( .A(n12793), .B(n14811), .S(n12606), .Z(n12573) );
  NAND2_X1 U14934 ( .A1(n12574), .A2(n12573), .ZN(n12580) );
  INV_X1 U14935 ( .A(n12575), .ZN(n12578) );
  INV_X1 U14936 ( .A(n12576), .ZN(n12577) );
  NAND2_X1 U14937 ( .A1(n12578), .A2(n12577), .ZN(n12579) );
  MUX2_X1 U14938 ( .A(n12792), .B(n14819), .S(n12606), .Z(n12584) );
  NAND2_X1 U14939 ( .A1(n12583), .A2(n12584), .ZN(n12582) );
  MUX2_X1 U14940 ( .A(n12792), .B(n14819), .S(n12694), .Z(n12581) );
  NAND2_X1 U14941 ( .A1(n12582), .A2(n12581), .ZN(n12588) );
  INV_X1 U14942 ( .A(n12583), .ZN(n12586) );
  INV_X1 U14943 ( .A(n12584), .ZN(n12585) );
  NAND2_X1 U14944 ( .A1(n12586), .A2(n12585), .ZN(n12587) );
  NAND2_X1 U14945 ( .A1(n12588), .A2(n12587), .ZN(n12591) );
  MUX2_X1 U14946 ( .A(n12791), .B(n12589), .S(n12694), .Z(n12592) );
  MUX2_X1 U14947 ( .A(n12791), .B(n12589), .S(n12606), .Z(n12590) );
  INV_X1 U14948 ( .A(n12592), .ZN(n12593) );
  MUX2_X1 U14949 ( .A(n14305), .B(n12594), .S(n12606), .Z(n12597) );
  INV_X1 U14950 ( .A(n12719), .ZN(n12694) );
  MUX2_X1 U14951 ( .A(n14305), .B(n12594), .S(n12694), .Z(n12595) );
  NAND2_X1 U14952 ( .A1(n12596), .A2(n12595), .ZN(n12598) );
  MUX2_X1 U14953 ( .A(n12790), .B(n12599), .S(n12694), .Z(n12602) );
  NAND2_X1 U14954 ( .A1(n12603), .A2(n12602), .ZN(n12601) );
  MUX2_X1 U14955 ( .A(n12790), .B(n12599), .S(n12606), .Z(n12600) );
  NAND2_X1 U14956 ( .A1(n12601), .A2(n12600), .ZN(n12605) );
  NAND2_X1 U14957 ( .A1(n12605), .A2(n12604), .ZN(n12609) );
  MUX2_X1 U14958 ( .A(n14307), .B(n13137), .S(n12606), .Z(n12610) );
  NAND2_X1 U14959 ( .A1(n12609), .A2(n12610), .ZN(n12608) );
  MUX2_X1 U14960 ( .A(n14307), .B(n13137), .S(n12694), .Z(n12607) );
  NAND2_X1 U14961 ( .A1(n12608), .A2(n12607), .ZN(n12614) );
  INV_X1 U14962 ( .A(n12609), .ZN(n12612) );
  INV_X1 U14963 ( .A(n12610), .ZN(n12611) );
  NAND2_X1 U14964 ( .A1(n12612), .A2(n12611), .ZN(n12613) );
  MUX2_X1 U14965 ( .A(n12789), .B(n14327), .S(n12694), .Z(n12616) );
  MUX2_X1 U14966 ( .A(n12789), .B(n14327), .S(n12606), .Z(n12615) );
  INV_X1 U14967 ( .A(n12616), .ZN(n12617) );
  MUX2_X1 U14968 ( .A(n13028), .B(n12618), .S(n12606), .Z(n12622) );
  NAND2_X1 U14969 ( .A1(n12621), .A2(n12622), .ZN(n12620) );
  MUX2_X1 U14970 ( .A(n13028), .B(n12618), .S(n12694), .Z(n12619) );
  NAND2_X1 U14971 ( .A1(n12620), .A2(n12619), .ZN(n12626) );
  INV_X1 U14972 ( .A(n12621), .ZN(n12624) );
  INV_X1 U14973 ( .A(n12622), .ZN(n12623) );
  NAND2_X1 U14974 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  MUX2_X1 U14975 ( .A(n12788), .B(n13045), .S(n12694), .Z(n12628) );
  MUX2_X1 U14976 ( .A(n12788), .B(n13045), .S(n12606), .Z(n12627) );
  MUX2_X1 U14977 ( .A(n13031), .B(n13114), .S(n12606), .Z(n12632) );
  MUX2_X1 U14978 ( .A(n13031), .B(n13114), .S(n12694), .Z(n12630) );
  NAND2_X1 U14979 ( .A1(n12631), .A2(n12630), .ZN(n12634) );
  NAND2_X1 U14980 ( .A1(n12634), .A2(n12633), .ZN(n12637) );
  MUX2_X1 U14981 ( .A(n13109), .B(n12787), .S(n12719), .Z(n12638) );
  NAND2_X1 U14982 ( .A1(n12637), .A2(n12638), .ZN(n12636) );
  MUX2_X1 U14983 ( .A(n12787), .B(n13109), .S(n12719), .Z(n12635) );
  INV_X1 U14984 ( .A(n12637), .ZN(n12640) );
  INV_X1 U14985 ( .A(n12638), .ZN(n12639) );
  MUX2_X1 U14986 ( .A(n12997), .B(n13105), .S(n12606), .Z(n12642) );
  MUX2_X1 U14987 ( .A(n12997), .B(n13105), .S(n12694), .Z(n12641) );
  INV_X1 U14988 ( .A(n12642), .ZN(n12643) );
  MUX2_X1 U14989 ( .A(n12945), .B(n13099), .S(n12694), .Z(n12646) );
  NAND2_X1 U14990 ( .A1(n12647), .A2(n12646), .ZN(n12645) );
  MUX2_X1 U14991 ( .A(n12945), .B(n13099), .S(n12528), .Z(n12644) );
  NAND2_X1 U14992 ( .A1(n12645), .A2(n12644), .ZN(n12649) );
  MUX2_X1 U14993 ( .A(n12786), .B(n13094), .S(n12528), .Z(n12653) );
  NAND2_X1 U14994 ( .A1(n12652), .A2(n12653), .ZN(n12651) );
  MUX2_X1 U14995 ( .A(n13094), .B(n12786), .S(n12528), .Z(n12650) );
  INV_X1 U14996 ( .A(n12652), .ZN(n12654) );
  MUX2_X1 U14997 ( .A(n13089), .B(n12944), .S(n12606), .Z(n12657) );
  MUX2_X1 U14998 ( .A(n12928), .B(n12915), .S(n12606), .Z(n12659) );
  MUX2_X1 U14999 ( .A(n12893), .B(n13084), .S(n12694), .Z(n12658) );
  MUX2_X1 U15000 ( .A(n12944), .B(n13089), .S(n12606), .Z(n12655) );
  INV_X1 U15001 ( .A(n12655), .ZN(n12656) );
  MUX2_X1 U15002 ( .A(n12912), .B(n12900), .S(n12719), .Z(n12697) );
  MUX2_X1 U15003 ( .A(n12785), .B(n13078), .S(n12694), .Z(n12696) );
  AOI22_X1 U15004 ( .A1(n12697), .A2(n12696), .B1(n12659), .B2(n12658), .ZN(
        n12660) );
  NAND2_X1 U15005 ( .A1(n12685), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12662) );
  INV_X1 U15006 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n12667) );
  NOR2_X1 U15007 ( .A1(n12668), .A2(n12667), .ZN(n12673) );
  INV_X1 U15008 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12847) );
  NOR2_X1 U15009 ( .A1(n9239), .A2(n12847), .ZN(n12672) );
  INV_X1 U15010 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n12669) );
  NOR2_X1 U15011 ( .A1(n12670), .A2(n12669), .ZN(n12671) );
  OR3_X1 U15012 ( .A1(n12673), .A2(n12672), .A3(n12671), .ZN(n12849) );
  NAND2_X1 U15013 ( .A1(n12849), .A2(n12694), .ZN(n12720) );
  OR2_X1 U15014 ( .A1(n12725), .A2(n12674), .ZN(n12770) );
  NAND4_X1 U15015 ( .A1(n12720), .A2(n12767), .A3(n12764), .A4(n12770), .ZN(
        n12675) );
  AND2_X1 U15016 ( .A1(n12675), .A2(n12783), .ZN(n12676) );
  AOI21_X1 U15017 ( .B1(n12853), .B2(n12719), .A(n12676), .ZN(n12708) );
  MUX2_X1 U15018 ( .A(n12784), .B(n13059), .S(n12719), .Z(n12677) );
  INV_X1 U15019 ( .A(n12677), .ZN(n12705) );
  MUX2_X1 U15020 ( .A(n13059), .B(n12784), .S(n12719), .Z(n12704) );
  OAI22_X1 U15021 ( .A1(n12707), .A2(n12708), .B1(n12705), .B2(n12704), .ZN(
        n12690) );
  MUX2_X1 U15022 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8042), .Z(n12681) );
  XNOR2_X1 U15023 ( .A(n12681), .B(SI_31_), .ZN(n12682) );
  NAND2_X1 U15024 ( .A1(n13473), .A2(n12684), .ZN(n12687) );
  NAND2_X1 U15025 ( .A1(n12685), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12686) );
  INV_X1 U15026 ( .A(n12851), .ZN(n13054) );
  INV_X1 U15027 ( .A(n12849), .ZN(n12688) );
  NAND2_X1 U15028 ( .A1(n12851), .A2(n12849), .ZN(n12689) );
  NAND2_X1 U15029 ( .A1(n12690), .A2(n6769), .ZN(n12710) );
  MUX2_X1 U15030 ( .A(n12692), .B(n13065), .S(n12691), .Z(n12701) );
  MUX2_X1 U15031 ( .A(n11425), .B(n12872), .S(n12719), .Z(n12700) );
  NAND2_X1 U15032 ( .A1(n12701), .A2(n12700), .ZN(n12693) );
  MUX2_X1 U15033 ( .A(n12695), .B(n13072), .S(n12694), .Z(n12712) );
  MUX2_X1 U15034 ( .A(n12894), .B(n12888), .S(n12719), .Z(n12711) );
  NOR2_X1 U15035 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  AOI21_X1 U15036 ( .B1(n12712), .B2(n12711), .A(n12698), .ZN(n12699) );
  INV_X1 U15037 ( .A(n12700), .ZN(n12703) );
  INV_X1 U15038 ( .A(n12701), .ZN(n12702) );
  AOI22_X1 U15039 ( .A1(n12705), .A2(n12704), .B1(n12703), .B2(n12702), .ZN(
        n12706) );
  AOI22_X1 U15040 ( .A1(n12710), .A2(n12709), .B1(n12708), .B2(n12707), .ZN(
        n12717) );
  INV_X1 U15041 ( .A(n12711), .ZN(n12714) );
  INV_X1 U15042 ( .A(n12712), .ZN(n12713) );
  NAND2_X1 U15043 ( .A1(n6764), .A2(n12719), .ZN(n12721) );
  NAND3_X1 U15044 ( .A1(n12722), .A2(n12721), .A3(n12720), .ZN(n12723) );
  INV_X1 U15045 ( .A(n12783), .ZN(n12726) );
  INV_X1 U15046 ( .A(n6559), .ZN(n12768) );
  NAND4_X1 U15047 ( .A1(n12729), .A2(n12728), .A3(n12768), .A4(n12727), .ZN(
        n12732) );
  NOR3_X1 U15048 ( .A1(n12732), .A2(n12731), .A3(n12730), .ZN(n12736) );
  NAND4_X1 U15049 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12739) );
  OR4_X1 U15050 ( .A1(n12740), .A2(n12739), .A3(n12738), .A4(n12737), .ZN(
        n12741) );
  NOR2_X1 U15051 ( .A1(n12742), .A2(n12741), .ZN(n12745) );
  NAND4_X1 U15052 ( .A1(n12746), .A2(n12745), .A3(n12744), .A4(n12743), .ZN(
        n12749) );
  OR4_X1 U15053 ( .A1(n12750), .A2(n12749), .A3(n12748), .A4(n12747), .ZN(
        n12751) );
  NOR2_X1 U15054 ( .A1(n12752), .A2(n12751), .ZN(n12753) );
  XNOR2_X1 U15055 ( .A(n13114), .B(n13031), .ZN(n13008) );
  NAND3_X1 U15056 ( .A1(n12996), .A2(n12753), .A3(n13008), .ZN(n12754) );
  NOR2_X1 U15057 ( .A1(n12974), .A2(n12754), .ZN(n12757) );
  NAND2_X1 U15058 ( .A1(n12756), .A2(n12755), .ZN(n12953) );
  NAND4_X1 U15059 ( .A1(n12937), .A2(n12961), .A3(n12757), .A4(n12953), .ZN(
        n12758) );
  NOR2_X1 U15060 ( .A1(n12908), .A2(n12758), .ZN(n12759) );
  XNOR2_X1 U15061 ( .A(n13078), .B(n12785), .ZN(n12901) );
  NAND2_X1 U15062 ( .A1(n12762), .A2(n12767), .ZN(n12763) );
  OAI211_X1 U15063 ( .C1(n12765), .C2(n12778), .A(n12764), .B(n12763), .ZN(
        n12766) );
  INV_X1 U15064 ( .A(n12766), .ZN(n12773) );
  NAND3_X1 U15065 ( .A1(n12768), .A2(n12842), .A3(n12767), .ZN(n12769) );
  NAND2_X1 U15066 ( .A1(n12770), .A2(n12769), .ZN(n12771) );
  OAI21_X1 U15067 ( .B1(n12774), .B2(n12773), .A(n12772), .ZN(n12775) );
  NOR2_X1 U15068 ( .A1(n12776), .A2(n12775), .ZN(n12782) );
  NOR3_X1 U15069 ( .A1(n12777), .A2(n6777), .A3(n13004), .ZN(n12780) );
  OAI21_X1 U15070 ( .B1(n12781), .B2(n12778), .A(P2_B_REG_SCAN_IN), .ZN(n12779) );
  OAI22_X1 U15071 ( .A1(n12782), .A2(n12781), .B1(n12780), .B2(n12779), .ZN(
        P2_U3328) );
  MUX2_X1 U15072 ( .A(n12849), .B(P2_DATAO_REG_31__SCAN_IN), .S(n12795), .Z(
        P2_U3562) );
  MUX2_X1 U15073 ( .A(n12783), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12795), .Z(
        P2_U3561) );
  MUX2_X1 U15074 ( .A(n12784), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12795), .Z(
        P2_U3560) );
  MUX2_X1 U15075 ( .A(n11425), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12795), .Z(
        P2_U3559) );
  MUX2_X1 U15076 ( .A(n12894), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12795), .Z(
        P2_U3558) );
  MUX2_X1 U15077 ( .A(n12785), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12795), .Z(
        P2_U3557) );
  MUX2_X1 U15078 ( .A(n12893), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12795), .Z(
        P2_U3556) );
  MUX2_X1 U15079 ( .A(n12944), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12795), .Z(
        P2_U3555) );
  MUX2_X1 U15080 ( .A(n12786), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12795), .Z(
        P2_U3554) );
  MUX2_X1 U15081 ( .A(n12945), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12795), .Z(
        P2_U3553) );
  MUX2_X1 U15082 ( .A(n12997), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12795), .Z(
        P2_U3552) );
  MUX2_X1 U15083 ( .A(n12787), .B(P2_DATAO_REG_20__SCAN_IN), .S(n12795), .Z(
        P2_U3551) );
  MUX2_X1 U15084 ( .A(n13031), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12804), .Z(
        P2_U3550) );
  MUX2_X1 U15085 ( .A(n12788), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12795), .Z(
        P2_U3549) );
  MUX2_X1 U15086 ( .A(n13028), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12795), .Z(
        P2_U3548) );
  MUX2_X1 U15087 ( .A(n12789), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12804), .Z(
        P2_U3547) );
  MUX2_X1 U15088 ( .A(n14307), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12795), .Z(
        P2_U3546) );
  MUX2_X1 U15089 ( .A(n12790), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12795), .Z(
        P2_U3545) );
  MUX2_X1 U15090 ( .A(n14305), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12804), .Z(
        P2_U3544) );
  MUX2_X1 U15091 ( .A(n12791), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12795), .Z(
        P2_U3543) );
  MUX2_X1 U15092 ( .A(n12792), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12804), .Z(
        P2_U3542) );
  MUX2_X1 U15093 ( .A(n12793), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12804), .Z(
        P2_U3541) );
  MUX2_X1 U15094 ( .A(n12794), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12795), .Z(
        P2_U3540) );
  MUX2_X1 U15095 ( .A(n12796), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12795), .Z(
        P2_U3539) );
  MUX2_X1 U15096 ( .A(n12797), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12804), .Z(
        P2_U3538) );
  MUX2_X1 U15097 ( .A(n12798), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12804), .Z(
        P2_U3537) );
  MUX2_X1 U15098 ( .A(n12799), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12804), .Z(
        P2_U3536) );
  MUX2_X1 U15099 ( .A(n12800), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12804), .Z(
        P2_U3535) );
  MUX2_X1 U15100 ( .A(n12801), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12804), .Z(
        P2_U3534) );
  MUX2_X1 U15101 ( .A(n12802), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12804), .Z(
        P2_U3533) );
  MUX2_X1 U15102 ( .A(n12803), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12804), .Z(
        P2_U3532) );
  MUX2_X1 U15103 ( .A(n12805), .B(P2_DATAO_REG_0__SCAN_IN), .S(n12804), .Z(
        P2_U3531) );
  OAI21_X1 U15104 ( .B1(n12808), .B2(n12807), .A(n12806), .ZN(n12809) );
  NAND2_X1 U15105 ( .A1(n12809), .A2(n14715), .ZN(n12818) );
  INV_X1 U15106 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U15107 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n12810)
         );
  OAI21_X1 U15108 ( .B1(n14722), .B2(n14396), .A(n12810), .ZN(n12811) );
  AOI21_X1 U15109 ( .B1(n12812), .B2(n14719), .A(n12811), .ZN(n12817) );
  OAI211_X1 U15110 ( .C1(n12815), .C2(n12814), .A(n12813), .B(n14655), .ZN(
        n12816) );
  NAND3_X1 U15111 ( .A1(n12818), .A2(n12817), .A3(n12816), .ZN(P2_U3225) );
  AOI21_X1 U15112 ( .B1(n12820), .B2(P2_REG1_REG_14__SCAN_IN), .A(n12819), 
        .ZN(n12821) );
  NOR2_X1 U15113 ( .A1(n12821), .A2(n12830), .ZN(n12822) );
  XNOR2_X1 U15114 ( .A(n12830), .B(n12821), .ZN(n14673) );
  NOR2_X1 U15115 ( .A1(n14672), .A2(n14673), .ZN(n14671) );
  NOR2_X1 U15116 ( .A1(n12822), .A2(n14671), .ZN(n14682) );
  XNOR2_X1 U15117 ( .A(n14689), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14681) );
  NOR2_X1 U15118 ( .A1(n14682), .A2(n14681), .ZN(n14680) );
  AOI21_X1 U15119 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n14689), .A(n14680), 
        .ZN(n14700) );
  XNOR2_X1 U15120 ( .A(n14703), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14699) );
  NOR2_X1 U15121 ( .A1(n14700), .A2(n14699), .ZN(n14698) );
  AOI21_X1 U15122 ( .B1(n14703), .B2(P2_REG1_REG_17__SCAN_IN), .A(n14698), 
        .ZN(n12823) );
  NOR2_X1 U15123 ( .A1(n12823), .A2(n12835), .ZN(n12824) );
  XNOR2_X1 U15124 ( .A(n12835), .B(n12823), .ZN(n14710) );
  NOR2_X1 U15125 ( .A1(n14709), .A2(n14710), .ZN(n14708) );
  NOR2_X1 U15126 ( .A1(n12824), .A2(n14708), .ZN(n12826) );
  INV_X1 U15127 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n12825) );
  XOR2_X1 U15128 ( .A(n12826), .B(n12825), .Z(n12839) );
  NOR2_X1 U15129 ( .A1(n12828), .A2(n12827), .ZN(n12829) );
  NOR2_X1 U15130 ( .A1(n12829), .A2(n12830), .ZN(n12831) );
  XNOR2_X1 U15131 ( .A(n12830), .B(n12829), .ZN(n14670) );
  NOR2_X1 U15132 ( .A1(n9102), .A2(n14670), .ZN(n14669) );
  NOR2_X1 U15133 ( .A1(n12831), .A2(n14669), .ZN(n14686) );
  XNOR2_X1 U15134 ( .A(n14689), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n14685) );
  NAND2_X1 U15135 ( .A1(n14689), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U15136 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n14703), .ZN(n12833) );
  OAI21_X1 U15137 ( .B1(n14703), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12833), 
        .ZN(n14696) );
  INV_X1 U15138 ( .A(n14696), .ZN(n12834) );
  NAND2_X1 U15139 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  INV_X1 U15140 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14712) );
  NAND2_X1 U15141 ( .A1(n14713), .A2(n14712), .ZN(n14711) );
  NAND2_X1 U15142 ( .A1(n12837), .A2(n14711), .ZN(n12838) );
  XNOR2_X1 U15143 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12838), .ZN(n12840) );
  AOI22_X1 U15144 ( .A1(n12839), .A2(n14655), .B1(n12840), .B2(n14715), .ZN(
        n12843) );
  INV_X1 U15145 ( .A(n12839), .ZN(n12841) );
  XNOR2_X1 U15146 ( .A(n12855), .B(n6764), .ZN(n12846) );
  NAND2_X1 U15147 ( .A1(n12846), .A2(n12913), .ZN(n13053) );
  NOR2_X1 U15148 ( .A1(n12979), .A2(n12847), .ZN(n12850) );
  NAND2_X1 U15149 ( .A1(n12849), .A2(n12848), .ZN(n13055) );
  NOR2_X1 U15150 ( .A1(n13051), .A2(n13055), .ZN(n12858) );
  AOI211_X1 U15151 ( .C1(n6764), .C2(n13044), .A(n12850), .B(n12858), .ZN(
        n12852) );
  OAI21_X1 U15152 ( .B1(n13053), .B2(n13047), .A(n12852), .ZN(P2_U3234) );
  OAI211_X1 U15153 ( .C1(n13057), .C2(n6892), .A(n12856), .B(n12913), .ZN(
        n13056) );
  NOR2_X1 U15154 ( .A1(n13057), .A2(n13018), .ZN(n12857) );
  AOI211_X1 U15155 ( .C1(n13051), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12858), 
        .B(n12857), .ZN(n12859) );
  OAI21_X1 U15156 ( .B1(n13047), .B2(n13056), .A(n12859), .ZN(P2_U3235) );
  OAI211_X1 U15157 ( .C1(n12862), .C2(n12861), .A(n12860), .B(n13026), .ZN(
        n12864) );
  OAI21_X1 U15158 ( .B1(n12867), .B2(n12866), .A(n12865), .ZN(n13069) );
  INV_X1 U15159 ( .A(n13069), .ZN(n12875) );
  OAI211_X1 U15160 ( .C1(n13065), .C2(n12882), .A(n12913), .B(n12868), .ZN(
        n13064) );
  INV_X1 U15161 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n12869) );
  OAI22_X1 U15162 ( .A1(n12870), .A2(n13041), .B1(n12869), .B2(n12979), .ZN(
        n12871) );
  AOI21_X1 U15163 ( .B1(n12872), .B2(n13044), .A(n12871), .ZN(n12873) );
  OAI21_X1 U15164 ( .B1(n13064), .B2(n13047), .A(n12873), .ZN(n12874) );
  AOI21_X1 U15165 ( .B1(n12875), .B2(n13049), .A(n12874), .ZN(n12876) );
  OAI21_X1 U15166 ( .B1(n13068), .B2(n13051), .A(n12876), .ZN(P2_U3237) );
  XNOR2_X1 U15167 ( .A(n12878), .B(n12877), .ZN(n12880) );
  AOI21_X1 U15168 ( .B1(n12880), .B2(n13026), .A(n12879), .ZN(n13076) );
  OAI21_X1 U15169 ( .B1(n13072), .B2(n12895), .A(n12913), .ZN(n12881) );
  OR2_X1 U15170 ( .A1(n6696), .A2(n12883), .ZN(n13071) );
  NAND3_X1 U15171 ( .A1(n13071), .A2(n13070), .A3(n13049), .ZN(n12890) );
  NAND2_X1 U15172 ( .A1(n12884), .A2(n13015), .ZN(n12885) );
  OAI21_X1 U15173 ( .B1(n12979), .B2(n12886), .A(n12885), .ZN(n12887) );
  AOI21_X1 U15174 ( .B1(n12888), .B2(n13044), .A(n12887), .ZN(n12889) );
  OAI211_X1 U15175 ( .C1(n13075), .C2(n13047), .A(n12890), .B(n12889), .ZN(
        n12891) );
  INV_X1 U15176 ( .A(n12891), .ZN(n12892) );
  OAI21_X1 U15177 ( .B1(n13076), .B2(n13051), .A(n12892), .ZN(P2_U3238) );
  INV_X1 U15178 ( .A(n12917), .ZN(n12896) );
  AOI211_X1 U15179 ( .C1(n13078), .C2(n12896), .A(n9183), .B(n12895), .ZN(
        n13077) );
  INV_X1 U15180 ( .A(n12897), .ZN(n12898) );
  AOI22_X1 U15181 ( .A1(n12898), .A2(n13015), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13051), .ZN(n12899) );
  OAI21_X1 U15182 ( .B1(n12900), .B2(n13018), .A(n12899), .ZN(n12904) );
  XOR2_X1 U15183 ( .A(n12902), .B(n12901), .Z(n13081) );
  NOR2_X1 U15184 ( .A1(n13081), .A2(n13002), .ZN(n12903) );
  AOI211_X1 U15185 ( .C1(n13077), .C2(n13023), .A(n12904), .B(n12903), .ZN(
        n12905) );
  OAI21_X1 U15186 ( .B1(n13080), .B2(n13051), .A(n12905), .ZN(P2_U3239) );
  XOR2_X1 U15187 ( .A(n12906), .B(n12908), .Z(n13086) );
  AOI21_X1 U15188 ( .B1(n12909), .B2(n12908), .A(n12907), .ZN(n12910) );
  OAI222_X1 U15189 ( .A1(n13006), .A2(n12912), .B1(n13004), .B2(n12911), .C1(
        n12977), .C2(n12910), .ZN(n13083) );
  OAI21_X1 U15190 ( .B1(n12915), .B2(n12914), .A(n12913), .ZN(n12916) );
  OR2_X1 U15191 ( .A1(n12917), .A2(n12916), .ZN(n13082) );
  AOI22_X1 U15192 ( .A1(n12918), .A2(n13015), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13051), .ZN(n12920) );
  NAND2_X1 U15193 ( .A1(n13084), .A2(n13044), .ZN(n12919) );
  OAI211_X1 U15194 ( .C1(n13082), .C2(n13047), .A(n12920), .B(n12919), .ZN(
        n12921) );
  AOI21_X1 U15195 ( .B1(n13083), .B2(n12979), .A(n12921), .ZN(n12922) );
  OAI21_X1 U15196 ( .B1(n13086), .B2(n13002), .A(n12922), .ZN(P2_U3240) );
  AOI21_X1 U15197 ( .B1(n12925), .B2(n12924), .A(n12923), .ZN(n12926) );
  OAI222_X1 U15198 ( .A1(n13006), .A2(n12928), .B1(n13004), .B2(n12927), .C1(
        n12977), .C2(n12926), .ZN(n12929) );
  INV_X1 U15199 ( .A(n12929), .ZN(n13091) );
  INV_X1 U15200 ( .A(n13089), .ZN(n12930) );
  XNOR2_X1 U15201 ( .A(n12930), .B(n12946), .ZN(n12931) );
  AND2_X1 U15202 ( .A1(n12931), .A2(n12913), .ZN(n13088) );
  NAND2_X1 U15203 ( .A1(n13089), .A2(n13044), .ZN(n12934) );
  AOI22_X1 U15204 ( .A1(n12932), .A2(n13015), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13051), .ZN(n12933) );
  NAND2_X1 U15205 ( .A1(n12934), .A2(n12933), .ZN(n12935) );
  AOI21_X1 U15206 ( .B1(n13088), .B2(n13023), .A(n12935), .ZN(n12941) );
  INV_X1 U15207 ( .A(n12936), .ZN(n12939) );
  NAND2_X1 U15208 ( .A1(n12938), .A2(n12937), .ZN(n13087) );
  NAND3_X1 U15209 ( .A1(n12939), .A2(n13049), .A3(n13087), .ZN(n12940) );
  OAI211_X1 U15210 ( .C1(n13091), .C2(n13051), .A(n12941), .B(n12940), .ZN(
        P2_U3241) );
  XOR2_X1 U15211 ( .A(n12942), .B(n12953), .Z(n12943) );
  AOI222_X1 U15212 ( .A1(n12945), .A2(n13029), .B1(n12944), .B2(n13030), .C1(
        n13026), .C2(n12943), .ZN(n13096) );
  INV_X1 U15213 ( .A(n12946), .ZN(n12947) );
  AOI211_X1 U15214 ( .C1(n13094), .C2(n12965), .A(n9183), .B(n12947), .ZN(
        n13093) );
  INV_X1 U15215 ( .A(n12948), .ZN(n12949) );
  AOI22_X1 U15216 ( .A1(n12949), .A2(n13015), .B1(n13051), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n12950) );
  OAI21_X1 U15217 ( .B1(n12951), .B2(n13018), .A(n12950), .ZN(n12955) );
  XOR2_X1 U15218 ( .A(n12953), .B(n12952), .Z(n13097) );
  NOR2_X1 U15219 ( .A1(n13097), .A2(n13002), .ZN(n12954) );
  AOI211_X1 U15220 ( .C1(n13093), .C2(n13023), .A(n12955), .B(n12954), .ZN(
        n12956) );
  OAI21_X1 U15221 ( .B1(n13096), .B2(n13051), .A(n12956), .ZN(P2_U3242) );
  OAI211_X1 U15222 ( .C1(n12958), .C2(n12961), .A(n12957), .B(n13026), .ZN(
        n12960) );
  NAND2_X1 U15223 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  NAND2_X1 U15224 ( .A1(n12964), .A2(n12963), .ZN(n13102) );
  INV_X1 U15225 ( .A(n13102), .ZN(n12971) );
  AOI21_X1 U15226 ( .B1(n13099), .B2(n12980), .A(n9183), .ZN(n12966) );
  AND2_X1 U15227 ( .A1(n12966), .A2(n12965), .ZN(n13098) );
  NAND2_X1 U15228 ( .A1(n13098), .A2(n13023), .ZN(n12969) );
  AOI22_X1 U15229 ( .A1(n13051), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n12967), 
        .B2(n13015), .ZN(n12968) );
  OAI211_X1 U15230 ( .C1(n6885), .C2(n13018), .A(n12969), .B(n12968), .ZN(
        n12970) );
  AOI21_X1 U15231 ( .B1(n12971), .B2(n13049), .A(n12970), .ZN(n12972) );
  OAI21_X1 U15232 ( .B1(n13101), .B2(n13051), .A(n12972), .ZN(P2_U3243) );
  XNOR2_X1 U15233 ( .A(n12973), .B(n12974), .ZN(n13107) );
  XNOR2_X1 U15234 ( .A(n6776), .B(n12974), .ZN(n12976) );
  OAI222_X1 U15235 ( .A1(n13006), .A2(n12978), .B1(n13004), .B2(n13007), .C1(
        n12977), .C2(n12976), .ZN(n13103) );
  NAND2_X1 U15236 ( .A1(n13103), .A2(n12979), .ZN(n12987) );
  INV_X1 U15237 ( .A(n12980), .ZN(n12981) );
  AOI211_X1 U15238 ( .C1(n13105), .C2(n12990), .A(n9183), .B(n12981), .ZN(
        n13104) );
  AOI22_X1 U15239 ( .A1(n13051), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n12982), 
        .B2(n13015), .ZN(n12983) );
  OAI21_X1 U15240 ( .B1(n12984), .B2(n13018), .A(n12983), .ZN(n12985) );
  AOI21_X1 U15241 ( .B1(n13104), .B2(n13023), .A(n12985), .ZN(n12986) );
  OAI211_X1 U15242 ( .C1(n13107), .C2(n13002), .A(n12987), .B(n12986), .ZN(
        P2_U3244) );
  XNOR2_X1 U15243 ( .A(n12988), .B(n12996), .ZN(n13112) );
  OR2_X1 U15244 ( .A1(n13013), .A2(n12993), .ZN(n12989) );
  AND3_X1 U15245 ( .A1(n12990), .A2(n12913), .A3(n12989), .ZN(n13108) );
  AOI22_X1 U15246 ( .A1(n13051), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n12991), 
        .B2(n13015), .ZN(n12992) );
  OAI21_X1 U15247 ( .B1(n12993), .B2(n13018), .A(n12992), .ZN(n13000) );
  OAI21_X1 U15248 ( .B1(n12996), .B2(n12995), .A(n12994), .ZN(n12998) );
  AOI222_X1 U15249 ( .A1(n13026), .A2(n12998), .B1(n12997), .B2(n13030), .C1(
        n13031), .C2(n13029), .ZN(n13111) );
  NOR2_X1 U15250 ( .A1(n13111), .A2(n13051), .ZN(n12999) );
  AOI211_X1 U15251 ( .C1(n13108), .C2(n13023), .A(n13000), .B(n12999), .ZN(
        n13001) );
  OAI21_X1 U15252 ( .B1(n13112), .B2(n13002), .A(n13001), .ZN(P2_U3245) );
  XNOR2_X1 U15253 ( .A(n13003), .B(n13008), .ZN(n13012) );
  OAI22_X1 U15254 ( .A1(n13007), .A2(n13006), .B1(n13005), .B2(n13004), .ZN(
        n13011) );
  XNOR2_X1 U15255 ( .A(n13009), .B(n13008), .ZN(n13117) );
  NOR2_X1 U15256 ( .A1(n13117), .A2(n9731), .ZN(n13010) );
  AOI211_X1 U15257 ( .C1(n13012), .C2(n13026), .A(n13011), .B(n13010), .ZN(
        n13116) );
  AOI211_X1 U15258 ( .C1(n13114), .C2(n13039), .A(n9183), .B(n13013), .ZN(
        n13113) );
  INV_X1 U15259 ( .A(n13014), .ZN(n13016) );
  AOI22_X1 U15260 ( .A1(n13051), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13016), 
        .B2(n13015), .ZN(n13017) );
  OAI21_X1 U15261 ( .B1(n13019), .B2(n13018), .A(n13017), .ZN(n13022) );
  NOR2_X1 U15262 ( .A1(n13117), .A2(n13020), .ZN(n13021) );
  AOI211_X1 U15263 ( .C1(n13113), .C2(n13023), .A(n13022), .B(n13021), .ZN(
        n13024) );
  OAI21_X1 U15264 ( .B1(n13116), .B2(n13051), .A(n13024), .ZN(P2_U3246) );
  XNOR2_X1 U15265 ( .A(n13025), .B(n13034), .ZN(n13027) );
  NAND2_X1 U15266 ( .A1(n13027), .A2(n13026), .ZN(n13033) );
  AOI22_X1 U15267 ( .A1(n13031), .A2(n13030), .B1(n13029), .B2(n13028), .ZN(
        n13032) );
  NAND2_X1 U15268 ( .A1(n13033), .A2(n13032), .ZN(n13123) );
  INV_X1 U15269 ( .A(n13123), .ZN(n13052) );
  NAND2_X1 U15270 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NAND2_X1 U15271 ( .A1(n13037), .A2(n13036), .ZN(n13118) );
  AOI21_X1 U15272 ( .B1(n13045), .B2(n13038), .A(n9183), .ZN(n13040) );
  NAND2_X1 U15273 ( .A1(n13040), .A2(n13039), .ZN(n13119) );
  OAI22_X1 U15274 ( .A1(n12979), .A2(n14712), .B1(n13042), .B2(n13041), .ZN(
        n13043) );
  AOI21_X1 U15275 ( .B1(n13045), .B2(n13044), .A(n13043), .ZN(n13046) );
  OAI21_X1 U15276 ( .B1(n13119), .B2(n13047), .A(n13046), .ZN(n13048) );
  AOI21_X1 U15277 ( .B1(n13118), .B2(n13049), .A(n13048), .ZN(n13050) );
  OAI21_X1 U15278 ( .B1(n13052), .B2(n13051), .A(n13050), .ZN(P2_U3247) );
  OAI211_X1 U15279 ( .C1(n13054), .C2(n14797), .A(n13053), .B(n13055), .ZN(
        n13142) );
  MUX2_X1 U15280 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13142), .S(n14842), .Z(
        P2_U3530) );
  OAI211_X1 U15281 ( .C1(n13057), .C2(n14797), .A(n13056), .B(n13055), .ZN(
        n13143) );
  MUX2_X1 U15282 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13143), .S(n14842), .Z(
        P2_U3529) );
  INV_X1 U15283 ( .A(n13059), .ZN(n13061) );
  OAI21_X1 U15284 ( .B1(n13061), .B2(n14797), .A(n13060), .ZN(n13062) );
  MUX2_X1 U15285 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13144), .S(n14842), .Z(
        P2_U3528) );
  OAI21_X1 U15286 ( .B1(n13065), .B2(n14797), .A(n13064), .ZN(n13066) );
  INV_X1 U15287 ( .A(n13066), .ZN(n13067) );
  OAI211_X1 U15288 ( .C1(n13140), .C2(n13069), .A(n13068), .B(n13067), .ZN(
        n13145) );
  MUX2_X1 U15289 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13145), .S(n14842), .Z(
        P2_U3527) );
  NAND3_X1 U15290 ( .A1(n13071), .A2(n13070), .A3(n14787), .ZN(n13074) );
  OR2_X1 U15291 ( .A1(n13072), .A2(n14797), .ZN(n13073) );
  NAND4_X1 U15292 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13146) );
  MUX2_X1 U15293 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13146), .S(n14842), .Z(
        P2_U3526) );
  AOI21_X1 U15294 ( .B1(n14818), .B2(n13078), .A(n13077), .ZN(n13079) );
  OAI211_X1 U15295 ( .C1(n13140), .C2(n13081), .A(n13080), .B(n13079), .ZN(
        n13147) );
  MUX2_X1 U15296 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13147), .S(n14842), .Z(
        P2_U3525) );
  OAI21_X1 U15297 ( .B1(n13140), .B2(n13086), .A(n13085), .ZN(n13148) );
  MUX2_X1 U15298 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13148), .S(n14842), .Z(
        P2_U3524) );
  NAND2_X1 U15299 ( .A1(n13087), .A2(n14787), .ZN(n13092) );
  AOI21_X1 U15300 ( .B1(n14818), .B2(n13089), .A(n13088), .ZN(n13090) );
  OAI211_X1 U15301 ( .C1(n12936), .C2(n13092), .A(n13091), .B(n13090), .ZN(
        n13149) );
  MUX2_X1 U15302 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13149), .S(n14842), .Z(
        P2_U3523) );
  AOI21_X1 U15303 ( .B1(n14818), .B2(n13094), .A(n13093), .ZN(n13095) );
  OAI211_X1 U15304 ( .C1(n13140), .C2(n13097), .A(n13096), .B(n13095), .ZN(
        n13150) );
  MUX2_X1 U15305 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13150), .S(n14842), .Z(
        P2_U3522) );
  AOI21_X1 U15306 ( .B1(n14818), .B2(n13099), .A(n13098), .ZN(n13100) );
  OAI211_X1 U15307 ( .C1(n13140), .C2(n13102), .A(n13101), .B(n13100), .ZN(
        n13151) );
  MUX2_X1 U15308 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13151), .S(n14842), .Z(
        P2_U3521) );
  AOI211_X1 U15309 ( .C1(n14818), .C2(n13105), .A(n13104), .B(n13103), .ZN(
        n13106) );
  OAI21_X1 U15310 ( .B1(n13140), .B2(n13107), .A(n13106), .ZN(n13152) );
  MUX2_X1 U15311 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13152), .S(n14842), .Z(
        P2_U3520) );
  AOI21_X1 U15312 ( .B1(n14818), .B2(n13109), .A(n13108), .ZN(n13110) );
  OAI211_X1 U15313 ( .C1(n13140), .C2(n13112), .A(n13111), .B(n13110), .ZN(
        n13153) );
  MUX2_X1 U15314 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13153), .S(n14842), .Z(
        P2_U3519) );
  AOI21_X1 U15315 ( .B1(n14818), .B2(n13114), .A(n13113), .ZN(n13115) );
  OAI211_X1 U15316 ( .C1(n14822), .C2(n13117), .A(n13116), .B(n13115), .ZN(
        n13154) );
  MUX2_X1 U15317 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13154), .S(n14842), .Z(
        P2_U3518) );
  AND2_X1 U15318 ( .A1(n13118), .A2(n14787), .ZN(n13122) );
  OAI21_X1 U15319 ( .B1(n13120), .B2(n14797), .A(n13119), .ZN(n13121) );
  MUX2_X1 U15320 ( .A(n13155), .B(P2_REG1_REG_18__SCAN_IN), .S(n14840), .Z(
        P2_U3517) );
  AND2_X1 U15321 ( .A1(n13124), .A2(n14787), .ZN(n13128) );
  OAI21_X1 U15322 ( .B1(n13126), .B2(n14797), .A(n13125), .ZN(n13127) );
  MUX2_X1 U15323 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13156), .S(n14842), .Z(
        P2_U3516) );
  INV_X1 U15324 ( .A(n14327), .ZN(n13131) );
  OAI21_X1 U15325 ( .B1(n13131), .B2(n14797), .A(n13130), .ZN(n13132) );
  AOI21_X1 U15326 ( .B1(n13133), .B2(n14787), .A(n13132), .ZN(n13134) );
  NAND2_X1 U15327 ( .A1(n13135), .A2(n13134), .ZN(n13157) );
  MUX2_X1 U15328 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13157), .S(n14842), .Z(
        P2_U3515) );
  AOI21_X1 U15329 ( .B1(n14818), .B2(n13137), .A(n13136), .ZN(n13138) );
  OAI211_X1 U15330 ( .C1(n13141), .C2(n13140), .A(n13139), .B(n13138), .ZN(
        n13158) );
  MUX2_X1 U15331 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13158), .S(n14842), .Z(
        P2_U3514) );
  MUX2_X1 U15332 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13142), .S(n14829), .Z(
        P2_U3498) );
  MUX2_X1 U15333 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13143), .S(n14829), .Z(
        P2_U3497) );
  MUX2_X1 U15334 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13145), .S(n14829), .Z(
        P2_U3495) );
  MUX2_X1 U15335 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13146), .S(n14829), .Z(
        P2_U3494) );
  MUX2_X1 U15336 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13147), .S(n14829), .Z(
        P2_U3493) );
  MUX2_X1 U15337 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13148), .S(n14829), .Z(
        P2_U3492) );
  MUX2_X1 U15338 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13149), .S(n14829), .Z(
        P2_U3491) );
  MUX2_X1 U15339 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13150), .S(n14829), .Z(
        P2_U3490) );
  MUX2_X1 U15340 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13151), .S(n14829), .Z(
        P2_U3489) );
  MUX2_X1 U15341 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13152), .S(n14829), .Z(
        P2_U3488) );
  MUX2_X1 U15342 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13153), .S(n14829), .Z(
        P2_U3487) );
  MUX2_X1 U15343 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13154), .S(n14829), .Z(
        P2_U3486) );
  MUX2_X1 U15344 ( .A(n13155), .B(P2_REG0_REG_18__SCAN_IN), .S(n14827), .Z(
        P2_U3484) );
  MUX2_X1 U15345 ( .A(n13156), .B(P2_REG0_REG_17__SCAN_IN), .S(n14827), .Z(
        P2_U3481) );
  MUX2_X1 U15346 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13157), .S(n14829), .Z(
        P2_U3478) );
  MUX2_X1 U15347 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13158), .S(n14829), .Z(
        P2_U3475) );
  INV_X1 U15348 ( .A(n13473), .ZN(n14037) );
  NAND3_X1 U15349 ( .A1(n13159), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13161) );
  OAI22_X1 U15350 ( .A1(n8808), .A2(n13161), .B1(n15354), .B2(n13160), .ZN(
        n13162) );
  INV_X1 U15351 ( .A(n13162), .ZN(n13163) );
  OAI21_X1 U15352 ( .B1(n14037), .B2(n13178), .A(n13163), .ZN(P2_U3296) );
  NAND2_X1 U15353 ( .A1(n13165), .A2(n13164), .ZN(n13167) );
  OAI211_X1 U15354 ( .C1(n13160), .C2(n13168), .A(n13167), .B(n13166), .ZN(
        P2_U3299) );
  INV_X1 U15355 ( .A(n13169), .ZN(n14042) );
  OAI222_X1 U15356 ( .A1(n13160), .A2(n13172), .B1(n13178), .B2(n14042), .C1(
        P2_U3088), .C2(n6777), .ZN(P2_U3300) );
  INV_X1 U15357 ( .A(n13173), .ZN(n14045) );
  INV_X1 U15358 ( .A(n13174), .ZN(n13175) );
  OAI222_X1 U15359 ( .A1(n13178), .A2(n14045), .B1(n13175), .B2(P2_U3088), 
        .C1(n15293), .C2(n13160), .ZN(P2_U3301) );
  INV_X1 U15360 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15367) );
  INV_X1 U15361 ( .A(n13176), .ZN(n14049) );
  OAI222_X1 U15362 ( .A1(n13160), .A2(n15367), .B1(n13178), .B2(n14049), .C1(
        P2_U3088), .C2(n13177), .ZN(P2_U3302) );
  INV_X1 U15363 ( .A(n13179), .ZN(n13180) );
  MUX2_X1 U15364 ( .A(n13180), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15365 ( .A(n13182), .B(n13181), .Z(n13188) );
  AOI22_X1 U15366 ( .A1(n14353), .A2(n13183), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13184) );
  OAI21_X1 U15367 ( .B1(n14369), .B2(n13185), .A(n13184), .ZN(n13186) );
  AOI21_X1 U15368 ( .B1(n13915), .B2(n9693), .A(n13186), .ZN(n13187) );
  OAI21_X1 U15369 ( .B1(n13188), .B2(n13286), .A(n13187), .ZN(P1_U3214) );
  XOR2_X1 U15370 ( .A(n13190), .B(n13189), .Z(n13196) );
  NAND2_X1 U15371 ( .A1(n13554), .A2(n13864), .ZN(n13192) );
  NAND2_X1 U15372 ( .A1(n13552), .A2(n13262), .ZN(n13191) );
  NAND2_X1 U15373 ( .A1(n13192), .A2(n13191), .ZN(n13938) );
  AOI22_X1 U15374 ( .A1(n14353), .A2(n13938), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13193) );
  OAI21_X1 U15375 ( .B1(n14369), .B2(n13783), .A(n13193), .ZN(n13194) );
  AOI21_X1 U15376 ( .B1(n13939), .B2(n9693), .A(n13194), .ZN(n13195) );
  OAI21_X1 U15377 ( .B1(n13196), .B2(n13286), .A(n13195), .ZN(P1_U3216) );
  INV_X1 U15378 ( .A(n14022), .ZN(n13205) );
  OAI211_X1 U15379 ( .C1(n13199), .C2(n13198), .A(n13197), .B(n14365), .ZN(
        n13204) );
  OR2_X1 U15380 ( .A1(n13400), .A2(n13686), .ZN(n13201) );
  NAND2_X1 U15381 ( .A1(n13558), .A2(n13864), .ZN(n13200) );
  AND2_X1 U15382 ( .A1(n13201), .A2(n13200), .ZN(n13844) );
  NAND2_X1 U15383 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13680)
         );
  OAI21_X1 U15384 ( .B1(n13844), .B2(n14360), .A(n13680), .ZN(n13202) );
  AOI21_X1 U15385 ( .B1(n13850), .B2(n13293), .A(n13202), .ZN(n13203) );
  OAI211_X1 U15386 ( .C1(n13205), .C2(n14362), .A(n13204), .B(n13203), .ZN(
        P1_U3219) );
  INV_X1 U15387 ( .A(n13206), .ZN(n13207) );
  AOI21_X1 U15388 ( .B1(n13209), .B2(n13208), .A(n13207), .ZN(n13215) );
  OR2_X1 U15389 ( .A1(n13400), .A2(n13542), .ZN(n13211) );
  NAND2_X1 U15390 ( .A1(n13554), .A2(n13262), .ZN(n13210) );
  NAND2_X1 U15391 ( .A1(n13211), .A2(n13210), .ZN(n13811) );
  AOI22_X1 U15392 ( .A1(n13811), .A2(n14353), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13212) );
  OAI21_X1 U15393 ( .B1(n14369), .B2(n13814), .A(n13212), .ZN(n13213) );
  AOI21_X1 U15394 ( .B1(n13950), .B2(n9693), .A(n13213), .ZN(n13214) );
  OAI21_X1 U15395 ( .B1(n13215), .B2(n13286), .A(n13214), .ZN(P1_U3223) );
  XOR2_X1 U15396 ( .A(n13217), .B(n13216), .Z(n13223) );
  NAND2_X1 U15397 ( .A1(n13550), .A2(n13262), .ZN(n13219) );
  NAND2_X1 U15398 ( .A1(n13552), .A2(n13864), .ZN(n13218) );
  NAND2_X1 U15399 ( .A1(n13219), .A2(n13218), .ZN(n13749) );
  AOI22_X1 U15400 ( .A1(n14353), .A2(n13749), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13220) );
  OAI21_X1 U15401 ( .B1(n14369), .B2(n13752), .A(n13220), .ZN(n13221) );
  AOI21_X1 U15402 ( .B1(n14007), .B2(n9693), .A(n13221), .ZN(n13222) );
  OAI21_X1 U15403 ( .B1(n13223), .B2(n13286), .A(n13222), .ZN(P1_U3225) );
  OAI21_X1 U15404 ( .B1(n13226), .B2(n13225), .A(n13224), .ZN(n13227) );
  NAND2_X1 U15405 ( .A1(n13227), .A2(n14365), .ZN(n13232) );
  INV_X1 U15406 ( .A(n13228), .ZN(n13881) );
  AND2_X1 U15407 ( .A1(n13559), .A2(n13864), .ZN(n13229) );
  AOI21_X1 U15408 ( .B1(n13558), .B2(n13262), .A(n13229), .ZN(n13880) );
  NAND2_X1 U15409 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14477)
         );
  OAI21_X1 U15410 ( .B1(n13880), .B2(n14360), .A(n14477), .ZN(n13230) );
  AOI21_X1 U15411 ( .B1(n13293), .B2(n13881), .A(n13230), .ZN(n13231) );
  OAI211_X1 U15412 ( .C1(n6880), .C2(n14362), .A(n13232), .B(n13231), .ZN(
        P1_U3228) );
  XOR2_X1 U15413 ( .A(n13234), .B(n13233), .Z(n13240) );
  NAND2_X1 U15414 ( .A1(n13551), .A2(n13262), .ZN(n13236) );
  NAND2_X1 U15415 ( .A1(n13553), .A2(n13864), .ZN(n13235) );
  NAND2_X1 U15416 ( .A1(n13236), .A2(n13235), .ZN(n13762) );
  AOI22_X1 U15417 ( .A1(n14353), .A2(n13762), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13237) );
  OAI21_X1 U15418 ( .B1(n14369), .B2(n13770), .A(n13237), .ZN(n13238) );
  AOI21_X1 U15419 ( .B1(n14011), .B2(n9693), .A(n13238), .ZN(n13239) );
  OAI21_X1 U15420 ( .B1(n13240), .B2(n13286), .A(n13239), .ZN(P1_U3229) );
  OAI211_X1 U15421 ( .C1(n13243), .C2(n13242), .A(n13241), .B(n14365), .ZN(
        n13249) );
  OR2_X1 U15422 ( .A1(n13271), .A2(n13542), .ZN(n13245) );
  NAND2_X1 U15423 ( .A1(n13555), .A2(n13262), .ZN(n13244) );
  AND2_X1 U15424 ( .A1(n13245), .A2(n13244), .ZN(n13955) );
  OAI22_X1 U15425 ( .A1(n13955), .A2(n14360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13246), .ZN(n13247) );
  AOI21_X1 U15426 ( .B1(n13826), .B2(n13293), .A(n13247), .ZN(n13248) );
  OAI211_X1 U15427 ( .C1(n13831), .C2(n14362), .A(n13249), .B(n13248), .ZN(
        P1_U3233) );
  OAI211_X1 U15428 ( .C1(n13251), .C2(n13250), .A(n14350), .B(n14365), .ZN(
        n13257) );
  NAND2_X1 U15429 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14426)
         );
  INV_X1 U15430 ( .A(n14426), .ZN(n13254) );
  NOR2_X1 U15431 ( .A1(n14369), .A2(n13252), .ZN(n13253) );
  AOI211_X1 U15432 ( .C1(n14353), .C2(n13255), .A(n13254), .B(n13253), .ZN(
        n13256) );
  OAI211_X1 U15433 ( .C1(n6875), .C2(n14362), .A(n13257), .B(n13256), .ZN(
        P1_U3234) );
  OAI21_X1 U15434 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(n13261) );
  NAND2_X1 U15435 ( .A1(n13261), .A2(n14365), .ZN(n13267) );
  INV_X1 U15436 ( .A(n13802), .ZN(n13265) );
  AOI22_X1 U15437 ( .A1(n13864), .A2(n13555), .B1(n13553), .B2(n13262), .ZN(
        n13796) );
  INV_X1 U15438 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13263) );
  OAI22_X1 U15439 ( .A1(n14360), .A2(n13796), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13263), .ZN(n13264) );
  AOI21_X1 U15440 ( .B1(n13293), .B2(n13265), .A(n13264), .ZN(n13266) );
  OAI211_X1 U15441 ( .C1(n14362), .C2(n13268), .A(n13267), .B(n13266), .ZN(
        P1_U3235) );
  XOR2_X1 U15442 ( .A(n13270), .B(n13269), .Z(n13278) );
  NOR2_X1 U15443 ( .A1(n14369), .A2(n13870), .ZN(n13276) );
  NOR2_X1 U15444 ( .A1(n13271), .A2(n13686), .ZN(n13863) );
  NAND2_X1 U15445 ( .A1(n13863), .A2(n14353), .ZN(n13272) );
  NAND2_X1 U15446 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14497)
         );
  OAI211_X1 U15447 ( .C1(n13274), .C2(n13273), .A(n13272), .B(n14497), .ZN(
        n13275) );
  AOI211_X1 U15448 ( .C1(n13873), .C2(n9693), .A(n13276), .B(n13275), .ZN(
        n13277) );
  OAI21_X1 U15449 ( .B1(n13278), .B2(n13286), .A(n13277), .ZN(P1_U3238) );
  XOR2_X1 U15450 ( .A(n13280), .B(n13279), .Z(n13287) );
  OAI22_X1 U15451 ( .A1(n13282), .A2(n13542), .B1(n13281), .B2(n13686), .ZN(
        n13736) );
  AOI22_X1 U15452 ( .A1(n14353), .A2(n13736), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13283) );
  OAI21_X1 U15453 ( .B1(n14369), .B2(n13730), .A(n13283), .ZN(n13284) );
  AOI21_X1 U15454 ( .B1(n13729), .B2(n9693), .A(n13284), .ZN(n13285) );
  OAI21_X1 U15455 ( .B1(n13287), .B2(n13286), .A(n13285), .ZN(P1_U3240) );
  OAI211_X1 U15456 ( .C1(n13290), .C2(n13289), .A(n13288), .B(n14365), .ZN(
        n13295) );
  NAND2_X1 U15457 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14450)
         );
  OAI21_X1 U15458 ( .B1(n14360), .B2(n14387), .A(n14450), .ZN(n13291) );
  AOI21_X1 U15459 ( .B1(n13293), .B2(n13292), .A(n13291), .ZN(n13294) );
  OAI211_X1 U15460 ( .C1(n13296), .C2(n14362), .A(n13295), .B(n13294), .ZN(
        P1_U3241) );
  MUX2_X1 U15461 ( .A(n13549), .B(n13915), .S(n6563), .Z(n13428) );
  INV_X1 U15462 ( .A(n13314), .ZN(n13298) );
  NAND2_X1 U15463 ( .A1(n13298), .A2(n13485), .ZN(n13306) );
  NAND3_X1 U15464 ( .A1(n13300), .A2(n13485), .A3(n13299), .ZN(n13305) );
  NAND3_X1 U15465 ( .A1(n13314), .A2(n13301), .A3(n6563), .ZN(n13304) );
  INV_X1 U15466 ( .A(n13299), .ZN(n13302) );
  NAND2_X1 U15467 ( .A1(n13302), .A2(n6563), .ZN(n13303) );
  NAND2_X1 U15468 ( .A1(n13310), .A2(n13307), .ZN(n13309) );
  NAND2_X1 U15469 ( .A1(n13313), .A2(n13312), .ZN(n13315) );
  MUX2_X1 U15470 ( .A(n13319), .B(n13318), .S(n6563), .Z(n13320) );
  MUX2_X1 U15471 ( .A(n13321), .B(n14565), .S(n13485), .Z(n13324) );
  MUX2_X1 U15472 ( .A(n13571), .B(n13322), .S(n6563), .Z(n13323) );
  MUX2_X1 U15473 ( .A(n13570), .B(n14571), .S(n6563), .Z(n13327) );
  MUX2_X1 U15474 ( .A(n13570), .B(n14571), .S(n13485), .Z(n13326) );
  INV_X1 U15475 ( .A(n13327), .ZN(n13328) );
  NAND2_X1 U15476 ( .A1(n6662), .A2(n13328), .ZN(n13329) );
  MUX2_X1 U15477 ( .A(n13569), .B(n13330), .S(n13485), .Z(n13332) );
  MUX2_X1 U15478 ( .A(n13569), .B(n13330), .S(n6563), .Z(n13331) );
  MUX2_X1 U15479 ( .A(n13568), .B(n13333), .S(n6563), .Z(n13337) );
  NAND2_X1 U15480 ( .A1(n13336), .A2(n13337), .ZN(n13335) );
  MUX2_X1 U15481 ( .A(n13568), .B(n13333), .S(n13485), .Z(n13334) );
  NAND2_X1 U15482 ( .A1(n13335), .A2(n13334), .ZN(n13341) );
  INV_X1 U15483 ( .A(n13336), .ZN(n13339) );
  INV_X1 U15484 ( .A(n13337), .ZN(n13338) );
  NAND2_X1 U15485 ( .A1(n13339), .A2(n13338), .ZN(n13340) );
  MUX2_X1 U15486 ( .A(n13567), .B(n14578), .S(n13485), .Z(n13343) );
  MUX2_X1 U15487 ( .A(n13567), .B(n14578), .S(n6563), .Z(n13342) );
  INV_X1 U15488 ( .A(n13343), .ZN(n13344) );
  MUX2_X1 U15489 ( .A(n13566), .B(n13345), .S(n6563), .Z(n13348) );
  MUX2_X1 U15490 ( .A(n13566), .B(n13345), .S(n13485), .Z(n13346) );
  INV_X1 U15491 ( .A(n13347), .ZN(n13350) );
  INV_X1 U15492 ( .A(n13348), .ZN(n13349) );
  NAND2_X1 U15493 ( .A1(n13350), .A2(n13349), .ZN(n13351) );
  MUX2_X1 U15494 ( .A(n13565), .B(n13352), .S(n13485), .Z(n13354) );
  MUX2_X1 U15495 ( .A(n13565), .B(n13352), .S(n6563), .Z(n13353) );
  MUX2_X1 U15496 ( .A(n13564), .B(n13355), .S(n6563), .Z(n13359) );
  NAND2_X1 U15497 ( .A1(n13358), .A2(n13359), .ZN(n13357) );
  MUX2_X1 U15498 ( .A(n13564), .B(n13355), .S(n13485), .Z(n13356) );
  INV_X1 U15499 ( .A(n13358), .ZN(n13361) );
  INV_X1 U15500 ( .A(n13359), .ZN(n13360) );
  NAND2_X1 U15501 ( .A1(n13361), .A2(n13360), .ZN(n13362) );
  MUX2_X1 U15502 ( .A(n13563), .B(n13363), .S(n13485), .Z(n13365) );
  MUX2_X1 U15503 ( .A(n13563), .B(n13363), .S(n6563), .Z(n13364) );
  MUX2_X1 U15504 ( .A(n13562), .B(n13366), .S(n6563), .Z(n13370) );
  NAND2_X1 U15505 ( .A1(n13369), .A2(n13370), .ZN(n13368) );
  MUX2_X1 U15506 ( .A(n13562), .B(n13366), .S(n13485), .Z(n13367) );
  INV_X1 U15507 ( .A(n13369), .ZN(n13371) );
  NAND2_X1 U15508 ( .A1(n13378), .A2(n13372), .ZN(n13375) );
  NAND2_X1 U15509 ( .A1(n13379), .A2(n13373), .ZN(n13374) );
  MUX2_X1 U15510 ( .A(n13375), .B(n13374), .S(n13485), .Z(n13376) );
  INV_X1 U15511 ( .A(n13378), .ZN(n13381) );
  INV_X1 U15512 ( .A(n13379), .ZN(n13380) );
  MUX2_X1 U15513 ( .A(n13381), .B(n13380), .S(n6563), .Z(n13382) );
  MUX2_X1 U15514 ( .A(n13559), .B(n13988), .S(n6563), .Z(n13386) );
  NAND2_X1 U15515 ( .A1(n13385), .A2(n13386), .ZN(n13384) );
  MUX2_X1 U15516 ( .A(n13559), .B(n13988), .S(n13485), .Z(n13383) );
  NOR2_X1 U15517 ( .A1(n13386), .A2(n13385), .ZN(n13390) );
  MUX2_X1 U15518 ( .A(n13388), .B(n13387), .S(n13485), .Z(n13389) );
  MUX2_X1 U15519 ( .A(n13865), .B(n13979), .S(n6563), .Z(n13391) );
  MUX2_X1 U15520 ( .A(n13558), .B(n13873), .S(n13485), .Z(n13395) );
  MUX2_X1 U15521 ( .A(n13398), .B(n13397), .S(n6563), .Z(n13399) );
  MUX2_X1 U15522 ( .A(n13400), .B(n13831), .S(n6563), .Z(n13402) );
  MUX2_X1 U15523 ( .A(n13556), .B(n14018), .S(n13485), .Z(n13401) );
  MUX2_X1 U15524 ( .A(n13555), .B(n13950), .S(n13485), .Z(n13405) );
  MUX2_X1 U15525 ( .A(n13555), .B(n13950), .S(n6563), .Z(n13403) );
  NAND2_X1 U15526 ( .A1(n13404), .A2(n13403), .ZN(n13406) );
  MUX2_X1 U15527 ( .A(n13554), .B(n13946), .S(n6563), .Z(n13408) );
  MUX2_X1 U15528 ( .A(n13554), .B(n13946), .S(n13485), .Z(n13407) );
  INV_X1 U15529 ( .A(n13408), .ZN(n13409) );
  MUX2_X1 U15530 ( .A(n13553), .B(n13939), .S(n13485), .Z(n13412) );
  MUX2_X1 U15531 ( .A(n13553), .B(n13939), .S(n6563), .Z(n13410) );
  INV_X1 U15532 ( .A(n13412), .ZN(n13413) );
  MUX2_X1 U15533 ( .A(n13552), .B(n14011), .S(n6563), .Z(n13416) );
  MUX2_X1 U15534 ( .A(n14011), .B(n13552), .S(n6563), .Z(n13414) );
  INV_X1 U15535 ( .A(n13416), .ZN(n13417) );
  MUX2_X1 U15536 ( .A(n13551), .B(n14007), .S(n13485), .Z(n13421) );
  NAND2_X1 U15537 ( .A1(n13420), .A2(n13421), .ZN(n13419) );
  MUX2_X1 U15538 ( .A(n13551), .B(n14007), .S(n6563), .Z(n13418) );
  INV_X1 U15539 ( .A(n13421), .ZN(n13422) );
  NAND2_X1 U15540 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  MUX2_X1 U15541 ( .A(n13550), .B(n13729), .S(n6563), .Z(n13426) );
  MUX2_X1 U15542 ( .A(n13729), .B(n13550), .S(n6563), .Z(n13425) );
  MUX2_X1 U15543 ( .A(n13549), .B(n13915), .S(n13485), .Z(n13427) );
  MUX2_X1 U15544 ( .A(n13430), .B(n13429), .S(n6563), .Z(n13432) );
  INV_X1 U15545 ( .A(n13430), .ZN(n13708) );
  MUX2_X1 U15546 ( .A(n13721), .B(n13708), .S(n6563), .Z(n13431) );
  OAI21_X1 U15547 ( .B1(n13433), .B2(n13432), .A(n13431), .ZN(n13460) );
  NAND2_X1 U15548 ( .A1(n13433), .A2(n13432), .ZN(n13459) );
  INV_X1 U15549 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13437) );
  NAND2_X1 U15550 ( .A1(n13434), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U15551 ( .A1(n13439), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n13435) );
  OAI211_X1 U15552 ( .C1(n13438), .C2(n13437), .A(n13436), .B(n13435), .ZN(
        n13687) );
  INV_X1 U15553 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15305) );
  NAND2_X1 U15554 ( .A1(n7991), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13441) );
  NAND2_X1 U15555 ( .A1(n13439), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n13440) );
  OAI211_X1 U15556 ( .C1(n13442), .C2(n15305), .A(n13441), .B(n13440), .ZN(
        n13705) );
  OAI21_X1 U15557 ( .B1(n13687), .B2(n13477), .A(n13705), .ZN(n13443) );
  INV_X1 U15558 ( .A(n13443), .ZN(n13448) );
  OR2_X1 U15559 ( .A1(n13445), .A2(n13444), .ZN(n13447) );
  NAND2_X1 U15560 ( .A1(n13474), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13446) );
  MUX2_X1 U15561 ( .A(n13448), .B(n13997), .S(n13485), .Z(n13464) );
  NAND2_X1 U15562 ( .A1(n13997), .A2(n6563), .ZN(n13453) );
  INV_X1 U15563 ( .A(n13687), .ZN(n13489) );
  OAI22_X1 U15564 ( .A1(n6563), .A2(n13489), .B1(n13450), .B2(n13449), .ZN(
        n13451) );
  NAND2_X1 U15565 ( .A1(n13451), .A2(n13705), .ZN(n13452) );
  AND2_X1 U15566 ( .A1(n13453), .A2(n13452), .ZN(n13469) );
  NAND2_X1 U15567 ( .A1(n13454), .A2(n13472), .ZN(n13456) );
  NAND2_X1 U15568 ( .A1(n13474), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13455) );
  MUX2_X1 U15569 ( .A(n13548), .B(n13905), .S(n6563), .Z(n13462) );
  INV_X1 U15570 ( .A(n13462), .ZN(n13457) );
  MUX2_X1 U15571 ( .A(n13905), .B(n13548), .S(n6563), .Z(n13461) );
  AOI22_X1 U15572 ( .A1(n13464), .A2(n13469), .B1(n13457), .B2(n13461), .ZN(
        n13458) );
  NAND3_X1 U15573 ( .A1(n13460), .A2(n13459), .A3(n13458), .ZN(n13471) );
  INV_X1 U15574 ( .A(n13461), .ZN(n13463) );
  AND2_X1 U15575 ( .A1(n13463), .A2(n13462), .ZN(n13467) );
  INV_X1 U15576 ( .A(n13469), .ZN(n13466) );
  INV_X1 U15577 ( .A(n13464), .ZN(n13465) );
  OAI21_X1 U15578 ( .B1(n13467), .B2(n13466), .A(n13465), .ZN(n13470) );
  INV_X1 U15579 ( .A(n13467), .ZN(n13468) );
  NAND2_X1 U15580 ( .A1(n13471), .A2(n7541), .ZN(n13491) );
  NAND2_X1 U15581 ( .A1(n13473), .A2(n13472), .ZN(n13476) );
  NAND2_X1 U15582 ( .A1(n13474), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n13475) );
  NOR2_X1 U15583 ( .A1(n13526), .A2(n13485), .ZN(n13531) );
  INV_X1 U15584 ( .A(n13297), .ZN(n13478) );
  NAND2_X1 U15585 ( .A1(n13478), .A2(n13477), .ZN(n13479) );
  NAND2_X1 U15586 ( .A1(n13480), .A2(n13479), .ZN(n13482) );
  NAND2_X1 U15587 ( .A1(n13482), .A2(n13481), .ZN(n13532) );
  NAND2_X1 U15588 ( .A1(n13484), .A2(n13483), .ZN(n13536) );
  NAND2_X1 U15589 ( .A1(n13532), .A2(n13536), .ZN(n13527) );
  NAND2_X1 U15590 ( .A1(n13526), .A2(n13485), .ZN(n13529) );
  NOR2_X1 U15591 ( .A1(n13529), .A2(n13687), .ZN(n13486) );
  AOI211_X1 U15592 ( .C1(n13531), .C2(n13687), .A(n13527), .B(n13486), .ZN(
        n13487) );
  INV_X1 U15593 ( .A(n13487), .ZN(n13488) );
  XNOR2_X1 U15594 ( .A(n13526), .B(n13489), .ZN(n13492) );
  NOR2_X1 U15595 ( .A1(n13492), .A2(n13532), .ZN(n13490) );
  XNOR2_X1 U15596 ( .A(n13997), .B(n13705), .ZN(n13523) );
  INV_X1 U15597 ( .A(n13492), .ZN(n13522) );
  NAND2_X1 U15598 ( .A1(n14530), .A2(n13493), .ZN(n13494) );
  NOR4_X1 U15599 ( .A1(n13496), .A2(n14502), .A3(n13495), .A4(n13494), .ZN(
        n13499) );
  NAND4_X1 U15600 ( .A1(n13500), .A2(n13499), .A3(n13498), .A4(n13497), .ZN(
        n13501) );
  NOR4_X1 U15601 ( .A1(n13504), .A2(n13503), .A3(n13502), .A4(n13501), .ZN(
        n13507) );
  NAND4_X1 U15602 ( .A1(n13508), .A2(n13507), .A3(n13506), .A4(n13505), .ZN(
        n13509) );
  NOR4_X1 U15603 ( .A1(n13891), .A2(n6984), .A3(n13510), .A4(n13509), .ZN(
        n13512) );
  NAND4_X1 U15604 ( .A1(n13513), .A2(n13512), .A3(n13511), .A4(n13862), .ZN(
        n13514) );
  NOR4_X1 U15605 ( .A1(n13795), .A2(n13825), .A3(n13808), .A4(n13514), .ZN(
        n13515) );
  NAND4_X1 U15606 ( .A1(n13516), .A2(n13515), .A3(n13778), .A4(n13760), .ZN(
        n13517) );
  NOR4_X1 U15607 ( .A1(n13519), .A2(n13518), .A3(n13734), .A4(n13517), .ZN(
        n13520) );
  XNOR2_X1 U15608 ( .A(n13905), .B(n13548), .ZN(n13699) );
  NAND3_X1 U15609 ( .A1(n13523), .A2(n13522), .A3(n13521), .ZN(n13524) );
  XOR2_X1 U15610 ( .A(n13525), .B(n13524), .Z(n13537) );
  NOR3_X1 U15611 ( .A1(n13994), .A2(n13687), .A3(n13527), .ZN(n13530) );
  NOR3_X1 U15612 ( .A1(n13529), .A2(n13687), .A3(n13532), .ZN(n13528) );
  AOI21_X1 U15613 ( .B1(n13530), .B2(n13529), .A(n13528), .ZN(n13535) );
  XOR2_X1 U15614 ( .A(n13532), .B(n13531), .Z(n13533) );
  NAND4_X1 U15615 ( .A1(n13533), .A2(n13994), .A3(n13687), .A4(n13536), .ZN(
        n13534) );
  OAI211_X1 U15616 ( .C1(n13537), .C2(n13536), .A(n13535), .B(n13534), .ZN(
        n13538) );
  INV_X1 U15617 ( .A(n13538), .ZN(n13539) );
  NOR3_X1 U15618 ( .A1(n13543), .A2(n14041), .A3(n13542), .ZN(n13545) );
  OAI21_X1 U15619 ( .B1(n13546), .B2(n13297), .A(P1_B_REG_SCAN_IN), .ZN(n13544) );
  OAI22_X1 U15620 ( .A1(n13547), .A2(n13546), .B1(n13545), .B2(n13544), .ZN(
        P1_U3242) );
  MUX2_X1 U15621 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13687), .S(n13591), .Z(
        P1_U3591) );
  MUX2_X1 U15622 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13705), .S(n13591), .Z(
        P1_U3590) );
  MUX2_X1 U15623 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13548), .S(n13591), .Z(
        P1_U3589) );
  MUX2_X1 U15624 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13708), .S(n13591), .Z(
        P1_U3588) );
  MUX2_X1 U15625 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13549), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15626 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13550), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15627 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13551), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15628 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13552), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15629 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13553), .S(n13591), .Z(
        P1_U3583) );
  MUX2_X1 U15630 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13554), .S(n13591), .Z(
        P1_U3582) );
  MUX2_X1 U15631 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13555), .S(n13591), .Z(
        P1_U3581) );
  MUX2_X1 U15632 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13556), .S(n13591), .Z(
        P1_U3580) );
  MUX2_X1 U15633 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13557), .S(n13591), .Z(
        P1_U3579) );
  MUX2_X1 U15634 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13558), .S(n13591), .Z(
        P1_U3578) );
  MUX2_X1 U15635 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13865), .S(n13591), .Z(
        P1_U3577) );
  MUX2_X1 U15636 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13559), .S(n13591), .Z(
        P1_U3576) );
  MUX2_X1 U15637 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13560), .S(n13591), .Z(
        P1_U3575) );
  MUX2_X1 U15638 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13561), .S(n13591), .Z(
        P1_U3574) );
  MUX2_X1 U15639 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13562), .S(n13591), .Z(
        P1_U3573) );
  MUX2_X1 U15640 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13563), .S(n13591), .Z(
        P1_U3572) );
  MUX2_X1 U15641 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13564), .S(n13591), .Z(
        P1_U3571) );
  MUX2_X1 U15642 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13565), .S(n13591), .Z(
        P1_U3570) );
  MUX2_X1 U15643 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13566), .S(n13591), .Z(
        P1_U3569) );
  MUX2_X1 U15644 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13567), .S(n13591), .Z(
        P1_U3568) );
  MUX2_X1 U15645 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13568), .S(n13591), .Z(
        P1_U3567) );
  MUX2_X1 U15646 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13569), .S(n13591), .Z(
        P1_U3566) );
  MUX2_X1 U15647 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13570), .S(n13591), .Z(
        P1_U3565) );
  MUX2_X1 U15648 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13571), .S(n13591), .Z(
        P1_U3564) );
  MUX2_X1 U15649 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13572), .S(n13591), .Z(
        P1_U3563) );
  MUX2_X1 U15650 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13573), .S(n13591), .Z(
        P1_U3562) );
  MUX2_X1 U15651 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13574), .S(n13591), .Z(
        P1_U3560) );
  OAI22_X1 U15652 ( .A1(n14499), .A2(n7224), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13575), .ZN(n13576) );
  AOI21_X1 U15653 ( .B1(n13577), .B2(n14493), .A(n13576), .ZN(n13585) );
  OAI211_X1 U15654 ( .C1(n13580), .C2(n13579), .A(n14483), .B(n13578), .ZN(
        n13584) );
  OAI211_X1 U15655 ( .C1(n13582), .C2(n13587), .A(n14468), .B(n13581), .ZN(
        n13583) );
  NAND3_X1 U15656 ( .A1(n13585), .A2(n13584), .A3(n13583), .ZN(P1_U3244) );
  MUX2_X1 U15657 ( .A(n13588), .B(n13587), .S(n13586), .Z(n13590) );
  NAND2_X1 U15658 ( .A1(n13590), .A2(n13589), .ZN(n13592) );
  OAI211_X1 U15659 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n13593), .A(n13592), .B(
        n13591), .ZN(n13632) );
  OAI22_X1 U15660 ( .A1(n14499), .A2(n14053), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13594), .ZN(n13595) );
  AOI21_X1 U15661 ( .B1(n13596), .B2(n14493), .A(n13595), .ZN(n13605) );
  OAI211_X1 U15662 ( .C1(n13599), .C2(n13598), .A(n14468), .B(n13597), .ZN(
        n13604) );
  OAI211_X1 U15663 ( .C1(n13602), .C2(n13601), .A(n14483), .B(n13600), .ZN(
        n13603) );
  NAND4_X1 U15664 ( .A1(n13632), .A2(n13605), .A3(n13604), .A4(n13603), .ZN(
        P1_U3245) );
  INV_X1 U15665 ( .A(n13606), .ZN(n13609) );
  INV_X1 U15666 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14107) );
  OAI21_X1 U15667 ( .B1(n14499), .B2(n14107), .A(n13607), .ZN(n13608) );
  AOI21_X1 U15668 ( .B1(n13609), .B2(n14493), .A(n13608), .ZN(n13618) );
  OAI211_X1 U15669 ( .C1(n13612), .C2(n13611), .A(n14468), .B(n13610), .ZN(
        n13617) );
  OAI211_X1 U15670 ( .C1(n13615), .C2(n13614), .A(n14483), .B(n13613), .ZN(
        n13616) );
  NAND3_X1 U15671 ( .A1(n13618), .A2(n13617), .A3(n13616), .ZN(P1_U3246) );
  OAI21_X1 U15672 ( .B1(n14499), .B2(n6774), .A(n13619), .ZN(n13620) );
  INV_X1 U15673 ( .A(n13620), .ZN(n13631) );
  NOR2_X1 U15674 ( .A1(n13622), .A2(n13621), .ZN(n13623) );
  NOR2_X1 U15675 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  AOI22_X1 U15676 ( .A1(n13626), .A2(n14493), .B1(n14483), .B2(n13625), .ZN(
        n13630) );
  OAI211_X1 U15677 ( .C1(n13628), .C2(n13627), .A(n14468), .B(n6815), .ZN(
        n13629) );
  NAND4_X1 U15678 ( .A1(n13632), .A2(n13631), .A3(n13630), .A4(n13629), .ZN(
        P1_U3247) );
  AOI21_X1 U15679 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n13642), .A(n13633), 
        .ZN(n13636) );
  MUX2_X1 U15680 ( .A(n10867), .B(P1_REG2_REG_12__SCAN_IN), .S(n13666), .Z(
        n13634) );
  INV_X1 U15681 ( .A(n13634), .ZN(n13635) );
  NAND2_X1 U15682 ( .A1(n13636), .A2(n13635), .ZN(n13665) );
  OAI21_X1 U15683 ( .B1(n13636), .B2(n13635), .A(n13665), .ZN(n13637) );
  NAND2_X1 U15684 ( .A1(n13637), .A2(n14468), .ZN(n13649) );
  AOI21_X1 U15685 ( .B1(n13639), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n13638), 
        .ZN(n13648) );
  MUX2_X1 U15686 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n13640), .S(n13666), .Z(
        n13644) );
  OAI21_X1 U15687 ( .B1(n13644), .B2(n13643), .A(n13652), .ZN(n13645) );
  NAND2_X1 U15688 ( .A1(n13645), .A2(n14483), .ZN(n13647) );
  NAND2_X1 U15689 ( .A1(n14493), .A2(n13666), .ZN(n13646) );
  NAND4_X1 U15690 ( .A1(n13649), .A2(n13648), .A3(n13647), .A4(n13646), .ZN(
        P1_U3255) );
  INV_X1 U15691 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13650) );
  XNOR2_X1 U15692 ( .A(n13671), .B(n13650), .ZN(n14467) );
  NAND2_X1 U15693 ( .A1(n14461), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n13657) );
  XNOR2_X1 U15694 ( .A(n14461), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14454) );
  MUX2_X1 U15695 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n13651), .S(n13667), .Z(
        n14430) );
  OAI21_X1 U15696 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n13666), .A(n13652), 
        .ZN(n14419) );
  MUX2_X1 U15697 ( .A(n13653), .B(P1_REG1_REG_13__SCAN_IN), .S(n14425), .Z(
        n14418) );
  NOR2_X1 U15698 ( .A1(n14419), .A2(n14418), .ZN(n14417) );
  NAND2_X1 U15699 ( .A1(n14430), .A2(n14431), .ZN(n14429) );
  OAI21_X1 U15700 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n13667), .A(n14429), 
        .ZN(n13654) );
  NAND2_X1 U15701 ( .A1(n14445), .A2(n13654), .ZN(n13655) );
  INV_X1 U15702 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U15703 ( .A1(n13655), .A2(n14442), .ZN(n14455) );
  NOR2_X1 U15704 ( .A1(n14454), .A2(n14455), .ZN(n14453) );
  INV_X1 U15705 ( .A(n14453), .ZN(n13656) );
  NAND2_X1 U15706 ( .A1(n13657), .A2(n13656), .ZN(n14466) );
  NAND2_X1 U15707 ( .A1(n14467), .A2(n14466), .ZN(n14465) );
  NAND2_X1 U15708 ( .A1(n13671), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n13658) );
  XNOR2_X1 U15709 ( .A(n13659), .B(n14491), .ZN(n14480) );
  NOR2_X1 U15710 ( .A1(n14479), .A2(n14480), .ZN(n14481) );
  NOR2_X1 U15711 ( .A1(n13659), .A2(n14491), .ZN(n13660) );
  NOR2_X1 U15712 ( .A1(n14481), .A2(n13660), .ZN(n13662) );
  INV_X1 U15713 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13883) );
  XNOR2_X1 U15714 ( .A(n13671), .B(n13883), .ZN(n14471) );
  NAND2_X1 U15715 ( .A1(n14461), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13670) );
  OAI21_X1 U15716 ( .B1(n14461), .B2(P1_REG2_REG_16__SCAN_IN), .A(n13670), 
        .ZN(n14457) );
  MUX2_X1 U15717 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n7806), .S(n13667), .Z(
        n13663) );
  INV_X1 U15718 ( .A(n13663), .ZN(n14434) );
  MUX2_X1 U15719 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11075), .S(n14425), .Z(
        n13664) );
  INV_X1 U15720 ( .A(n13664), .ZN(n14421) );
  OAI21_X1 U15721 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n13666), .A(n13665), 
        .ZN(n14422) );
  NOR2_X1 U15722 ( .A1(n14421), .A2(n14422), .ZN(n14420) );
  NAND2_X1 U15723 ( .A1(n13668), .A2(n14445), .ZN(n13669) );
  NAND2_X1 U15724 ( .A1(n14447), .A2(n7840), .ZN(n14446) );
  NAND2_X1 U15725 ( .A1(n14471), .A2(n14470), .ZN(n14469) );
  NAND2_X1 U15726 ( .A1(n13671), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13672) );
  NOR2_X1 U15727 ( .A1(n13673), .A2(n14491), .ZN(n13674) );
  INV_X1 U15728 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14485) );
  XNOR2_X1 U15729 ( .A(n13673), .B(n14491), .ZN(n14486) );
  NOR2_X1 U15730 ( .A1(n14485), .A2(n14486), .ZN(n14487) );
  NOR2_X1 U15731 ( .A1(n13674), .A2(n14487), .ZN(n13675) );
  XNOR2_X1 U15732 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13675), .ZN(n13677) );
  AOI22_X1 U15733 ( .A1(n13678), .A2(n14483), .B1(n13677), .B2(n14468), .ZN(
        n13679) );
  NOR2_X1 U15734 ( .A1(n13997), .A2(n13703), .ZN(n13682) );
  XNOR2_X1 U15735 ( .A(n13994), .B(n13682), .ZN(n13683) );
  NOR2_X2 U15736 ( .A1(n13683), .A2(n13884), .ZN(n13898) );
  NAND2_X1 U15737 ( .A1(n13898), .A2(n14517), .ZN(n13689) );
  NOR2_X1 U15738 ( .A1(n14041), .A2(n13684), .ZN(n13685) );
  NOR2_X1 U15739 ( .A1(n13686), .A2(n13685), .ZN(n13704) );
  AND2_X1 U15740 ( .A1(n13687), .A2(n13704), .ZN(n13897) );
  INV_X1 U15741 ( .A(n13897), .ZN(n13901) );
  NOR2_X1 U15742 ( .A1(n14521), .A2(n13901), .ZN(n13692) );
  AOI21_X1 U15743 ( .B1(n14521), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13692), 
        .ZN(n13688) );
  OAI211_X1 U15744 ( .C1(n13994), .C2(n14376), .A(n13689), .B(n13688), .ZN(
        P1_U3263) );
  XNOR2_X1 U15745 ( .A(n13690), .B(n13997), .ZN(n13691) );
  NAND2_X1 U15746 ( .A1(n13691), .A2(n14513), .ZN(n13902) );
  AOI21_X1 U15747 ( .B1(n14521), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13692), 
        .ZN(n13694) );
  NAND2_X1 U15748 ( .A1(n13997), .A2(n14512), .ZN(n13693) );
  OAI211_X1 U15749 ( .C1(n13902), .C2(n13888), .A(n13694), .B(n13693), .ZN(
        P1_U3264) );
  XNOR2_X1 U15750 ( .A(n13696), .B(n13699), .ZN(n13913) );
  NAND2_X1 U15751 ( .A1(n13698), .A2(n13697), .ZN(n13700) );
  XNOR2_X1 U15752 ( .A(n13700), .B(n13699), .ZN(n13911) );
  NAND2_X1 U15753 ( .A1(n13905), .A2(n13701), .ZN(n13702) );
  NAND3_X1 U15754 ( .A1(n13703), .A2(n14513), .A3(n13702), .ZN(n13909) );
  NAND2_X1 U15755 ( .A1(n13705), .A2(n13704), .ZN(n13906) );
  OAI22_X1 U15756 ( .A1(n13707), .A2(n13906), .B1(n14508), .B2(n13706), .ZN(
        n13710) );
  NAND2_X1 U15757 ( .A1(n13708), .A2(n13864), .ZN(n13907) );
  NOR2_X1 U15758 ( .A1(n14521), .A2(n13907), .ZN(n13709) );
  AOI211_X1 U15759 ( .C1(n14521), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13710), 
        .B(n13709), .ZN(n13712) );
  NAND2_X1 U15760 ( .A1(n13905), .A2(n14512), .ZN(n13711) );
  OAI211_X1 U15761 ( .C1(n13909), .C2(n13888), .A(n13712), .B(n13711), .ZN(
        n13713) );
  AOI21_X1 U15762 ( .B1(n13911), .B2(n14532), .A(n13713), .ZN(n13714) );
  OAI21_X1 U15763 ( .B1(n13913), .B2(n13895), .A(n13714), .ZN(P1_U3356) );
  OR2_X1 U15764 ( .A1(n13715), .A2(n14521), .ZN(n13723) );
  OAI22_X1 U15765 ( .A1(n14536), .A2(n13717), .B1(n13716), .B2(n14508), .ZN(
        n13720) );
  NOR2_X1 U15766 ( .A1(n13718), .A2(n13888), .ZN(n13719) );
  AOI211_X1 U15767 ( .C1(n14512), .C2(n13721), .A(n13720), .B(n13719), .ZN(
        n13722) );
  OAI211_X1 U15768 ( .C1(n13895), .C2(n13724), .A(n13723), .B(n13722), .ZN(
        P1_U3265) );
  XOR2_X1 U15769 ( .A(n13725), .B(n13734), .Z(n13921) );
  INV_X1 U15770 ( .A(n13921), .ZN(n13741) );
  INV_X1 U15771 ( .A(n13727), .ZN(n13728) );
  AOI211_X1 U15772 ( .C1(n13729), .C2(n13751), .A(n13884), .B(n13728), .ZN(
        n13920) );
  INV_X1 U15773 ( .A(n13730), .ZN(n13731) );
  AOI22_X1 U15774 ( .A1(n14521), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13731), 
        .B2(n14528), .ZN(n13732) );
  OAI21_X1 U15775 ( .B1(n14004), .B2(n14376), .A(n13732), .ZN(n13733) );
  AOI21_X1 U15776 ( .B1(n13920), .B2(n14517), .A(n13733), .ZN(n13740) );
  XNOR2_X1 U15777 ( .A(n13735), .B(n13734), .ZN(n13738) );
  INV_X1 U15778 ( .A(n13736), .ZN(n13737) );
  OAI21_X1 U15779 ( .B1(n13738), .B2(n14505), .A(n13737), .ZN(n13919) );
  NAND2_X1 U15780 ( .A1(n13919), .A2(n14536), .ZN(n13739) );
  OAI211_X1 U15781 ( .C1(n13741), .C2(n13895), .A(n13740), .B(n13739), .ZN(
        P1_U3267) );
  OAI21_X1 U15782 ( .B1(n13743), .B2(n13744), .A(n13742), .ZN(n13928) );
  NOR2_X1 U15783 ( .A1(n13928), .A2(n13895), .ZN(n13758) );
  NAND2_X1 U15784 ( .A1(n13745), .A2(n13744), .ZN(n13746) );
  NAND2_X1 U15785 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  NAND2_X1 U15786 ( .A1(n13748), .A2(n14585), .ZN(n13926) );
  INV_X1 U15787 ( .A(n13749), .ZN(n13924) );
  AOI21_X1 U15788 ( .B1(n13926), .B2(n13924), .A(n14521), .ZN(n13757) );
  NAND2_X1 U15789 ( .A1(n13769), .A2(n14007), .ZN(n13750) );
  NAND3_X1 U15790 ( .A1(n13751), .A2(n14513), .A3(n13750), .ZN(n13925) );
  INV_X1 U15791 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n13753) );
  OAI22_X1 U15792 ( .A1(n14536), .A2(n13753), .B1(n13752), .B2(n14508), .ZN(
        n13754) );
  AOI21_X1 U15793 ( .B1(n14007), .B2(n14512), .A(n13754), .ZN(n13755) );
  OAI21_X1 U15794 ( .B1(n13925), .B2(n13888), .A(n13755), .ZN(n13756) );
  OR3_X1 U15795 ( .A1(n13758), .A2(n13757), .A3(n13756), .ZN(P1_U3268) );
  OAI211_X1 U15796 ( .C1(n13761), .C2(n13760), .A(n13759), .B(n14585), .ZN(
        n13764) );
  INV_X1 U15797 ( .A(n13762), .ZN(n13763) );
  AND2_X1 U15798 ( .A1(n13764), .A2(n13763), .ZN(n13934) );
  OAI21_X1 U15799 ( .B1(n13767), .B2(n13766), .A(n13765), .ZN(n13931) );
  AOI21_X1 U15800 ( .B1(n13781), .B2(n14011), .A(n13884), .ZN(n13768) );
  NAND2_X1 U15801 ( .A1(n13769), .A2(n13768), .ZN(n13932) );
  INV_X1 U15802 ( .A(n13770), .ZN(n13771) );
  AOI22_X1 U15803 ( .A1(n14521), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13771), 
        .B2(n14528), .ZN(n13773) );
  NAND2_X1 U15804 ( .A1(n14011), .A2(n14512), .ZN(n13772) );
  OAI211_X1 U15805 ( .C1(n13932), .C2(n13888), .A(n13773), .B(n13772), .ZN(
        n13774) );
  AOI21_X1 U15806 ( .B1(n13931), .B2(n13775), .A(n13774), .ZN(n13776) );
  OAI21_X1 U15807 ( .B1(n13934), .B2(n14521), .A(n13776), .ZN(P1_U3269) );
  XNOR2_X1 U15808 ( .A(n13777), .B(n13778), .ZN(n13943) );
  XNOR2_X1 U15809 ( .A(n13779), .B(n13778), .ZN(n13940) );
  NAND2_X1 U15810 ( .A1(n13940), .A2(n14532), .ZN(n13790) );
  AOI21_X1 U15811 ( .B1(n13798), .B2(n13939), .A(n13884), .ZN(n13782) );
  AND2_X1 U15812 ( .A1(n13782), .A2(n13781), .ZN(n13937) );
  NAND2_X1 U15813 ( .A1(n13939), .A2(n14512), .ZN(n13787) );
  NOR2_X1 U15814 ( .A1(n14508), .A2(n13783), .ZN(n13784) );
  AOI21_X1 U15815 ( .B1(n14536), .B2(n13938), .A(n13784), .ZN(n13786) );
  NAND2_X1 U15816 ( .A1(n14521), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n13785) );
  NAND3_X1 U15817 ( .A1(n13787), .A2(n13786), .A3(n13785), .ZN(n13788) );
  AOI21_X1 U15818 ( .B1(n13937), .B2(n14517), .A(n13788), .ZN(n13789) );
  OAI211_X1 U15819 ( .C1(n13943), .C2(n13895), .A(n13790), .B(n13789), .ZN(
        P1_U3270) );
  XOR2_X1 U15820 ( .A(n13791), .B(n13795), .Z(n13948) );
  INV_X1 U15821 ( .A(n13792), .ZN(n13793) );
  AOI21_X1 U15822 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n13797) );
  OAI21_X1 U15823 ( .B1(n13797), .B2(n14505), .A(n13796), .ZN(n13944) );
  NAND2_X1 U15824 ( .A1(n13944), .A2(n14536), .ZN(n13805) );
  AOI21_X1 U15825 ( .B1(n13946), .B2(n6607), .A(n13884), .ZN(n13799) );
  AND2_X1 U15826 ( .A1(n13799), .A2(n13798), .ZN(n13945) );
  NAND2_X1 U15827 ( .A1(n13946), .A2(n14512), .ZN(n13801) );
  NAND2_X1 U15828 ( .A1(n14521), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n13800) );
  OAI211_X1 U15829 ( .C1(n14508), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        n13803) );
  AOI21_X1 U15830 ( .B1(n13945), .B2(n14517), .A(n13803), .ZN(n13804) );
  OAI211_X1 U15831 ( .C1(n13948), .C2(n13895), .A(n13805), .B(n13804), .ZN(
        P1_U3271) );
  NAND3_X1 U15832 ( .A1(n13806), .A2(n13808), .A3(n13807), .ZN(n13809) );
  AND3_X1 U15833 ( .A1(n13810), .A2(n14585), .A3(n13809), .ZN(n13812) );
  NOR2_X1 U15834 ( .A1(n13812), .A2(n13811), .ZN(n13952) );
  INV_X1 U15835 ( .A(n6607), .ZN(n13813) );
  AOI211_X1 U15836 ( .C1(n13950), .C2(n13830), .A(n13884), .B(n13813), .ZN(
        n13949) );
  INV_X1 U15837 ( .A(n13950), .ZN(n13817) );
  INV_X1 U15838 ( .A(n13814), .ZN(n13815) );
  AOI22_X1 U15839 ( .A1(n14521), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13815), 
        .B2(n14528), .ZN(n13816) );
  OAI21_X1 U15840 ( .B1(n13817), .B2(n14376), .A(n13816), .ZN(n13823) );
  INV_X1 U15841 ( .A(n13818), .ZN(n13819) );
  AOI21_X1 U15842 ( .B1(n13821), .B2(n13820), .A(n13819), .ZN(n13953) );
  NOR2_X1 U15843 ( .A1(n13953), .A2(n13895), .ZN(n13822) );
  AOI211_X1 U15844 ( .C1(n13949), .C2(n14517), .A(n13823), .B(n13822), .ZN(
        n13824) );
  OAI21_X1 U15845 ( .B1(n14521), .B2(n13952), .A(n13824), .ZN(P1_U3272) );
  NAND2_X1 U15846 ( .A1(n6665), .A2(n13825), .ZN(n13954) );
  NAND3_X1 U15847 ( .A1(n13954), .A2(n14532), .A3(n13806), .ZN(n13838) );
  INV_X1 U15848 ( .A(n13955), .ZN(n13827) );
  AOI22_X1 U15849 ( .A1(n13827), .A2(n14536), .B1(n13826), .B2(n14528), .ZN(
        n13828) );
  OAI21_X1 U15850 ( .B1(n13829), .B2(n14536), .A(n13828), .ZN(n13833) );
  OAI211_X1 U15851 ( .C1(n13849), .C2(n13831), .A(n14513), .B(n13830), .ZN(
        n13956) );
  NOR2_X1 U15852 ( .A1(n13956), .A2(n13888), .ZN(n13832) );
  AOI211_X1 U15853 ( .C1(n14512), .C2(n14018), .A(n13833), .B(n13832), .ZN(
        n13837) );
  NAND2_X1 U15854 ( .A1(n13835), .A2(n13834), .ZN(n13957) );
  NAND3_X1 U15855 ( .A1(n13958), .A2(n13957), .A3(n14533), .ZN(n13836) );
  NAND3_X1 U15856 ( .A1(n13838), .A2(n13837), .A3(n13836), .ZN(P1_U3273) );
  XNOR2_X1 U15857 ( .A(n13839), .B(n13840), .ZN(n13964) );
  INV_X1 U15858 ( .A(n13964), .ZN(n13858) );
  NAND2_X1 U15859 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  NAND2_X1 U15860 ( .A1(n13843), .A2(n13842), .ZN(n13846) );
  INV_X1 U15861 ( .A(n13844), .ZN(n13845) );
  AOI21_X1 U15862 ( .B1(n13846), .B2(n14585), .A(n13845), .ZN(n13967) );
  INV_X1 U15863 ( .A(n13967), .ZN(n13856) );
  NAND2_X1 U15864 ( .A1(n14022), .A2(n6558), .ZN(n13847) );
  NAND2_X1 U15865 ( .A1(n13847), .A2(n14513), .ZN(n13848) );
  OR2_X1 U15866 ( .A1(n13849), .A2(n13848), .ZN(n13965) );
  INV_X1 U15867 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n13852) );
  INV_X1 U15868 ( .A(n13850), .ZN(n13851) );
  OAI22_X1 U15869 ( .A1(n14536), .A2(n13852), .B1(n13851), .B2(n14508), .ZN(
        n13853) );
  AOI21_X1 U15870 ( .B1(n14022), .B2(n14512), .A(n13853), .ZN(n13854) );
  OAI21_X1 U15871 ( .B1(n13965), .B2(n13888), .A(n13854), .ZN(n13855) );
  AOI21_X1 U15872 ( .B1(n13856), .B2(n14536), .A(n13855), .ZN(n13857) );
  OAI21_X1 U15873 ( .B1(n13858), .B2(n13895), .A(n13857), .ZN(P1_U3274) );
  XNOR2_X1 U15874 ( .A(n13859), .B(n13862), .ZN(n13972) );
  INV_X1 U15875 ( .A(n13972), .ZN(n13878) );
  OAI211_X1 U15876 ( .C1(n13862), .C2(n13861), .A(n13860), .B(n14585), .ZN(
        n13868) );
  INV_X1 U15877 ( .A(n13863), .ZN(n13867) );
  NAND2_X1 U15878 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  NAND3_X1 U15879 ( .A1(n13868), .A2(n13867), .A3(n13866), .ZN(n13869) );
  AOI21_X1 U15880 ( .B1(n13972), .B2(n14557), .A(n13869), .ZN(n13974) );
  OAI21_X1 U15881 ( .B1(n13870), .B2(n14508), .A(n13974), .ZN(n13871) );
  NAND2_X1 U15882 ( .A1(n13871), .A2(n14536), .ZN(n13876) );
  AOI21_X1 U15883 ( .B1(n13873), .B2(n13886), .A(n13884), .ZN(n13872) );
  AND2_X1 U15884 ( .A1(n13872), .A2(n6558), .ZN(n13971) );
  INV_X1 U15885 ( .A(n13873), .ZN(n14029) );
  OAI22_X1 U15886 ( .A1(n14029), .A2(n14376), .B1(n14485), .B2(n14536), .ZN(
        n13874) );
  AOI21_X1 U15887 ( .B1(n14517), .B2(n13971), .A(n13874), .ZN(n13875) );
  OAI211_X1 U15888 ( .C1(n13878), .C2(n13877), .A(n13876), .B(n13875), .ZN(
        P1_U3275) );
  XNOR2_X1 U15889 ( .A(n13879), .B(n13891), .ZN(n13977) );
  INV_X1 U15890 ( .A(n13977), .ZN(n13896) );
  INV_X1 U15891 ( .A(n13880), .ZN(n13978) );
  AOI22_X1 U15892 ( .A1(n13978), .A2(n14536), .B1(n13881), .B2(n14528), .ZN(
        n13882) );
  OAI21_X1 U15893 ( .B1(n13883), .B2(n14536), .A(n13882), .ZN(n13890) );
  AOI21_X1 U15894 ( .B1(n13979), .B2(n13885), .A(n13884), .ZN(n13887) );
  NAND2_X1 U15895 ( .A1(n13887), .A2(n13886), .ZN(n13982) );
  NOR2_X1 U15896 ( .A1(n13982), .A2(n13888), .ZN(n13889) );
  AOI211_X1 U15897 ( .C1(n14512), .C2(n13979), .A(n13890), .B(n13889), .ZN(
        n13894) );
  NAND2_X1 U15898 ( .A1(n13892), .A2(n13891), .ZN(n13980) );
  NAND3_X1 U15899 ( .A1(n13981), .A2(n13980), .A3(n14532), .ZN(n13893) );
  OAI211_X1 U15900 ( .C1(n13896), .C2(n13895), .A(n13894), .B(n13893), .ZN(
        P1_U3276) );
  INV_X1 U15901 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n13899) );
  NOR2_X1 U15902 ( .A1(n13898), .A2(n13897), .ZN(n13992) );
  MUX2_X1 U15903 ( .A(n13899), .B(n13992), .S(n14600), .Z(n13900) );
  OAI21_X1 U15904 ( .B1(n13994), .B2(n13976), .A(n13900), .ZN(P1_U3559) );
  NAND2_X1 U15905 ( .A1(n13902), .A2(n13901), .ZN(n13995) );
  MUX2_X1 U15906 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n13995), .S(n14600), .Z(
        n13903) );
  AOI21_X1 U15907 ( .B1(n13969), .B2(n13997), .A(n13903), .ZN(n13904) );
  INV_X1 U15908 ( .A(n13904), .ZN(P1_U3558) );
  NAND2_X1 U15909 ( .A1(n13905), .A2(n14549), .ZN(n13908) );
  NAND4_X1 U15910 ( .A1(n13909), .A2(n13908), .A3(n13907), .A4(n13906), .ZN(
        n13910) );
  OAI21_X1 U15911 ( .B1(n13913), .B2(n13991), .A(n13912), .ZN(n13999) );
  MUX2_X1 U15912 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n13999), .S(n14597), .Z(
        P1_U3557) );
  AOI21_X1 U15913 ( .B1(n13915), .B2(n14549), .A(n13914), .ZN(n13916) );
  OAI211_X1 U15914 ( .C1(n13918), .C2(n14553), .A(n13917), .B(n13916), .ZN(
        n14000) );
  MUX2_X1 U15915 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14000), .S(n14600), .Z(
        P1_U3555) );
  INV_X1 U15916 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n13922) );
  AOI211_X1 U15917 ( .C1(n14590), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        n14001) );
  MUX2_X1 U15918 ( .A(n13922), .B(n14001), .S(n14597), .Z(n13923) );
  OAI21_X1 U15919 ( .B1(n14004), .B2(n13976), .A(n13923), .ZN(P1_U3554) );
  AND2_X1 U15920 ( .A1(n13925), .A2(n13924), .ZN(n13927) );
  OAI211_X1 U15921 ( .C1(n13928), .C2(n13991), .A(n13927), .B(n13926), .ZN(
        n14005) );
  MUX2_X1 U15922 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14005), .S(n14600), .Z(
        n13929) );
  AOI21_X1 U15923 ( .B1(n13969), .B2(n14007), .A(n13929), .ZN(n13930) );
  INV_X1 U15924 ( .A(n13930), .ZN(P1_U3553) );
  NAND2_X1 U15925 ( .A1(n13931), .A2(n14590), .ZN(n13933) );
  NAND3_X1 U15926 ( .A1(n13934), .A2(n13933), .A3(n13932), .ZN(n14009) );
  MUX2_X1 U15927 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14009), .S(n14600), .Z(
        n13935) );
  AOI21_X1 U15928 ( .B1(n13969), .B2(n14011), .A(n13935), .ZN(n13936) );
  INV_X1 U15929 ( .A(n13936), .ZN(P1_U3552) );
  AOI211_X1 U15930 ( .C1(n13939), .C2(n14549), .A(n13938), .B(n13937), .ZN(
        n13942) );
  NAND2_X1 U15931 ( .A1(n13940), .A2(n14585), .ZN(n13941) );
  OAI211_X1 U15932 ( .C1(n13943), .C2(n13991), .A(n13942), .B(n13941), .ZN(
        n14013) );
  MUX2_X1 U15933 ( .A(n14013), .B(P1_REG1_REG_23__SCAN_IN), .S(n14598), .Z(
        P1_U3551) );
  AOI211_X1 U15934 ( .C1(n13946), .C2(n14549), .A(n13945), .B(n13944), .ZN(
        n13947) );
  OAI21_X1 U15935 ( .B1(n13991), .B2(n13948), .A(n13947), .ZN(n14014) );
  MUX2_X1 U15936 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14014), .S(n14600), .Z(
        P1_U3550) );
  AOI21_X1 U15937 ( .B1(n13950), .B2(n14549), .A(n13949), .ZN(n13951) );
  OAI211_X1 U15938 ( .C1(n13953), .C2(n13991), .A(n13952), .B(n13951), .ZN(
        n14015) );
  MUX2_X1 U15939 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14015), .S(n14600), .Z(
        P1_U3549) );
  NAND3_X1 U15940 ( .A1(n13954), .A2(n14585), .A3(n13806), .ZN(n13961) );
  AND2_X1 U15941 ( .A1(n13956), .A2(n13955), .ZN(n13960) );
  NAND3_X1 U15942 ( .A1(n13958), .A2(n13957), .A3(n14590), .ZN(n13959) );
  NAND3_X1 U15943 ( .A1(n13961), .A2(n13960), .A3(n13959), .ZN(n14016) );
  MUX2_X1 U15944 ( .A(n14016), .B(P1_REG1_REG_20__SCAN_IN), .S(n14598), .Z(
        n13962) );
  AOI21_X1 U15945 ( .B1(n13969), .B2(n14018), .A(n13962), .ZN(n13963) );
  INV_X1 U15946 ( .A(n13963), .ZN(P1_U3548) );
  NAND2_X1 U15947 ( .A1(n13964), .A2(n14590), .ZN(n13966) );
  NAND3_X1 U15948 ( .A1(n13967), .A2(n13966), .A3(n13965), .ZN(n14020) );
  MUX2_X1 U15949 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14020), .S(n14597), .Z(
        n13968) );
  AOI21_X1 U15950 ( .B1(n13969), .B2(n14022), .A(n13968), .ZN(n13970) );
  INV_X1 U15951 ( .A(n13970), .ZN(P1_U3547) );
  AOI21_X1 U15952 ( .B1(n13972), .B2(n14576), .A(n13971), .ZN(n13973) );
  AND2_X1 U15953 ( .A1(n13974), .A2(n13973), .ZN(n14025) );
  MUX2_X1 U15954 ( .A(n14479), .B(n14025), .S(n14597), .Z(n13975) );
  OAI21_X1 U15955 ( .B1(n14029), .B2(n13976), .A(n13975), .ZN(P1_U3546) );
  NAND2_X1 U15956 ( .A1(n13977), .A2(n14590), .ZN(n13985) );
  AOI21_X1 U15957 ( .B1(n13979), .B2(n14549), .A(n13978), .ZN(n13984) );
  NAND3_X1 U15958 ( .A1(n13981), .A2(n14585), .A3(n13980), .ZN(n13983) );
  NAND4_X1 U15959 ( .A1(n13985), .A2(n13984), .A3(n13983), .A4(n13982), .ZN(
        n14030) );
  MUX2_X1 U15960 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14030), .S(n14597), .Z(
        P1_U3545) );
  AOI211_X1 U15961 ( .C1(n13988), .C2(n14549), .A(n13987), .B(n13986), .ZN(
        n13989) );
  OAI21_X1 U15962 ( .B1(n13991), .B2(n13990), .A(n13989), .ZN(n14031) );
  MUX2_X1 U15963 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14031), .S(n14597), .Z(
        P1_U3544) );
  INV_X1 U15964 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n13993) );
  MUX2_X1 U15965 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n13995), .S(n8150), .Z(
        n13996) );
  AOI21_X1 U15966 ( .B1(n14023), .B2(n13997), .A(n13996), .ZN(n13998) );
  INV_X1 U15967 ( .A(n13998), .ZN(P1_U3526) );
  MUX2_X1 U15968 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n13999), .S(n8150), .Z(
        P1_U3525) );
  MUX2_X1 U15969 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14000), .S(n8150), .Z(
        P1_U3523) );
  INV_X1 U15970 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14002) );
  MUX2_X1 U15971 ( .A(n14002), .B(n14001), .S(n8150), .Z(n14003) );
  OAI21_X1 U15972 ( .B1(n14004), .B2(n14028), .A(n14003), .ZN(P1_U3522) );
  MUX2_X1 U15973 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14005), .S(n8150), .Z(
        n14006) );
  AOI21_X1 U15974 ( .B1(n14023), .B2(n14007), .A(n14006), .ZN(n14008) );
  INV_X1 U15975 ( .A(n14008), .ZN(P1_U3521) );
  MUX2_X1 U15976 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14009), .S(n8150), .Z(
        n14010) );
  AOI21_X1 U15977 ( .B1(n14023), .B2(n14011), .A(n14010), .ZN(n14012) );
  INV_X1 U15978 ( .A(n14012), .ZN(P1_U3520) );
  MUX2_X1 U15979 ( .A(n14013), .B(P1_REG0_REG_23__SCAN_IN), .S(n14577), .Z(
        P1_U3519) );
  MUX2_X1 U15980 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14014), .S(n8150), .Z(
        P1_U3518) );
  MUX2_X1 U15981 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14015), .S(n8150), .Z(
        P1_U3517) );
  MUX2_X1 U15982 ( .A(n14016), .B(P1_REG0_REG_20__SCAN_IN), .S(n14577), .Z(
        n14017) );
  AOI21_X1 U15983 ( .B1(n14023), .B2(n14018), .A(n14017), .ZN(n14019) );
  INV_X1 U15984 ( .A(n14019), .ZN(P1_U3516) );
  MUX2_X1 U15985 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14020), .S(n8150), .Z(
        n14021) );
  AOI21_X1 U15986 ( .B1(n14023), .B2(n14022), .A(n14021), .ZN(n14024) );
  INV_X1 U15987 ( .A(n14024), .ZN(P1_U3515) );
  INV_X1 U15988 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14026) );
  MUX2_X1 U15989 ( .A(n14026), .B(n14025), .S(n8150), .Z(n14027) );
  OAI21_X1 U15990 ( .B1(n14029), .B2(n14028), .A(n14027), .ZN(P1_U3513) );
  MUX2_X1 U15991 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14030), .S(n8150), .Z(
        P1_U3510) );
  MUX2_X1 U15992 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14031), .S(n8150), .Z(
        P1_U3507) );
  NOR4_X1 U15993 ( .A1(n14032), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14033), .A4(
        P1_U3086), .ZN(n14034) );
  AOI21_X1 U15994 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14035), .A(n14034), 
        .ZN(n14036) );
  OAI21_X1 U15995 ( .B1(n14037), .B2(n14043), .A(n14036), .ZN(P1_U3324) );
  OAI222_X1 U15996 ( .A1(n14040), .A2(P1_U3086), .B1(n14043), .B2(n14039), 
        .C1(n14038), .C2(n14047), .ZN(P1_U3326) );
  OAI222_X1 U15997 ( .A1(n14047), .A2(n15299), .B1(n14043), .B2(n14042), .C1(
        P1_U3086), .C2(n14041), .ZN(P1_U3328) );
  OAI222_X1 U15998 ( .A1(n14047), .A2(n14046), .B1(n14043), .B2(n14045), .C1(
        n14044), .C2(P1_U3086), .ZN(P1_U3329) );
  OAI222_X1 U15999 ( .A1(n14047), .A2(n15366), .B1(n14043), .B2(n14049), .C1(
        P1_U3086), .C2(n14048), .ZN(P1_U3330) );
  MUX2_X1 U16000 ( .A(n13297), .B(n14050), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16001 ( .A(n14051), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16002 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14723) );
  INV_X1 U16003 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14428) );
  XOR2_X1 U16004 ( .A(n14898), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14139) );
  INV_X1 U16005 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14879) );
  INV_X1 U16006 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14075) );
  INV_X1 U16007 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14072) );
  XOR2_X1 U16008 ( .A(n14072), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14130) );
  INV_X1 U16009 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15211) );
  NAND2_X1 U16010 ( .A1(n14100), .A2(n14099), .ZN(n14052) );
  XOR2_X1 U16011 ( .A(n14053), .B(P3_ADDR_REG_2__SCAN_IN), .Z(n14098) );
  NOR2_X1 U16012 ( .A1(n14054), .A2(n15220), .ZN(n14056) );
  NOR2_X1 U16013 ( .A1(n14060), .A2(n14059), .ZN(n14062) );
  XNOR2_X1 U16014 ( .A(n14060), .B(n14059), .ZN(n14110) );
  NOR2_X1 U16015 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14116), .ZN(n14064) );
  INV_X1 U16016 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14063) );
  NOR2_X1 U16017 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14065), .ZN(n14067) );
  XNOR2_X1 U16018 ( .A(n14065), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14121) );
  NOR2_X1 U16019 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n14068), .ZN(n14070) );
  NAND2_X1 U16020 ( .A1(n14130), .A2(n14129), .ZN(n14071) );
  XNOR2_X1 U16021 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14073), .ZN(n14093) );
  XNOR2_X1 U16022 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n14076), .ZN(n14135) );
  NAND2_X1 U16023 ( .A1(n14139), .A2(n14138), .ZN(n14078) );
  INV_X1 U16024 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U16025 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14915), .ZN(n14079) );
  INV_X1 U16026 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14441) );
  NAND2_X1 U16027 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n14441), .ZN(n14080) );
  INV_X1 U16028 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14937) );
  INV_X1 U16029 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15350) );
  OR2_X1 U16030 ( .A1(n15350), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U16031 ( .A1(n14141), .A2(n14081), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n15350), .ZN(n14082) );
  NOR2_X1 U16032 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14082), .ZN(n14084) );
  INV_X1 U16033 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14210) );
  INV_X1 U16034 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14464) );
  XOR2_X1 U16035 ( .A(n14464), .B(n14082), .Z(n14144) );
  NOR2_X1 U16036 ( .A1(n14210), .A2(n14144), .ZN(n14083) );
  NOR2_X1 U16037 ( .A1(n14084), .A2(n14083), .ZN(n14085) );
  NOR2_X1 U16038 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14085), .ZN(n14087) );
  INV_X1 U16039 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14228) );
  INV_X1 U16040 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15318) );
  XOR2_X1 U16041 ( .A(n15318), .B(n14085), .Z(n14147) );
  NOR2_X1 U16042 ( .A1(n14228), .A2(n14147), .ZN(n14086) );
  NOR2_X1 U16043 ( .A1(n14087), .A2(n14086), .ZN(n14181) );
  INV_X1 U16044 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14500) );
  XNOR2_X1 U16045 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n14500), .ZN(n14180) );
  XNOR2_X1 U16046 ( .A(n14181), .B(n14180), .ZN(n14178) );
  INV_X1 U16047 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14679) );
  XNOR2_X1 U16048 ( .A(n14937), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14088) );
  XNOR2_X1 U16049 ( .A(n14089), .B(n14088), .ZN(n14408) );
  XOR2_X1 U16050 ( .A(n14915), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14091) );
  XNOR2_X1 U16051 ( .A(n14091), .B(n14090), .ZN(n14403) );
  XOR2_X1 U16052 ( .A(n14093), .B(n14092), .Z(n14134) );
  INV_X1 U16053 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14132) );
  XOR2_X1 U16054 ( .A(n15151), .B(n14094), .Z(n14128) );
  INV_X1 U16055 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14625) );
  OR2_X1 U16056 ( .A1(n14625), .A2(n14096), .ZN(n14109) );
  XOR2_X1 U16057 ( .A(n14096), .B(n14625), .Z(n15389) );
  INV_X1 U16058 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14105) );
  XNOR2_X1 U16059 ( .A(n14097), .B(n14098), .ZN(n14151) );
  XNOR2_X1 U16060 ( .A(n14100), .B(n14099), .ZN(n14101) );
  NAND2_X1 U16061 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14101), .ZN(n14103) );
  AOI21_X1 U16062 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14850), .A(n14100), .ZN(
        n15392) );
  INV_X1 U16063 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15391) );
  NOR2_X1 U16064 ( .A1(n15392), .A2(n15391), .ZN(n15401) );
  XOR2_X1 U16065 ( .A(n14101), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15400) );
  NAND2_X1 U16066 ( .A1(n15401), .A2(n15400), .ZN(n14102) );
  NAND2_X1 U16067 ( .A1(n14103), .A2(n14102), .ZN(n14152) );
  NAND2_X1 U16068 ( .A1(n14151), .A2(n14152), .ZN(n14104) );
  NOR2_X1 U16069 ( .A1(n14151), .A2(n14152), .ZN(n14150) );
  AOI21_X1 U16070 ( .B1(n14105), .B2(n14104), .A(n14150), .ZN(n15396) );
  XOR2_X1 U16071 ( .A(n14107), .B(n14106), .Z(n15397) );
  NOR2_X1 U16072 ( .A1(n15396), .A2(n15397), .ZN(n14108) );
  NAND2_X1 U16073 ( .A1(n15396), .A2(n15397), .ZN(n15395) );
  OAI21_X1 U16074 ( .B1(n14108), .B2(n15398), .A(n15395), .ZN(n15388) );
  XOR2_X1 U16075 ( .A(n15321), .B(n14110), .Z(n14111) );
  NOR2_X1 U16076 ( .A1(n14112), .A2(n14111), .ZN(n14114) );
  XNOR2_X1 U16077 ( .A(n14112), .B(n14111), .ZN(n15390) );
  NOR2_X1 U16078 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15390), .ZN(n14113) );
  NAND2_X1 U16079 ( .A1(n14115), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14120) );
  INV_X1 U16080 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14638) );
  XOR2_X1 U16081 ( .A(n14116), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14118) );
  XOR2_X1 U16082 ( .A(n14118), .B(n14117), .Z(n14159) );
  NAND2_X1 U16083 ( .A1(n14160), .A2(n14159), .ZN(n14119) );
  NAND2_X1 U16084 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14123), .ZN(n14126) );
  XOR2_X1 U16085 ( .A(n14122), .B(n14121), .Z(n15394) );
  XNOR2_X1 U16086 ( .A(n14130), .B(n14129), .ZN(n14167) );
  NAND2_X1 U16087 ( .A1(n14168), .A2(n14167), .ZN(n14131) );
  NOR2_X1 U16088 ( .A1(n14168), .A2(n14167), .ZN(n14166) );
  NOR2_X1 U16089 ( .A1(n14134), .A2(n14133), .ZN(n14171) );
  XOR2_X1 U16090 ( .A(n14136), .B(n14135), .Z(n14394) );
  NAND2_X1 U16091 ( .A1(n14395), .A2(n14394), .ZN(n14393) );
  XNOR2_X1 U16092 ( .A(n14139), .B(n14138), .ZN(n14399) );
  INV_X1 U16093 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U16094 ( .A1(n14400), .A2(n14399), .ZN(n14398) );
  INV_X1 U16095 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14668) );
  NAND2_X1 U16096 ( .A1(n14408), .A2(n14407), .ZN(n14140) );
  XOR2_X1 U16097 ( .A(n15350), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14142) );
  XNOR2_X1 U16098 ( .A(n14142), .B(n14141), .ZN(n14411) );
  NAND2_X1 U16099 ( .A1(n14412), .A2(n14411), .ZN(n14143) );
  XNOR2_X1 U16100 ( .A(n14210), .B(n14144), .ZN(n14146) );
  NOR2_X1 U16101 ( .A1(n14145), .A2(n14146), .ZN(n14415) );
  XOR2_X1 U16102 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14147), .Z(n14175) );
  INV_X1 U16103 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14706) );
  XNOR2_X1 U16104 ( .A(n14178), .B(n14177), .ZN(n14179) );
  XOR2_X1 U16105 ( .A(n14723), .B(n14179), .Z(SUB_1596_U62) );
  AOI21_X1 U16106 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14148) );
  OAI21_X1 U16107 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14148), 
        .ZN(U28) );
  AOI21_X1 U16108 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14149) );
  OAI21_X1 U16109 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14149), 
        .ZN(U29) );
  AOI21_X1 U16110 ( .B1(n14152), .B2(n14151), .A(n14150), .ZN(n14153) );
  XOR2_X1 U16111 ( .A(n14153), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  OR2_X1 U16112 ( .A1(n14155), .A2(n14154), .ZN(n14157) );
  NAND2_X1 U16113 ( .A1(n14161), .A2(SI_13_), .ZN(n14156) );
  AND2_X1 U16114 ( .A1(n14157), .A2(n14156), .ZN(n14158) );
  OAI21_X1 U16115 ( .B1(P3_U3151), .B2(n14916), .A(n14158), .ZN(P3_U3282) );
  XOR2_X1 U16116 ( .A(n14160), .B(n14159), .Z(SUB_1596_U57) );
  AOI22_X1 U16117 ( .A1(n14163), .A2(n14162), .B1(SI_16_), .B2(n14161), .ZN(
        n14164) );
  OAI21_X1 U16118 ( .B1(P3_U3151), .B2(n14211), .A(n14164), .ZN(P3_U3279) );
  XNOR2_X1 U16119 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14165), .ZN(SUB_1596_U55)
         );
  AOI21_X1 U16120 ( .B1(n14168), .B2(n14167), .A(n14166), .ZN(n14169) );
  XOR2_X1 U16121 ( .A(n14169), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  NOR2_X1 U16122 ( .A1(n14171), .A2(n14170), .ZN(n14172) );
  XOR2_X1 U16123 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14172), .Z(SUB_1596_U70)
         );
  OAI21_X1 U16124 ( .B1(n14175), .B2(n14174), .A(n14173), .ZN(n14176) );
  XOR2_X1 U16125 ( .A(n14176), .B(n14706), .Z(SUB_1596_U63) );
  NOR2_X1 U16126 ( .A1(n14181), .A2(n14180), .ZN(n14182) );
  AOI21_X1 U16127 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14500), .A(n14182), 
        .ZN(n14183) );
  XOR2_X1 U16128 ( .A(n14183), .B(P3_ADDR_REG_19__SCAN_IN), .Z(n14184) );
  AOI22_X1 U16129 ( .A1(n14866), .A2(n14185), .B1(n14860), .B2(
        P3_ADDR_REG_15__SCAN_IN), .ZN(n14199) );
  OAI21_X1 U16130 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14187), .A(n14186), 
        .ZN(n14191) );
  XNOR2_X1 U16131 ( .A(n14189), .B(n14188), .ZN(n14190) );
  AOI22_X1 U16132 ( .A1(n14191), .A2(n14929), .B1(n14893), .B2(n14190), .ZN(
        n14198) );
  NAND2_X1 U16133 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P3_U3151), .ZN(n14197)
         );
  OAI221_X1 U16134 ( .B1(n14195), .B2(n14194), .C1(n14195), .C2(n14193), .A(
        n14192), .ZN(n14196) );
  NAND4_X1 U16135 ( .A1(n14199), .A2(n14198), .A3(n14197), .A4(n14196), .ZN(
        P3_U3197) );
  AOI21_X1 U16136 ( .B1(n6649), .B2(n14201), .A(n14200), .ZN(n14217) );
  OAI21_X1 U16137 ( .B1(n14204), .B2(n14203), .A(n14202), .ZN(n14205) );
  AND2_X1 U16138 ( .A1(n14205), .A2(n14929), .ZN(n14214) );
  OAI211_X1 U16139 ( .C1(n14208), .C2(n14207), .A(n14206), .B(n14893), .ZN(
        n14209) );
  INV_X1 U16140 ( .A(n14209), .ZN(n14213) );
  OAI22_X1 U16141 ( .A1(n14939), .A2(n14211), .B1(n14210), .B2(n14936), .ZN(
        n14212) );
  NOR4_X1 U16142 ( .A1(n14215), .A2(n14214), .A3(n14213), .A4(n14212), .ZN(
        n14216) );
  OAI21_X1 U16143 ( .B1(n14217), .B2(n14945), .A(n14216), .ZN(P3_U3198) );
  AOI21_X1 U16144 ( .B1(n14220), .B2(n14219), .A(n14218), .ZN(n14235) );
  OAI21_X1 U16145 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14222), .A(n14221), 
        .ZN(n14223) );
  AND2_X1 U16146 ( .A1(n14929), .A2(n14223), .ZN(n14232) );
  OAI21_X1 U16147 ( .B1(n14225), .B2(n14224), .A(n14893), .ZN(n14227) );
  NOR2_X1 U16148 ( .A1(n14227), .A2(n14226), .ZN(n14231) );
  OAI22_X1 U16149 ( .A1(n14939), .A2(n14229), .B1(n14228), .B2(n14936), .ZN(
        n14230) );
  NOR4_X1 U16150 ( .A1(n14233), .A2(n14232), .A3(n14231), .A4(n14230), .ZN(
        n14234) );
  OAI21_X1 U16151 ( .B1(n14235), .B2(n14945), .A(n14234), .ZN(P3_U3199) );
  AOI21_X1 U16152 ( .B1(n14238), .B2(n14237), .A(n14236), .ZN(n14252) );
  NOR2_X1 U16153 ( .A1(n14939), .A2(n14239), .ZN(n14240) );
  AOI211_X1 U16154 ( .C1(n14860), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n14241), 
        .B(n14240), .ZN(n14251) );
  OAI21_X1 U16155 ( .B1(n14244), .B2(n14243), .A(n14242), .ZN(n14249) );
  OAI21_X1 U16156 ( .B1(n14247), .B2(n14246), .A(n14245), .ZN(n14248) );
  AOI22_X1 U16157 ( .A1(n14249), .A2(n14929), .B1(n14893), .B2(n14248), .ZN(
        n14250) );
  OAI211_X1 U16158 ( .C1(n14252), .C2(n14945), .A(n14251), .B(n14250), .ZN(
        P3_U3200) );
  AOI22_X1 U16159 ( .A1(n14285), .A2(n14253), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15018), .ZN(n14254) );
  NAND2_X1 U16160 ( .A1(n14255), .A2(n14254), .ZN(P3_U3203) );
  XNOR2_X1 U16161 ( .A(n14256), .B(n14264), .ZN(n14257) );
  NAND2_X1 U16162 ( .A1(n14257), .A2(n14982), .ZN(n14261) );
  AOI22_X1 U16163 ( .A1(n14980), .A2(n14259), .B1(n14258), .B2(n14977), .ZN(
        n14260) );
  NAND2_X1 U16164 ( .A1(n14261), .A2(n14260), .ZN(n14291) );
  OAI22_X1 U16165 ( .A1(n14263), .A2(n14995), .B1(n15010), .B2(n14262), .ZN(
        n14271) );
  INV_X1 U16166 ( .A(n14264), .ZN(n14265) );
  XNOR2_X1 U16167 ( .A(n14266), .B(n14265), .ZN(n14289) );
  OR2_X1 U16168 ( .A1(n14267), .A2(n14988), .ZN(n14287) );
  OAI22_X1 U16169 ( .A1(n14289), .A2(n14269), .B1(n14287), .B2(n14268), .ZN(
        n14270) );
  AOI211_X1 U16170 ( .C1(n14995), .C2(n14291), .A(n14271), .B(n14270), .ZN(
        n14272) );
  INV_X1 U16171 ( .A(n14272), .ZN(P3_U3221) );
  INV_X1 U16172 ( .A(n14995), .ZN(n15018) );
  XOR2_X1 U16173 ( .A(n14273), .B(n14278), .Z(n14276) );
  AOI222_X1 U16174 ( .A1(n14982), .A2(n14276), .B1(n14275), .B2(n14980), .C1(
        n14274), .C2(n14977), .ZN(n14292) );
  AOI22_X1 U16175 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n15018), .B1(n14991), 
        .B2(n14277), .ZN(n14283) );
  XNOR2_X1 U16176 ( .A(n14279), .B(n14278), .ZN(n14295) );
  NOR2_X1 U16177 ( .A1(n14280), .A2(n14988), .ZN(n14294) );
  AOI22_X1 U16178 ( .A1(n14295), .A2(n14281), .B1(n14294), .B2(n14992), .ZN(
        n14282) );
  OAI211_X1 U16179 ( .C1(n15018), .C2(n14292), .A(n14283), .B(n14282), .ZN(
        P3_U3222) );
  AOI21_X1 U16180 ( .B1(n14285), .B2(n15043), .A(n14284), .ZN(n14297) );
  INV_X1 U16181 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U16182 ( .A1(n15072), .A2(n14297), .B1(n14286), .B2(n8777), .ZN(
        P3_U3489) );
  OAI21_X1 U16183 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n14290) );
  NOR2_X1 U16184 ( .A1(n14291), .A2(n14290), .ZN(n14298) );
  AOI22_X1 U16185 ( .A1(n15072), .A2(n14298), .B1(n15274), .B2(n8777), .ZN(
        P3_U3471) );
  INV_X1 U16186 ( .A(n14292), .ZN(n14293) );
  AOI211_X1 U16187 ( .C1(n15054), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        n14299) );
  INV_X1 U16188 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U16189 ( .A1(n15072), .A2(n14299), .B1(n14296), .B2(n8777), .ZN(
        P3_U3470) );
  AOI22_X1 U16190 ( .A1(n15056), .A2(n8695), .B1(n14297), .B2(n15055), .ZN(
        P3_U3457) );
  AOI22_X1 U16191 ( .A1(n15056), .A2(n8429), .B1(n14298), .B2(n15055), .ZN(
        P3_U3426) );
  AOI22_X1 U16192 ( .A1(n15056), .A2(n8407), .B1(n14299), .B2(n15055), .ZN(
        P3_U3423) );
  NAND2_X1 U16193 ( .A1(n14301), .A2(n14300), .ZN(n14303) );
  AOI21_X1 U16194 ( .B1(n14304), .B2(n14303), .A(n14302), .ZN(n14312) );
  AOI22_X1 U16195 ( .A1(n14308), .A2(n14307), .B1(n14306), .B2(n14305), .ZN(
        n14309) );
  OAI21_X1 U16196 ( .B1(n14333), .B2(n14310), .A(n14309), .ZN(n14311) );
  NOR2_X1 U16197 ( .A1(n14312), .A2(n14311), .ZN(n14314) );
  OAI211_X1 U16198 ( .C1(n14331), .C2(n14315), .A(n14314), .B(n14313), .ZN(
        P2_U3187) );
  INV_X1 U16199 ( .A(n14316), .ZN(n14320) );
  INV_X1 U16200 ( .A(n14317), .ZN(n14319) );
  AOI21_X1 U16201 ( .B1(n14320), .B2(n14319), .A(n14318), .ZN(n14323) );
  OAI21_X1 U16202 ( .B1(n14323), .B2(n14322), .A(n14321), .ZN(n14324) );
  AOI222_X1 U16203 ( .A1(n14328), .A2(n14327), .B1(n14326), .B2(n14325), .C1(
        n14324), .C2(n9282), .ZN(n14329) );
  NAND2_X1 U16204 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14690)
         );
  OAI211_X1 U16205 ( .C1(n14331), .C2(n14330), .A(n14329), .B(n14690), .ZN(
        P2_U3198) );
  OAI21_X1 U16206 ( .B1(n14333), .B2(n14797), .A(n14332), .ZN(n14336) );
  INV_X1 U16207 ( .A(n14334), .ZN(n14335) );
  AOI211_X1 U16208 ( .C1(n14337), .C2(n14787), .A(n14336), .B(n14335), .ZN(
        n14345) );
  AOI22_X1 U16209 ( .A1(n14842), .A2(n14345), .B1(n10923), .B2(n14840), .ZN(
        P2_U3513) );
  AND2_X1 U16210 ( .A1(n14338), .A2(n14787), .ZN(n14342) );
  OAI21_X1 U16211 ( .B1(n14340), .B2(n14797), .A(n14339), .ZN(n14341) );
  NOR3_X1 U16212 ( .A1(n14343), .A2(n14342), .A3(n14341), .ZN(n14347) );
  AOI22_X1 U16213 ( .A1(n14842), .A2(n14347), .B1(n10919), .B2(n14840), .ZN(
        P2_U3512) );
  INV_X1 U16214 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14344) );
  AOI22_X1 U16215 ( .A1(n14829), .A2(n14345), .B1(n14344), .B2(n14827), .ZN(
        P2_U3472) );
  INV_X1 U16216 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U16217 ( .A1(n14829), .A2(n14347), .B1(n14346), .B2(n14827), .ZN(
        P2_U3469) );
  AOI21_X1 U16218 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n14351) );
  OR2_X1 U16219 ( .A1(n6697), .A2(n14351), .ZN(n14352) );
  AOI222_X1 U16220 ( .A1(n9693), .A2(n14370), .B1(n14354), .B2(n14353), .C1(
        n14352), .C2(n14365), .ZN(n14355) );
  NAND2_X1 U16221 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14439)
         );
  OAI211_X1 U16222 ( .C1(n14369), .C2(n14372), .A(n14355), .B(n14439), .ZN(
        P1_U3215) );
  AND2_X1 U16223 ( .A1(n13288), .A2(n14356), .ZN(n14359) );
  OAI21_X1 U16224 ( .B1(n14359), .B2(n14358), .A(n14357), .ZN(n14366) );
  OAI22_X1 U16225 ( .A1(n14363), .A2(n14362), .B1(n14361), .B2(n14360), .ZN(
        n14364) );
  AOI21_X1 U16226 ( .B1(n14366), .B2(n14365), .A(n14364), .ZN(n14367) );
  NAND2_X1 U16227 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14462)
         );
  OAI211_X1 U16228 ( .C1(n14369), .C2(n14368), .A(n14367), .B(n14462), .ZN(
        P1_U3226) );
  INV_X1 U16229 ( .A(n14370), .ZN(n14377) );
  NAND2_X1 U16230 ( .A1(n14371), .A2(n14517), .ZN(n14375) );
  INV_X1 U16231 ( .A(n14372), .ZN(n14373) );
  AOI22_X1 U16232 ( .A1(n14521), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n14373), 
        .B2(n14528), .ZN(n14374) );
  OAI211_X1 U16233 ( .C1(n14377), .C2(n14376), .A(n14375), .B(n14374), .ZN(
        n14378) );
  AOI21_X1 U16234 ( .B1(n14379), .B2(n14533), .A(n14378), .ZN(n14380) );
  OAI21_X1 U16235 ( .B1(n14521), .B2(n14381), .A(n14380), .ZN(P1_U3279) );
  NAND3_X1 U16236 ( .A1(n14383), .A2(n14382), .A3(n14585), .ZN(n14388) );
  NAND2_X1 U16237 ( .A1(n14384), .A2(n14549), .ZN(n14385) );
  NAND4_X1 U16238 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14389) );
  AOI21_X1 U16239 ( .B1(n14390), .B2(n14590), .A(n14389), .ZN(n14392) );
  AOI22_X1 U16240 ( .A1(n14600), .A2(n14392), .B1(n14443), .B2(n14598), .ZN(
        P1_U3543) );
  INV_X1 U16241 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U16242 ( .A1(n8150), .A2(n14392), .B1(n14391), .B2(n14577), .ZN(
        P1_U3504) );
  OAI21_X1 U16243 ( .B1(n14395), .B2(n14394), .A(n14393), .ZN(n14397) );
  XOR2_X1 U16244 ( .A(n14397), .B(n14396), .Z(SUB_1596_U69) );
  OAI21_X1 U16245 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n14401) );
  XOR2_X1 U16246 ( .A(n14401), .B(n14654), .Z(SUB_1596_U68) );
  OAI21_X1 U16247 ( .B1(n14404), .B2(n14403), .A(n14402), .ZN(n14405) );
  XOR2_X1 U16248 ( .A(n14405), .B(n14668), .Z(SUB_1596_U67) );
  AOI21_X1 U16249 ( .B1(n14408), .B2(n14407), .A(n14406), .ZN(n14409) );
  XOR2_X1 U16250 ( .A(n14409), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16251 ( .B1(n14412), .B2(n14411), .A(n14410), .ZN(n14413) );
  XOR2_X1 U16252 ( .A(n14413), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  INV_X1 U16253 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14692) );
  NOR2_X1 U16254 ( .A1(n14415), .A2(n14414), .ZN(n14416) );
  XNOR2_X1 U16255 ( .A(n14692), .B(n14416), .ZN(SUB_1596_U64) );
  AOI211_X1 U16256 ( .C1(n14419), .C2(n14418), .A(n14417), .B(n14452), .ZN(
        n14424) );
  AOI211_X1 U16257 ( .C1(n14422), .C2(n14421), .A(n14420), .B(n14488), .ZN(
        n14423) );
  AOI211_X1 U16258 ( .C1(n14493), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        n14427) );
  OAI211_X1 U16259 ( .C1(n14428), .C2(n14499), .A(n14427), .B(n14426), .ZN(
        P1_U3256) );
  OAI21_X1 U16260 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14438) );
  NOR2_X1 U16261 ( .A1(n14432), .A2(n14475), .ZN(n14437) );
  AOI211_X1 U16262 ( .C1(n14435), .C2(n14434), .A(n14488), .B(n14433), .ZN(
        n14436) );
  AOI211_X1 U16263 ( .C1(n14483), .C2(n14438), .A(n14437), .B(n14436), .ZN(
        n14440) );
  OAI211_X1 U16264 ( .C1(n14441), .C2(n14499), .A(n14440), .B(n14439), .ZN(
        P1_U3257) );
  OAI21_X1 U16265 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14449) );
  OAI21_X1 U16266 ( .B1(n14447), .B2(n7840), .A(n14446), .ZN(n14448) );
  AOI222_X1 U16267 ( .A1(n14449), .A2(n14483), .B1(n6747), .B2(n14493), .C1(
        n14448), .C2(n14468), .ZN(n14451) );
  OAI211_X1 U16268 ( .C1(n15350), .C2(n14499), .A(n14451), .B(n14450), .ZN(
        P1_U3258) );
  AOI211_X1 U16269 ( .C1(n14455), .C2(n14454), .A(n14453), .B(n14452), .ZN(
        n14460) );
  AOI211_X1 U16270 ( .C1(n14458), .C2(n14457), .A(n14456), .B(n14488), .ZN(
        n14459) );
  AOI211_X1 U16271 ( .C1(n14493), .C2(n14461), .A(n14460), .B(n14459), .ZN(
        n14463) );
  OAI211_X1 U16272 ( .C1(n14464), .C2(n14499), .A(n14463), .B(n14462), .ZN(
        P1_U3259) );
  OAI211_X1 U16273 ( .C1(n14467), .C2(n14466), .A(n14465), .B(n14483), .ZN(
        n14473) );
  OAI211_X1 U16274 ( .C1(n14471), .C2(n14470), .A(n14469), .B(n14468), .ZN(
        n14472) );
  OAI211_X1 U16275 ( .C1(n14475), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        n14476) );
  INV_X1 U16276 ( .A(n14476), .ZN(n14478) );
  OAI211_X1 U16277 ( .C1(n15318), .C2(n14499), .A(n14478), .B(n14477), .ZN(
        P1_U3260) );
  NAND2_X1 U16278 ( .A1(n14480), .A2(n14479), .ZN(n14484) );
  INV_X1 U16279 ( .A(n14481), .ZN(n14482) );
  NAND3_X1 U16280 ( .A1(n14484), .A2(n14483), .A3(n14482), .ZN(n14496) );
  NAND2_X1 U16281 ( .A1(n14486), .A2(n14485), .ZN(n14490) );
  NOR2_X1 U16282 ( .A1(n14488), .A2(n14487), .ZN(n14489) );
  NAND2_X1 U16283 ( .A1(n14490), .A2(n14489), .ZN(n14495) );
  INV_X1 U16284 ( .A(n14491), .ZN(n14492) );
  NAND2_X1 U16285 ( .A1(n14493), .A2(n14492), .ZN(n14494) );
  OAI211_X1 U16286 ( .C1(n14500), .C2(n14499), .A(n14498), .B(n14497), .ZN(
        P1_U3261) );
  XNOR2_X1 U16287 ( .A(n14501), .B(n14502), .ZN(n14563) );
  XNOR2_X1 U16288 ( .A(n14503), .B(n14502), .ZN(n14506) );
  OAI21_X1 U16289 ( .B1(n14506), .B2(n14505), .A(n14504), .ZN(n14507) );
  AOI21_X1 U16290 ( .B1(n14557), .B2(n14563), .A(n14507), .ZN(n14560) );
  OAI22_X1 U16291 ( .A1(n14536), .A2(n14509), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14508), .ZN(n14510) );
  AOI21_X1 U16292 ( .B1(n14512), .B2(n14511), .A(n14510), .ZN(n14520) );
  OAI211_X1 U16293 ( .C1(n14515), .C2(n14559), .A(n14514), .B(n14513), .ZN(
        n14558) );
  INV_X1 U16294 ( .A(n14558), .ZN(n14516) );
  AOI22_X1 U16295 ( .A1(n14518), .A2(n14563), .B1(n14517), .B2(n14516), .ZN(
        n14519) );
  OAI211_X1 U16296 ( .C1(n14521), .C2(n14560), .A(n14520), .B(n14519), .ZN(
        P1_U3290) );
  AOI21_X1 U16297 ( .B1(n14524), .B2(n14523), .A(n14522), .ZN(n14527) );
  OAI21_X1 U16298 ( .B1(n14527), .B2(n14526), .A(n14525), .ZN(n14529) );
  AOI22_X1 U16299 ( .A1(n14536), .A2(n14529), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n14528), .ZN(n14535) );
  INV_X1 U16300 ( .A(n14530), .ZN(n14531) );
  OAI21_X1 U16301 ( .B1(n14533), .B2(n14532), .A(n14531), .ZN(n14534) );
  OAI211_X1 U16302 ( .C1(n14536), .C2(n7574), .A(n14535), .B(n14534), .ZN(
        P1_U3293) );
  AND2_X1 U16303 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14537), .ZN(P1_U3294) );
  AND2_X1 U16304 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14537), .ZN(P1_U3295) );
  AND2_X1 U16305 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14537), .ZN(P1_U3296) );
  AND2_X1 U16306 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14537), .ZN(P1_U3297) );
  AND2_X1 U16307 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14537), .ZN(P1_U3298) );
  AND2_X1 U16308 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14537), .ZN(P1_U3299) );
  AND2_X1 U16309 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14537), .ZN(P1_U3300) );
  NOR2_X1 U16310 ( .A1(n14538), .A2(n15363), .ZN(P1_U3301) );
  AND2_X1 U16311 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14537), .ZN(P1_U3302) );
  AND2_X1 U16312 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14537), .ZN(P1_U3303) );
  AND2_X1 U16313 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14537), .ZN(P1_U3304) );
  AND2_X1 U16314 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14537), .ZN(P1_U3305) );
  AND2_X1 U16315 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14537), .ZN(P1_U3306) );
  AND2_X1 U16316 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14537), .ZN(P1_U3307) );
  AND2_X1 U16317 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14537), .ZN(P1_U3308) );
  NOR2_X1 U16318 ( .A1(n14538), .A2(n15360), .ZN(P1_U3309) );
  NOR2_X1 U16319 ( .A1(n14538), .A2(n15259), .ZN(P1_U3310) );
  NOR2_X1 U16320 ( .A1(n14538), .A2(n15300), .ZN(P1_U3311) );
  AND2_X1 U16321 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14537), .ZN(P1_U3312) );
  AND2_X1 U16322 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14537), .ZN(P1_U3313) );
  AND2_X1 U16323 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14537), .ZN(P1_U3314) );
  AND2_X1 U16324 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14537), .ZN(P1_U3315) );
  INV_X1 U16325 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15286) );
  NOR2_X1 U16326 ( .A1(n14538), .A2(n15286), .ZN(P1_U3316) );
  INV_X1 U16327 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15137) );
  NOR2_X1 U16328 ( .A1(n14538), .A2(n15137), .ZN(P1_U3317) );
  AND2_X1 U16329 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14537), .ZN(P1_U3318) );
  AND2_X1 U16330 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14537), .ZN(P1_U3319) );
  AND2_X1 U16331 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14537), .ZN(P1_U3320) );
  INV_X1 U16332 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15141) );
  NOR2_X1 U16333 ( .A1(n14538), .A2(n15141), .ZN(P1_U3321) );
  AND2_X1 U16334 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14537), .ZN(P1_U3322) );
  INV_X1 U16335 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15205) );
  NOR2_X1 U16336 ( .A1(n14538), .A2(n15205), .ZN(P1_U3323) );
  INV_X1 U16337 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U16338 ( .A1(n8150), .A2(n14540), .B1(n14539), .B2(n14577), .ZN(
        P1_U3459) );
  INV_X1 U16339 ( .A(n14541), .ZN(n14542) );
  OAI21_X1 U16340 ( .B1(n14543), .B2(n14582), .A(n14542), .ZN(n14546) );
  INV_X1 U16341 ( .A(n14544), .ZN(n14545) );
  AOI211_X1 U16342 ( .C1(n14576), .C2(n14547), .A(n14546), .B(n14545), .ZN(
        n14592) );
  AOI22_X1 U16343 ( .A1(n8150), .A2(n14592), .B1(n7585), .B2(n14577), .ZN(
        P1_U3462) );
  AOI21_X1 U16344 ( .B1(n14550), .B2(n14549), .A(n14548), .ZN(n14551) );
  OAI211_X1 U16345 ( .C1(n14554), .C2(n14553), .A(n14552), .B(n14551), .ZN(
        n14555) );
  AOI21_X1 U16346 ( .B1(n14557), .B2(n14556), .A(n14555), .ZN(n14593) );
  AOI22_X1 U16347 ( .A1(n8150), .A2(n14593), .B1(n7599), .B2(n14577), .ZN(
        P1_U3465) );
  OAI21_X1 U16348 ( .B1(n14559), .B2(n14582), .A(n14558), .ZN(n14562) );
  INV_X1 U16349 ( .A(n14560), .ZN(n14561) );
  AOI211_X1 U16350 ( .C1(n14576), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14594) );
  AOI22_X1 U16351 ( .A1(n8150), .A2(n14594), .B1(n7614), .B2(n14577), .ZN(
        P1_U3468) );
  OAI21_X1 U16352 ( .B1(n14565), .B2(n14582), .A(n14564), .ZN(n14567) );
  AOI211_X1 U16353 ( .C1(n14568), .C2(n14590), .A(n14567), .B(n14566), .ZN(
        n14595) );
  INV_X1 U16354 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14569) );
  AOI22_X1 U16355 ( .A1(n8150), .A2(n14595), .B1(n14569), .B2(n14577), .ZN(
        P1_U3471) );
  INV_X1 U16356 ( .A(n14570), .ZN(n14575) );
  OAI21_X1 U16357 ( .B1(n6874), .B2(n14582), .A(n14572), .ZN(n14574) );
  AOI211_X1 U16358 ( .C1(n14576), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14596) );
  INV_X1 U16359 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U16360 ( .A1(n8150), .A2(n14596), .B1(n15239), .B2(n14577), .ZN(
        P1_U3474) );
  INV_X1 U16361 ( .A(n14578), .ZN(n14583) );
  INV_X1 U16362 ( .A(n14579), .ZN(n14580) );
  OAI211_X1 U16363 ( .C1(n14583), .C2(n14582), .A(n14581), .B(n14580), .ZN(
        n14588) );
  AND3_X1 U16364 ( .A1(n14586), .A2(n14585), .A3(n14584), .ZN(n14587) );
  AOI211_X1 U16365 ( .C1(n14590), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14599) );
  INV_X1 U16366 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U16367 ( .A1(n8150), .A2(n14599), .B1(n14591), .B2(n14577), .ZN(
        P1_U3483) );
  AOI22_X1 U16368 ( .A1(n14597), .A2(n14592), .B1(n7586), .B2(n14598), .ZN(
        P1_U3529) );
  AOI22_X1 U16369 ( .A1(n14597), .A2(n14593), .B1(n7598), .B2(n14598), .ZN(
        P1_U3530) );
  AOI22_X1 U16370 ( .A1(n14597), .A2(n14594), .B1(n9606), .B2(n14598), .ZN(
        P1_U3531) );
  AOI22_X1 U16371 ( .A1(n14600), .A2(n14595), .B1(n7635), .B2(n14598), .ZN(
        P1_U3532) );
  AOI22_X1 U16372 ( .A1(n14597), .A2(n14596), .B1(n9608), .B2(n14598), .ZN(
        P1_U3533) );
  AOI22_X1 U16373 ( .A1(n14600), .A2(n14599), .B1(n9667), .B2(n14598), .ZN(
        P1_U3536) );
  NOR2_X1 U16374 ( .A1(n14601), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16375 ( .A1(n14601), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14612) );
  OAI211_X1 U16376 ( .C1(n14604), .C2(n14603), .A(n14715), .B(n14602), .ZN(
        n14609) );
  OAI211_X1 U16377 ( .C1(n14607), .C2(n14606), .A(n14655), .B(n14605), .ZN(
        n14608) );
  OAI211_X1 U16378 ( .C1(n14621), .C2(n8859), .A(n14609), .B(n14608), .ZN(
        n14610) );
  INV_X1 U16379 ( .A(n14610), .ZN(n14611) );
  NAND2_X1 U16380 ( .A1(n14612), .A2(n14611), .ZN(P2_U3215) );
  OAI211_X1 U16381 ( .C1(n14614), .C2(n14613), .A(n14715), .B(n6908), .ZN(
        n14619) );
  OAI211_X1 U16382 ( .C1(n14617), .C2(n14616), .A(n14655), .B(n14615), .ZN(
        n14618) );
  OAI211_X1 U16383 ( .C1(n14621), .C2(n14620), .A(n14619), .B(n14618), .ZN(
        n14622) );
  INV_X1 U16384 ( .A(n14622), .ZN(n14624) );
  OAI211_X1 U16385 ( .C1(n14722), .C2(n14625), .A(n14624), .B(n14623), .ZN(
        P2_U3218) );
  OAI211_X1 U16386 ( .C1(n14628), .C2(n14627), .A(n14655), .B(n14626), .ZN(
        n14629) );
  INV_X1 U16387 ( .A(n14629), .ZN(n14634) );
  AOI211_X1 U16388 ( .C1(n14632), .C2(n14631), .A(n14695), .B(n14630), .ZN(
        n14633) );
  AOI211_X1 U16389 ( .C1(n14719), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14637) );
  OAI211_X1 U16390 ( .C1(n14722), .C2(n14638), .A(n14637), .B(n14636), .ZN(
        P2_U3220) );
  INV_X1 U16391 ( .A(n14639), .ZN(n14641) );
  OAI21_X1 U16392 ( .B1(n14641), .B2(n14640), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14642) );
  OAI21_X1 U16393 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_12__SCAN_IN), 
        .A(n14642), .ZN(n14653) );
  OAI21_X1 U16394 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n14651) );
  NAND2_X1 U16395 ( .A1(n14647), .A2(n14646), .ZN(n14648) );
  AOI21_X1 U16396 ( .B1(n14649), .B2(n14648), .A(n14707), .ZN(n14650) );
  AOI21_X1 U16397 ( .B1(n14651), .B2(n14715), .A(n14650), .ZN(n14652) );
  OAI211_X1 U16398 ( .C1(n14654), .C2(n14722), .A(n14653), .B(n14652), .ZN(
        P2_U3226) );
  OAI211_X1 U16399 ( .C1(n14658), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14659) );
  INV_X1 U16400 ( .A(n14659), .ZN(n14664) );
  AOI211_X1 U16401 ( .C1(n14662), .C2(n14661), .A(n14695), .B(n14660), .ZN(
        n14663) );
  AOI211_X1 U16402 ( .C1(n14719), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14667) );
  NAND2_X1 U16403 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14666)
         );
  OAI211_X1 U16404 ( .C1(n14668), .C2(n14722), .A(n14667), .B(n14666), .ZN(
        P2_U3227) );
  AOI211_X1 U16405 ( .C1(n14670), .C2(n9102), .A(n14669), .B(n14695), .ZN(
        n14675) );
  AOI211_X1 U16406 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14707), .ZN(
        n14674) );
  AOI211_X1 U16407 ( .C1(n14719), .C2(n14676), .A(n14675), .B(n14674), .ZN(
        n14678) );
  NAND2_X1 U16408 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14677)
         );
  OAI211_X1 U16409 ( .C1(n14679), .C2(n14722), .A(n14678), .B(n14677), .ZN(
        P2_U3229) );
  AOI211_X1 U16410 ( .C1(n14682), .C2(n14681), .A(n14707), .B(n14680), .ZN(
        n14688) );
  INV_X1 U16411 ( .A(n14683), .ZN(n14684) );
  AOI211_X1 U16412 ( .C1(n14686), .C2(n14685), .A(n14695), .B(n14684), .ZN(
        n14687) );
  AOI211_X1 U16413 ( .C1(n14719), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        n14691) );
  OAI211_X1 U16414 ( .C1(n14692), .C2(n14722), .A(n14691), .B(n14690), .ZN(
        P2_U3230) );
  INV_X1 U16415 ( .A(n14693), .ZN(n14697) );
  AOI211_X1 U16416 ( .C1(n14697), .C2(n14696), .A(n14695), .B(n14694), .ZN(
        n14702) );
  AOI211_X1 U16417 ( .C1(n14700), .C2(n14699), .A(n14707), .B(n14698), .ZN(
        n14701) );
  AOI211_X1 U16418 ( .C1(n14719), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14705) );
  OAI211_X1 U16419 ( .C1(n14706), .C2(n14722), .A(n14705), .B(n14704), .ZN(
        P2_U3231) );
  AOI211_X1 U16420 ( .C1(n14710), .C2(n14709), .A(n14708), .B(n14707), .ZN(
        n14717) );
  OAI21_X1 U16421 ( .B1(n14713), .B2(n14712), .A(n14711), .ZN(n14714) );
  AND2_X1 U16422 ( .A1(n14715), .A2(n14714), .ZN(n14716) );
  AOI211_X1 U16423 ( .C1(n14719), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14721) );
  OAI211_X1 U16424 ( .C1(n14723), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        P2_U3232) );
  INV_X1 U16425 ( .A(n14751), .ZN(n14753) );
  INV_X1 U16426 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15196) );
  NOR2_X1 U16427 ( .A1(n14749), .A2(n15196), .ZN(P2_U3266) );
  INV_X1 U16428 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15164) );
  NOR2_X1 U16429 ( .A1(n14749), .A2(n15164), .ZN(P2_U3267) );
  INV_X1 U16430 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14725) );
  NOR2_X1 U16431 ( .A1(n14749), .A2(n14725), .ZN(P2_U3268) );
  INV_X1 U16432 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14726) );
  NOR2_X1 U16433 ( .A1(n14746), .A2(n14726), .ZN(P2_U3269) );
  INV_X1 U16434 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14727) );
  NOR2_X1 U16435 ( .A1(n14746), .A2(n14727), .ZN(P2_U3270) );
  INV_X1 U16436 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14728) );
  NOR2_X1 U16437 ( .A1(n14746), .A2(n14728), .ZN(P2_U3271) );
  INV_X1 U16438 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14729) );
  NOR2_X1 U16439 ( .A1(n14746), .A2(n14729), .ZN(P2_U3272) );
  INV_X1 U16440 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14730) );
  NOR2_X1 U16441 ( .A1(n14746), .A2(n14730), .ZN(P2_U3273) );
  INV_X1 U16442 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15194) );
  NOR2_X1 U16443 ( .A1(n14746), .A2(n15194), .ZN(P2_U3274) );
  INV_X1 U16444 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14731) );
  NOR2_X1 U16445 ( .A1(n14746), .A2(n14731), .ZN(P2_U3275) );
  INV_X1 U16446 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14732) );
  NOR2_X1 U16447 ( .A1(n14746), .A2(n14732), .ZN(P2_U3276) );
  INV_X1 U16448 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14733) );
  NOR2_X1 U16449 ( .A1(n14746), .A2(n14733), .ZN(P2_U3277) );
  INV_X1 U16450 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15266) );
  NOR2_X1 U16451 ( .A1(n14749), .A2(n15266), .ZN(P2_U3278) );
  INV_X1 U16452 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14734) );
  NOR2_X1 U16453 ( .A1(n14749), .A2(n14734), .ZN(P2_U3279) );
  INV_X1 U16454 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U16455 ( .A1(n14749), .A2(n15333), .ZN(P2_U3280) );
  INV_X1 U16456 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14735) );
  NOR2_X1 U16457 ( .A1(n14749), .A2(n14735), .ZN(P2_U3281) );
  INV_X1 U16458 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15306) );
  NOR2_X1 U16459 ( .A1(n14749), .A2(n15306), .ZN(P2_U3282) );
  INV_X1 U16460 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U16461 ( .A1(n14749), .A2(n14736), .ZN(P2_U3283) );
  INV_X1 U16462 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14737) );
  NOR2_X1 U16463 ( .A1(n14749), .A2(n14737), .ZN(P2_U3284) );
  INV_X1 U16464 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14738) );
  NOR2_X1 U16465 ( .A1(n14749), .A2(n14738), .ZN(P2_U3285) );
  INV_X1 U16466 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14739) );
  NOR2_X1 U16467 ( .A1(n14749), .A2(n14739), .ZN(P2_U3286) );
  INV_X1 U16468 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14740) );
  NOR2_X1 U16469 ( .A1(n14749), .A2(n14740), .ZN(P2_U3287) );
  INV_X1 U16470 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15325) );
  NOR2_X1 U16471 ( .A1(n14749), .A2(n15325), .ZN(P2_U3288) );
  INV_X1 U16472 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14741) );
  NOR2_X1 U16473 ( .A1(n14749), .A2(n14741), .ZN(P2_U3289) );
  INV_X1 U16474 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14742) );
  NOR2_X1 U16475 ( .A1(n14749), .A2(n14742), .ZN(P2_U3290) );
  INV_X1 U16476 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14743) );
  NOR2_X1 U16477 ( .A1(n14746), .A2(n14743), .ZN(P2_U3291) );
  INV_X1 U16478 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14744) );
  NOR2_X1 U16479 ( .A1(n14749), .A2(n14744), .ZN(P2_U3292) );
  INV_X1 U16480 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14745) );
  NOR2_X1 U16481 ( .A1(n14746), .A2(n14745), .ZN(P2_U3293) );
  INV_X1 U16482 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14747) );
  NOR2_X1 U16483 ( .A1(n14749), .A2(n14747), .ZN(P2_U3294) );
  INV_X1 U16484 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14748) );
  NOR2_X1 U16485 ( .A1(n14749), .A2(n14748), .ZN(P2_U3295) );
  AOI22_X1 U16486 ( .A1(n14751), .A2(n14750), .B1(n15260), .B2(n14753), .ZN(
        P2_U3416) );
  AOI21_X1 U16487 ( .B1(n15273), .B2(n14753), .A(n14752), .ZN(P2_U3417) );
  INV_X1 U16488 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U16489 ( .A1(n14829), .A2(n14755), .B1(n14754), .B2(n14827), .ZN(
        P2_U3430) );
  OAI21_X1 U16490 ( .B1(n14757), .B2(n14797), .A(n14756), .ZN(n14759) );
  AOI211_X1 U16491 ( .C1(n14802), .C2(n14760), .A(n14759), .B(n14758), .ZN(
        n14830) );
  INV_X1 U16492 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14761) );
  AOI22_X1 U16493 ( .A1(n14829), .A2(n14830), .B1(n14761), .B2(n14827), .ZN(
        P2_U3436) );
  OAI21_X1 U16494 ( .B1(n14763), .B2(n14797), .A(n14762), .ZN(n14766) );
  INV_X1 U16495 ( .A(n14764), .ZN(n14765) );
  AOI211_X1 U16496 ( .C1(n14787), .C2(n14767), .A(n14766), .B(n14765), .ZN(
        n14831) );
  INV_X1 U16497 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U16498 ( .A1(n14829), .A2(n14831), .B1(n15319), .B2(n14827), .ZN(
        P2_U3439) );
  OAI21_X1 U16499 ( .B1(n14769), .B2(n14797), .A(n14768), .ZN(n14772) );
  INV_X1 U16500 ( .A(n14770), .ZN(n14771) );
  AOI211_X1 U16501 ( .C1(n14787), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14832) );
  AOI22_X1 U16502 ( .A1(n14829), .A2(n14832), .B1(n8918), .B2(n14827), .ZN(
        P2_U3442) );
  OAI211_X1 U16503 ( .C1(n14776), .C2(n14797), .A(n14775), .B(n14774), .ZN(
        n14779) );
  AOI21_X1 U16504 ( .B1(n9731), .B2(n14822), .A(n14777), .ZN(n14778) );
  NOR2_X1 U16505 ( .A1(n14779), .A2(n14778), .ZN(n14834) );
  AOI22_X1 U16506 ( .A1(n14829), .A2(n14834), .B1(n8933), .B2(n14827), .ZN(
        P2_U3445) );
  AOI21_X1 U16507 ( .B1(n9731), .B2(n14822), .A(n14780), .ZN(n14785) );
  NOR2_X1 U16508 ( .A1(n14781), .A2(n14797), .ZN(n14782) );
  NOR4_X1 U16509 ( .A1(n14785), .A2(n14784), .A3(n14783), .A4(n14782), .ZN(
        n14835) );
  INV_X1 U16510 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U16511 ( .A1(n14829), .A2(n14835), .B1(n14786), .B2(n14827), .ZN(
        P2_U3448) );
  AND2_X1 U16512 ( .A1(n14788), .A2(n14787), .ZN(n14793) );
  OAI21_X1 U16513 ( .B1(n14790), .B2(n14797), .A(n14789), .ZN(n14791) );
  NOR3_X1 U16514 ( .A1(n14793), .A2(n14792), .A3(n14791), .ZN(n14836) );
  INV_X1 U16515 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14794) );
  AOI22_X1 U16516 ( .A1(n14829), .A2(n14836), .B1(n14794), .B2(n14827), .ZN(
        P2_U3451) );
  INV_X1 U16517 ( .A(n14795), .ZN(n14801) );
  OAI21_X1 U16518 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14800) );
  AOI211_X1 U16519 ( .C1(n14802), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        n14837) );
  AOI22_X1 U16520 ( .A1(n14829), .A2(n14837), .B1(n8985), .B2(n14827), .ZN(
        P2_U3454) );
  NAND2_X1 U16521 ( .A1(n14803), .A2(n14818), .ZN(n14805) );
  OAI211_X1 U16522 ( .C1(n14806), .C2(n14822), .A(n14805), .B(n14804), .ZN(
        n14809) );
  NOR2_X1 U16523 ( .A1(n14806), .A2(n9731), .ZN(n14808) );
  NOR3_X1 U16524 ( .A1(n14809), .A2(n14808), .A3(n14807), .ZN(n14838) );
  INV_X1 U16525 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U16526 ( .A1(n14829), .A2(n14838), .B1(n14810), .B2(n14827), .ZN(
        P2_U3457) );
  NAND2_X1 U16527 ( .A1(n14811), .A2(n14818), .ZN(n14813) );
  OAI211_X1 U16528 ( .C1(n14814), .C2(n14822), .A(n14813), .B(n14812), .ZN(
        n14817) );
  NOR2_X1 U16529 ( .A1(n14814), .A2(n9731), .ZN(n14816) );
  NOR3_X1 U16530 ( .A1(n14817), .A2(n14816), .A3(n14815), .ZN(n14839) );
  AOI22_X1 U16531 ( .A1(n14829), .A2(n14839), .B1(n9020), .B2(n14827), .ZN(
        P2_U3460) );
  NAND2_X1 U16532 ( .A1(n14819), .A2(n14818), .ZN(n14821) );
  OAI211_X1 U16533 ( .C1(n14823), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        n14826) );
  NOR2_X1 U16534 ( .A1(n14823), .A2(n9731), .ZN(n14825) );
  NOR3_X1 U16535 ( .A1(n14826), .A2(n14825), .A3(n14824), .ZN(n14841) );
  INV_X1 U16536 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14828) );
  AOI22_X1 U16537 ( .A1(n14829), .A2(n14841), .B1(n14828), .B2(n14827), .ZN(
        P2_U3463) );
  AOI22_X1 U16538 ( .A1(n14842), .A2(n14830), .B1(n8887), .B2(n14840), .ZN(
        P2_U3501) );
  AOI22_X1 U16539 ( .A1(n14842), .A2(n14831), .B1(n8903), .B2(n14840), .ZN(
        P2_U3502) );
  AOI22_X1 U16540 ( .A1(n14842), .A2(n14832), .B1(n9578), .B2(n14840), .ZN(
        P2_U3503) );
  AOI22_X1 U16541 ( .A1(n14842), .A2(n14834), .B1(n14833), .B2(n14840), .ZN(
        P2_U3504) );
  AOI22_X1 U16542 ( .A1(n14842), .A2(n14835), .B1(n8950), .B2(n14840), .ZN(
        P2_U3505) );
  AOI22_X1 U16543 ( .A1(n14842), .A2(n14836), .B1(n8968), .B2(n14840), .ZN(
        P2_U3506) );
  AOI22_X1 U16544 ( .A1(n14842), .A2(n14837), .B1(n8989), .B2(n14840), .ZN(
        P2_U3507) );
  AOI22_X1 U16545 ( .A1(n14842), .A2(n14838), .B1(n9936), .B2(n14840), .ZN(
        P2_U3508) );
  AOI22_X1 U16546 ( .A1(n14842), .A2(n14839), .B1(n9935), .B2(n14840), .ZN(
        P2_U3509) );
  AOI22_X1 U16547 ( .A1(n14842), .A2(n14841), .B1(n9039), .B2(n14840), .ZN(
        P2_U3510) );
  NOR2_X1 U16548 ( .A1(P3_U3897), .A2(n14860), .ZN(P3_U3150) );
  AOI22_X1 U16549 ( .A1(n14866), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n14849) );
  NOR2_X1 U16550 ( .A1(n14843), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14846) );
  NAND3_X1 U16551 ( .A1(n14945), .A2(n14844), .A3(n14933), .ZN(n14845) );
  OAI21_X1 U16552 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(n14848) );
  OAI211_X1 U16553 ( .C1(n14850), .C2(n14936), .A(n14849), .B(n14848), .ZN(
        P3_U3182) );
  AOI21_X1 U16554 ( .B1(n14853), .B2(n14852), .A(n14851), .ZN(n14869) );
  OAI21_X1 U16555 ( .B1(n14856), .B2(n14855), .A(n14854), .ZN(n14857) );
  AND2_X1 U16556 ( .A1(n14857), .A2(n14929), .ZN(n14858) );
  AOI211_X1 U16557 ( .C1(P3_ADDR_REG_10__SCAN_IN), .C2(n14860), .A(n14859), 
        .B(n14858), .ZN(n14868) );
  OAI21_X1 U16558 ( .B1(n14863), .B2(n14862), .A(n14861), .ZN(n14864) );
  AOI22_X1 U16559 ( .A1(n14866), .A2(n14865), .B1(n14893), .B2(n14864), .ZN(
        n14867) );
  OAI211_X1 U16560 ( .C1(n14869), .C2(n14945), .A(n14868), .B(n14867), .ZN(
        P3_U3192) );
  AOI21_X1 U16561 ( .B1(n14872), .B2(n14871), .A(n14870), .ZN(n14886) );
  OAI21_X1 U16562 ( .B1(n14874), .B2(P3_REG1_REG_11__SCAN_IN), .A(n14873), 
        .ZN(n14875) );
  AND2_X1 U16563 ( .A1(n14875), .A2(n14929), .ZN(n14883) );
  XOR2_X1 U16564 ( .A(n14877), .B(n14876), .Z(n14878) );
  NOR2_X1 U16565 ( .A1(n14878), .A2(n14933), .ZN(n14882) );
  OAI22_X1 U16566 ( .A1(n14939), .A2(n14880), .B1(n14879), .B2(n14936), .ZN(
        n14881) );
  NOR4_X1 U16567 ( .A1(n14884), .A2(n14883), .A3(n14882), .A4(n14881), .ZN(
        n14885) );
  OAI21_X1 U16568 ( .B1(n14886), .B2(n14945), .A(n14885), .ZN(P3_U3193) );
  AOI21_X1 U16569 ( .B1(n6722), .B2(n14888), .A(n14887), .ZN(n14905) );
  OAI21_X1 U16570 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14892) );
  AND2_X1 U16571 ( .A1(n14892), .A2(n14929), .ZN(n14902) );
  OAI211_X1 U16572 ( .C1(n14896), .C2(n14895), .A(n14894), .B(n14893), .ZN(
        n14897) );
  INV_X1 U16573 ( .A(n14897), .ZN(n14901) );
  OAI22_X1 U16574 ( .A1(n14939), .A2(n14899), .B1(n14898), .B2(n14936), .ZN(
        n14900) );
  NOR4_X1 U16575 ( .A1(n14903), .A2(n14902), .A3(n14901), .A4(n14900), .ZN(
        n14904) );
  OAI21_X1 U16576 ( .B1(n14905), .B2(n14945), .A(n14904), .ZN(P3_U3194) );
  AOI21_X1 U16577 ( .B1(n11248), .B2(n14907), .A(n14906), .ZN(n14922) );
  OAI21_X1 U16578 ( .B1(n14909), .B2(P3_REG1_REG_13__SCAN_IN), .A(n14908), 
        .ZN(n14910) );
  AND2_X1 U16579 ( .A1(n14929), .A2(n14910), .ZN(n14919) );
  NAND2_X1 U16580 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  AOI21_X1 U16581 ( .B1(n14914), .B2(n14913), .A(n14933), .ZN(n14918) );
  OAI22_X1 U16582 ( .A1(n14939), .A2(n14916), .B1(n14915), .B2(n14936), .ZN(
        n14917) );
  NOR4_X1 U16583 ( .A1(n14920), .A2(n14919), .A3(n14918), .A4(n14917), .ZN(
        n14921) );
  OAI21_X1 U16584 ( .B1(n14922), .B2(n14945), .A(n14921), .ZN(P3_U3195) );
  AOI21_X1 U16585 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14946) );
  AND2_X1 U16586 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n14943) );
  OAI21_X1 U16587 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n14930) );
  AND2_X1 U16588 ( .A1(n14930), .A2(n14929), .ZN(n14942) );
  INV_X1 U16589 ( .A(n14931), .ZN(n14932) );
  AOI211_X1 U16590 ( .C1(n14935), .C2(n14934), .A(n14933), .B(n14932), .ZN(
        n14941) );
  OAI22_X1 U16591 ( .A1(n14939), .A2(n14938), .B1(n14937), .B2(n14936), .ZN(
        n14940) );
  NOR4_X1 U16592 ( .A1(n14943), .A2(n14942), .A3(n14941), .A4(n14940), .ZN(
        n14944) );
  OAI21_X1 U16593 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(P3_U3196) );
  XNOR2_X1 U16594 ( .A(n14947), .B(n14949), .ZN(n14954) );
  INV_X1 U16595 ( .A(n14954), .ZN(n15046) );
  OAI21_X1 U16596 ( .B1(n6719), .B2(n14949), .A(n14948), .ZN(n14950) );
  NAND2_X1 U16597 ( .A1(n14950), .A2(n14982), .ZN(n14953) );
  AOI22_X1 U16598 ( .A1(n14980), .A2(n14964), .B1(n14951), .B2(n14977), .ZN(
        n14952) );
  OAI211_X1 U16599 ( .C1(n15038), .C2(n14954), .A(n14953), .B(n14952), .ZN(
        n15044) );
  AOI21_X1 U16600 ( .B1(n15003), .B2(n15046), .A(n15044), .ZN(n14959) );
  AND2_X1 U16601 ( .A1(n14955), .A2(n15043), .ZN(n15045) );
  AOI22_X1 U16602 ( .A1(n14992), .A2(n15045), .B1(n14991), .B2(n14956), .ZN(
        n14957) );
  OAI221_X1 U16603 ( .B1(n15018), .B2(n14959), .C1(n14995), .C2(n14958), .A(
        n14957), .ZN(P3_U3225) );
  AND2_X1 U16604 ( .A1(n14960), .A2(n15043), .ZN(n15034) );
  AOI22_X1 U16605 ( .A1(n14992), .A2(n15034), .B1(n14991), .B2(n14961), .ZN(
        n14973) );
  OAI21_X1 U16606 ( .B1(n14963), .B2(n14966), .A(n14962), .ZN(n15035) );
  INV_X1 U16607 ( .A(n15035), .ZN(n14970) );
  AOI22_X1 U16608 ( .A1(n14980), .A2(n14965), .B1(n14964), .B2(n14977), .ZN(
        n14969) );
  OAI211_X1 U16609 ( .C1(n6720), .C2(n8337), .A(n14982), .B(n14967), .ZN(
        n14968) );
  OAI211_X1 U16610 ( .C1(n14970), .C2(n15038), .A(n14969), .B(n14968), .ZN(
        n15033) );
  AOI22_X1 U16611 ( .A1(n15033), .A2(n14995), .B1(n14971), .B2(n15035), .ZN(
        n14972) );
  OAI211_X1 U16612 ( .C1(n14974), .C2(n14995), .A(n14973), .B(n14972), .ZN(
        P3_U3227) );
  OAI21_X1 U16613 ( .B1(n14976), .B2(n8753), .A(n14975), .ZN(n15024) );
  INV_X1 U16614 ( .A(n15024), .ZN(n14987) );
  AOI22_X1 U16615 ( .A1(n14980), .A2(n14979), .B1(n14978), .B2(n14977), .ZN(
        n14986) );
  OAI211_X1 U16616 ( .C1(n14984), .C2(n14983), .A(n14982), .B(n14981), .ZN(
        n14985) );
  OAI211_X1 U16617 ( .C1(n14987), .C2(n15038), .A(n14986), .B(n14985), .ZN(
        n15022) );
  AOI21_X1 U16618 ( .B1(n15003), .B2(n15024), .A(n15022), .ZN(n14996) );
  NOR2_X1 U16619 ( .A1(n14989), .A2(n14988), .ZN(n15023) );
  AOI22_X1 U16620 ( .A1(n14992), .A2(n15023), .B1(n14991), .B2(n14990), .ZN(
        n14993) );
  OAI221_X1 U16621 ( .B1(n15018), .B2(n14996), .C1(n14995), .C2(n14994), .A(
        n14993), .ZN(P3_U3230) );
  INV_X1 U16622 ( .A(n14997), .ZN(n15002) );
  OAI22_X1 U16623 ( .A1(n14999), .A2(n14998), .B1(n15010), .B2(n15247), .ZN(
        n15001) );
  AOI211_X1 U16624 ( .C1(n15003), .C2(n15002), .A(n15001), .B(n15000), .ZN(
        n15004) );
  AOI22_X1 U16625 ( .A1(n15018), .A2(n15005), .B1(n15004), .B2(n14995), .ZN(
        P3_U3231) );
  INV_X1 U16626 ( .A(n15006), .ZN(n15007) );
  AOI21_X1 U16627 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15017) );
  OAI22_X1 U16628 ( .A1(n15013), .A2(n15012), .B1(n15011), .B2(n15010), .ZN(
        n15014) );
  INV_X1 U16629 ( .A(n15014), .ZN(n15015) );
  OAI221_X1 U16630 ( .B1(n15018), .B2(n15017), .C1(n14995), .C2(n15016), .A(
        n15015), .ZN(P3_U3232) );
  INV_X1 U16631 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U16632 ( .A1(n15056), .A2(n15020), .B1(n15019), .B2(n15055), .ZN(
        P3_U3393) );
  AOI22_X1 U16633 ( .A1(n15056), .A2(n8263), .B1(n15021), .B2(n15055), .ZN(
        P3_U3396) );
  AOI211_X1 U16634 ( .C1(n15049), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        n15058) );
  AOI22_X1 U16635 ( .A1(n15056), .A2(n8269), .B1(n15058), .B2(n15055), .ZN(
        P3_U3399) );
  AOI211_X1 U16636 ( .C1(n15027), .C2(n15049), .A(n15026), .B(n15025), .ZN(
        n15059) );
  AOI22_X1 U16637 ( .A1(n15056), .A2(n8283), .B1(n15059), .B2(n15055), .ZN(
        P3_U3402) );
  INV_X1 U16638 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15032) );
  INV_X1 U16639 ( .A(n15028), .ZN(n15031) );
  AOI211_X1 U16640 ( .C1(n15031), .C2(n15049), .A(n15030), .B(n15029), .ZN(
        n15061) );
  AOI22_X1 U16641 ( .A1(n15056), .A2(n15032), .B1(n15061), .B2(n15055), .ZN(
        P3_U3405) );
  AOI211_X1 U16642 ( .C1(n15049), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        n15063) );
  AOI22_X1 U16643 ( .A1(n15056), .A2(n8319), .B1(n15063), .B2(n15055), .ZN(
        P3_U3408) );
  AOI21_X1 U16644 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15041) );
  INV_X1 U16645 ( .A(n15039), .ZN(n15040) );
  AOI211_X1 U16646 ( .C1(n15043), .C2(n15042), .A(n15041), .B(n15040), .ZN(
        n15065) );
  AOI22_X1 U16647 ( .A1(n15056), .A2(n8341), .B1(n15065), .B2(n15055), .ZN(
        P3_U3411) );
  AOI211_X1 U16648 ( .C1(n15046), .C2(n15049), .A(n15045), .B(n15044), .ZN(
        n15067) );
  AOI22_X1 U16649 ( .A1(n15056), .A2(n8357), .B1(n15067), .B2(n15055), .ZN(
        P3_U3414) );
  AOI211_X1 U16650 ( .C1(n15050), .C2(n15049), .A(n15048), .B(n15047), .ZN(
        n15069) );
  AOI22_X1 U16651 ( .A1(n15056), .A2(n8371), .B1(n15069), .B2(n15055), .ZN(
        P3_U3417) );
  AOI211_X1 U16652 ( .C1(n15054), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15071) );
  AOI22_X1 U16653 ( .A1(n15056), .A2(n8389), .B1(n15071), .B2(n15055), .ZN(
        P3_U3420) );
  INV_X1 U16654 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U16655 ( .A1(n15072), .A2(n15058), .B1(n15057), .B2(n8777), .ZN(
        P3_U3462) );
  AOI22_X1 U16656 ( .A1(n15072), .A2(n15059), .B1(n10279), .B2(n8777), .ZN(
        P3_U3463) );
  INV_X1 U16657 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15060) );
  AOI22_X1 U16658 ( .A1(n15072), .A2(n15061), .B1(n15060), .B2(n8777), .ZN(
        P3_U3464) );
  AOI22_X1 U16659 ( .A1(n15072), .A2(n15063), .B1(n15062), .B2(n8777), .ZN(
        P3_U3465) );
  INV_X1 U16660 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15064) );
  AOI22_X1 U16661 ( .A1(n15072), .A2(n15065), .B1(n15064), .B2(n8777), .ZN(
        P3_U3466) );
  AOI22_X1 U16662 ( .A1(n15072), .A2(n15067), .B1(n15066), .B2(n8777), .ZN(
        P3_U3467) );
  INV_X1 U16663 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15068) );
  AOI22_X1 U16664 ( .A1(n15072), .A2(n15069), .B1(n15068), .B2(n8777), .ZN(
        P3_U3468) );
  AOI22_X1 U16665 ( .A1(n15072), .A2(n15071), .B1(n15070), .B2(n8777), .ZN(
        P3_U3469) );
  NAND2_X1 U16666 ( .A1(n15073), .A2(n15075), .ZN(n15074) );
  OAI21_X1 U16667 ( .B1(n15075), .B2(P3_D_REG_1__SCAN_IN), .A(n15074), .ZN(
        n15387) );
  INV_X1 U16668 ( .A(keyinput108), .ZN(n15076) );
  NOR4_X1 U16669 ( .A1(keyinput62), .A2(keyinput70), .A3(keyinput63), .A4(
        n15076), .ZN(n15078) );
  INV_X1 U16670 ( .A(keyinput115), .ZN(n15077) );
  NAND4_X1 U16671 ( .A1(keyinput9), .A2(keyinput13), .A3(n15078), .A4(n15077), 
        .ZN(n15089) );
  NAND4_X1 U16672 ( .A1(keyinput2), .A2(keyinput110), .A3(keyinput67), .A4(
        keyinput44), .ZN(n15088) );
  NOR3_X1 U16673 ( .A1(keyinput46), .A2(keyinput52), .A3(keyinput30), .ZN(
        n15079) );
  NAND2_X1 U16674 ( .A1(keyinput91), .A2(n15079), .ZN(n15087) );
  INV_X1 U16675 ( .A(keyinput39), .ZN(n15080) );
  NOR4_X1 U16676 ( .A1(keyinput3), .A2(keyinput82), .A3(keyinput68), .A4(
        n15080), .ZN(n15085) );
  NOR4_X1 U16677 ( .A1(keyinput96), .A2(keyinput73), .A3(keyinput11), .A4(
        keyinput43), .ZN(n15084) );
  INV_X1 U16678 ( .A(keyinput105), .ZN(n15081) );
  NOR4_X1 U16679 ( .A1(keyinput113), .A2(keyinput47), .A3(keyinput49), .A4(
        n15081), .ZN(n15083) );
  AND4_X1 U16680 ( .A1(keyinput27), .A2(keyinput94), .A3(keyinput38), .A4(
        keyinput14), .ZN(n15082) );
  NAND4_X1 U16681 ( .A1(n15085), .A2(n15084), .A3(n15083), .A4(n15082), .ZN(
        n15086) );
  NOR4_X1 U16682 ( .A1(n15089), .A2(n15088), .A3(n15087), .A4(n15086), .ZN(
        n15135) );
  NOR2_X1 U16683 ( .A1(keyinput23), .A2(keyinput104), .ZN(n15090) );
  NAND3_X1 U16684 ( .A1(keyinput121), .A2(keyinput10), .A3(n15090), .ZN(n15097) );
  NOR2_X1 U16685 ( .A1(keyinput120), .A2(keyinput71), .ZN(n15091) );
  NAND3_X1 U16686 ( .A1(keyinput119), .A2(keyinput18), .A3(n15091), .ZN(n15096) );
  NOR2_X1 U16687 ( .A1(keyinput4), .A2(keyinput78), .ZN(n15092) );
  NAND3_X1 U16688 ( .A1(keyinput29), .A2(keyinput21), .A3(n15092), .ZN(n15095)
         );
  INV_X1 U16689 ( .A(keyinput122), .ZN(n15093) );
  NAND4_X1 U16690 ( .A1(keyinput36), .A2(keyinput85), .A3(keyinput114), .A4(
        n15093), .ZN(n15094) );
  NOR4_X1 U16691 ( .A1(n15097), .A2(n15096), .A3(n15095), .A4(n15094), .ZN(
        n15134) );
  NAND4_X1 U16692 ( .A1(keyinput64), .A2(keyinput72), .A3(keyinput74), .A4(
        keyinput83), .ZN(n15104) );
  NOR2_X1 U16693 ( .A1(keyinput17), .A2(keyinput117), .ZN(n15098) );
  NAND3_X1 U16694 ( .A1(keyinput97), .A2(keyinput40), .A3(n15098), .ZN(n15103)
         );
  INV_X1 U16695 ( .A(keyinput1), .ZN(n15099) );
  NAND4_X1 U16696 ( .A1(keyinput37), .A2(keyinput123), .A3(keyinput86), .A4(
        n15099), .ZN(n15102) );
  NOR2_X1 U16697 ( .A1(keyinput54), .A2(keyinput25), .ZN(n15100) );
  NAND3_X1 U16698 ( .A1(keyinput5), .A2(keyinput56), .A3(n15100), .ZN(n15101)
         );
  NOR4_X1 U16699 ( .A1(n15104), .A2(n15103), .A3(n15102), .A4(n15101), .ZN(
        n15133) );
  INV_X1 U16700 ( .A(keyinput76), .ZN(n15105) );
  NOR4_X1 U16701 ( .A1(keyinput24), .A2(keyinput22), .A3(keyinput66), .A4(
        n15105), .ZN(n15111) );
  NAND3_X1 U16702 ( .A1(keyinput92), .A2(keyinput112), .A3(keyinput12), .ZN(
        n15106) );
  NOR2_X1 U16703 ( .A1(keyinput84), .A2(n15106), .ZN(n15110) );
  NAND2_X1 U16704 ( .A1(keyinput8), .A2(keyinput42), .ZN(n15107) );
  NOR3_X1 U16705 ( .A1(keyinput99), .A2(keyinput116), .A3(n15107), .ZN(n15109)
         );
  NOR4_X1 U16706 ( .A1(keyinput126), .A2(keyinput51), .A3(keyinput32), .A4(
        keyinput75), .ZN(n15108) );
  NAND4_X1 U16707 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15131) );
  NOR4_X1 U16708 ( .A1(keyinput7), .A2(keyinput31), .A3(keyinput33), .A4(
        keyinput89), .ZN(n15117) );
  INV_X1 U16709 ( .A(keyinput59), .ZN(n15112) );
  NOR4_X1 U16710 ( .A1(keyinput50), .A2(keyinput125), .A3(keyinput6), .A4(
        n15112), .ZN(n15116) );
  NOR4_X1 U16711 ( .A1(keyinput107), .A2(keyinput15), .A3(keyinput0), .A4(
        keyinput101), .ZN(n15115) );
  NAND3_X1 U16712 ( .A1(keyinput26), .A2(keyinput34), .A3(keyinput61), .ZN(
        n15113) );
  NOR2_X1 U16713 ( .A1(keyinput57), .A2(n15113), .ZN(n15114) );
  NAND4_X1 U16714 ( .A1(n15117), .A2(n15116), .A3(n15115), .A4(n15114), .ZN(
        n15130) );
  AND4_X1 U16715 ( .A1(keyinput16), .A2(keyinput127), .A3(keyinput58), .A4(
        keyinput93), .ZN(n15122) );
  NOR4_X1 U16716 ( .A1(keyinput28), .A2(keyinput124), .A3(keyinput35), .A4(
        keyinput98), .ZN(n15121) );
  NOR4_X1 U16717 ( .A1(keyinput95), .A2(keyinput65), .A3(keyinput55), .A4(
        keyinput106), .ZN(n15120) );
  INV_X1 U16718 ( .A(keyinput118), .ZN(n15118) );
  NOR4_X1 U16719 ( .A1(keyinput87), .A2(keyinput79), .A3(keyinput45), .A4(
        n15118), .ZN(n15119) );
  NAND4_X1 U16720 ( .A1(n15122), .A2(n15121), .A3(n15120), .A4(n15119), .ZN(
        n15129) );
  AND4_X1 U16721 ( .A1(keyinput20), .A2(keyinput77), .A3(keyinput19), .A4(
        keyinput69), .ZN(n15127) );
  NOR4_X1 U16722 ( .A1(keyinput111), .A2(keyinput48), .A3(keyinput90), .A4(
        keyinput41), .ZN(n15126) );
  INV_X1 U16723 ( .A(keyinput100), .ZN(n15123) );
  NOR4_X1 U16724 ( .A1(keyinput88), .A2(keyinput81), .A3(keyinput109), .A4(
        n15123), .ZN(n15125) );
  AND4_X1 U16725 ( .A1(keyinput103), .A2(keyinput53), .A3(keyinput80), .A4(
        keyinput102), .ZN(n15124) );
  NAND4_X1 U16726 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        n15128) );
  NOR4_X1 U16727 ( .A1(n15131), .A2(n15130), .A3(n15129), .A4(n15128), .ZN(
        n15132) );
  NAND4_X1 U16728 ( .A1(n15135), .A2(n15134), .A3(n15133), .A4(n15132), .ZN(
        n15384) );
  AOI22_X1 U16729 ( .A1(n15138), .A2(keyinput6), .B1(keyinput7), .B2(n15137), 
        .ZN(n15136) );
  OAI221_X1 U16730 ( .B1(n15138), .B2(keyinput6), .C1(n15137), .C2(keyinput7), 
        .A(n15136), .ZN(n15149) );
  AOI22_X1 U16731 ( .A1(n15141), .A2(keyinput125), .B1(keyinput50), .B2(n15140), .ZN(n15139) );
  OAI221_X1 U16732 ( .B1(n15141), .B2(keyinput125), .C1(n15140), .C2(
        keyinput50), .A(n15139), .ZN(n15148) );
  AOI22_X1 U16733 ( .A1(P2_U3088), .A2(keyinput31), .B1(keyinput33), .B2(
        n15143), .ZN(n15142) );
  OAI221_X1 U16734 ( .B1(P2_U3088), .B2(keyinput31), .C1(n15143), .C2(
        keyinput33), .A(n15142), .ZN(n15147) );
  XNOR2_X1 U16735 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput12), .ZN(n15145)
         );
  XNOR2_X1 U16736 ( .A(keyinput89), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n15144) );
  NAND2_X1 U16737 ( .A1(n15145), .A2(n15144), .ZN(n15146) );
  NOR4_X1 U16738 ( .A1(n15149), .A2(n15148), .A3(n15147), .A4(n15146), .ZN(
        n15192) );
  AOI22_X1 U16739 ( .A1(n15152), .A2(keyinput92), .B1(n15151), .B2(keyinput24), 
        .ZN(n15150) );
  OAI221_X1 U16740 ( .B1(n15152), .B2(keyinput92), .C1(n15151), .C2(keyinput24), .A(n15150), .ZN(n15161) );
  AOI22_X1 U16741 ( .A1(n9623), .A2(keyinput84), .B1(n15154), .B2(keyinput112), 
        .ZN(n15153) );
  OAI221_X1 U16742 ( .B1(n9623), .B2(keyinput84), .C1(n15154), .C2(keyinput112), .A(n15153), .ZN(n15160) );
  XOR2_X1 U16743 ( .A(n11441), .B(keyinput34), .Z(n15158) );
  XNOR2_X1 U16744 ( .A(SI_9_), .B(keyinput22), .ZN(n15157) );
  XNOR2_X1 U16745 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput76), .ZN(n15156) );
  XNOR2_X1 U16746 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput66), .ZN(n15155) );
  NAND4_X1 U16747 ( .A1(n15158), .A2(n15157), .A3(n15156), .A4(n15155), .ZN(
        n15159) );
  NOR3_X1 U16748 ( .A1(n15161), .A2(n15160), .A3(n15159), .ZN(n15191) );
  AOI22_X1 U16749 ( .A1(n15164), .A2(keyinput101), .B1(keyinput126), .B2(
        n15163), .ZN(n15162) );
  OAI221_X1 U16750 ( .B1(n15164), .B2(keyinput101), .C1(n15163), .C2(
        keyinput126), .A(n15162), .ZN(n15173) );
  AOI22_X1 U16751 ( .A1(n8989), .A2(keyinput26), .B1(keyinput107), .B2(n15166), 
        .ZN(n15165) );
  OAI221_X1 U16752 ( .B1(n8989), .B2(keyinput26), .C1(n15166), .C2(keyinput107), .A(n15165), .ZN(n15172) );
  XOR2_X1 U16753 ( .A(n12886), .B(keyinput0), .Z(n15170) );
  XNOR2_X1 U16754 ( .A(P2_REG0_REG_27__SCAN_IN), .B(keyinput57), .ZN(n15169)
         );
  XNOR2_X1 U16755 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput61), .ZN(n15168) );
  XNOR2_X1 U16756 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput15), .ZN(n15167) );
  NAND4_X1 U16757 ( .A1(n15170), .A2(n15169), .A3(n15168), .A4(n15167), .ZN(
        n15171) );
  NOR3_X1 U16758 ( .A1(n15173), .A2(n15172), .A3(n15171), .ZN(n15190) );
  AOI22_X1 U16759 ( .A1(n15176), .A2(keyinput116), .B1(keyinput32), .B2(n15175), .ZN(n15174) );
  OAI221_X1 U16760 ( .B1(n15176), .B2(keyinput116), .C1(n15175), .C2(
        keyinput32), .A(n15174), .ZN(n15188) );
  AOI22_X1 U16761 ( .A1(n15179), .A2(keyinput99), .B1(n15178), .B2(keyinput8), 
        .ZN(n15177) );
  OAI221_X1 U16762 ( .B1(n15179), .B2(keyinput99), .C1(n15178), .C2(keyinput8), 
        .A(n15177), .ZN(n15187) );
  AOI22_X1 U16763 ( .A1(n15182), .A2(keyinput51), .B1(keyinput42), .B2(n15181), 
        .ZN(n15180) );
  OAI221_X1 U16764 ( .B1(n15182), .B2(keyinput51), .C1(n15181), .C2(keyinput42), .A(n15180), .ZN(n15186) );
  XNOR2_X1 U16765 ( .A(P3_IR_REG_24__SCAN_IN), .B(keyinput111), .ZN(n15184) );
  XNOR2_X1 U16766 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput75), .ZN(n15183)
         );
  NAND2_X1 U16767 ( .A1(n15184), .A2(n15183), .ZN(n15185) );
  NOR4_X1 U16768 ( .A1(n15188), .A2(n15187), .A3(n15186), .A4(n15185), .ZN(
        n15189) );
  NAND4_X1 U16769 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15382) );
  AOI22_X1 U16770 ( .A1(n15195), .A2(keyinput69), .B1(n15194), .B2(keyinput103), .ZN(n15193) );
  OAI221_X1 U16771 ( .B1(n15195), .B2(keyinput69), .C1(n15194), .C2(
        keyinput103), .A(n15193), .ZN(n15201) );
  XNOR2_X1 U16772 ( .A(n15196), .B(keyinput19), .ZN(n15200) );
  XNOR2_X1 U16773 ( .A(n15197), .B(keyinput77), .ZN(n15199) );
  XOR2_X1 U16774 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput41), .Z(n15198) );
  OR4_X1 U16775 ( .A1(n15201), .A2(n15200), .A3(n15199), .A4(n15198), .ZN(
        n15208) );
  INV_X1 U16776 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U16777 ( .A1(n15204), .A2(keyinput48), .B1(keyinput20), .B2(n15203), 
        .ZN(n15202) );
  OAI221_X1 U16778 ( .B1(n15204), .B2(keyinput48), .C1(n15203), .C2(keyinput20), .A(n15202), .ZN(n15207) );
  XNOR2_X1 U16779 ( .A(n15205), .B(keyinput90), .ZN(n15206) );
  NOR3_X1 U16780 ( .A1(n15208), .A2(n15207), .A3(n15206), .ZN(n15257) );
  AOI22_X1 U16781 ( .A1(n15211), .A2(keyinput53), .B1(n15210), .B2(keyinput88), 
        .ZN(n15209) );
  OAI221_X1 U16782 ( .B1(n15211), .B2(keyinput53), .C1(n15210), .C2(keyinput88), .A(n15209), .ZN(n15215) );
  XOR2_X1 U16783 ( .A(SI_3_), .B(keyinput100), .Z(n15214) );
  XNOR2_X1 U16784 ( .A(n15212), .B(keyinput102), .ZN(n15213) );
  OR3_X1 U16785 ( .A1(n15215), .A2(n15214), .A3(n15213), .ZN(n15223) );
  AOI22_X1 U16786 ( .A1(n15217), .A2(keyinput109), .B1(keyinput28), .B2(n14509), .ZN(n15216) );
  OAI221_X1 U16787 ( .B1(n15217), .B2(keyinput109), .C1(n14509), .C2(
        keyinput28), .A(n15216), .ZN(n15222) );
  AOI22_X1 U16788 ( .A1(n15220), .A2(keyinput81), .B1(n15219), .B2(keyinput80), 
        .ZN(n15218) );
  OAI221_X1 U16789 ( .B1(n15220), .B2(keyinput81), .C1(n15219), .C2(keyinput80), .A(n15218), .ZN(n15221) );
  NOR3_X1 U16790 ( .A1(n15223), .A2(n15222), .A3(n15221), .ZN(n15256) );
  AOI22_X1 U16791 ( .A1(n15226), .A2(keyinput124), .B1(n15225), .B2(keyinput16), .ZN(n15224) );
  OAI221_X1 U16792 ( .B1(n15226), .B2(keyinput124), .C1(n15225), .C2(
        keyinput16), .A(n15224), .ZN(n15227) );
  INV_X1 U16793 ( .A(n15227), .ZN(n15231) );
  XOR2_X1 U16794 ( .A(keyinput35), .B(n15228), .Z(n15230) );
  XNOR2_X1 U16795 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput127), .ZN(n15229)
         );
  NAND3_X1 U16796 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(n15237) );
  AOI22_X1 U16797 ( .A1(n15233), .A2(keyinput93), .B1(keyinput118), .B2(n7598), 
        .ZN(n15232) );
  OAI221_X1 U16798 ( .B1(n15233), .B2(keyinput93), .C1(n7598), .C2(keyinput118), .A(n15232), .ZN(n15236) );
  AOI22_X1 U16799 ( .A1(n11033), .A2(keyinput98), .B1(keyinput58), .B2(n9565), 
        .ZN(n15234) );
  OAI221_X1 U16800 ( .B1(n11033), .B2(keyinput98), .C1(n9565), .C2(keyinput58), 
        .A(n15234), .ZN(n15235) );
  NOR3_X1 U16801 ( .A1(n15237), .A2(n15236), .A3(n15235), .ZN(n15255) );
  AOI22_X1 U16802 ( .A1(n15240), .A2(keyinput9), .B1(keyinput106), .B2(n15239), 
        .ZN(n15238) );
  OAI221_X1 U16803 ( .B1(n15240), .B2(keyinput9), .C1(n15239), .C2(keyinput106), .A(n15238), .ZN(n15253) );
  AOI22_X1 U16804 ( .A1(n15243), .A2(keyinput45), .B1(keyinput95), .B2(n15242), 
        .ZN(n15241) );
  OAI221_X1 U16805 ( .B1(n15243), .B2(keyinput45), .C1(n15242), .C2(keyinput95), .A(n15241), .ZN(n15252) );
  AOI22_X1 U16806 ( .A1(n15246), .A2(keyinput65), .B1(n15245), .B2(keyinput55), 
        .ZN(n15244) );
  OAI221_X1 U16807 ( .B1(n15246), .B2(keyinput65), .C1(n15245), .C2(keyinput55), .A(n15244), .ZN(n15251) );
  INV_X1 U16808 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15247) );
  XOR2_X1 U16809 ( .A(n15247), .B(keyinput79), .Z(n15249) );
  XNOR2_X1 U16810 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput87), .ZN(n15248) );
  NAND2_X1 U16811 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  NOR4_X1 U16812 ( .A1(n15253), .A2(n15252), .A3(n15251), .A4(n15250), .ZN(
        n15254) );
  NAND4_X1 U16813 ( .A1(n15257), .A2(n15256), .A3(n15255), .A4(n15254), .ZN(
        n15381) );
  AOI22_X1 U16814 ( .A1(n15260), .A2(keyinput5), .B1(keyinput25), .B2(n15259), 
        .ZN(n15258) );
  OAI221_X1 U16815 ( .B1(n15260), .B2(keyinput5), .C1(n15259), .C2(keyinput25), 
        .A(n15258), .ZN(n15270) );
  AOI22_X1 U16816 ( .A1(n15262), .A2(keyinput86), .B1(keyinput119), .B2(n8407), 
        .ZN(n15261) );
  OAI221_X1 U16817 ( .B1(n15262), .B2(keyinput86), .C1(n8407), .C2(keyinput119), .A(n15261), .ZN(n15269) );
  XNOR2_X1 U16818 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput1), .ZN(n15265)
         );
  XNOR2_X1 U16819 ( .A(SI_5_), .B(keyinput37), .ZN(n15264) );
  XNOR2_X1 U16820 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput123), .ZN(n15263)
         );
  NAND3_X1 U16821 ( .A1(n15265), .A2(n15264), .A3(n15263), .ZN(n15268) );
  XNOR2_X1 U16822 ( .A(n15266), .B(keyinput56), .ZN(n15267) );
  NOR4_X1 U16823 ( .A1(n15270), .A2(n15269), .A3(n15268), .A4(n15267), .ZN(
        n15316) );
  AOI22_X1 U16824 ( .A1(n9618), .A2(keyinput83), .B1(keyinput40), .B2(n10491), 
        .ZN(n15271) );
  OAI221_X1 U16825 ( .B1(n9618), .B2(keyinput83), .C1(n10491), .C2(keyinput40), 
        .A(n15271), .ZN(n15283) );
  AOI22_X1 U16826 ( .A1(n15274), .A2(keyinput97), .B1(n15273), .B2(keyinput64), 
        .ZN(n15272) );
  OAI221_X1 U16827 ( .B1(n15274), .B2(keyinput97), .C1(n15273), .C2(keyinput64), .A(n15272), .ZN(n15282) );
  AOI22_X1 U16828 ( .A1(n15277), .A2(keyinput72), .B1(n15276), .B2(keyinput74), 
        .ZN(n15275) );
  OAI221_X1 U16829 ( .B1(n15277), .B2(keyinput72), .C1(n15276), .C2(keyinput74), .A(n15275), .ZN(n15281) );
  XNOR2_X1 U16830 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput117), .ZN(n15279)
         );
  XNOR2_X1 U16831 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput54), .ZN(n15278) );
  NAND2_X1 U16832 ( .A1(n15279), .A2(n15278), .ZN(n15280) );
  NOR4_X1 U16833 ( .A1(n15283), .A2(n15282), .A3(n15281), .A4(n15280), .ZN(
        n15315) );
  AOI22_X1 U16834 ( .A1(n15286), .A2(keyinput122), .B1(n15285), .B2(keyinput29), .ZN(n15284) );
  OAI221_X1 U16835 ( .B1(n15286), .B2(keyinput122), .C1(n15285), .C2(
        keyinput29), .A(n15284), .ZN(n15297) );
  AOI22_X1 U16836 ( .A1(n15289), .A2(keyinput36), .B1(n15288), .B2(keyinput114), .ZN(n15287) );
  OAI221_X1 U16837 ( .B1(n15289), .B2(keyinput36), .C1(n15288), .C2(
        keyinput114), .A(n15287), .ZN(n15296) );
  AOI22_X1 U16838 ( .A1(n9515), .A2(keyinput21), .B1(n10923), .B2(keyinput59), 
        .ZN(n15290) );
  OAI221_X1 U16839 ( .B1(n9515), .B2(keyinput21), .C1(n10923), .C2(keyinput59), 
        .A(n15290), .ZN(n15295) );
  AOI22_X1 U16840 ( .A1(n15293), .A2(keyinput78), .B1(keyinput4), .B2(n15292), 
        .ZN(n15291) );
  OAI221_X1 U16841 ( .B1(n15293), .B2(keyinput78), .C1(n15292), .C2(keyinput4), 
        .A(n15291), .ZN(n15294) );
  NOR4_X1 U16842 ( .A1(n15297), .A2(n15296), .A3(n15295), .A4(n15294), .ZN(
        n15314) );
  AOI22_X1 U16843 ( .A1(n15300), .A2(keyinput71), .B1(n15299), .B2(keyinput120), .ZN(n15298) );
  OAI221_X1 U16844 ( .B1(n15300), .B2(keyinput71), .C1(n15299), .C2(
        keyinput120), .A(n15298), .ZN(n15312) );
  AOI22_X1 U16845 ( .A1(n15303), .A2(keyinput18), .B1(keyinput23), .B2(n15302), 
        .ZN(n15301) );
  OAI221_X1 U16846 ( .B1(n15303), .B2(keyinput18), .C1(n15302), .C2(keyinput23), .A(n15301), .ZN(n15311) );
  AOI22_X1 U16847 ( .A1(n15306), .A2(keyinput121), .B1(keyinput104), .B2(
        n15305), .ZN(n15304) );
  OAI221_X1 U16848 ( .B1(n15306), .B2(keyinput121), .C1(n15305), .C2(
        keyinput104), .A(n15304), .ZN(n15310) );
  XNOR2_X1 U16849 ( .A(P3_REG1_REG_22__SCAN_IN), .B(keyinput10), .ZN(n15308)
         );
  XNOR2_X1 U16850 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput85), .ZN(n15307) );
  NAND2_X1 U16851 ( .A1(n15308), .A2(n15307), .ZN(n15309) );
  NOR4_X1 U16852 ( .A1(n15312), .A2(n15311), .A3(n15310), .A4(n15309), .ZN(
        n15313) );
  NAND4_X1 U16853 ( .A1(n15316), .A2(n15315), .A3(n15314), .A4(n15313), .ZN(
        n15380) );
  AOI22_X1 U16854 ( .A1(n15319), .A2(keyinput52), .B1(keyinput96), .B2(n15318), 
        .ZN(n15317) );
  OAI221_X1 U16855 ( .B1(n15319), .B2(keyinput52), .C1(n15318), .C2(keyinput96), .A(n15317), .ZN(n15331) );
  INV_X1 U16856 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U16857 ( .A1(n15322), .A2(keyinput91), .B1(keyinput2), .B2(n15321), 
        .ZN(n15320) );
  OAI221_X1 U16858 ( .B1(n15322), .B2(keyinput91), .C1(n15321), .C2(keyinput2), 
        .A(n15320), .ZN(n15330) );
  INV_X1 U16859 ( .A(keyinput110), .ZN(n15324) );
  AOI22_X1 U16860 ( .A1(n15325), .A2(keyinput67), .B1(P3_WR_REG_SCAN_IN), .B2(
        n15324), .ZN(n15323) );
  OAI221_X1 U16861 ( .B1(n15325), .B2(keyinput67), .C1(n15324), .C2(
        P3_WR_REG_SCAN_IN), .A(n15323), .ZN(n15329) );
  XNOR2_X1 U16862 ( .A(P3_REG1_REG_1__SCAN_IN), .B(keyinput44), .ZN(n15327) );
  XNOR2_X1 U16863 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput30), .ZN(n15326)
         );
  NAND2_X1 U16864 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  NOR4_X1 U16865 ( .A1(n15331), .A2(n15330), .A3(n15329), .A4(n15328), .ZN(
        n15378) );
  AOI22_X1 U16866 ( .A1(n15334), .A2(keyinput13), .B1(n15333), .B2(keyinput108), .ZN(n15332) );
  OAI221_X1 U16867 ( .B1(n15334), .B2(keyinput13), .C1(n15333), .C2(
        keyinput108), .A(n15332), .ZN(n15345) );
  INV_X1 U16868 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n15337) );
  AOI22_X1 U16869 ( .A1(n15337), .A2(keyinput62), .B1(n15336), .B2(keyinput70), 
        .ZN(n15335) );
  OAI221_X1 U16870 ( .B1(n15337), .B2(keyinput62), .C1(n15336), .C2(keyinput70), .A(n15335), .ZN(n15344) );
  AOI22_X1 U16871 ( .A1(n13575), .A2(keyinput63), .B1(n15339), .B2(keyinput46), 
        .ZN(n15338) );
  OAI221_X1 U16872 ( .B1(n13575), .B2(keyinput63), .C1(n15339), .C2(keyinput46), .A(n15338), .ZN(n15343) );
  INV_X1 U16873 ( .A(keyinput60), .ZN(n15341) );
  XNOR2_X1 U16874 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput115), .ZN(n15340) );
  OAI21_X1 U16875 ( .B1(P3_REG0_REG_20__SCAN_IN), .B2(n15341), .A(n15340), 
        .ZN(n15342) );
  NOR4_X1 U16876 ( .A1(n15345), .A2(n15344), .A3(n15343), .A4(n15342), .ZN(
        n15377) );
  AOI22_X1 U16877 ( .A1(n15391), .A2(keyinput14), .B1(n15347), .B2(keyinput105), .ZN(n15346) );
  OAI221_X1 U16878 ( .B1(n15391), .B2(keyinput14), .C1(n15347), .C2(
        keyinput105), .A(n15346), .ZN(n15358) );
  AOI22_X1 U16879 ( .A1(n15350), .A2(keyinput94), .B1(n15349), .B2(keyinput38), 
        .ZN(n15348) );
  OAI221_X1 U16880 ( .B1(n15350), .B2(keyinput94), .C1(n15349), .C2(keyinput38), .A(n15348), .ZN(n15357) );
  AOI22_X1 U16881 ( .A1(n15352), .A2(keyinput49), .B1(n9849), .B2(keyinput17), 
        .ZN(n15351) );
  OAI221_X1 U16882 ( .B1(n15352), .B2(keyinput49), .C1(n9849), .C2(keyinput17), 
        .A(n15351), .ZN(n15356) );
  AOI22_X1 U16883 ( .A1(n15354), .A2(keyinput47), .B1(n10739), .B2(keyinput113), .ZN(n15353) );
  OAI221_X1 U16884 ( .B1(n15354), .B2(keyinput47), .C1(n10739), .C2(
        keyinput113), .A(n15353), .ZN(n15355) );
  NOR4_X1 U16885 ( .A1(n15358), .A2(n15357), .A3(n15356), .A4(n15355), .ZN(
        n15376) );
  AOI22_X1 U16886 ( .A1(n15361), .A2(keyinput68), .B1(keyinput27), .B2(n15360), 
        .ZN(n15359) );
  OAI221_X1 U16887 ( .B1(n15361), .B2(keyinput68), .C1(n15360), .C2(keyinput27), .A(n15359), .ZN(n15374) );
  AOI22_X1 U16888 ( .A1(n15364), .A2(keyinput73), .B1(keyinput11), .B2(n15363), 
        .ZN(n15362) );
  OAI221_X1 U16889 ( .B1(n15364), .B2(keyinput73), .C1(n15363), .C2(keyinput11), .A(n15362), .ZN(n15373) );
  AOI22_X1 U16890 ( .A1(n15367), .A2(keyinput43), .B1(n15366), .B2(keyinput3), 
        .ZN(n15365) );
  OAI221_X1 U16891 ( .B1(n15367), .B2(keyinput43), .C1(n15366), .C2(keyinput3), 
        .A(n15365), .ZN(n15372) );
  XOR2_X1 U16892 ( .A(n15368), .B(keyinput82), .Z(n15370) );
  XNOR2_X1 U16893 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput39), .ZN(n15369) );
  NAND2_X1 U16894 ( .A1(n15370), .A2(n15369), .ZN(n15371) );
  NOR4_X1 U16895 ( .A1(n15374), .A2(n15373), .A3(n15372), .A4(n15371), .ZN(
        n15375) );
  NAND4_X1 U16896 ( .A1(n15378), .A2(n15377), .A3(n15376), .A4(n15375), .ZN(
        n15379) );
  NOR4_X1 U16897 ( .A1(n15382), .A2(n15381), .A3(n15380), .A4(n15379), .ZN(
        n15383) );
  OAI221_X1 U16898 ( .B1(n15385), .B2(keyinput60), .C1(n15385), .C2(n15384), 
        .A(n15383), .ZN(n15386) );
  XOR2_X1 U16899 ( .A(n15387), .B(n15386), .Z(P3_U3377) );
  XOR2_X1 U16900 ( .A(n15389), .B(n15388), .Z(SUB_1596_U59) );
  XNOR2_X1 U16901 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15390), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16902 ( .B1(n15392), .B2(n15391), .A(n15401), .ZN(SUB_1596_U53) );
  XOR2_X1 U16903 ( .A(n15394), .B(n15393), .Z(SUB_1596_U56) );
  OAI21_X1 U16904 ( .B1(n15397), .B2(n15396), .A(n15395), .ZN(n15399) );
  XOR2_X1 U16905 ( .A(n15399), .B(n15398), .Z(SUB_1596_U60) );
  XOR2_X1 U16906 ( .A(n15401), .B(n15400), .Z(SUB_1596_U5) );
  AND3_X1 U9853 ( .A1(n7564), .A2(n7563), .A3(n7562), .ZN(n8124) );
  NAND2_X1 U7371 ( .A1(n7584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7582) );
  INV_X2 U7321 ( .A(n7980), .ZN(n13439) );
  BUF_X2 U7323 ( .A(n8917), .Z(n11430) );
  NAND2_X2 U7338 ( .A1(n6970), .A2(n6969), .ZN(n13485) );
  NOR2_X1 U7359 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7282) );
  OR2_X1 U7369 ( .A1(n11591), .A2(n7035), .ZN(n7034) );
  INV_X2 U7379 ( .A(n13474), .ZN(n7790) );
  AND4_X1 U7381 ( .A1(n7278), .A2(n7277), .A3(n7276), .A4(n7275), .ZN(n7279)
         );
  CLKBUF_X1 U7507 ( .A(n8277), .Z(n11764) );
  NAND2_X2 U7628 ( .A1(n14041), .A2(n8115), .ZN(n9506) );
  CLKBUF_X1 U9212 ( .A(n8832), .Z(n6559) );
  AND2_X1 U9377 ( .A1(n7489), .A2(n7488), .ZN(n15407) );
endmodule

