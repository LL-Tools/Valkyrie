

module b20_C_gen_AntiSAT_k_128_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276;

  AND3_X1 U4852 ( .A1(n4785), .A2(n4787), .A3(n8484), .ZN(n8488) );
  NOR2_X1 U4853 ( .A1(n4403), .A2(n8304), .ZN(n8313) );
  AND2_X1 U4854 ( .A1(n7531), .A2(n7530), .ZN(n9417) );
  INV_X1 U4855 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n9827) );
  INV_X1 U4856 ( .A(n9140), .ZN(n9316) );
  NAND2_X1 U4857 ( .A1(n5641), .A2(n5640), .ZN(n9347) );
  CLKBUF_X2 U4858 ( .A(n5039), .Z(n7645) );
  CLKBUF_X2 U4859 ( .A(n5025), .Z(n6498) );
  CLKBUF_X2 U4860 ( .A(n5673), .Z(n5503) );
  CLKBUF_X1 U4861 ( .A(n5961), .Z(n6308) );
  INV_X1 U4862 ( .A(n5077), .ZN(n5118) );
  CLKBUF_X2 U4863 ( .A(n5088), .Z(n5664) );
  CLKBUF_X3 U4864 ( .A(n5094), .Z(n4352) );
  OR2_X2 U4865 ( .A1(n5758), .A2(n5893), .ZN(n5040) );
  CLKBUF_X2 U4866 ( .A(n5994), .Z(n4353) );
  NAND2_X1 U4867 ( .A1(n4960), .A2(n5857), .ZN(n4974) );
  XNOR2_X1 U4868 ( .A(n4991), .B(n4990), .ZN(n4996) );
  AND2_X1 U4869 ( .A1(n5949), .A2(n8856), .ZN(n5973) );
  INV_X1 U4870 ( .A(n5489), .ZN(n5886) );
  NAND2_X1 U4871 ( .A1(n9471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4991) );
  XNOR2_X1 U4872 ( .A(n4940), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5489) );
  INV_X1 U4875 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4876 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4933) );
  INV_X1 U4877 ( .A(n5118), .ZN(n5492) );
  NOR2_X1 U4878 ( .A1(n8436), .A2(n4566), .ZN(n8459) );
  INV_X1 U4879 ( .A(n8290), .ZN(n8297) );
  OR2_X1 U4881 ( .A1(n8438), .A2(n4788), .ZN(n4787) );
  INV_X1 U4882 ( .A(n5994), .ZN(n6204) );
  AND2_X1 U4883 ( .A1(n7161), .A2(n5260), .ZN(n5264) );
  OR2_X1 U4884 ( .A1(n5831), .A2(n4675), .ZN(n4465) );
  NAND2_X1 U4885 ( .A1(n4391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4971) );
  INV_X1 U4887 ( .A(n9347), .ZN(n8900) );
  INV_X2 U4888 ( .A(n5040), .ZN(n6478) );
  AND2_X1 U4889 ( .A1(n5266), .A2(n5242), .ZN(n4924) );
  AND2_X1 U4890 ( .A1(n5717), .A2(n5716), .ZN(n9327) );
  OR2_X1 U4891 ( .A1(n4392), .A2(n4474), .ZN(n9315) );
  NAND2_X1 U4892 ( .A1(n4643), .A2(n4499), .ZN(n6579) );
  NAND2_X1 U4893 ( .A1(n5787), .A2(n5786), .ZN(n7504) );
  XNOR2_X1 U4895 ( .A(n5164), .B(n10198), .ZN(n5162) );
  CLKBUF_X3 U4896 ( .A(n5267), .Z(n7525) );
  INV_X1 U4897 ( .A(n6673), .ZN(n6674) );
  NAND2_X1 U4898 ( .A1(n5689), .A2(n5688), .ZN(n9140) );
  BUF_X1 U4899 ( .A(n9011), .Z(n4349) );
  INV_X1 U4900 ( .A(n9148), .ZN(n5883) );
  AND2_X2 U4901 ( .A1(n4902), .A2(n4977), .ZN(n4900) );
  NOR2_X2 U4902 ( .A1(n4969), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4902) );
  NOR2_X4 U4903 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5041) );
  OR2_X1 U4904 ( .A1(n8523), .A2(n8283), .ZN(n4856) );
  INV_X2 U4905 ( .A(n6845), .ZN(n6687) );
  NAND2_X2 U4906 ( .A1(n6302), .A2(n6303), .ZN(n5970) );
  OR2_X2 U4907 ( .A1(n5560), .A2(n5559), .ZN(n4912) );
  OAI21_X2 U4908 ( .B1(n5533), .B2(n5534), .A(n5537), .ZN(n5560) );
  NOR2_X4 U4909 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5109) );
  NAND4_X1 U4910 ( .A1(n5093), .A2(n5092), .A3(n5091), .A4(n5090), .ZN(n9011)
         );
  AOI21_X4 U4911 ( .B1(n7140), .B2(n5264), .A(n4923), .ZN(n7313) );
  NAND2_X2 U4912 ( .A1(n7139), .A2(n7142), .ZN(n7140) );
  NAND2_X4 U4913 ( .A1(n5727), .A2(n4973), .ZN(n6395) );
  XNOR2_X2 U4914 ( .A(n4964), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5727) );
  AOI21_X2 U4915 ( .B1(n9549), .B2(n8224), .A(n6325), .ZN(n8677) );
  NAND2_X2 U4916 ( .A1(n8694), .A2(n8219), .ZN(n9549) );
  AOI211_X2 U4917 ( .C1(n7637), .C2(n7636), .A(n7635), .B(n7702), .ZN(n7640)
         );
  AOI21_X2 U4918 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8397), .A(n8396), .ZN(
        n8420) );
  XNOR2_X1 U4920 ( .A(n5982), .B(n5981), .ZN(n6420) );
  INV_X1 U4921 ( .A(n5118), .ZN(n4351) );
  INV_X1 U4922 ( .A(n4696), .ZN(n5077) );
  INV_X1 U4923 ( .A(n5118), .ZN(n5711) );
  OAI21_X1 U4924 ( .B1(n4975), .B2(n4974), .A(n6395), .ZN(n4696) );
  NAND2_X2 U4925 ( .A1(n4820), .A2(n4819), .ZN(n5063) );
  OR2_X2 U4926 ( .A1(n8846), .A2(n8847), .ZN(n5939) );
  AND2_X1 U4927 ( .A1(n5040), .A2(n7525), .ZN(n5094) );
  NAND2_X2 U4928 ( .A1(n5564), .A2(n5563), .ZN(n9222) );
  AND2_X1 U4929 ( .A1(n6343), .A2(n6342), .ZN(n7877) );
  NOR2_X2 U4930 ( .A1(n9127), .A2(n9316), .ZN(n7724) );
  AND2_X1 U4931 ( .A1(n5883), .A2(n9159), .ZN(n7708) );
  NAND2_X2 U4932 ( .A1(n7705), .A2(n7719), .ZN(n9163) );
  INV_X1 U4933 ( .A(n9355), .ZN(n9375) );
  INV_X1 U4934 ( .A(n6319), .ZN(n9917) );
  NAND2_X1 U4935 ( .A1(n8154), .A2(n8155), .ZN(n6319) );
  NAND2_X1 U4936 ( .A1(n5206), .A2(n5205), .ZN(n5236) );
  INV_X1 U4937 ( .A(n7105), .ZN(n6994) );
  OR2_X1 U4938 ( .A1(n5986), .A2(n9930), .ZN(n8154) );
  OR2_X1 U4939 ( .A1(n7745), .A2(n5310), .ZN(n5005) );
  OAI211_X1 U4940 ( .C1(n5995), .C2(n6455), .A(n4639), .B(n4410), .ZN(n6845)
         );
  CLKBUF_X1 U4941 ( .A(n5811), .Z(n9013) );
  NAND2_X1 U4942 ( .A1(n5117), .A2(n5116), .ZN(n9770) );
  INV_X1 U4943 ( .A(n7654), .ZN(n7660) );
  INV_X1 U4944 ( .A(n5094), .ZN(n5212) );
  OR2_X1 U4945 ( .A1(n5989), .A2(n6402), .ZN(n5956) );
  CLKBUF_X2 U4947 ( .A(n6303), .Z(n8473) );
  OAI21_X1 U4948 ( .B1(n4963), .B2(n4962), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4964) );
  NAND2_X1 U4949 ( .A1(n7877), .A2(n6345), .ZN(n6392) );
  OAI21_X1 U4950 ( .B1(n8116), .B2(n4363), .A(n4373), .ZN(n4846) );
  INV_X1 U4951 ( .A(n8152), .ZN(n8309) );
  AND2_X1 U4952 ( .A1(n4502), .A2(n7657), .ZN(n7658) );
  OR2_X1 U4953 ( .A1(n7653), .A2(n9084), .ZN(n7651) );
  OR2_X1 U4954 ( .A1(n7653), .A2(n9421), .ZN(n4502) );
  AOI21_X1 U4955 ( .B1(n8305), .B2(n8306), .A(n8304), .ZN(n8314) );
  MUX2_X1 U4956 ( .A(n7642), .B(n7641), .S(n7654), .Z(n7644) );
  OR2_X1 U4957 ( .A1(n8703), .A2(n8117), .ZN(n8298) );
  OR2_X1 U4958 ( .A1(n9123), .A2(n4875), .ZN(n4874) );
  AOI21_X1 U4959 ( .B1(n8845), .B2(n8115), .A(n8114), .ZN(n8763) );
  NAND2_X1 U4960 ( .A1(n7647), .A2(n7646), .ZN(n9084) );
  NAND2_X1 U4961 ( .A1(n5854), .A2(n5853), .ZN(n5897) );
  NAND2_X1 U4962 ( .A1(n4471), .A2(n5840), .ZN(n9162) );
  NAND2_X1 U4963 ( .A1(n8461), .A2(n4786), .ZN(n4785) );
  OR2_X1 U4964 ( .A1(n9118), .A2(n9327), .ZN(n7728) );
  NAND2_X1 U4965 ( .A1(n4472), .A2(n4400), .ZN(n9192) );
  NAND2_X1 U4966 ( .A1(n6256), .A2(n6255), .ZN(n8712) );
  NAND2_X1 U4967 ( .A1(n5708), .A2(n5707), .ZN(n5781) );
  NAND2_X1 U4968 ( .A1(n6248), .A2(n6247), .ZN(n8784) );
  NAND2_X2 U4969 ( .A1(n5606), .A2(n5605), .ZN(n9187) );
  NAND2_X1 U4970 ( .A1(n4740), .A2(n4737), .ZN(n8053) );
  NOR2_X1 U4971 ( .A1(n7881), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U4972 ( .A1(n5586), .A2(n5585), .ZN(n9203) );
  NAND2_X1 U4973 ( .A1(n4888), .A2(n4886), .ZN(n7438) );
  NAND2_X1 U4974 ( .A1(n4792), .A2(n4791), .ZN(n8343) );
  OR2_X1 U4975 ( .A1(n7411), .A2(n7363), .ZN(n4792) );
  NOR2_X1 U4976 ( .A1(n7412), .A2(n10001), .ZN(n7411) );
  NAND2_X1 U4977 ( .A1(n7096), .A2(n5822), .ZN(n7051) );
  NAND2_X1 U4978 ( .A1(n4473), .A2(n4398), .ZN(n7096) );
  XNOR2_X1 U4979 ( .A(n7362), .B(n7386), .ZN(n7412) );
  AND2_X1 U4980 ( .A1(n7361), .A2(n7360), .ZN(n7362) );
  OR2_X1 U4981 ( .A1(n9736), .A2(n9735), .ZN(n4473) );
  NAND2_X1 U4982 ( .A1(n4563), .A2(n4562), .ZN(n7361) );
  NAND2_X1 U4983 ( .A1(n4894), .A2(n4895), .ZN(n7203) );
  OR2_X1 U4984 ( .A1(n7126), .A2(n7127), .ZN(n4563) );
  NOR2_X1 U4985 ( .A1(n7187), .A2(n4918), .ZN(n7190) );
  OR2_X1 U4986 ( .A1(n5508), .A2(n5507), .ZN(n5510) );
  XNOR2_X1 U4987 ( .A(n7124), .B(n7125), .ZN(n7079) );
  OAI21_X1 U4988 ( .B1(n7076), .B2(n4796), .A(n4795), .ZN(n7124) );
  NAND2_X1 U4989 ( .A1(n4797), .A2(n7077), .ZN(n4796) );
  NAND2_X1 U4990 ( .A1(n5357), .A2(n5356), .ZN(n7433) );
  NAND2_X1 U4991 ( .A1(n5406), .A2(n5405), .ZN(n5430) );
  NOR2_X1 U4992 ( .A1(n9996), .A2(n6913), .ZN(n7076) );
  NAND2_X1 U4993 ( .A1(n5246), .A2(n5245), .ZN(n9788) );
  XNOR2_X1 U4994 ( .A(n4569), .B(n7060), .ZN(n6913) );
  AND3_X2 U4995 ( .A1(n6391), .A2(n6390), .A3(n6617), .ZN(n10003) );
  NAND2_X1 U4996 ( .A1(n9885), .A2(n6912), .ZN(n4569) );
  OR2_X1 U4997 ( .A1(n9883), .A2(n9884), .ZN(n9885) );
  NAND2_X1 U4998 ( .A1(n5236), .A2(n4364), .ZN(n4527) );
  NAND2_X1 U4999 ( .A1(n5006), .A2(n5005), .ZN(n5020) );
  NAND2_X1 U5000 ( .A1(n6609), .A2(n6687), .ZN(n8161) );
  AND2_X1 U5001 ( .A1(n8175), .A2(n8183), .ZN(n8172) );
  NOR2_X1 U5002 ( .A1(n9861), .A2(n9993), .ZN(n9860) );
  NAND2_X1 U5003 ( .A1(n6679), .A2(n6678), .ZN(n6712) );
  NOR2_X2 U5004 ( .A1(n8456), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U5005 ( .A1(n9737), .A2(n5861), .ZN(n9812) );
  AND2_X1 U5006 ( .A1(n5136), .A2(n5135), .ZN(n7544) );
  AND2_X1 U5007 ( .A1(n6909), .A2(n4437), .ZN(n6910) );
  NOR2_X1 U5008 ( .A1(n9014), .A2(n6755), .ZN(n6524) );
  AND3_X1 U5009 ( .A1(n5985), .A2(n5984), .A3(n5983), .ZN(n9930) );
  CLKBUF_X1 U5010 ( .A(n5863), .Z(n9014) );
  INV_X1 U5011 ( .A(n6579), .ZN(n7745) );
  AND3_X1 U5012 ( .A1(n4387), .A2(n4526), .A3(n4525), .ZN(n4524) );
  NAND4_X1 U5013 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n9012)
         );
  XNOR2_X1 U5014 ( .A(n6353), .B(n6352), .ZN(n7806) );
  AND4_X2 U5015 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n9923)
         );
  AND4_X1 U5016 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n9921)
         );
  CLKBUF_X1 U5017 ( .A(n5975), .Z(n4356) );
  XNOR2_X1 U5018 ( .A(n6203), .B(n6202), .ZN(n8482) );
  NAND2_X1 U5019 ( .A1(n6357), .A2(n6356), .ZN(n6362) );
  NAND2_X1 U5020 ( .A1(n5970), .A2(n5064), .ZN(n5995) );
  OR2_X1 U5021 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  INV_X1 U5022 ( .A(n5002), .ZN(n6795) );
  NAND2_X1 U5023 ( .A1(n4939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U5024 ( .A1(n5933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  OR2_X1 U5025 ( .A1(n7669), .A2(n4909), .ZN(n5002) );
  XNOR2_X1 U5026 ( .A(n5942), .B(n5941), .ZN(n8856) );
  OR2_X1 U5027 ( .A1(n4957), .A2(n4956), .ZN(n4958) );
  NAND2_X1 U5028 ( .A1(n9908), .A2(n7077), .ZN(n4795) );
  NAND2_X2 U5029 ( .A1(n7525), .A2(P1_U3086), .ZN(n6469) );
  MUX2_X1 U5030 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5932), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5934) );
  NAND2_X1 U5031 ( .A1(n4989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4978) );
  OR2_X1 U5032 ( .A1(n4992), .A2(n4945), .ZN(n4994) );
  XNOR2_X1 U5033 ( .A(n4953), .B(n4954), .ZN(n7669) );
  NAND2_X1 U5034 ( .A1(n4776), .A2(n6417), .ZN(n9851) );
  NAND2_X1 U5035 ( .A1(n4938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5511) );
  OR2_X1 U5036 ( .A1(n6561), .A2(n6402), .ZN(n4776) );
  OR2_X1 U5037 ( .A1(n4955), .A2(n4945), .ZN(n4953) );
  OAI21_X1 U5038 ( .B1(n5064), .B2(n5066), .A(n5065), .ZN(n5098) );
  NAND2_X1 U5039 ( .A1(n4470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4980) );
  OAI21_X1 U5040 ( .B1(n6437), .B2(n6416), .A(n6417), .ZN(n6561) );
  AND2_X1 U5041 ( .A1(n4758), .A2(n5980), .ZN(n4483) );
  NOR2_X1 U5042 ( .A1(n5926), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4872) );
  AND3_X1 U5043 ( .A1(n4941), .A2(n4961), .A3(n4948), .ZN(n4968) );
  AND2_X1 U5044 ( .A1(n6007), .A2(n5916), .ZN(n4758) );
  AND2_X1 U5045 ( .A1(n4981), .A2(n4976), .ZN(n4977) );
  INV_X1 U5046 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6377) );
  INV_X1 U5047 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4757) );
  INV_X1 U5048 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5931) );
  INV_X1 U5049 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4990) );
  INV_X1 U5050 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4948) );
  INV_X2 U5051 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5981) );
  INV_X1 U5052 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6185) );
  NOR2_X1 U5053 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4934) );
  NOR2_X1 U5054 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4936) );
  XNOR2_X2 U5055 ( .A(n5232), .B(n5233), .ZN(n7139) );
  XNOR2_X2 U5056 ( .A(n5397), .B(n5398), .ZN(n8859) );
  NAND2_X2 U5057 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  NAND4_X2 U5058 ( .A1(n5001), .A2(n5000), .A3(n4999), .A4(n4998), .ZN(n5811)
         );
  OAI21_X1 U5059 ( .B1(n8975), .B2(n5724), .A(n5725), .ZN(n5726) );
  CLKBUF_X2 U5060 ( .A(n5986), .Z(n4354) );
  INV_X2 U5061 ( .A(n9923), .ZN(n6609) );
  XNOR2_X1 U5062 ( .A(n4978), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5758) );
  OR2_X1 U5063 ( .A1(n4996), .A2(n4995), .ZN(n5088) );
  AND2_X1 U5064 ( .A1(n4995), .A2(n4996), .ZN(n5058) );
  NAND4_X2 U5065 ( .A1(n5041), .A2(n4889), .A3(n5109), .A4(n4932), .ZN(n5182)
         );
  NOR2_X2 U5066 ( .A1(n5940), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8846) );
  XNOR2_X2 U5067 ( .A(n4971), .B(n4970), .ZN(n7408) );
  CLKBUF_X1 U5068 ( .A(n5893), .Z(n4358) );
  XNOR2_X1 U5069 ( .A(n4982), .B(n4981), .ZN(n5893) );
  NAND2_X1 U5070 ( .A1(n6302), .A2(n6303), .ZN(n4359) );
  NAND2_X1 U5071 ( .A1(n6302), .A2(n6303), .ZN(n4360) );
  NAND2_X1 U5072 ( .A1(n9476), .A2(n4995), .ZN(n4361) );
  NAND2_X4 U5073 ( .A1(n9476), .A2(n4995), .ZN(n5089) );
  OAI21_X2 U5074 ( .B1(n8642), .B2(n6328), .A(n8235), .ZN(n8633) );
  NAND2_X2 U5075 ( .A1(n6327), .A2(n8231), .ZN(n8642) );
  AOI21_X2 U5076 ( .B1(n8499), .B2(n8500), .A(n6336), .ZN(n8106) );
  XNOR2_X2 U5077 ( .A(n5939), .B(n5938), .ZN(n5949) );
  NOR2_X2 U5078 ( .A1(n8897), .A2(n8896), .ZN(n8895) );
  NAND2_X1 U5079 ( .A1(n4359), .A2(n7525), .ZN(n5994) );
  XNOR2_X2 U5080 ( .A(n5930), .B(n5929), .ZN(n6302) );
  NAND2_X1 U5081 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NOR2_X1 U5082 ( .A1(n8424), .A2(n8750), .ZN(n4566) );
  AOI21_X1 U5083 ( .B1(n4602), .B2(n8144), .A(n4405), .ZN(n4600) );
  INV_X1 U5084 ( .A(n4839), .ZN(n4838) );
  OAI21_X1 U5085 ( .B1(n4841), .B2(n4840), .A(n5376), .ZN(n4839) );
  NOR2_X1 U5086 ( .A1(n8432), .A2(n4802), .ZN(n8445) );
  NOR2_X1 U5087 ( .A1(n8424), .A2(n8652), .ZN(n4802) );
  INV_X1 U5088 ( .A(n8482), .ZN(n8472) );
  NAND2_X1 U5089 ( .A1(n5839), .A2(n4679), .ZN(n4471) );
  NOR2_X1 U5090 ( .A1(n4412), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U5091 ( .A1(n4509), .A2(n4508), .ZN(n7571) );
  NAND2_X1 U5092 ( .A1(n4515), .A2(n8993), .ZN(n4508) );
  NAND2_X1 U5093 ( .A1(n4510), .A2(n9398), .ZN(n4509) );
  OR2_X1 U5094 ( .A1(n4515), .A2(n8993), .ZN(n4510) );
  NAND2_X1 U5095 ( .A1(n7604), .A2(n7771), .ZN(n4523) );
  NAND2_X1 U5096 ( .A1(n8276), .A2(n4534), .ZN(n4533) );
  AND2_X1 U5097 ( .A1(n8525), .A2(n8281), .ZN(n4535) );
  NAND2_X1 U5098 ( .A1(n4381), .A2(n6511), .ZN(n4727) );
  INV_X1 U5099 ( .A(n4619), .ZN(n4618) );
  OAI21_X1 U5100 ( .B1(n4366), .B2(n4362), .A(n4395), .ZN(n4619) );
  AND2_X1 U5101 ( .A1(n4710), .A2(n4712), .ZN(n4709) );
  INV_X1 U5102 ( .A(n8888), .ZN(n4710) );
  NOR2_X1 U5103 ( .A1(n4388), .A2(n4735), .ZN(n4734) );
  NOR2_X1 U5104 ( .A1(n4919), .A2(n4736), .ZN(n4735) );
  INV_X1 U5105 ( .A(n4764), .ZN(n4761) );
  NAND2_X1 U5106 ( .A1(n9850), .A2(n6421), .ZN(n4784) );
  NAND2_X1 U5107 ( .A1(n9878), .A2(n6934), .ZN(n7066) );
  NOR2_X1 U5108 ( .A1(n7079), .A2(n6067), .ZN(n7126) );
  OR2_X1 U5109 ( .A1(n8291), .A2(n8503), .ZN(n8293) );
  INV_X1 U5110 ( .A(n4598), .ZN(n4596) );
  AOI21_X1 U5111 ( .B1(n4599), .B2(n8501), .A(n4603), .ZN(n4598) );
  INV_X1 U5112 ( .A(n4600), .ZN(n4599) );
  INV_X1 U5113 ( .A(n8133), .ZN(n4633) );
  OR2_X1 U5114 ( .A1(n8774), .A2(n8504), .ZN(n8287) );
  OR2_X1 U5115 ( .A1(n7911), .A2(n6333), .ZN(n8274) );
  AND2_X1 U5116 ( .A1(n4859), .A2(n8259), .ZN(n4858) );
  OR2_X1 U5117 ( .A1(n8260), .A2(n4860), .ZN(n4859) );
  OR2_X1 U5118 ( .A1(n8735), .A2(n8614), .ZN(n8258) );
  OR2_X1 U5119 ( .A1(n8814), .A2(n8031), .ZN(n8251) );
  NOR2_X1 U5120 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5921) );
  NOR2_X1 U5121 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5920) );
  NOR2_X1 U5122 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5919) );
  OR2_X1 U5123 ( .A1(n7504), .A2(n9317), .ZN(n7633) );
  NOR2_X1 U5124 ( .A1(n5351), .A2(n4842), .ZN(n4841) );
  INV_X1 U5125 ( .A(n5323), .ZN(n4842) );
  AND2_X1 U5126 ( .A1(n4771), .A2(n4770), .ZN(n4769) );
  INV_X1 U5127 ( .A(n8028), .ZN(n4770) );
  OR2_X1 U5128 ( .A1(n4773), .A2(n4385), .ZN(n4771) );
  INV_X4 U5129 ( .A(n6712), .ZN(n7961) );
  AND2_X1 U5130 ( .A1(n8308), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5131 ( .A1(n8307), .A2(n8313), .ZN(n8308) );
  CLKBUF_X1 U5132 ( .A(n5974), .Z(n6157) );
  XNOR2_X1 U5133 ( .A(n6910), .B(n6930), .ZN(n9861) );
  XNOR2_X1 U5134 ( .A(n8420), .B(n8421), .ZN(n8398) );
  NAND2_X1 U5135 ( .A1(n8416), .A2(n8417), .ZN(n8434) );
  OR2_X1 U5136 ( .A1(n8438), .A2(n8745), .ZN(n4790) );
  OR2_X1 U5137 ( .A1(n6268), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U5138 ( .A1(n6224), .A2(n5947), .ZN(n6233) );
  AND2_X1 U5139 ( .A1(n6341), .A2(n6623), .ZN(n9919) );
  XNOR2_X1 U5140 ( .A(n8512), .B(n8153), .ZN(n8501) );
  OAI21_X1 U5141 ( .B1(n8526), .B2(n4601), .A(n4600), .ZN(n8502) );
  OR2_X1 U5142 ( .A1(n8050), .A2(n7947), .ZN(n8265) );
  INV_X1 U5143 ( .A(n5995), .ZN(n8115) );
  NAND2_X1 U5144 ( .A1(n8118), .A2(n6301), .ZN(n8671) );
  NAND2_X1 U5145 ( .A1(n6361), .A2(n6360), .ZN(n6387) );
  OR2_X1 U5146 ( .A1(n4365), .A2(n8847), .ZN(n6152) );
  NAND2_X1 U5147 ( .A1(n7658), .A2(n4818), .ZN(n4814) );
  INV_X1 U5148 ( .A(n5089), .ZN(n5794) );
  NAND2_X1 U5149 ( .A1(n9192), .A2(n5837), .ZN(n5839) );
  NAND2_X1 U5150 ( .A1(n9238), .A2(n4884), .ZN(n4883) );
  NOR2_X1 U5151 ( .A1(n9227), .A2(n4885), .ZN(n4884) );
  AOI21_X1 U5152 ( .B1(n4674), .B2(n4467), .A(n4445), .ZN(n4466) );
  INV_X1 U5153 ( .A(n4677), .ZN(n4467) );
  NAND2_X1 U5154 ( .A1(n9398), .A2(n8993), .ZN(n7774) );
  AND3_X1 U5155 ( .A1(n6395), .A2(n6479), .A3(P1_STATE_REG_SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U5156 ( .A(n4501), .B(n5436), .ZN(n6662) );
  NAND2_X1 U5157 ( .A1(n4834), .A2(n5435), .ZN(n4501) );
  INV_X1 U5158 ( .A(n8528), .ZN(n8504) );
  OR2_X1 U5159 ( .A1(n8360), .A2(n8361), .ZN(n4808) );
  INV_X1 U5160 ( .A(n8358), .ZN(n8359) );
  XNOR2_X1 U5161 ( .A(n8445), .B(n8460), .ZN(n8433) );
  INV_X1 U5162 ( .A(n8192), .ZN(n4556) );
  OR2_X1 U5163 ( .A1(n7603), .A2(n7660), .ZN(n4522) );
  NAND2_X1 U5164 ( .A1(n7607), .A2(n7654), .ZN(n4520) );
  OR2_X1 U5165 ( .A1(n7570), .A2(n7660), .ZN(n7597) );
  AOI21_X1 U5166 ( .B1(n4561), .B2(n8227), .A(n8226), .ZN(n4560) );
  OAI21_X1 U5167 ( .B1(n8223), .B2(n8222), .A(n4414), .ZN(n4561) );
  NAND2_X1 U5168 ( .A1(n4559), .A2(n4558), .ZN(n4557) );
  INV_X1 U5169 ( .A(n8230), .ZN(n4558) );
  INV_X1 U5170 ( .A(n8543), .ZN(n4534) );
  NAND2_X1 U5171 ( .A1(n8249), .A2(n8297), .ZN(n4542) );
  NOR2_X1 U5172 ( .A1(n4541), .A2(n8252), .ZN(n4540) );
  INV_X1 U5173 ( .A(n8255), .ZN(n4541) );
  NAND2_X1 U5174 ( .A1(n8255), .A2(n4407), .ZN(n4538) );
  NOR2_X1 U5175 ( .A1(n8254), .A2(n8290), .ZN(n4539) );
  NAND2_X1 U5176 ( .A1(n4529), .A2(n8289), .ZN(n8306) );
  NAND2_X1 U5177 ( .A1(n5980), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6438) );
  INV_X1 U5178 ( .A(n8789), .ZN(n6333) );
  OR2_X1 U5179 ( .A1(n7295), .A2(n4701), .ZN(n4700) );
  INV_X1 U5180 ( .A(n5347), .ZN(n4701) );
  NOR2_X1 U5181 ( .A1(n9245), .A2(n9386), .ZN(n4651) );
  INV_X1 U5182 ( .A(n5373), .ZN(n5375) );
  INV_X1 U5183 ( .A(n7909), .ZN(n4736) );
  NAND2_X1 U5184 ( .A1(n6677), .A2(n8310), .ZN(n6678) );
  NAND2_X1 U5185 ( .A1(n6675), .A2(n4921), .ZN(n6679) );
  AND2_X1 U5186 ( .A1(n4850), .A2(n4849), .ZN(n4848) );
  INV_X1 U5187 ( .A(n8298), .ZN(n4850) );
  NAND2_X1 U5188 ( .A1(n4422), .A2(n8763), .ZN(n4847) );
  NAND2_X1 U5189 ( .A1(n6434), .A2(n4801), .ZN(n9836) );
  NAND2_X1 U5190 ( .A1(n4350), .A2(n6435), .ZN(n6434) );
  OR2_X1 U5191 ( .A1(n4350), .A2(n6435), .ZN(n4801) );
  AND2_X1 U5192 ( .A1(n7384), .A2(n7383), .ZN(n7385) );
  NAND2_X1 U5193 ( .A1(n8343), .A2(n8342), .ZN(n8374) );
  INV_X1 U5194 ( .A(n8425), .ZN(n4780) );
  INV_X1 U5195 ( .A(n8398), .ZN(n4568) );
  INV_X1 U5196 ( .A(n6078), .ZN(n4622) );
  NOR2_X1 U5197 ( .A1(n6323), .A2(n4624), .ZN(n4623) );
  INV_X1 U5198 ( .A(n6066), .ZN(n4624) );
  NOR2_X1 U5199 ( .A1(n6012), .A2(n4638), .ZN(n4637) );
  INV_X1 U5200 ( .A(n5998), .ZN(n4638) );
  INV_X1 U5201 ( .A(n8310), .ZN(n8299) );
  OAI21_X1 U5202 ( .B1(n6358), .B2(n4381), .A(n4725), .ZN(n6672) );
  INV_X1 U5203 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5204 ( .B1(n7806), .B2(n4381), .A(n6511), .ZN(n4726) );
  AND2_X1 U5205 ( .A1(n8265), .A2(n8264), .ZN(n8575) );
  OR2_X1 U5206 ( .A1(n8802), .A2(n8570), .ZN(n8259) );
  AOI21_X1 U5207 ( .B1(n4618), .B2(n4362), .A(n4416), .ZN(n4617) );
  OR2_X1 U5208 ( .A1(n8749), .A2(n8094), .ZN(n8235) );
  NAND2_X1 U5209 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  INV_X1 U5210 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4983) );
  INV_X1 U5211 ( .A(n5531), .ZN(n4714) );
  AND2_X1 U5212 ( .A1(n4708), .A2(n4498), .ZN(n4497) );
  NAND2_X1 U5213 ( .A1(n4709), .A2(n5526), .ZN(n4498) );
  NAND2_X1 U5214 ( .A1(n9425), .A2(n9327), .ZN(n4694) );
  AND2_X1 U5215 ( .A1(n4694), .A2(n4692), .ZN(n4684) );
  NOR2_X1 U5216 ( .A1(n7504), .A2(n9118), .ZN(n4659) );
  NAND2_X1 U5217 ( .A1(n5882), .A2(n8900), .ZN(n7719) );
  NAND2_X1 U5218 ( .A1(n9187), .A2(n5880), .ZN(n7704) );
  NOR2_X1 U5219 ( .A1(n9285), .A2(n9280), .ZN(n9255) );
  OR2_X1 U5220 ( .A1(n8961), .A2(n7317), .ZN(n7574) );
  OR2_X1 U5221 ( .A1(n9788), .A2(n9741), .ZN(n7563) );
  INV_X1 U5222 ( .A(n5866), .ZN(n4891) );
  OR2_X1 U5223 ( .A1(n5089), .A2(n9029), .ZN(n5008) );
  OAI21_X1 U5224 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(n7524) );
  OR2_X1 U5225 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  XNOR2_X1 U5226 ( .A(n7514), .B(n7513), .ZN(n7517) );
  NAND2_X1 U5227 ( .A1(n4963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4957) );
  AND2_X1 U5228 ( .A1(n4723), .A2(n4426), .ZN(n4722) );
  AND2_X1 U5229 ( .A1(n4911), .A2(n5435), .ZN(n4833) );
  INV_X1 U5230 ( .A(SI_12_), .ZN(n5325) );
  INV_X1 U5231 ( .A(n5321), .ZN(n4526) );
  AOI21_X1 U5232 ( .B1(n4924), .B2(n4831), .A(n4830), .ZN(n4829) );
  INV_X1 U5233 ( .A(n5237), .ZN(n4831) );
  INV_X1 U5234 ( .A(n5266), .ZN(n4830) );
  INV_X1 U5235 ( .A(n4924), .ZN(n4832) );
  INV_X1 U5236 ( .A(SI_10_), .ZN(n5268) );
  AOI21_X1 U5237 ( .B1(n7924), .B2(n4755), .A(n7959), .ZN(n4754) );
  INV_X1 U5238 ( .A(n8075), .ZN(n4755) );
  INV_X1 U5239 ( .A(n4754), .ZN(n4752) );
  INV_X1 U5240 ( .A(n8686), .ZN(n8680) );
  AND2_X1 U5241 ( .A1(n4765), .A2(n4766), .ZN(n4764) );
  NAND2_X1 U5242 ( .A1(n6980), .A2(n6833), .ZN(n4765) );
  NAND2_X1 U5243 ( .A1(n4774), .A2(n4446), .ZN(n4773) );
  NAND2_X1 U5244 ( .A1(n7952), .A2(n4775), .ZN(n4774) );
  INV_X1 U5245 ( .A(n7900), .ZN(n4775) );
  AND2_X1 U5246 ( .A1(n7880), .A2(n7879), .ZN(n7881) );
  AND3_X1 U5247 ( .A1(n6245), .A2(n6244), .A3(n6243), .ZN(n7911) );
  OR2_X1 U5248 ( .A1(n6308), .A2(n6016), .ZN(n6017) );
  NAND2_X1 U5249 ( .A1(n4781), .A2(n4783), .ZN(n4782) );
  NOR2_X1 U5250 ( .A1(n9847), .A2(n4408), .ZN(n6534) );
  NAND2_X1 U5251 ( .A1(n4784), .A2(n6536), .ZN(n6423) );
  NAND3_X1 U5252 ( .A1(n4782), .A2(P2_REG1_REG_3__SCAN_IN), .A3(n6423), .ZN(
        n6544) );
  XNOR2_X1 U5253 ( .A(n6931), .B(n6930), .ZN(n9863) );
  NOR2_X1 U5254 ( .A1(n9860), .A2(n6911), .ZN(n9883) );
  NOR2_X1 U5255 ( .A1(n9856), .A2(n6921), .ZN(n9875) );
  NAND2_X1 U5256 ( .A1(n9875), .A2(n9876), .ZN(n9874) );
  XNOR2_X1 U5257 ( .A(n7066), .B(n7060), .ZN(n6935) );
  INV_X1 U5258 ( .A(n7066), .ZN(n7067) );
  NOR2_X1 U5259 ( .A1(n6935), .A2(n7184), .ZN(n7069) );
  INV_X1 U5260 ( .A(n9904), .ZN(n7070) );
  INV_X1 U5261 ( .A(n4569), .ZN(n7073) );
  INV_X1 U5262 ( .A(n7128), .ZN(n4562) );
  OAI21_X1 U5263 ( .B1(n7115), .B2(n4491), .A(n4490), .ZN(n7418) );
  NAND2_X1 U5264 ( .A1(n4492), .A2(n7370), .ZN(n4490) );
  NAND2_X1 U5265 ( .A1(n4493), .A2(n4492), .ZN(n4491) );
  INV_X1 U5266 ( .A(n7420), .ZN(n4492) );
  NOR2_X1 U5267 ( .A1(n8362), .A2(n8421), .ZN(n4581) );
  NAND2_X1 U5268 ( .A1(n8362), .A2(n4584), .ZN(n4582) );
  OR2_X1 U5269 ( .A1(n8421), .A2(n4805), .ZN(n4585) );
  AND2_X1 U5270 ( .A1(n8421), .A2(n4805), .ZN(n4584) );
  NAND2_X1 U5271 ( .A1(n8414), .A2(n8415), .ZN(n8416) );
  OR2_X1 U5272 ( .A1(n8145), .A2(n8144), .ZN(n8525) );
  NAND2_X1 U5273 ( .A1(n7236), .A2(n4623), .ZN(n7324) );
  OR2_X1 U5274 ( .A1(n8331), .A2(n9962), .ZN(n8199) );
  NAND2_X1 U5275 ( .A1(n7174), .A2(n8192), .ZN(n4845) );
  AND2_X1 U5276 ( .A1(n8310), .A2(n8472), .ZN(n6844) );
  OR2_X1 U5277 ( .A1(n5989), .A2(n5960), .ZN(n5965) );
  NAND2_X1 U5278 ( .A1(n6386), .A2(n8297), .ZN(n6774) );
  AOI21_X1 U5279 ( .B1(n4854), .B2(n8283), .A(n4852), .ZN(n4851) );
  INV_X1 U5280 ( .A(n8287), .ZN(n4852) );
  OR2_X1 U5281 ( .A1(n8784), .A2(n8326), .ZN(n6254) );
  INV_X1 U5282 ( .A(n6238), .ZN(n4611) );
  OR2_X1 U5283 ( .A1(n8795), .A2(n8327), .ZN(n4609) );
  OR2_X1 U5284 ( .A1(n4614), .A2(n6238), .ZN(n4610) );
  INV_X1 U5285 ( .A(n8687), .ZN(n9922) );
  AOI21_X1 U5286 ( .B1(n8588), .B2(n8567), .A(n8575), .ZN(n8569) );
  OR2_X1 U5287 ( .A1(n8271), .A2(n8141), .ZN(n8560) );
  INV_X1 U5288 ( .A(n8258), .ZN(n4863) );
  NOR2_X1 U5289 ( .A1(n8252), .A2(n8119), .ZN(n4865) );
  NAND2_X1 U5290 ( .A1(n6312), .A2(n8290), .ZN(n9920) );
  NAND2_X1 U5291 ( .A1(n6329), .A2(n4867), .ZN(n4866) );
  NOR2_X1 U5292 ( .A1(n8242), .A2(n4868), .ZN(n4867) );
  INV_X1 U5293 ( .A(n8245), .ZN(n4868) );
  OR2_X1 U5294 ( .A1(n8826), .A2(n8650), .ZN(n8245) );
  OR2_X1 U5295 ( .A1(n8757), .A2(n8659), .ZN(n4627) );
  AND2_X1 U5296 ( .A1(n6685), .A2(n8290), .ZN(n8687) );
  INV_X1 U5297 ( .A(n9920), .ZN(n8684) );
  NOR2_X1 U5298 ( .A1(n6625), .A2(n8843), .ZN(n6631) );
  NOR2_X1 U5299 ( .A1(n6617), .A2(n6379), .ZN(n6636) );
  NAND2_X1 U5300 ( .A1(n4729), .A2(n6359), .ZN(n6477) );
  AND2_X1 U5301 ( .A1(n6619), .A2(n6513), .ZN(n6637) );
  NOR2_X1 U5302 ( .A1(n4871), .A2(n4413), .ZN(n4870) );
  INV_X1 U5303 ( .A(n4871), .ZN(n4482) );
  AND2_X1 U5304 ( .A1(n4872), .A2(n5931), .ZN(n4479) );
  AND2_X1 U5305 ( .A1(n5924), .A2(n4756), .ZN(n4480) );
  INV_X1 U5306 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6352) );
  INV_X1 U5307 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U5308 ( .A1(n6351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U5309 ( .A1(n6296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  NOR2_X1 U5310 ( .A1(n4374), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4544) );
  OR2_X1 U5311 ( .A1(n6294), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6296) );
  AND2_X1 U5312 ( .A1(n5915), .A2(n5981), .ZN(n4759) );
  NAND2_X1 U5313 ( .A1(n4957), .A2(n4956), .ZN(n5741) );
  OR2_X1 U5314 ( .A1(n5683), .A2(n5682), .ZN(n5763) );
  NAND2_X1 U5315 ( .A1(n5493), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U5316 ( .A1(n5414), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5441) );
  INV_X1 U5317 ( .A(n8905), .ZN(n4720) );
  INV_X1 U5318 ( .A(n8990), .ZN(n4721) );
  OR2_X1 U5319 ( .A1(n5610), .A2(n5609), .ZN(n5635) );
  INV_X1 U5320 ( .A(n8940), .ZN(n4706) );
  INV_X1 U5321 ( .A(n8921), .ZN(n4704) );
  INV_X1 U5322 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5358) );
  OR2_X1 U5323 ( .A1(n5333), .A2(n5332), .ZN(n5359) );
  OAI21_X1 U5324 ( .B1(n4696), .B2(n7745), .A(n5003), .ZN(n5004) );
  AND2_X1 U5325 ( .A1(n4959), .A2(n7746), .ZN(n7735) );
  AND2_X1 U5326 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  NAND2_X1 U5327 ( .A1(n9421), .A2(n7654), .ZN(n7656) );
  INV_X1 U5328 ( .A(n5025), .ZN(n5518) );
  INV_X1 U5329 ( .A(n5058), .ZN(n5888) );
  AND2_X1 U5330 ( .A1(n7633), .A2(n7638), .ZN(n7694) );
  AND2_X1 U5331 ( .A1(n7694), .A2(n4881), .ZN(n4880) );
  NAND2_X1 U5332 ( .A1(n7693), .A2(n7636), .ZN(n4881) );
  NAND2_X1 U5333 ( .A1(n9110), .A2(n7636), .ZN(n4876) );
  NOR2_X1 U5334 ( .A1(n9127), .A2(n9146), .ZN(n9126) );
  NOR2_X1 U5335 ( .A1(n7708), .A2(n4904), .ZN(n4903) );
  INV_X1 U5336 ( .A(n7705), .ZN(n4904) );
  AND2_X1 U5337 ( .A1(n7620), .A2(n7704), .ZN(n9173) );
  INV_X1 U5338 ( .A(n9210), .ZN(n4472) );
  AND2_X1 U5339 ( .A1(n9209), .A2(n7608), .ZN(n4882) );
  NAND2_X1 U5340 ( .A1(n4469), .A2(n4468), .ZN(n9228) );
  OR2_X1 U5341 ( .A1(n9245), .A2(n9265), .ZN(n4468) );
  NAND2_X1 U5342 ( .A1(n4465), .A2(n4464), .ZN(n4469) );
  AND2_X1 U5343 ( .A1(n4466), .A2(n4436), .ZN(n4464) );
  AND2_X1 U5344 ( .A1(n7777), .A2(n7782), .ZN(n9240) );
  NAND2_X1 U5345 ( .A1(n9298), .A2(n4898), .ZN(n4897) );
  NOR2_X1 U5346 ( .A1(n7689), .A2(n4899), .ZN(n4898) );
  INV_X1 U5347 ( .A(n7774), .ZN(n4899) );
  NOR2_X1 U5348 ( .A1(n5833), .A2(n4678), .ZN(n4677) );
  INV_X1 U5349 ( .A(n5830), .ZN(n4678) );
  AND2_X1 U5350 ( .A1(n7776), .A2(n7599), .ZN(n9263) );
  NAND2_X1 U5351 ( .A1(n7438), .A2(n7764), .ZN(n9299) );
  OR2_X1 U5352 ( .A1(n9807), .A2(n7400), .ZN(n7575) );
  OR2_X1 U5353 ( .A1(n7208), .A2(n9807), .ZN(n7285) );
  AOI21_X1 U5354 ( .B1(n4663), .B2(n4665), .A(n4411), .ZN(n4661) );
  OR2_X1 U5355 ( .A1(n5301), .A2(n5300), .ZN(n5303) );
  NAND2_X1 U5356 ( .A1(n5281), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5333) );
  INV_X1 U5357 ( .A(n5303), .ZN(n5281) );
  INV_X1 U5358 ( .A(n5871), .ZN(n4896) );
  NAND2_X1 U5359 ( .A1(n6896), .A2(n5821), .ZN(n9736) );
  OR2_X1 U5360 ( .A1(n7536), .A2(n7537), .ZN(n7543) );
  OR2_X1 U5361 ( .A1(n6804), .A2(n9770), .ZN(n6822) );
  OR2_X1 U5362 ( .A1(n5811), .A2(n6579), .ZN(n5812) );
  NOR2_X1 U5363 ( .A1(n6579), .A2(n6556), .ZN(n6589) );
  XNOR2_X1 U5364 ( .A(n5814), .B(n5813), .ZN(n6587) );
  OR2_X1 U5365 ( .A1(n6519), .A2(n4909), .ZN(n9291) );
  NAND2_X1 U5366 ( .A1(n4987), .A2(n7525), .ZN(n4646) );
  NAND2_X1 U5367 ( .A1(n5064), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4645) );
  INV_X1 U5368 ( .A(n5040), .ZN(n4500) );
  AND2_X1 U5369 ( .A1(n5769), .A2(n5768), .ZN(n9317) );
  AND2_X1 U5370 ( .A1(n6749), .A2(n5856), .ZN(n9806) );
  INV_X1 U5371 ( .A(n9738), .ZN(n9796) );
  INV_X1 U5372 ( .A(n9746), .ZN(n9331) );
  AND2_X1 U5373 ( .A1(n5729), .A2(n7451), .ZN(n6485) );
  NOR2_X1 U5374 ( .A1(n4673), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4671) );
  INV_X1 U5375 ( .A(n5182), .ZN(n4672) );
  XNOR2_X1 U5376 ( .A(n5781), .B(n5780), .ZN(n7480) );
  NAND2_X1 U5377 ( .A1(n4420), .A2(n4527), .ZN(n5322) );
  AND2_X1 U5378 ( .A1(n4443), .A2(n4824), .ZN(n4823) );
  AND3_X1 U5379 ( .A1(n5953), .A2(n5952), .A3(n5951), .ZN(n7947) );
  AND4_X1 U5380 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n7458)
         );
  AND4_X1 U5381 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n8614)
         );
  AOI21_X1 U5382 ( .B1(n4744), .B2(n4743), .A(n4447), .ZN(n4742) );
  AND3_X1 U5383 ( .A1(n6237), .A2(n6236), .A3(n6235), .ZN(n8571) );
  NAND2_X1 U5384 ( .A1(n5936), .A2(n5935), .ZN(n8050) );
  INV_X1 U5385 ( .A(n8093), .ZN(n8066) );
  INV_X1 U5386 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5929) );
  AND2_X1 U5387 ( .A1(n8113), .A2(n6291), .ZN(n8503) );
  NAND2_X1 U5388 ( .A1(n6275), .A2(n6274), .ZN(n8528) );
  INV_X1 U5389 ( .A(n7911), .ZN(n8561) );
  INV_X1 U5390 ( .A(n7947), .ZN(n8590) );
  INV_X1 U5391 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U5392 ( .A1(n4565), .A2(n6422), .ZN(n6909) );
  NAND2_X1 U5393 ( .A1(n6423), .A2(n6544), .ZN(n4565) );
  NOR2_X1 U5394 ( .A1(n7115), .A2(n7114), .ZN(n7369) );
  INV_X1 U5395 ( .A(n4806), .ZN(n8389) );
  OR2_X1 U5396 ( .A1(n8408), .A2(n8409), .ZN(n4804) );
  INV_X1 U5397 ( .A(n8423), .ZN(n4778) );
  AND2_X1 U5398 ( .A1(n4804), .A2(n4803), .ZN(n8432) );
  INV_X1 U5399 ( .A(n8410), .ZN(n4803) );
  NAND2_X1 U5400 ( .A1(n8442), .A2(n6411), .ZN(n4573) );
  NOR2_X1 U5401 ( .A1(n8441), .A2(n4572), .ZN(n4571) );
  NOR2_X1 U5402 ( .A1(n9841), .A2(n8439), .ZN(n4572) );
  NOR2_X1 U5403 ( .A1(n8433), .A2(n8638), .ZN(n8446) );
  NAND2_X1 U5404 ( .A1(n4790), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U5405 ( .A1(n8438), .A2(n8745), .ZN(n4575) );
  NAND2_X1 U5406 ( .A1(n4785), .A2(n4787), .ZN(n8485) );
  NAND2_X1 U5407 ( .A1(n4593), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5408 ( .A1(n8447), .A2(n4593), .ZN(n4591) );
  INV_X1 U5409 ( .A(n8448), .ZN(n4593) );
  NAND2_X1 U5410 ( .A1(n4485), .A2(n8476), .ZN(n4484) );
  NAND2_X1 U5411 ( .A1(n4486), .A2(n9871), .ZN(n4485) );
  NAND2_X1 U5412 ( .A1(n8457), .A2(P2_U3893), .ZN(n4486) );
  INV_X1 U5413 ( .A(n4488), .ZN(n4487) );
  OAI21_X1 U5414 ( .B1(n8457), .B2(n4379), .A(n4489), .ZN(n4488) );
  AOI21_X1 U5415 ( .B1(n9900), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8458), .ZN(
        n4489) );
  NAND2_X1 U5416 ( .A1(n8490), .A2(n8489), .ZN(n4794) );
  INV_X1 U5417 ( .A(n4793), .ZN(n4586) );
  OAI21_X1 U5418 ( .B1(n4927), .B2(n9857), .A(n8491), .ZN(n4793) );
  NOR2_X1 U5419 ( .A1(n6280), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8492) );
  AOI21_X1 U5420 ( .B1(n6316), .B2(n8671), .A(n6315), .ZN(n6343) );
  NAND2_X1 U5421 ( .A1(n6279), .A2(n6278), .ZN(n8512) );
  NAND2_X1 U5422 ( .A1(n6215), .A2(n6214), .ZN(n8735) );
  NAND2_X1 U5423 ( .A1(n5439), .A2(n5438), .ZN(n9398) );
  NAND2_X1 U5424 ( .A1(n6662), .A2(n4352), .ZN(n5439) );
  INV_X1 U5425 ( .A(n9002), .ZN(n8971) );
  AND4_X1 U5426 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n8993)
         );
  NAND2_X1 U5427 ( .A1(n5669), .A2(n5668), .ZN(n9159) );
  OR2_X1 U5428 ( .A1(n9149), .A2(n5664), .ZN(n5669) );
  CLKBUF_X1 U5429 ( .A(n5897), .Z(n9090) );
  AOI21_X1 U5430 ( .B1(n4687), .B2(n4688), .A(n7693), .ZN(n4474) );
  NAND2_X1 U5431 ( .A1(n5776), .A2(n6554), .ZN(n9753) );
  AND2_X2 U5432 ( .A1(n5911), .A2(n5910), .ZN(n9826) );
  NAND2_X1 U5433 ( .A1(n9816), .A2(n9806), .ZN(n9466) );
  INV_X1 U5434 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4945) );
  AOI21_X1 U5435 ( .B1(n7562), .B2(n7561), .A(n7560), .ZN(n7578) );
  INV_X1 U5436 ( .A(n7764), .ZN(n4515) );
  INV_X1 U5437 ( .A(n7765), .ZN(n4505) );
  OR2_X1 U5438 ( .A1(n7567), .A2(n7575), .ZN(n4511) );
  NOR2_X1 U5439 ( .A1(n7567), .A2(n4507), .ZN(n4506) );
  NOR2_X1 U5440 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  INV_X1 U5441 ( .A(n7582), .ZN(n4513) );
  NOR2_X1 U5442 ( .A1(n7572), .A2(n7654), .ZN(n7595) );
  NAND2_X1 U5443 ( .A1(n8197), .A2(n4409), .ZN(n4552) );
  NAND2_X1 U5444 ( .A1(n4521), .A2(n4406), .ZN(n4518) );
  NAND2_X1 U5445 ( .A1(n7605), .A2(n7660), .ZN(n4519) );
  NAND2_X1 U5446 ( .A1(n7717), .A2(n7660), .ZN(n7617) );
  OAI21_X1 U5447 ( .B1(n4560), .B2(n4557), .A(n8234), .ZN(n8240) );
  AOI22_X1 U5448 ( .A1(n8263), .A2(n8290), .B1(n4418), .B2(n4537), .ZN(n4536)
         );
  NAND2_X1 U5449 ( .A1(n4532), .A2(n4528), .ZN(n4530) );
  INV_X1 U5450 ( .A(n4532), .ZN(n4531) );
  AOI21_X1 U5451 ( .B1(n8451), .B2(n8452), .A(n4476), .ZN(n8454) );
  AND2_X1 U5452 ( .A1(n8450), .A2(n8460), .ZN(n4476) );
  NAND2_X1 U5453 ( .A1(n8336), .A2(n6994), .ZN(n8174) );
  NAND2_X1 U5454 ( .A1(n4863), .A2(n8256), .ZN(n4860) );
  NOR2_X1 U5455 ( .A1(n8260), .A2(n4862), .ZN(n4861) );
  INV_X1 U5456 ( .A(n8256), .ZN(n4862) );
  NOR2_X1 U5457 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5918) );
  INV_X1 U5458 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4821) );
  AOI21_X1 U5459 ( .B1(n4709), .B2(n4715), .A(n4396), .ZN(n4708) );
  NOR2_X1 U5460 ( .A1(n9234), .A2(n4650), .ZN(n4649) );
  INV_X1 U5461 ( .A(n4651), .ZN(n4650) );
  NAND2_X1 U5462 ( .A1(n5851), .A2(n5850), .ZN(n7514) );
  AOI21_X1 U5463 ( .B1(n5534), .B2(n5537), .A(SI_20_), .ZN(n4836) );
  INV_X1 U5464 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U5465 ( .A1(n4419), .A2(n5350), .ZN(n4840) );
  AND2_X1 U5466 ( .A1(n4829), .A2(n5293), .ZN(n4364) );
  INV_X1 U5467 ( .A(SI_11_), .ZN(n10099) );
  INV_X1 U5468 ( .A(SI_9_), .ZN(n10088) );
  INV_X1 U5469 ( .A(SI_26_), .ZN(n10090) );
  INV_X1 U5470 ( .A(n8313), .ZN(n4549) );
  NAND2_X1 U5471 ( .A1(n9836), .A2(n9835), .ZN(n9834) );
  OAI21_X1 U5472 ( .B1(n9836), .B2(n4800), .A(n4799), .ZN(n6443) );
  INV_X1 U5473 ( .A(n6439), .ZN(n4800) );
  AOI21_X1 U5474 ( .B1(n4798), .B2(n6439), .A(n4783), .ZN(n4799) );
  AND2_X1 U5475 ( .A1(n6928), .A2(n4812), .ZN(n6931) );
  NAND2_X1 U5476 ( .A1(n6929), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4812) );
  OAI211_X1 U5477 ( .C1(n6935), .C2(n4376), .A(n4590), .B(n4452), .ZN(n7116)
         );
  INV_X1 U5478 ( .A(n7114), .ZN(n4493) );
  NAND2_X1 U5479 ( .A1(n6174), .A2(n6173), .ZN(n6190) );
  OR2_X1 U5480 ( .A1(n9978), .A2(n8680), .ZN(n8211) );
  NAND2_X1 U5481 ( .A1(n7153), .A2(n4386), .ZN(n7177) );
  NOR2_X1 U5482 ( .A1(n4855), .A2(n8284), .ZN(n4854) );
  INV_X1 U5483 ( .A(n8288), .ZN(n4855) );
  AND2_X1 U5484 ( .A1(n8140), .A2(n8552), .ZN(n8272) );
  OR2_X1 U5485 ( .A1(n8784), .A2(n8549), .ZN(n8279) );
  NAND2_X1 U5486 ( .A1(n5931), .A2(n5927), .ZN(n5937) );
  INV_X1 U5487 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U5488 ( .A1(n5924), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U5489 ( .A1(n6298), .A2(n5925), .ZN(n6350) );
  NAND2_X1 U5490 ( .A1(n4365), .A2(n6169), .ZN(n6180) );
  INV_X1 U5491 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6169) );
  OR2_X1 U5492 ( .A1(n6117), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6118) );
  INV_X1 U5493 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5917) );
  AOI21_X1 U5494 ( .B1(n4369), .B2(n4701), .A(n4399), .ZN(n4697) );
  NOR2_X1 U5495 ( .A1(n9090), .A2(n4658), .ZN(n4657) );
  INV_X1 U5496 ( .A(n4659), .ZN(n4658) );
  INV_X1 U5497 ( .A(n5838), .ZN(n4680) );
  NOR2_X1 U5498 ( .A1(n9203), .A2(n9218), .ZN(n9182) );
  OR2_X1 U5499 ( .A1(n9398), .A2(n8993), .ZN(n7770) );
  NAND2_X1 U5500 ( .A1(n4655), .A2(n9467), .ZN(n4654) );
  INV_X1 U5501 ( .A(n4656), .ZN(n4655) );
  OR2_X1 U5502 ( .A1(n7344), .A2(n7433), .ZN(n4656) );
  INV_X1 U5503 ( .A(n4664), .ZN(n4663) );
  OAI21_X1 U5504 ( .B1(n7679), .B2(n4665), .A(n7201), .ZN(n4664) );
  INV_X1 U5505 ( .A(n5823), .ZN(n4665) );
  OR2_X1 U5506 ( .A1(n7678), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U5507 ( .A1(n6882), .A2(n7674), .ZN(n6898) );
  OR2_X1 U5508 ( .A1(n4361), .A2(n7812), .ZN(n5001) );
  NAND2_X1 U5509 ( .A1(n9255), .A2(n4647), .ZN(n9218) );
  NOR2_X1 U5510 ( .A1(n4648), .A2(n9222), .ZN(n4647) );
  INV_X1 U5511 ( .A(n4649), .ZN(n4648) );
  NAND2_X1 U5512 ( .A1(n9255), .A2(n4649), .ZN(n9231) );
  CLKBUF_X1 U5513 ( .A(n5748), .Z(n5856) );
  NAND2_X1 U5514 ( .A1(n5679), .A2(n5678), .ZN(n5704) );
  OAI21_X1 U5515 ( .B1(n5584), .B2(n5583), .A(n5582), .ZN(n5600) );
  INV_X1 U5516 ( .A(n5580), .ZN(n5581) );
  INV_X1 U5517 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4954) );
  INV_X1 U5518 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4942) );
  INV_X1 U5519 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4943) );
  NOR2_X1 U5520 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4723) );
  NAND2_X1 U5521 ( .A1(n5433), .A2(n5432), .ZN(n4834) );
  NAND2_X1 U5522 ( .A1(n4364), .A2(n5235), .ZN(n4525) );
  NAND2_X1 U5523 ( .A1(n5177), .A2(n4826), .ZN(n4824) );
  INV_X1 U5524 ( .A(n5165), .ZN(n4826) );
  NAND2_X1 U5525 ( .A1(n5267), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5106) );
  INV_X1 U5526 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5066) );
  INV_X1 U5527 ( .A(SI_28_), .ZN(n10201) );
  INV_X1 U5528 ( .A(SI_21_), .ZN(n10199) );
  INV_X1 U5529 ( .A(SI_13_), .ZN(n10210) );
  INV_X1 U5530 ( .A(SI_15_), .ZN(n10188) );
  INV_X1 U5531 ( .A(SI_24_), .ZN(n10184) );
  INV_X1 U5532 ( .A(SI_22_), .ZN(n10123) );
  INV_X1 U5533 ( .A(SI_25_), .ZN(n10114) );
  NAND2_X1 U5534 ( .A1(n7908), .A2(n4919), .ZN(n4733) );
  NAND2_X1 U5535 ( .A1(n6069), .A2(n6068), .ZN(n6087) );
  INV_X1 U5536 ( .A(n4929), .ZN(n4743) );
  NOR2_X1 U5537 ( .A1(n6146), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U5538 ( .A1(n4732), .A2(n4730), .ZN(n8020) );
  AND2_X1 U5539 ( .A1(n7914), .A2(n4731), .ZN(n4730) );
  NAND2_X1 U5540 ( .A1(n4734), .A2(n4736), .ZN(n4731) );
  XNOR2_X1 U5541 ( .A(n7961), .B(n9930), .ZN(n6734) );
  NAND2_X1 U5542 ( .A1(n4370), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5543 ( .A1(n4746), .A2(n4929), .ZN(n4745) );
  INV_X1 U5544 ( .A(n7931), .ZN(n4746) );
  INV_X1 U5545 ( .A(n4846), .ZN(n4551) );
  OAI21_X1 U5546 ( .B1(n8303), .B2(n8302), .A(n8307), .ZN(n4550) );
  NAND2_X1 U5547 ( .A1(n5980), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U5548 ( .A1(n6572), .A2(n6405), .ZN(n9845) );
  AND2_X1 U5549 ( .A1(n9845), .A2(n9844), .ZN(n9847) );
  OR2_X1 U5550 ( .A1(n6539), .A2(n6401), .ZN(n6537) );
  NOR2_X1 U5551 ( .A1(n9863), .A2(n6016), .ZN(n9862) );
  OR2_X1 U5552 ( .A1(n9880), .A2(n9881), .ZN(n9878) );
  NAND2_X1 U5553 ( .A1(n9874), .A2(n6922), .ZN(n6924) );
  NAND2_X1 U5554 ( .A1(n6924), .A2(n6923), .ZN(n7062) );
  INV_X1 U5555 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7255) );
  XNOR2_X1 U5556 ( .A(n7116), .B(n7078), .ZN(n7071) );
  NOR2_X1 U5557 ( .A1(n7071), .A2(n7327), .ZN(n7118) );
  NAND2_X1 U5558 ( .A1(n4579), .A2(n4578), .ZN(n7384) );
  INV_X1 U5559 ( .A(n7366), .ZN(n4791) );
  NAND2_X1 U5560 ( .A1(n4810), .A2(n4809), .ZN(n8347) );
  INV_X1 U5561 ( .A(n4576), .ZN(n4810) );
  OR2_X1 U5562 ( .A1(n7414), .A2(n7368), .ZN(n4811) );
  XNOR2_X1 U5563 ( .A(n8358), .B(n8364), .ZN(n8348) );
  NOR2_X1 U5564 ( .A1(n7418), .A2(n7373), .ZN(n8339) );
  NAND2_X1 U5565 ( .A1(n8347), .A2(n8346), .ZN(n8358) );
  INV_X1 U5566 ( .A(n4779), .ZN(n8422) );
  NAND2_X1 U5567 ( .A1(n8397), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U5568 ( .A1(n4777), .A2(n4567), .ZN(n8436) );
  NAND2_X1 U5569 ( .A1(n8423), .A2(n4780), .ZN(n4777) );
  NAND2_X1 U5570 ( .A1(n4568), .A2(n4380), .ZN(n4567) );
  OR2_X1 U5571 ( .A1(n8398), .A2(n8752), .ZN(n4779) );
  NAND2_X1 U5572 ( .A1(n8434), .A2(n4477), .ZN(n8451) );
  NAND2_X1 U5573 ( .A1(n4478), .A2(n8424), .ZN(n4477) );
  INV_X1 U5574 ( .A(n8435), .ZN(n4478) );
  OR2_X1 U5575 ( .A1(n8463), .A2(n8745), .ZN(n4788) );
  INV_X1 U5576 ( .A(n8463), .ZN(n4786) );
  AOI21_X1 U5577 ( .B1(n4597), .B2(n4371), .A(n4596), .ZN(n6292) );
  NOR2_X1 U5578 ( .A1(n6249), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6258) );
  AND2_X1 U5579 ( .A1(n6332), .A2(n8265), .ZN(n4864) );
  OR2_X1 U5580 ( .A1(n6233), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6241) );
  AND4_X1 U5581 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n8570)
         );
  AND2_X1 U5582 ( .A1(n6222), .A2(n5946), .ZN(n6224) );
  NOR2_X1 U5583 ( .A1(n6207), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6222) );
  INV_X1 U5584 ( .A(n8132), .ZN(n4629) );
  INV_X1 U5585 ( .A(n6115), .ZN(n4630) );
  INV_X1 U5586 ( .A(n4632), .ZN(n4631) );
  INV_X1 U5587 ( .A(n8659), .ZN(n9559) );
  INV_X1 U5588 ( .A(n8222), .ZN(n8691) );
  OR2_X1 U5589 ( .A1(n6087), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6097) );
  OR2_X1 U5590 ( .A1(n6097), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6108) );
  OAI21_X1 U5591 ( .B1(n7236), .B2(n4622), .A(n4620), .ZN(n6093) );
  INV_X1 U5592 ( .A(n4621), .ZN(n4620) );
  OAI21_X1 U5593 ( .B1(n4623), .B2(n4622), .A(n7347), .ZN(n4621) );
  NOR2_X1 U5594 ( .A1(n8127), .A2(n4844), .ZN(n4843) );
  INV_X1 U5595 ( .A(n8199), .ZN(n4844) );
  AND2_X1 U5596 ( .A1(n8199), .A2(n8194), .ZN(n7243) );
  INV_X1 U5597 ( .A(n7243), .ZN(n6063) );
  NOR2_X1 U5598 ( .A1(n6038), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6052) );
  AND4_X1 U5599 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n7194)
         );
  AOI21_X1 U5600 ( .B1(n4636), .B2(n4635), .A(n4417), .ZN(n7155) );
  AND2_X1 U5601 ( .A1(n4433), .A2(n6011), .ZN(n4635) );
  OR2_X1 U5602 ( .A1(n6026), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6038) );
  INV_X1 U5603 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U5604 ( .A1(n4636), .A2(n6011), .ZN(n7024) );
  NAND2_X1 U5605 ( .A1(n7028), .A2(n8124), .ZN(n7150) );
  NAND2_X1 U5606 ( .A1(n5999), .A2(n5998), .ZN(n7014) );
  NAND2_X1 U5607 ( .A1(n6608), .A2(n6788), .ZN(n6761) );
  NAND2_X1 U5608 ( .A1(n6286), .A2(n6285), .ZN(n8291) );
  INV_X1 U5609 ( .A(n8501), .ZN(n8500) );
  NAND2_X1 U5610 ( .A1(n4606), .A2(n4605), .ZN(n8537) );
  OR2_X1 U5611 ( .A1(n4607), .A2(n6246), .ZN(n4605) );
  AND2_X1 U5612 ( .A1(n4368), .A2(n4442), .ZN(n4607) );
  AND2_X1 U5613 ( .A1(n6232), .A2(n6231), .ZN(n7910) );
  NAND2_X1 U5614 ( .A1(n4616), .A2(n4617), .ZN(n8598) );
  NAND2_X1 U5615 ( .A1(n4616), .A2(n4394), .ZN(n8600) );
  INV_X1 U5616 ( .A(n8597), .ZN(n4615) );
  AND2_X1 U5617 ( .A1(n8258), .A2(n8256), .ZN(n8597) );
  AOI21_X1 U5618 ( .B1(n6168), .B2(n4366), .A(n4362), .ZN(n8612) );
  AND2_X1 U5619 ( .A1(n4869), .A2(n8251), .ZN(n8610) );
  OR2_X1 U5620 ( .A1(n8242), .A2(n8119), .ZN(n8625) );
  AND2_X1 U5621 ( .A1(n6168), .A2(n6167), .ZN(n8634) );
  AND2_X1 U5622 ( .A1(n8235), .A2(n8236), .ZN(n8646) );
  AND2_X1 U5623 ( .A1(n6080), .A2(n6079), .ZN(n6083) );
  INV_X1 U5624 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5916) );
  AND3_X1 U5625 ( .A1(n4759), .A2(n5980), .A3(n6007), .ZN(n6021) );
  OR2_X1 U5626 ( .A1(n7006), .A2(n7005), .ZN(n4475) );
  AND2_X1 U5627 ( .A1(n5702), .A2(n5701), .ZN(n5724) );
  INV_X1 U5628 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5220) );
  OR2_X1 U5629 ( .A1(n5221), .A2(n5220), .ZN(n5249) );
  AND2_X1 U5630 ( .A1(n4713), .A2(n5556), .ZN(n4712) );
  NAND2_X1 U5631 ( .A1(n4714), .A2(n5553), .ZN(n4713) );
  INV_X1 U5632 ( .A(n5553), .ZN(n4715) );
  INV_X1 U5633 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5332) );
  OR2_X1 U5634 ( .A1(n5441), .A2(n5440), .ZN(n5464) );
  OAI21_X1 U5635 ( .B1(n8939), .B2(n8943), .A(n8867), .ZN(n8922) );
  CLKBUF_X1 U5636 ( .A(n7140), .Z(n7141) );
  NAND2_X1 U5637 ( .A1(n5015), .A2(n4908), .ZN(n6552) );
  OR2_X1 U5638 ( .A1(n8876), .A2(n5526), .ZN(n5532) );
  NOR2_X1 U5639 ( .A1(n8941), .A2(n8940), .ZN(n8939) );
  NAND2_X1 U5640 ( .A1(n5565), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5610) );
  OR2_X1 U5641 ( .A1(n5515), .A2(n5514), .ZN(n5517) );
  NAND2_X1 U5642 ( .A1(n5462), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5515) );
  INV_X1 U5643 ( .A(n5464), .ZN(n5462) );
  NAND2_X1 U5644 ( .A1(n8989), .A2(n8990), .ZN(n8988) );
  NAND2_X1 U5645 ( .A1(n4503), .A2(n7652), .ZN(n7659) );
  AND2_X1 U5646 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  AND2_X1 U5647 ( .A1(n9417), .A2(n9076), .ZN(n7790) );
  AND2_X1 U5648 ( .A1(n9701), .A2(n7827), .ZN(n9706) );
  AND3_X1 U5649 ( .A1(n5891), .A2(n5890), .A3(n5889), .ZN(n7664) );
  AOI21_X1 U5650 ( .B1(n4880), .B2(n4878), .A(n7639), .ZN(n4877) );
  INV_X1 U5651 ( .A(n7636), .ZN(n4878) );
  NAND2_X1 U5652 ( .A1(n4683), .A2(n4694), .ZN(n4682) );
  INV_X1 U5653 ( .A(n4685), .ZN(n4683) );
  AND2_X1 U5654 ( .A1(n5793), .A2(n5764), .ZN(n9100) );
  NOR2_X1 U5655 ( .A1(n4690), .A2(n4689), .ZN(n4688) );
  NOR2_X1 U5656 ( .A1(n9429), .A2(n9316), .ZN(n4689) );
  NOR2_X1 U5657 ( .A1(n5844), .A2(n4691), .ZN(n4690) );
  NAND2_X1 U5658 ( .A1(n5843), .A2(n5842), .ZN(n4691) );
  NOR2_X1 U5659 ( .A1(n5844), .A2(n4693), .ZN(n4692) );
  INV_X1 U5660 ( .A(n5842), .ZN(n4693) );
  NOR2_X1 U5661 ( .A1(n9111), .A2(n4686), .ZN(n4685) );
  INV_X1 U5662 ( .A(n4688), .ZN(n4686) );
  OR2_X1 U5663 ( .A1(n7708), .A2(n7665), .ZN(n9143) );
  NAND2_X1 U5664 ( .A1(n9145), .A2(n5883), .ZN(n9146) );
  NAND2_X1 U5665 ( .A1(n5881), .A2(n7704), .ZN(n9156) );
  NOR2_X1 U5666 ( .A1(n9163), .A2(n4906), .ZN(n4905) );
  INV_X1 U5667 ( .A(n7704), .ZN(n4906) );
  NAND2_X1 U5668 ( .A1(n9255), .A2(n9261), .ZN(n9256) );
  INV_X1 U5669 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U5670 ( .B1(n5825), .B2(n4669), .A(n5827), .ZN(n4668) );
  NOR2_X1 U5671 ( .A1(n7686), .A2(n4887), .ZN(n4886) );
  INV_X1 U5672 ( .A(n7591), .ZN(n4887) );
  NAND2_X1 U5673 ( .A1(n4888), .A2(n7591), .ZN(n7436) );
  NAND2_X1 U5674 ( .A1(n5385), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5416) );
  OR2_X1 U5675 ( .A1(n5359), .A2(n5358), .ZN(n5387) );
  NOR2_X1 U5676 ( .A1(n7285), .A2(n7433), .ZN(n7341) );
  AND4_X1 U5677 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n8956)
         );
  AND2_X1 U5678 ( .A1(n4375), .A2(n7318), .ZN(n4640) );
  AND2_X1 U5679 ( .A1(n5873), .A2(n7049), .ZN(n4894) );
  NAND2_X1 U5680 ( .A1(n6901), .A2(n4367), .ZN(n9760) );
  NAND2_X1 U5681 ( .A1(n6901), .A2(n6970), .ZN(n9759) );
  AND4_X1 U5682 ( .A1(n5195), .A2(n5194), .A3(n5193), .A4(n5192), .ZN(n9739)
         );
  NOR2_X1 U5683 ( .A1(n6822), .A2(n7541), .ZN(n6890) );
  NAND2_X1 U5684 ( .A1(n6645), .A2(n5817), .ZN(n6793) );
  NAND2_X1 U5685 ( .A1(n4891), .A2(n7751), .ZN(n4890) );
  XNOR2_X1 U5686 ( .A(n6813), .B(n9012), .ZN(n7671) );
  NAND4_X1 U5687 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n5863)
         );
  NAND2_X1 U5688 ( .A1(n5413), .A2(n5412), .ZN(n7443) );
  NOR2_X1 U5689 ( .A1(n4916), .A2(n4907), .ZN(n5116) );
  NOR2_X1 U5690 ( .A1(n5907), .A2(n5906), .ZN(n5911) );
  INV_X1 U5691 ( .A(n9805), .ZN(n9740) );
  INV_X1 U5692 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4695) );
  INV_X1 U5693 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4993) );
  OAI21_X1 U5694 ( .B1(n7524), .B2(n7523), .A(n7522), .ZN(n7529) );
  XNOR2_X1 U5695 ( .A(n7524), .B(n7523), .ZN(n8101) );
  NAND2_X1 U5696 ( .A1(n4958), .A2(n5741), .ZN(n5747) );
  NAND2_X1 U5697 ( .A1(n4837), .A2(n5350), .ZN(n5374) );
  NAND2_X1 U5698 ( .A1(n5324), .A2(n4841), .ZN(n4837) );
  OR2_X1 U5699 ( .A1(n5295), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5326) );
  OAI21_X1 U5700 ( .B1(n5238), .B2(n4832), .A(n4829), .ZN(n5294) );
  INV_X1 U5701 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U5702 ( .A1(n7925), .A2(n7924), .ZN(n7960) );
  NAND2_X1 U5703 ( .A1(n4772), .A2(n7900), .ZN(n7951) );
  NAND2_X1 U5704 ( .A1(n8064), .A2(n8065), .ZN(n4772) );
  NOR2_X1 U5705 ( .A1(n7962), .A2(n4752), .ZN(n4749) );
  OAI22_X1 U5706 ( .A1(n4752), .A2(n4751), .B1(n7962), .B2(n4754), .ZN(n4750)
         );
  NOR2_X1 U5707 ( .A1(n7962), .A2(n7924), .ZN(n4751) );
  NAND2_X1 U5708 ( .A1(n7924), .A2(n7962), .ZN(n4753) );
  AOI21_X1 U5709 ( .B1(n4769), .B2(n4773), .A(n4451), .ZN(n4768) );
  INV_X1 U5710 ( .A(n8685), .ZN(n7981) );
  NAND2_X1 U5711 ( .A1(n6834), .A2(n6980), .ZN(n4763) );
  AND4_X1 U5712 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n8094)
         );
  NOR2_X1 U5713 ( .A1(n6834), .A2(n6833), .ZN(n6982) );
  INV_X1 U5714 ( .A(n8627), .ZN(n8031) );
  AOI21_X1 U5715 ( .B1(n8064), .B2(n4385), .A(n4773), .ZN(n8027) );
  INV_X1 U5716 ( .A(n8054), .ZN(n4738) );
  INV_X1 U5717 ( .A(n7881), .ZN(n4739) );
  INV_X1 U5718 ( .A(n8334), .ZN(n7044) );
  INV_X1 U5719 ( .A(n8091), .ZN(n8070) );
  AND2_X1 U5720 ( .A1(n6635), .A2(n6634), .ZN(n8082) );
  OR2_X1 U5721 ( .A1(n6629), .A2(n6685), .ZN(n8093) );
  NAND2_X1 U5722 ( .A1(n6639), .A2(n9553), .ZN(n8080) );
  INV_X1 U5723 ( .A(n8080), .ZN(n8099) );
  NAND2_X1 U5724 ( .A1(n4745), .A2(n4744), .ZN(n8087) );
  INV_X1 U5725 ( .A(n8082), .ZN(n8088) );
  XNOR2_X1 U5726 ( .A(n6300), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8319) );
  INV_X1 U5727 ( .A(n8153), .ZN(n8517) );
  NAND2_X1 U5728 ( .A1(n6264), .A2(n6263), .ZN(n8538) );
  INV_X1 U5729 ( .A(n8571), .ZN(n8327) );
  INV_X1 U5730 ( .A(n8614), .ZN(n8589) );
  INV_X1 U5731 ( .A(n7458), .ZN(n8330) );
  INV_X1 U5732 ( .A(n7194), .ZN(n8333) );
  INV_X1 U5733 ( .A(n9921), .ZN(n8336) );
  NAND2_X1 U5734 ( .A1(n6574), .A2(n6573), .ZN(n6572) );
  NAND2_X1 U5735 ( .A1(n4782), .A2(n6423), .ZN(n6542) );
  OR2_X1 U5736 ( .A1(n7069), .A2(n7068), .ZN(n9902) );
  NOR2_X1 U5737 ( .A1(n7076), .A2(n7075), .ZN(n9907) );
  INV_X1 U5738 ( .A(n4563), .ZN(n7129) );
  AND2_X1 U5739 ( .A1(n6431), .A2(n6430), .ZN(n9871) );
  NOR2_X1 U5740 ( .A1(n7369), .A2(n7370), .ZN(n7419) );
  INV_X1 U5741 ( .A(n4792), .ZN(n7367) );
  OAI211_X1 U5742 ( .C1(n4808), .C2(n4583), .A(n4459), .B(n4580), .ZN(n8390)
         );
  INV_X1 U5743 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5744 ( .A(n8474), .ZN(n4589) );
  OR2_X1 U5745 ( .A1(n6281), .A2(n8492), .ZN(n8511) );
  NAND2_X1 U5746 ( .A1(n6154), .A2(n6153), .ZN(n8749) );
  NAND2_X1 U5747 ( .A1(n6132), .A2(n6131), .ZN(n8757) );
  NAND2_X1 U5748 ( .A1(n7324), .A2(n6078), .ZN(n7350) );
  AND3_X1 U5749 ( .A1(n6050), .A2(n6049), .A3(n6048), .ZN(n9957) );
  NAND2_X1 U5750 ( .A1(n6787), .A2(n8673), .ZN(n8695) );
  INV_X1 U5751 ( .A(n9934), .ZN(n9553) );
  INV_X1 U5752 ( .A(n8667), .ZN(n8698) );
  INV_X1 U5753 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6435) );
  INV_X1 U5754 ( .A(n9562), .ZN(n9936) );
  INV_X1 U5755 ( .A(n8695), .ZN(n8664) );
  NAND2_X1 U5756 ( .A1(n10003), .A2(n9985), .ZN(n8736) );
  AND2_X1 U5757 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U5758 ( .A1(n7875), .A2(n6344), .ZN(n6345) );
  INV_X1 U5759 ( .A(n8291), .ZN(n7872) );
  OAI21_X1 U5760 ( .B1(n8508), .B2(n9928), .A(n8507), .ZN(n8767) );
  NOR2_X1 U5761 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  NOR2_X1 U5762 ( .A1(n8504), .A2(n9922), .ZN(n8505) );
  NAND2_X1 U5763 ( .A1(n6267), .A2(n6266), .ZN(n8774) );
  AND2_X1 U5764 ( .A1(n6240), .A2(n6239), .ZN(n8789) );
  NAND2_X1 U5765 ( .A1(n4608), .A2(n4368), .ZN(n8547) );
  NAND2_X1 U5766 ( .A1(n8569), .A2(n4611), .ZN(n4608) );
  INV_X1 U5767 ( .A(n7910), .ZN(n8795) );
  NOR2_X1 U5768 ( .A1(n8569), .A2(n4612), .ZN(n8559) );
  NAND2_X1 U5769 ( .A1(n8577), .A2(n8265), .ZN(n8558) );
  OR2_X1 U5770 ( .A1(n8731), .A2(n8730), .ZN(n8799) );
  NAND2_X1 U5771 ( .A1(n6221), .A2(n6220), .ZN(n8802) );
  OAI21_X1 U5772 ( .B1(n8596), .B2(n4863), .A(n8256), .ZN(n8583) );
  NAND2_X1 U5773 ( .A1(n6206), .A2(n6205), .ZN(n8814) );
  NAND2_X1 U5774 ( .A1(n6189), .A2(n6188), .ZN(n8820) );
  NAND2_X1 U5775 ( .A1(n6172), .A2(n6171), .ZN(n8826) );
  NAND2_X1 U5776 ( .A1(n6145), .A2(n6144), .ZN(n8837) );
  INV_X1 U5777 ( .A(n8807), .ZN(n8836) );
  INV_X1 U5778 ( .A(n7265), .ZN(n7492) );
  INV_X1 U5779 ( .A(n6387), .ZN(n8844) );
  AND2_X1 U5780 ( .A1(n6731), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6513) );
  INV_X1 U5781 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5938) );
  INV_X1 U5782 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U5783 ( .A1(n6346), .A2(n6349), .ZN(n7455) );
  NAND2_X1 U5784 ( .A1(n6357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6353) );
  INV_X1 U5785 ( .A(n8319), .ZN(n7235) );
  NAND2_X1 U5786 ( .A1(n6297), .A2(n6296), .ZN(n8310) );
  INV_X1 U5787 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6202) );
  INV_X1 U5788 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U5789 ( .A1(n4595), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5790 ( .A1(n5980), .A2(n5981), .ZN(n4595) );
  NAND2_X1 U5791 ( .A1(n4564), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5982) );
  INV_X1 U5792 ( .A(n5980), .ZN(n4564) );
  CLKBUF_X1 U5793 ( .A(n6437), .Z(n6568) );
  XNOR2_X1 U5794 ( .A(n5742), .B(n4961), .ZN(n6479) );
  NAND2_X1 U5795 ( .A1(n5491), .A2(n5490), .ZN(n9245) );
  NAND2_X1 U5796 ( .A1(n6277), .A2(n4352), .ZN(n5787) );
  NAND2_X1 U5797 ( .A1(n4711), .A2(n4712), .ZN(n8889) );
  OR2_X1 U5798 ( .A1(n5532), .A2(n4715), .ZN(n4711) );
  NAND2_X1 U5799 ( .A1(n8988), .A2(n5429), .ZN(n8906) );
  NAND2_X1 U5800 ( .A1(n8989), .A2(n4719), .ZN(n4718) );
  INV_X1 U5801 ( .A(n4717), .ZN(n4716) );
  NOR2_X1 U5802 ( .A1(n4720), .A2(n4721), .ZN(n4719) );
  OAI211_X1 U5803 ( .C1(n4705), .C2(n8941), .A(n4702), .B(n4703), .ZN(n8924)
         );
  NAND2_X1 U5804 ( .A1(n4707), .A2(n4704), .ZN(n4703) );
  NAND2_X1 U5805 ( .A1(n4707), .A2(n4393), .ZN(n4705) );
  NAND2_X1 U5806 ( .A1(n7304), .A2(n4352), .ZN(n4813) );
  NAND2_X1 U5807 ( .A1(n5532), .A2(n5531), .ZN(n8933) );
  XNOR2_X1 U5808 ( .A(n5370), .B(n5371), .ZN(n7399) );
  NAND2_X1 U5809 ( .A1(n7294), .A2(n7295), .ZN(n4699) );
  NAND2_X1 U5810 ( .A1(n5755), .A2(n7802), .ZN(n8980) );
  INV_X1 U5811 ( .A(n8975), .ZN(n8979) );
  AND2_X1 U5812 ( .A1(n5777), .A2(n9753), .ZN(n9002) );
  AND2_X1 U5813 ( .A1(n5774), .A2(n5749), .ZN(n8991) );
  NAND2_X1 U5814 ( .A1(n5616), .A2(n5615), .ZN(n9356) );
  INV_X1 U5815 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6508) );
  AND4_X1 U5816 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n7317)
         );
  INV_X1 U5817 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6504) );
  INV_X1 U5818 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6501) );
  AND4_X1 U5819 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n7536)
         );
  NAND2_X1 U5820 ( .A1(n4879), .A2(n7636), .ZN(n7501) );
  NAND2_X1 U5821 ( .A1(n4876), .A2(n4880), .ZN(n7500) );
  OR2_X1 U5822 ( .A1(n9110), .A2(n7693), .ZN(n4879) );
  OAI21_X1 U5823 ( .B1(n9144), .B2(n5843), .A(n5842), .ZN(n9122) );
  NAND2_X1 U5824 ( .A1(n5839), .A2(n5838), .ZN(n9174) );
  AND2_X1 U5825 ( .A1(n4883), .A2(n7608), .ZN(n9207) );
  NAND2_X1 U5826 ( .A1(n4465), .A2(n4466), .ZN(n9237) );
  AND2_X1 U5827 ( .A1(n4897), .A2(n7602), .ZN(n9264) );
  NAND2_X1 U5828 ( .A1(n4676), .A2(n5832), .ZN(n9254) );
  NAND2_X1 U5829 ( .A1(n5831), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5830 ( .A1(n9298), .A2(n7774), .ZN(n9270) );
  NAND2_X1 U5831 ( .A1(n5831), .A2(n5830), .ZN(n9274) );
  NAND2_X1 U5832 ( .A1(n5461), .A2(n5460), .ZN(n9285) );
  NAND2_X1 U5833 ( .A1(n7290), .A2(n7684), .ZN(n4670) );
  AND4_X1 U5834 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n7296)
         );
  NAND2_X1 U5835 ( .A1(n5331), .A2(n5330), .ZN(n9807) );
  NAND2_X1 U5836 ( .A1(n7051), .A2(n7679), .ZN(n4662) );
  AND4_X1 U5837 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n9741)
         );
  AND2_X1 U5838 ( .A1(n4473), .A2(n9733), .ZN(n7097) );
  INV_X1 U5839 ( .A(n9770), .ZN(n6806) );
  OR2_X1 U5840 ( .A1(n5088), .A2(n9034), .ZN(n5028) );
  OR2_X1 U5841 ( .A1(n5025), .A2(n7840), .ZN(n5026) );
  OR2_X1 U5842 ( .A1(n9295), .A2(n6748), .ZN(n9756) );
  NAND2_X1 U5843 ( .A1(n6747), .A2(n9753), .ZN(n9251) );
  INV_X1 U5844 ( .A(n9282), .ZN(n9764) );
  INV_X1 U5845 ( .A(n9756), .ZN(n9286) );
  INV_X1 U5846 ( .A(n9291), .ZN(n9761) );
  INV_X1 U5847 ( .A(n7544), .ZN(n7541) );
  NAND2_X1 U5848 ( .A1(n4500), .A2(n9018), .ZN(n4499) );
  NAND2_X1 U5849 ( .A1(n4646), .A2(n4645), .ZN(n4644) );
  AND2_X1 U5850 ( .A1(n9312), .A2(n9311), .ZN(n9418) );
  INV_X1 U5851 ( .A(n7504), .ZN(n9098) );
  NAND2_X1 U5852 ( .A1(n9315), .A2(n9812), .ZN(n9322) );
  INV_X1 U5853 ( .A(n9127), .ZN(n9429) );
  INV_X1 U5854 ( .A(n5882), .ZN(n9436) );
  INV_X1 U5855 ( .A(n9203), .ZN(n9444) );
  INV_X1 U5856 ( .A(n7443), .ZN(n9467) );
  NAND2_X1 U5857 ( .A1(n5279), .A2(n5278), .ZN(n8961) );
  NAND2_X1 U5858 ( .A1(n5039), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5046) );
  AND2_X2 U5859 ( .A1(n5911), .A2(n6745), .ZN(n9816) );
  NAND2_X1 U5860 ( .A1(n6486), .A2(n6554), .ZN(n9768) );
  INV_X1 U5861 ( .A(n7669), .ZN(n7746) );
  OR2_X1 U5862 ( .A1(n4949), .A2(n4948), .ZN(n4950) );
  NOR2_X1 U5863 ( .A1(n7525), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9479) );
  INV_X1 U5864 ( .A(n4808), .ZN(n8363) );
  INV_X1 U5865 ( .A(n4804), .ZN(n8411) );
  AOI21_X1 U5866 ( .B1(n4574), .B2(n8489), .A(n4570), .ZN(n8443) );
  NAND2_X1 U5867 ( .A1(n4573), .A2(n4571), .ZN(n4570) );
  AND2_X1 U5868 ( .A1(n4487), .A2(n4484), .ZN(n8466) );
  NAND2_X1 U5869 ( .A1(n4587), .A2(n4404), .ZN(P2_U3201) );
  NAND2_X1 U5870 ( .A1(n4588), .A2(n9838), .ZN(n4587) );
  XNOR2_X1 U5871 ( .A(n8471), .B(n4589), .ZN(n4588) );
  OR2_X1 U5872 ( .A1(n5898), .A2(n9406), .ZN(n4915) );
  OR2_X1 U5873 ( .A1(n5898), .A2(n9466), .ZN(n4914) );
  NOR2_X1 U5874 ( .A1(n6199), .A2(n6198), .ZN(n4362) );
  OR2_X1 U5875 ( .A1(n4848), .A2(n8118), .ZN(n4363) );
  INV_X2 U5876 ( .A(n5173), .ZN(n5310) );
  XNOR2_X1 U5877 ( .A(n6293), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U5878 ( .A1(n4483), .A2(n4756), .ZN(n6046) );
  AND2_X1 U5879 ( .A1(n4425), .A2(n4483), .ZN(n4365) );
  AND2_X1 U5880 ( .A1(n4745), .A2(n4747), .ZN(n7933) );
  AND2_X1 U5881 ( .A1(n6200), .A2(n6167), .ZN(n4366) );
  INV_X1 U5882 ( .A(n8763), .ZN(n4849) );
  AND2_X1 U5883 ( .A1(n6970), .A2(n4642), .ZN(n4367) );
  AND2_X1 U5884 ( .A1(n4610), .A2(n4609), .ZN(n4368) );
  AND2_X1 U5885 ( .A1(n4700), .A2(n7399), .ZN(n4369) );
  AND2_X1 U5886 ( .A1(n7038), .A2(n7037), .ZN(n4370) );
  AND2_X1 U5887 ( .A1(n4602), .A2(n8501), .ZN(n4371) );
  NAND3_X1 U5888 ( .A1(n4758), .A2(n4427), .A3(n5980), .ZN(n4372) );
  OR2_X1 U5889 ( .A1(n4847), .A2(n8118), .ZN(n4373) );
  OR2_X1 U5890 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4374) );
  AND2_X1 U5891 ( .A1(n4367), .A2(n4641), .ZN(n4375) );
  INV_X1 U5892 ( .A(n8145), .ZN(n4604) );
  BUF_X1 U5893 ( .A(n5489), .Z(n7662) );
  NAND2_X1 U5894 ( .A1(n7070), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4376) );
  AND2_X1 U5895 ( .A1(n4763), .A2(n4764), .ZN(n4377) );
  OR2_X1 U5896 ( .A1(n7285), .A2(n4656), .ZN(n4378) );
  OR2_X1 U5897 ( .A1(n9857), .A2(n8476), .ZN(n4379) );
  AND2_X1 U5898 ( .A1(n4780), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5899 ( .A1(n6359), .A2(n4728), .ZN(n4381) );
  NAND2_X1 U5900 ( .A1(n7563), .A2(n7573), .ZN(n4382) );
  AND2_X1 U5901 ( .A1(n5040), .A2(n5064), .ZN(n5039) );
  AND2_X1 U5902 ( .A1(n9238), .A2(n7782), .ZN(n4383) );
  AND2_X1 U5903 ( .A1(n4733), .A2(n7909), .ZN(n4384) );
  NAND4_X1 U5904 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n5986)
         );
  AND2_X1 U5905 ( .A1(n7952), .A2(n8065), .ZN(n4385) );
  INV_X1 U5906 ( .A(n6930), .ZN(n9870) );
  INV_X1 U5907 ( .A(n7782), .ZN(n4885) );
  AND2_X1 U5908 ( .A1(n8193), .A2(n6037), .ZN(n4386) );
  NAND2_X1 U5909 ( .A1(n4853), .A2(n4851), .ZN(n8499) );
  NAND2_X1 U5910 ( .A1(n5324), .A2(n5323), .ZN(n5352) );
  NAND2_X1 U5911 ( .A1(n4827), .A2(n5165), .ZN(n5178) );
  NAND2_X1 U5912 ( .A1(n5950), .A2(n8856), .ZN(n5961) );
  AND2_X1 U5913 ( .A1(n4828), .A2(n5270), .ZN(n4387) );
  AND2_X1 U5914 ( .A1(n7943), .A2(n8571), .ZN(n4388) );
  INV_X1 U5915 ( .A(n9084), .ZN(n9421) );
  AND2_X1 U5916 ( .A1(n5177), .A2(n5162), .ZN(n4389) );
  AND4_X1 U5917 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n4390)
         );
  OR2_X1 U5918 ( .A1(n5410), .A2(n4969), .ZN(n4391) );
  NAND2_X1 U5919 ( .A1(n5660), .A2(n5659), .ZN(n9148) );
  AND2_X1 U5920 ( .A1(n4687), .A2(n4685), .ZN(n4392) );
  NAND2_X1 U5921 ( .A1(n5540), .A2(n5539), .ZN(n9234) );
  AND2_X1 U5922 ( .A1(n8867), .A2(n4706), .ZN(n4393) );
  AND2_X1 U5923 ( .A1(n4617), .A2(n4615), .ZN(n4394) );
  OR2_X1 U5924 ( .A1(n8814), .A2(n8627), .ZN(n4395) );
  AND2_X1 U5925 ( .A1(n5579), .A2(n5578), .ZN(n4396) );
  NOR2_X1 U5926 ( .A1(n8446), .A2(n8447), .ZN(n4397) );
  NAND2_X1 U5927 ( .A1(n5513), .A2(n5512), .ZN(n9386) );
  INV_X1 U5928 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4981) );
  AND2_X1 U5929 ( .A1(n4382), .A2(n9733), .ZN(n4398) );
  AND2_X1 U5930 ( .A1(n5372), .A2(n5371), .ZN(n4399) );
  INV_X1 U5931 ( .A(n5826), .ZN(n4669) );
  NAND2_X1 U5932 ( .A1(n9222), .A2(n9355), .ZN(n4400) );
  OR2_X1 U5933 ( .A1(n7659), .A2(n7658), .ZN(n4401) );
  AND2_X1 U5934 ( .A1(n4779), .A2(n4778), .ZN(n4402) );
  OR2_X1 U5935 ( .A1(n8306), .A2(n8305), .ZN(n4403) );
  OAI21_X1 U5936 ( .B1(n8276), .B2(n8277), .A(n4534), .ZN(n4528) );
  AND2_X1 U5937 ( .A1(n4794), .A2(n4586), .ZN(n4404) );
  AND2_X1 U5938 ( .A1(n8774), .A2(n8528), .ZN(n4405) );
  AND2_X1 U5939 ( .A1(n4520), .A2(n4519), .ZN(n4406) );
  NAND2_X1 U5940 ( .A1(n8258), .A2(n8251), .ZN(n4407) );
  AND2_X1 U5941 ( .A1(n6407), .A2(n4350), .ZN(n4408) );
  AND2_X1 U5942 ( .A1(n4556), .A2(n8297), .ZN(n4409) );
  OR2_X1 U5943 ( .A1(n4360), .A2(n6568), .ZN(n4410) );
  NOR2_X1 U5944 ( .A1(n8961), .A2(n7298), .ZN(n4411) );
  AND2_X1 U5945 ( .A1(n8814), .A2(n8031), .ZN(n8252) );
  INV_X1 U5946 ( .A(n8252), .ZN(n4869) );
  AND2_X1 U5947 ( .A1(n9187), .A2(n9356), .ZN(n4412) );
  OR2_X1 U5948 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(n5937), .ZN(n4413) );
  INV_X1 U5949 ( .A(n4481), .ZN(n6347) );
  AND2_X1 U5950 ( .A1(n8220), .A2(n8221), .ZN(n4414) );
  AND2_X1 U5951 ( .A1(n7728), .A2(n7636), .ZN(n9111) );
  INV_X1 U5952 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4970) );
  INV_X1 U5953 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5925) );
  OR2_X1 U5954 ( .A1(n6392), .A2(n10004), .ZN(n4415) );
  INV_X1 U5955 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6181) );
  NOR2_X1 U5956 ( .A1(n6213), .A2(n8031), .ZN(n4416) );
  AND2_X1 U5957 ( .A1(n7044), .A2(n9948), .ZN(n4417) );
  AND2_X1 U5958 ( .A1(n4539), .A2(n4538), .ZN(n4418) );
  OR2_X1 U5959 ( .A1(n5375), .A2(n10210), .ZN(n4419) );
  AND2_X1 U5960 ( .A1(n4387), .A2(n4525), .ZN(n4420) );
  INV_X1 U5961 ( .A(n4602), .ZN(n4601) );
  AND2_X1 U5962 ( .A1(n4604), .A2(n6276), .ZN(n4602) );
  OR2_X1 U5963 ( .A1(n8763), .A2(n8494), .ZN(n4421) );
  NAND2_X1 U5964 ( .A1(n8766), .A2(n8315), .ZN(n4422) );
  AND2_X1 U5965 ( .A1(n4856), .A2(n8282), .ZN(n4423) );
  AND2_X1 U5966 ( .A1(n7684), .A2(n5826), .ZN(n4424) );
  AND2_X1 U5967 ( .A1(n4756), .A2(n4390), .ZN(n4425) );
  AND3_X1 U5968 ( .A1(n4943), .A2(n4942), .A3(n4941), .ZN(n4426) );
  AND3_X1 U5969 ( .A1(n4757), .A2(n5981), .A3(n5915), .ZN(n4427) );
  NAND2_X1 U5970 ( .A1(n5383), .A2(n5382), .ZN(n7344) );
  NAND2_X1 U5971 ( .A1(n9158), .A2(n7705), .ZN(n9138) );
  AND2_X1 U5972 ( .A1(n4707), .A2(n8867), .ZN(n4428) );
  AND2_X1 U5973 ( .A1(n4896), .A2(n7674), .ZN(n4429) );
  NOR2_X1 U5974 ( .A1(n4885), .A2(n4522), .ZN(n4430) );
  AND2_X1 U5975 ( .A1(n4877), .A2(n4873), .ZN(n4431) );
  AND2_X1 U5976 ( .A1(n4806), .A2(n4805), .ZN(n4432) );
  NAND2_X1 U5977 ( .A1(n8334), .A2(n6985), .ZN(n4433) );
  AND2_X1 U5978 ( .A1(n8197), .A2(n6321), .ZN(n4434) );
  AND2_X1 U5979 ( .A1(n4657), .A2(n9421), .ZN(n4435) );
  NAND2_X1 U5980 ( .A1(n9245), .A2(n9265), .ZN(n4436) );
  NAND2_X1 U5981 ( .A1(n6929), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4437) );
  AND2_X1 U5982 ( .A1(n4530), .A2(n8286), .ZN(n4438) );
  AND2_X1 U5983 ( .A1(n9263), .A2(n7602), .ZN(n4439) );
  AND2_X1 U5984 ( .A1(n4790), .A2(n4789), .ZN(n4440) );
  AND2_X1 U5985 ( .A1(n4613), .A2(n4611), .ZN(n4441) );
  NAND2_X1 U5986 ( .A1(n8789), .A2(n7911), .ZN(n4442) );
  INV_X1 U5987 ( .A(n4614), .ZN(n4612) );
  NAND2_X1 U5988 ( .A1(n8729), .A2(n7947), .ZN(n4614) );
  NAND2_X1 U5989 ( .A1(n5180), .A2(SI_6_), .ZN(n4443) );
  INV_X1 U5990 ( .A(n4675), .ZN(n4674) );
  NAND2_X1 U5991 ( .A1(n4926), .A2(n5832), .ZN(n4675) );
  INV_X1 U5992 ( .A(n6246), .ZN(n4613) );
  AND2_X1 U5993 ( .A1(n6333), .A2(n8561), .ZN(n6246) );
  INV_X1 U5994 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4941) );
  INV_X1 U5995 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4956) );
  INV_X1 U5996 ( .A(n5973), .ZN(n6040) );
  NAND2_X1 U5997 ( .A1(n8161), .A2(n8169), .ZN(n6757) );
  OR2_X1 U5998 ( .A1(n7462), .A2(n7463), .ZN(n4740) );
  AND2_X1 U5999 ( .A1(n5747), .A2(n7662), .ZN(n7654) );
  XNOR2_X1 U6000 ( .A(n7517), .B(SI_29_), .ZN(n8852) );
  AND2_X1 U6001 ( .A1(n9255), .A2(n4651), .ZN(n4444) );
  NAND2_X1 U6002 ( .A1(n4741), .A2(n4742), .ZN(n7997) );
  AND2_X2 U6003 ( .A1(n6673), .A2(n8319), .ZN(n8290) );
  NAND2_X1 U6004 ( .A1(n4866), .A2(n8247), .ZN(n8609) );
  NAND2_X1 U6005 ( .A1(n6329), .A2(n8245), .ZN(n8621) );
  NAND2_X1 U6006 ( .A1(n4463), .A2(n5824), .ZN(n7290) );
  NAND2_X1 U6007 ( .A1(n4662), .A2(n5823), .ZN(n7200) );
  NAND2_X1 U6008 ( .A1(n4670), .A2(n5825), .ZN(n7339) );
  NAND2_X1 U6009 ( .A1(n4699), .A2(n5347), .ZN(n7398) );
  AND2_X1 U6010 ( .A1(n9386), .A2(n9242), .ZN(n4445) );
  AOI21_X1 U6011 ( .B1(n4632), .B2(n4630), .A(n4629), .ZN(n4628) );
  OR2_X1 U6012 ( .A1(n7901), .A2(n8627), .ZN(n4446) );
  AND2_X1 U6013 ( .A1(n7889), .A2(n8669), .ZN(n4447) );
  NAND2_X1 U6014 ( .A1(n8757), .A2(n8659), .ZN(n4448) );
  INV_X1 U6015 ( .A(n9145), .ZN(n9164) );
  NOR2_X1 U6016 ( .A1(n9183), .A2(n5882), .ZN(n9145) );
  OR2_X1 U6017 ( .A1(n8084), .A2(n8085), .ZN(n4449) );
  NAND2_X1 U6018 ( .A1(n4811), .A2(n4577), .ZN(n4450) );
  AND2_X1 U6019 ( .A1(n7903), .A2(n8614), .ZN(n4451) );
  NAND2_X1 U6020 ( .A1(n9893), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4452) );
  AND2_X1 U6021 ( .A1(n8644), .A2(n8643), .ZN(n8657) );
  INV_X1 U6022 ( .A(n8657), .ZN(n4559) );
  AND2_X1 U6023 ( .A1(n7236), .A2(n6066), .ZN(n4453) );
  NOR2_X1 U6024 ( .A1(n4928), .A2(n4449), .ZN(n4744) );
  AND2_X1 U6025 ( .A1(n4740), .A2(n4739), .ZN(n4454) );
  INV_X2 U6026 ( .A(n9988), .ZN(n9986) );
  XNOR2_X1 U6027 ( .A(n4980), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7451) );
  NOR3_X1 U6028 ( .A1(n7285), .A2(n9398), .A3(n4654), .ZN(n4652) );
  INV_X1 U6029 ( .A(n8362), .ZN(n4807) );
  NAND2_X1 U6030 ( .A1(n4660), .A2(n4661), .ZN(n7221) );
  AND2_X1 U6031 ( .A1(n6901), .A2(n4375), .ZN(n4455) );
  NAND2_X1 U6032 ( .A1(n4845), .A2(n8199), .ZN(n7331) );
  NOR2_X1 U6033 ( .A1(n6982), .A2(n6981), .ZN(n4456) );
  NOR2_X1 U6034 ( .A1(n9907), .A2(n9908), .ZN(n4457) );
  INV_X1 U6035 ( .A(n4653), .ZN(n9292) );
  NOR2_X1 U6036 ( .A1(n7285), .A2(n4654), .ZN(n4653) );
  OR2_X1 U6037 ( .A1(n7118), .A2(n7119), .ZN(n4579) );
  AND2_X1 U6038 ( .A1(n9902), .A2(n7070), .ZN(n4458) );
  AND2_X1 U6039 ( .A1(n4582), .A2(n4585), .ZN(n4459) );
  AND2_X1 U6040 ( .A1(n7153), .A2(n6037), .ZN(n4460) );
  AND2_X1 U6041 ( .A1(n4895), .A2(n5873), .ZN(n4461) );
  INV_X1 U6042 ( .A(n7138), .ZN(n4642) );
  AND4_X1 U6043 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n6317)
         );
  AND3_X1 U6044 ( .A1(n4952), .A2(n4951), .A3(n4950), .ZN(n4909) );
  OR2_X2 U6045 ( .A1(n6619), .A2(n6628), .ZN(n8456) );
  INV_X1 U6046 ( .A(n9788), .ZN(n4641) );
  INV_X1 U6047 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4961) );
  INV_X1 U6048 ( .A(n7120), .ZN(n4578) );
  AND2_X1 U6049 ( .A1(n8346), .A2(n7389), .ZN(n4462) );
  XNOR2_X1 U6050 ( .A(n4594), .B(n5915), .ZN(n6536) );
  INV_X1 U6051 ( .A(n6536), .ZN(n4783) );
  NAND2_X1 U6052 ( .A1(n4992), .A2(n4993), .ZN(n9471) );
  INV_X1 U6053 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4728) );
  INV_X1 U6054 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4822) );
  INV_X2 U6055 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6056 ( .A1(n7598), .A2(n9273), .ZN(n7604) );
  NAND2_X1 U6057 ( .A1(n5238), .A2(n5237), .ZN(n5265) );
  NAND2_X1 U6058 ( .A1(n4523), .A2(n4430), .ZN(n4521) );
  NAND2_X1 U6059 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  NOR2_X1 U6060 ( .A1(n4518), .A2(n7606), .ZN(n7613) );
  AOI21_X1 U6061 ( .B1(n7566), .B2(n4506), .A(n4504), .ZN(n4516) );
  NAND2_X1 U6062 ( .A1(n7651), .A2(n7650), .ZN(n4503) );
  NAND2_X1 U6063 ( .A1(n7290), .A2(n4424), .ZN(n4666) );
  NAND2_X1 U6064 ( .A1(n7221), .A2(n7222), .ZN(n4463) );
  INV_X1 U6065 ( .A(n4901), .ZN(n5410) );
  NAND2_X1 U6066 ( .A1(n4902), .A2(n4901), .ZN(n4470) );
  AND2_X2 U6067 ( .A1(n4672), .A2(n4671), .ZN(n4901) );
  NAND2_X1 U6068 ( .A1(n6793), .A2(n6797), .ZN(n6792) );
  NAND2_X1 U6069 ( .A1(n6646), .A2(n7671), .ZN(n6645) );
  OAI21_X2 U6070 ( .B1(n7004), .B2(n5176), .A(n4475), .ZN(n6966) );
  NAND2_X2 U6071 ( .A1(n5153), .A2(n6943), .ZN(n7004) );
  NAND4_X1 U6072 ( .A1(n4483), .A2(n4480), .A3(n4390), .A4(n4479), .ZN(n6346)
         );
  NAND3_X1 U6073 ( .A1(n4425), .A2(n4483), .A3(n4482), .ZN(n4481) );
  NAND2_X1 U6074 ( .A1(n4495), .A2(n5086), .ZN(n6692) );
  NAND2_X1 U6075 ( .A1(n4495), .A2(n4494), .ZN(n6694) );
  AND2_X1 U6076 ( .A1(n5124), .A2(n5086), .ZN(n4494) );
  NAND2_X1 U6077 ( .A1(n6657), .A2(n6658), .ZN(n4495) );
  NAND2_X1 U6078 ( .A1(n8876), .A2(n4709), .ZN(n4496) );
  NAND2_X1 U6079 ( .A1(n4496), .A2(n4497), .ZN(n5598) );
  INV_X1 U6080 ( .A(n7766), .ZN(n4517) );
  AOI21_X1 U6081 ( .B1(n4511), .B2(n4517), .A(n4505), .ZN(n4504) );
  NAND2_X1 U6082 ( .A1(n4512), .A2(n7765), .ZN(n4507) );
  INV_X1 U6083 ( .A(n7583), .ZN(n4514) );
  AOI21_X1 U6084 ( .B1(n4516), .B2(n7770), .A(n7571), .ZN(n7568) );
  NAND2_X2 U6085 ( .A1(n4524), .A2(n4527), .ZN(n5324) );
  OR2_X1 U6086 ( .A1(n5236), .A2(n5235), .ZN(n5238) );
  OAI21_X1 U6087 ( .B1(n8278), .B2(n4531), .A(n4438), .ZN(n4529) );
  AND2_X1 U6088 ( .A1(n4535), .A2(n4533), .ZN(n4532) );
  NAND2_X1 U6089 ( .A1(n8250), .A2(n8290), .ZN(n4543) );
  NAND2_X1 U6090 ( .A1(n4543), .A2(n4542), .ZN(n8257) );
  INV_X1 U6091 ( .A(n4536), .ZN(n8270) );
  NAND3_X1 U6092 ( .A1(n4543), .A2(n4542), .A3(n4540), .ZN(n4537) );
  NAND2_X1 U6093 ( .A1(n6182), .A2(n4544), .ZN(n6294) );
  NAND2_X1 U6094 ( .A1(n4545), .A2(n4421), .ZN(n8316) );
  NAND4_X1 U6095 ( .A1(n4551), .A2(n4550), .A3(n4546), .A4(n8309), .ZN(n4545)
         );
  NAND2_X1 U6096 ( .A1(n4549), .A2(n4548), .ZN(n4547) );
  AOI21_X1 U6097 ( .B1(n8768), .B2(n8314), .A(n8312), .ZN(n4548) );
  NAND3_X1 U6098 ( .A1(n8207), .A2(n4552), .A3(n4553), .ZN(n8215) );
  NAND3_X1 U6099 ( .A1(n4555), .A2(n4554), .A3(n4434), .ZN(n4553) );
  NAND2_X1 U6100 ( .A1(n8190), .A2(n8290), .ZN(n4554) );
  NAND2_X1 U6101 ( .A1(n8191), .A2(n8297), .ZN(n4555) );
  NAND2_X1 U6102 ( .A1(n4577), .A2(n7414), .ZN(n4809) );
  OAI21_X1 U6103 ( .B1(n7387), .B2(P2_REG2_REG_11__SCAN_IN), .A(n4462), .ZN(
        n4576) );
  INV_X1 U6104 ( .A(n7387), .ZN(n4577) );
  NAND2_X1 U6105 ( .A1(n4808), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U6106 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  NOR2_X1 U6107 ( .A1(n8390), .A2(n8662), .ZN(n8408) );
  NAND2_X1 U6108 ( .A1(n7068), .A2(n7070), .ZN(n4590) );
  OAI21_X1 U6109 ( .B1(n8433), .B2(n4592), .A(n4591), .ZN(n8470) );
  INV_X1 U6110 ( .A(n8526), .ZN(n4597) );
  AOI21_X1 U6111 ( .B1(n8526), .B2(n8143), .A(n8145), .ZN(n8516) );
  AND2_X1 U6112 ( .A1(n8512), .A2(n8517), .ZN(n4603) );
  NAND2_X1 U6113 ( .A1(n8569), .A2(n4441), .ZN(n4606) );
  NAND2_X1 U6114 ( .A1(n6168), .A2(n4618), .ZN(n4616) );
  NAND3_X1 U6115 ( .A1(n4626), .A2(n4627), .A3(n4625), .ZN(n8658) );
  NAND3_X1 U6116 ( .A1(n4628), .A2(n4448), .A3(n4631), .ZN(n4625) );
  NAND3_X1 U6117 ( .A1(n7475), .A2(n4448), .A3(n4628), .ZN(n4626) );
  OAI21_X1 U6118 ( .B1(n7475), .B2(n4631), .A(n4628), .ZN(n8668) );
  OAI21_X1 U6119 ( .B1(n7475), .B2(n6116), .A(n6115), .ZN(n9556) );
  AOI21_X1 U6120 ( .B1(n6116), .B2(n6115), .A(n4633), .ZN(n4632) );
  NAND2_X1 U6121 ( .A1(n7177), .A2(n6051), .ZN(n7237) );
  INV_X1 U6122 ( .A(n7237), .ZN(n6064) );
  INV_X1 U6123 ( .A(n4634), .ZN(n4756) );
  NAND4_X1 U6124 ( .A1(n5917), .A2(n4757), .A3(n5981), .A4(n5915), .ZN(n4634)
         );
  NAND2_X1 U6125 ( .A1(n5999), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U6126 ( .A1(n6204), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U6127 ( .B1(n6392), .B2(n9988), .A(n4920), .ZN(n6383) );
  NAND2_X1 U6128 ( .A1(n4640), .A2(n6901), .ZN(n7209) );
  NAND2_X1 U6129 ( .A1(n4644), .A2(n5040), .ZN(n4643) );
  INV_X1 U6130 ( .A(n4652), .ZN(n9280) );
  AND2_X1 U6131 ( .A1(n9126), .A2(n4659), .ZN(n5899) );
  NAND2_X1 U6132 ( .A1(n9126), .A2(n4657), .ZN(n9079) );
  NAND2_X1 U6133 ( .A1(n4435), .A2(n9126), .ZN(n9080) );
  NAND2_X1 U6134 ( .A1(n9126), .A2(n9425), .ZN(n9112) );
  NAND2_X1 U6135 ( .A1(n7051), .A2(n4663), .ZN(n4660) );
  NAND2_X1 U6136 ( .A1(n4666), .A2(n4667), .ZN(n7442) );
  NAND4_X1 U6137 ( .A1(n4935), .A2(n4936), .A3(n4934), .A4(n4933), .ZN(n4673)
         );
  NOR2_X2 U6138 ( .A1(n5182), .A2(n4673), .ZN(n4937) );
  INV_X1 U6139 ( .A(n4937), .ZN(n5408) );
  NAND2_X1 U6140 ( .A1(n9144), .A2(n4684), .ZN(n4681) );
  NAND2_X1 U6141 ( .A1(n4681), .A2(n4682), .ZN(n7499) );
  NAND2_X1 U6142 ( .A1(n9144), .A2(n4692), .ZN(n4687) );
  NAND2_X1 U6143 ( .A1(n4901), .A2(n4900), .ZN(n4989) );
  AND3_X2 U6144 ( .A1(n4901), .A2(n4900), .A3(n4695), .ZN(n4992) );
  OAI21_X2 U6145 ( .B1(n9228), .B2(n5834), .A(n5835), .ZN(n9210) );
  NAND2_X1 U6146 ( .A1(n6897), .A2(n7533), .ZN(n6896) );
  NOR2_X2 U6147 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4889) );
  NAND3_X1 U6148 ( .A1(n5808), .A2(n5810), .A3(n5809), .ZN(P1_U3220) );
  NAND2_X2 U6149 ( .A1(n4974), .A2(n6395), .ZN(n5790) );
  NAND2_X2 U6150 ( .A1(n4975), .A2(n6395), .ZN(n5673) );
  NAND2_X1 U6151 ( .A1(n7294), .A2(n4369), .ZN(n4698) );
  NAND2_X2 U6152 ( .A1(n4698), .A2(n4697), .ZN(n5397) );
  NAND2_X1 U6153 ( .A1(n8943), .A2(n4428), .ZN(n4702) );
  NOR2_X1 U6154 ( .A1(n8924), .A2(n5652), .ZN(n8897) );
  INV_X1 U6155 ( .A(n8920), .ZN(n4707) );
  NAND2_X1 U6156 ( .A1(n4718), .A2(n4716), .ZN(n8913) );
  OAI21_X2 U6157 ( .B1(n5429), .B2(n4720), .A(n5455), .ZN(n4717) );
  NAND2_X1 U6158 ( .A1(n4937), .A2(n4723), .ZN(n4944) );
  NAND2_X1 U6160 ( .A1(n4727), .A2(n4724), .ZN(n6675) );
  NAND3_X1 U6161 ( .A1(n6358), .A2(n7806), .A3(n6511), .ZN(n4724) );
  NAND2_X1 U6162 ( .A1(n6358), .A2(n7806), .ZN(n4729) );
  NAND2_X1 U6163 ( .A1(n7908), .A2(n4734), .ZN(n4732) );
  XNOR2_X1 U6164 ( .A(n7878), .B(n8329), .ZN(n7462) );
  INV_X1 U6165 ( .A(n4740), .ZN(n7882) );
  NAND2_X1 U6166 ( .A1(n7931), .A2(n4744), .ZN(n4741) );
  INV_X1 U6167 ( .A(n4928), .ZN(n4747) );
  NAND2_X1 U6168 ( .A1(n7921), .A2(n4749), .ZN(n4748) );
  OAI211_X1 U6169 ( .C1(n7921), .C2(n4753), .A(n4750), .B(n4748), .ZN(n7967)
         );
  NAND2_X1 U6170 ( .A1(n7921), .A2(n8075), .ZN(n7925) );
  NAND3_X1 U6171 ( .A1(n4758), .A2(n4759), .A3(n5980), .ZN(n6032) );
  NAND2_X1 U6172 ( .A1(n4762), .A2(n4760), .ZN(n7187) );
  NAND3_X1 U6173 ( .A1(n4370), .A2(n6980), .A3(n6834), .ZN(n4762) );
  INV_X1 U6174 ( .A(n6983), .ZN(n4766) );
  NAND2_X1 U6175 ( .A1(n8064), .A2(n4769), .ZN(n4767) );
  NAND2_X1 U6176 ( .A1(n4767), .A2(n4768), .ZN(n7968) );
  XNOR2_X1 U6177 ( .A(n5958), .B(n5959), .ZN(n6437) );
  INV_X1 U6178 ( .A(n4784), .ZN(n4781) );
  INV_X1 U6179 ( .A(n8461), .ZN(n4789) );
  INV_X1 U6180 ( .A(n7075), .ZN(n4797) );
  INV_X1 U6181 ( .A(n9835), .ZN(n4798) );
  NAND2_X1 U6182 ( .A1(n9834), .A2(n6439), .ZN(n6440) );
  INV_X1 U6183 ( .A(n4811), .ZN(n7413) );
  NAND2_X2 U6184 ( .A1(n4813), .A2(n5632), .ZN(n5882) );
  XNOR2_X2 U6185 ( .A(n5654), .B(n5653), .ZN(n7304) );
  NAND2_X2 U6186 ( .A1(n5631), .A2(n5630), .ZN(n5654) );
  NAND2_X1 U6187 ( .A1(n7659), .A2(n4818), .ZN(n4815) );
  NAND3_X1 U6188 ( .A1(n4815), .A2(n4922), .A3(n4814), .ZN(n4817) );
  AOI21_X1 U6189 ( .B1(n4816), .B2(n7741), .A(n7740), .ZN(n7795) );
  NAND2_X1 U6190 ( .A1(n4817), .A2(n7737), .ZN(n4816) );
  INV_X1 U6191 ( .A(n7663), .ZN(n4818) );
  NAND3_X1 U6192 ( .A1(n10228), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4819) );
  NAND3_X1 U6193 ( .A1(n4983), .A2(n4822), .A3(n4821), .ZN(n4820) );
  NAND2_X1 U6194 ( .A1(n5163), .A2(n4389), .ZN(n4825) );
  NAND2_X1 U6195 ( .A1(n4825), .A2(n4823), .ZN(n5203) );
  NAND2_X1 U6196 ( .A1(n5163), .A2(n5162), .ZN(n4827) );
  NAND3_X1 U6197 ( .A1(n4829), .A2(n4832), .A3(n5293), .ZN(n4828) );
  NAND2_X1 U6198 ( .A1(n4834), .A2(n4833), .ZN(n5486) );
  NAND2_X1 U6199 ( .A1(n5533), .A2(n5537), .ZN(n4835) );
  NAND2_X1 U6200 ( .A1(n4835), .A2(n4836), .ZN(n5558) );
  OAI21_X2 U6201 ( .B1(n5324), .B2(n4840), .A(n4838), .ZN(n5402) );
  NAND2_X1 U6202 ( .A1(n4845), .A2(n4843), .ZN(n7330) );
  NAND2_X1 U6203 ( .A1(n8523), .A2(n4854), .ZN(n4853) );
  NAND2_X1 U6204 ( .A1(n8596), .A2(n4861), .ZN(n4857) );
  NAND2_X1 U6205 ( .A1(n4857), .A2(n4858), .ZN(n8576) );
  NAND2_X1 U6206 ( .A1(n8577), .A2(n4864), .ZN(n8553) );
  NAND2_X1 U6207 ( .A1(n8553), .A2(n8272), .ZN(n6334) );
  NAND3_X1 U6208 ( .A1(n5915), .A2(n5980), .A3(n5981), .ZN(n6006) );
  NAND2_X1 U6209 ( .A1(n4866), .A2(n4865), .ZN(n6331) );
  AND2_X1 U6210 ( .A1(n4365), .A2(n5924), .ZN(n6298) );
  NAND2_X1 U6211 ( .A1(n4365), .A2(n4870), .ZN(n5940) );
  AND2_X1 U6212 ( .A1(n9123), .A2(n7711), .ZN(n9110) );
  NAND2_X1 U6213 ( .A1(n4874), .A2(n4431), .ZN(n5885) );
  NAND2_X1 U6214 ( .A1(n4880), .A2(n7785), .ZN(n4873) );
  INV_X1 U6215 ( .A(n4880), .ZN(n4875) );
  NAND2_X1 U6216 ( .A1(n4883), .A2(n4882), .ZN(n9206) );
  NAND2_X1 U6217 ( .A1(n7280), .A2(n7590), .ZN(n4888) );
  NAND3_X1 U6218 ( .A1(n5109), .A2(n4889), .A3(n5041), .ZN(n5167) );
  NAND3_X1 U6219 ( .A1(n4892), .A2(n5867), .A3(n4890), .ZN(n6798) );
  NAND3_X1 U6220 ( .A1(n6585), .A2(n7667), .A3(n7751), .ZN(n4892) );
  NAND2_X1 U6221 ( .A1(n4893), .A2(n5866), .ZN(n6644) );
  NAND2_X1 U6222 ( .A1(n6585), .A2(n7667), .ZN(n4893) );
  NAND2_X1 U6223 ( .A1(n6882), .A2(n4429), .ZN(n4895) );
  NAND2_X1 U6224 ( .A1(n4897), .A2(n4439), .ZN(n9262) );
  NAND2_X1 U6225 ( .A1(n5881), .A2(n4905), .ZN(n9158) );
  NAND2_X1 U6226 ( .A1(n9158), .A2(n4903), .ZN(n5884) );
  NAND2_X1 U6227 ( .A1(n5152), .A2(n5151), .ZN(n6943) );
  INV_X1 U6228 ( .A(n5149), .ZN(n5152) );
  OR2_X1 U6229 ( .A1(n5025), .A2(n7841), .ZN(n5000) );
  INV_X1 U6230 ( .A(n4995), .ZN(n9480) );
  NAND2_X1 U6232 ( .A1(n6355), .A2(n6354), .ZN(n6357) );
  OR2_X1 U6233 ( .A1(n6477), .A2(n6373), .ZN(n6614) );
  OR2_X1 U6234 ( .A1(n6477), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6361) );
  NAND2_X2 U6235 ( .A1(n7701), .A2(n7712), .ZN(n7697) );
  XNOR2_X1 U6236 ( .A(n5032), .B(n4984), .ZN(n5031) );
  AND2_X1 U6237 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  NAND2_X2 U6238 ( .A1(n5785), .A2(n5784), .ZN(n5847) );
  NAND2_X1 U6239 ( .A1(n4996), .A2(n9480), .ZN(n5025) );
  AND2_X1 U6240 ( .A1(n6387), .A2(n6672), .ZN(n6772) );
  NAND2_X1 U6241 ( .A1(n5064), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6242 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  NAND2_X1 U6243 ( .A1(n7461), .A2(n7460), .ZN(n7878) );
  NAND2_X1 U6244 ( .A1(n5862), .A2(n6527), .ZN(n6526) );
  AOI21_X2 U6245 ( .B1(n5486), .B2(n5485), .A(n4925), .ZN(n5508) );
  OAI22_X2 U6246 ( .A1(n9162), .A2(n5841), .B1(n8900), .B2(n9436), .ZN(n9144)
         );
  NAND2_X1 U6247 ( .A1(n6317), .A2(n6788), .ZN(n8159) );
  AND2_X1 U6248 ( .A1(n6478), .A2(n9587), .ZN(n4907) );
  INV_X1 U6249 ( .A(n5899), .ZN(n7503) );
  OR2_X1 U6250 ( .A1(n6395), .A2(n5014), .ZN(n4908) );
  INV_X1 U6251 ( .A(n6314), .ZN(n6315) );
  XNOR2_X1 U6252 ( .A(n8106), .B(n6338), .ZN(n7875) );
  INV_X1 U6253 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6173) );
  INV_X1 U6254 ( .A(n7074), .ZN(n7060) );
  OR2_X1 U6255 ( .A1(n7872), .A2(n8807), .ZN(n4910) );
  OR2_X1 U6256 ( .A1(n5457), .A2(n10213), .ZN(n4911) );
  OR2_X1 U6257 ( .A1(n7872), .A2(n8736), .ZN(n4913) );
  AND2_X1 U6258 ( .A1(n5039), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4916) );
  OR2_X1 U6259 ( .A1(n9425), .A2(n9002), .ZN(n4917) );
  AND2_X1 U6260 ( .A1(n7186), .A2(n8333), .ZN(n4918) );
  OR2_X1 U6261 ( .A1(n8045), .A2(n8590), .ZN(n4919) );
  OR2_X1 U6262 ( .A1(n9986), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4920) );
  AND2_X1 U6263 ( .A1(n6674), .A2(n8299), .ZN(n4921) );
  OR2_X1 U6264 ( .A1(n5886), .A2(n7746), .ZN(n4922) );
  NOR2_X1 U6265 ( .A1(n5263), .A2(n7163), .ZN(n4923) );
  NOR2_X1 U6266 ( .A1(n5484), .A2(n5483), .ZN(n4925) );
  INV_X1 U6267 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6068) );
  INV_X1 U6268 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6121) );
  AND2_X1 U6269 ( .A1(n5064), .A2(n9827), .ZN(n7495) );
  NAND2_X2 U6270 ( .A1(n6786), .A2(n9553), .ZN(n9562) );
  INV_X1 U6271 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5036) );
  INV_X1 U6272 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5107) );
  OR2_X1 U6273 ( .A1(n9386), .A2(n9242), .ZN(n4926) );
  NAND2_X1 U6274 ( .A1(n6844), .A2(n7235), .ZN(n9969) );
  INV_X1 U6275 ( .A(n9969), .ZN(n6344) );
  INV_X1 U6276 ( .A(n7786), .ZN(n7652) );
  XNOR2_X1 U6277 ( .A(n8479), .B(n8478), .ZN(n4927) );
  NAND2_X1 U6278 ( .A1(n6350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6376) );
  NOR2_X1 U6279 ( .A1(n7887), .A2(n7932), .ZN(n4928) );
  NOR2_X1 U6280 ( .A1(n8037), .A2(n7887), .ZN(n4929) );
  OR2_X1 U6281 ( .A1(n7884), .A2(n9558), .ZN(n4930) );
  AND2_X1 U6282 ( .A1(n8113), .A2(n8112), .ZN(n8315) );
  OR2_X1 U6283 ( .A1(n7920), .A2(n8538), .ZN(n4931) );
  NOR2_X1 U6284 ( .A1(n7593), .A2(n7654), .ZN(n7594) );
  NOR2_X1 U6285 ( .A1(n7595), .A2(n7594), .ZN(n7596) );
  NAND2_X1 U6286 ( .A1(n7597), .A2(n7596), .ZN(n7598) );
  NAND2_X1 U6287 ( .A1(n7703), .A2(n7654), .ZN(n7616) );
  NAND2_X1 U6288 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  MUX2_X1 U6289 ( .A(n7719), .B(n7705), .S(n7654), .Z(n7623) );
  NAND2_X1 U6290 ( .A1(n7620), .A2(n7615), .ZN(n7703) );
  NAND2_X1 U6291 ( .A1(n9084), .A2(n7660), .ZN(n7648) );
  NAND2_X1 U6292 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  AND4_X1 U6293 ( .A1(n5923), .A2(n5922), .A3(n6181), .A4(n6185), .ZN(n5924)
         );
  NOR2_X1 U6294 ( .A1(n9417), .A2(n7664), .ZN(n7655) );
  OR2_X1 U6295 ( .A1(n8774), .A2(n8528), .ZN(n6276) );
  INV_X1 U6296 ( .A(SI_19_), .ZN(n10223) );
  INV_X1 U6297 ( .A(n7039), .ZN(n7037) );
  INV_X1 U6298 ( .A(n8856), .ZN(n5943) );
  INV_X1 U6299 ( .A(n5937), .ZN(n5928) );
  INV_X1 U6300 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5300) );
  XNOR2_X1 U6301 ( .A(n5004), .B(n5788), .ZN(n5022) );
  INV_X1 U6302 ( .A(n5517), .ZN(n5493) );
  NAND2_X1 U6303 ( .A1(n4956), .A2(n4961), .ZN(n4962) );
  INV_X1 U6304 ( .A(SI_23_), .ZN(n10214) );
  INV_X1 U6305 ( .A(SI_16_), .ZN(n10213) );
  INV_X1 U6306 ( .A(SI_8_), .ZN(n10116) );
  INV_X1 U6307 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10119) );
  OR2_X1 U6308 ( .A1(n6133), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U6309 ( .A1(n6347), .A2(n5928), .ZN(n5933) );
  NOR2_X1 U6310 ( .A1(n8378), .A2(n8377), .ZN(n8382) );
  INV_X1 U6311 ( .A(n9909), .ZN(n8489) );
  NAND2_X1 U6312 ( .A1(n8536), .A2(n6254), .ZN(n8526) );
  OR2_X1 U6313 ( .A1(n6190), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6207) );
  NOR2_X1 U6314 ( .A1(n6108), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6122) );
  NOR2_X1 U6315 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6013) );
  INV_X1 U6316 ( .A(n5567), .ZN(n5565) );
  OR2_X1 U6317 ( .A1(n8976), .A2(n8977), .ZN(n5698) );
  OR2_X1 U6318 ( .A1(n5662), .A2(n5661), .ZN(n5683) );
  OR2_X1 U6319 ( .A1(n5542), .A2(n5541), .ZN(n5567) );
  INV_X1 U6320 ( .A(n9090), .ZN(n5898) );
  XNOR2_X1 U6321 ( .A(n5811), .B(n7745), .ZN(n5862) );
  NAND2_X1 U6322 ( .A1(n5886), .A2(n7740), .ZN(n5748) );
  OR2_X1 U6323 ( .A1(n7209), .A2(n8961), .ZN(n7208) );
  INV_X1 U6324 ( .A(SI_27_), .ZN(n10065) );
  INV_X1 U6325 ( .A(SI_20_), .ZN(n5559) );
  INV_X1 U6326 ( .A(SI_17_), .ZN(n10182) );
  INV_X1 U6327 ( .A(SI_14_), .ZN(n10231) );
  NAND2_X1 U6328 ( .A1(n5063), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5035) );
  AND2_X1 U6329 ( .A1(n6052), .A2(n7255), .ZN(n6069) );
  AND2_X1 U6330 ( .A1(n6155), .A2(n10119), .ZN(n6174) );
  AND2_X1 U6331 ( .A1(n7268), .A2(n7267), .ZN(n7266) );
  INV_X1 U6332 ( .A(n8636), .ZN(n7955) );
  OR2_X1 U6333 ( .A1(n6241), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6249) );
  INV_X1 U6334 ( .A(n6672), .ZN(n6776) );
  NOR2_X1 U6335 ( .A1(n9969), .A2(n6673), .ZN(n6638) );
  AND3_X1 U6336 ( .A1(n6062), .A2(n6061), .A3(n6060), .ZN(n9962) );
  AND2_X1 U6337 ( .A1(n8176), .A2(n8182), .ZN(n8124) );
  INV_X1 U6338 ( .A(n8671), .ZN(n9928) );
  INV_X1 U6339 ( .A(n7455), .ZN(n6359) );
  AND2_X1 U6340 ( .A1(n6083), .A2(n6082), .ZN(n6104) );
  NOR2_X1 U6341 ( .A1(n4972), .A2(n7408), .ZN(n4973) );
  INV_X1 U6342 ( .A(n9159), .ZN(n9326) );
  INV_X1 U6343 ( .A(n7739), .ZN(n7741) );
  AND2_X1 U6344 ( .A1(n5763), .A2(n5684), .ZN(n9128) );
  INV_X1 U6345 ( .A(n5664), .ZN(n5798) );
  NAND2_X1 U6346 ( .A1(n7836), .A2(n9025), .ZN(n9721) );
  AND2_X1 U6347 ( .A1(n9705), .A2(n7829), .ZN(n9720) );
  AND2_X1 U6348 ( .A1(n7615), .A2(n7614), .ZN(n9195) );
  INV_X1 U6349 ( .A(n4909), .ZN(n7740) );
  AND2_X1 U6350 ( .A1(n7663), .A2(n7661), .ZN(n9746) );
  AND2_X1 U6351 ( .A1(n6686), .A2(n6685), .ZN(n8091) );
  OR2_X1 U6352 ( .A1(n6733), .A2(n6732), .ZN(n8096) );
  AOI21_X1 U6353 ( .B1(n8540), .B2(n4357), .A(n6253), .ZN(n8549) );
  AND4_X1 U6354 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n8650)
         );
  AND4_X1 U6355 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n9558)
         );
  NAND2_X1 U6356 ( .A1(n6375), .A2(n6374), .ZN(n6619) );
  INV_X1 U6357 ( .A(n9871), .ZN(n9896) );
  AND2_X1 U6358 ( .A1(n8211), .A2(n8212), .ZN(n8130) );
  AND2_X1 U6359 ( .A1(n6638), .A2(n6637), .ZN(n9934) );
  INV_X1 U6360 ( .A(n8736), .ZN(n8753) );
  NAND2_X1 U6361 ( .A1(n8844), .A2(n6776), .ZN(n6617) );
  INV_X1 U6362 ( .A(n9967), .ZN(n9985) );
  NAND2_X1 U6363 ( .A1(n6674), .A2(n7235), .ZN(n9967) );
  OR2_X1 U6364 ( .A1(n9919), .A2(n6344), .ZN(n9980) );
  NOR2_X1 U6365 ( .A1(n6084), .A2(n6104), .ZN(n7382) );
  INV_X1 U6366 ( .A(n8994), .ZN(n8985) );
  AND4_X1 U6367 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n7400)
         );
  INV_X1 U6368 ( .A(n9721), .ZN(n9712) );
  INV_X1 U6369 ( .A(n9307), .ZN(n9275) );
  AND2_X1 U6370 ( .A1(n5746), .A2(n9470), .ZN(n5910) );
  AND2_X1 U6371 ( .A1(n7654), .A2(n7740), .ZN(n9787) );
  INV_X1 U6372 ( .A(n5910), .ZN(n6745) );
  AND2_X1 U6373 ( .A1(n5329), .A2(n5354), .ZN(n9635) );
  AND2_X1 U6374 ( .A1(n5216), .A2(n5243), .ZN(n9521) );
  INV_X1 U6375 ( .A(n5970), .ZN(n6399) );
  INV_X1 U6376 ( .A(n8096), .ZN(n8040) );
  INV_X1 U6377 ( .A(n8315), .ZN(n8494) );
  INV_X1 U6378 ( .A(n8094), .ZN(n8660) );
  OR2_X1 U6379 ( .A1(P2_U3150), .A2(n6429), .ZN(n9841) );
  INV_X1 U6380 ( .A(n6411), .ZN(n9857) );
  NAND2_X1 U6381 ( .A1(n6433), .A2(n6432), .ZN(n9905) );
  NAND2_X1 U6382 ( .A1(n9562), .A2(n9561), .ZN(n8667) );
  NAND2_X1 U6383 ( .A1(n10003), .A2(n9980), .ZN(n8756) );
  INV_X1 U6384 ( .A(n10003), .ZN(n10004) );
  XOR2_X1 U6385 ( .A(n8515), .B(n4423), .Z(n8777) );
  OR2_X1 U6386 ( .A1(n9988), .A2(n9974), .ZN(n8840) );
  OR2_X1 U6387 ( .A1(n9988), .A2(n9967), .ZN(n8807) );
  AND2_X1 U6388 ( .A1(n6382), .A2(n6381), .ZN(n9988) );
  NAND2_X1 U6389 ( .A1(n6637), .A2(n6477), .ZN(n6510) );
  INV_X1 U6390 ( .A(n8380), .ZN(n8397) );
  INV_X1 U6391 ( .A(n7125), .ZN(n7078) );
  INV_X1 U6392 ( .A(n7344), .ZN(n9409) );
  INV_X1 U6393 ( .A(n8980), .ZN(n8996) );
  INV_X1 U6394 ( .A(n8991), .ZN(n8973) );
  INV_X1 U6395 ( .A(n9327), .ZN(n9131) );
  INV_X1 U6396 ( .A(n8993), .ZN(n9271) );
  INV_X1 U6397 ( .A(n7296), .ZN(n9804) );
  INV_X1 U6398 ( .A(n9593), .ZN(n9732) );
  OR2_X1 U6399 ( .A1(n9295), .A2(n7662), .ZN(n9282) );
  OR2_X1 U6400 ( .A1(n9295), .A2(n6796), .ZN(n9307) );
  NAND2_X1 U6401 ( .A1(n9826), .A2(n9806), .ZN(n9406) );
  INV_X1 U6402 ( .A(n9826), .ZN(n9824) );
  INV_X1 U6403 ( .A(n9118), .ZN(n9425) );
  INV_X1 U6404 ( .A(n9234), .ZN(n9452) );
  INV_X1 U6405 ( .A(n9816), .ZN(n9814) );
  INV_X1 U6406 ( .A(n8456), .ZN(P2_U3893) );
  AND2_X2 U6407 ( .A1(n6396), .A2(n6479), .ZN(P1_U3973) );
  INV_X2 U6408 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U6409 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4935) );
  NAND2_X1 U6410 ( .A1(n4944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6411 ( .A1(n5459), .A2(n4943), .ZN(n4938) );
  NAND2_X1 U6412 ( .A1(n5511), .A2(n4942), .ZN(n4939) );
  AND2_X2 U6413 ( .A1(n4946), .A2(n4948), .ZN(n4955) );
  INV_X1 U6414 ( .A(n4955), .ZN(n4952) );
  NAND2_X1 U6415 ( .A1(n4948), .A2(n4945), .ZN(n4951) );
  INV_X1 U6416 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6417 ( .A1(n4947), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6418 ( .A1(n5748), .A2(n5002), .ZN(n4960) );
  NAND2_X1 U6419 ( .A1(n4955), .A2(n4954), .ZN(n4963) );
  INV_X1 U6420 ( .A(n5747), .ZN(n4959) );
  NAND2_X2 U6421 ( .A1(n4959), .A2(n5886), .ZN(n5857) );
  NOR2_X1 U6422 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4967) );
  NOR2_X1 U6423 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4966) );
  NOR2_X1 U6424 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4965) );
  NAND4_X1 U6425 ( .A1(n4968), .A2(n4967), .A3(n4966), .A4(n4965), .ZN(n4969)
         );
  INV_X1 U6426 ( .A(n7451), .ZN(n4972) );
  INV_X1 U6428 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6429 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n4979) );
  NAND2_X1 U6430 ( .A1(n4980), .A2(n4979), .ZN(n4982) );
  INV_X4 U6431 ( .A(n5064), .ZN(n5267) );
  MUX2_X1 U6432 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5063), .Z(n5032) );
  INV_X1 U6433 ( .A(SI_1_), .ZN(n4984) );
  NAND3_X1 U6434 ( .A1(n5267), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4986) );
  AND2_X1 U6435 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6436 ( .A1(n5064), .A2(n4985), .ZN(n5968) );
  NAND2_X1 U6437 ( .A1(n4986), .A2(n5968), .ZN(n5030) );
  XNOR2_X1 U6438 ( .A(n5031), .B(n5030), .ZN(n6455) );
  INV_X1 U6439 ( .A(n6455), .ZN(n4987) );
  NAND2_X1 U6440 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4988) );
  XNOR2_X1 U6441 ( .A(n4988), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9018) );
  INV_X1 U6442 ( .A(n4996), .ZN(n9476) );
  XNOR2_X2 U6443 ( .A(n4994), .B(n4993), .ZN(n4995) );
  INV_X1 U6444 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7812) );
  INV_X1 U6445 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U6446 ( .A1(n5058), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4999) );
  INV_X1 U6447 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n4997) );
  OR2_X1 U6448 ( .A1(n5088), .A2(n4997), .ZN(n4998) );
  AND2_X2 U6449 ( .A1(n6395), .A2(n6795), .ZN(n5173) );
  NAND2_X1 U6450 ( .A1(n5811), .A2(n5173), .ZN(n5003) );
  INV_X4 U6451 ( .A(n5673), .ZN(n5788) );
  INV_X4 U6452 ( .A(n5790), .ZN(n5694) );
  NAND2_X1 U6453 ( .A1(n5811), .A2(n5694), .ZN(n5006) );
  XNOR2_X1 U6454 ( .A(n5022), .B(n5020), .ZN(n6577) );
  NAND2_X1 U6455 ( .A1(n5058), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5010) );
  INV_X1 U6456 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6751) );
  OR2_X1 U6457 ( .A1(n5088), .A2(n6751), .ZN(n5009) );
  INV_X1 U6458 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9029) );
  INV_X1 U6459 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5014) );
  OR2_X1 U6460 ( .A1(n5025), .A2(n5014), .ZN(n5007) );
  NAND2_X1 U6461 ( .A1(n5863), .A2(n5173), .ZN(n5013) );
  NAND2_X1 U6462 ( .A1(n7525), .A2(SI_0_), .ZN(n5011) );
  XNOR2_X1 U6463 ( .A(n5011), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9483) );
  MUX2_X1 U6464 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9483), .S(n5040), .Z(n6556) );
  NAND2_X1 U6465 ( .A1(n5077), .A2(n6556), .ZN(n5012) );
  NAND2_X1 U6466 ( .A1(n5013), .A2(n5012), .ZN(n5018) );
  INV_X1 U6467 ( .A(n5018), .ZN(n5015) );
  NAND2_X1 U6468 ( .A1(n5863), .A2(n5694), .ZN(n5017) );
  INV_X1 U6469 ( .A(n6395), .ZN(n5754) );
  AOI22_X1 U6470 ( .A1(n5173), .A2(n6556), .B1(n5754), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6471 ( .A1(n5017), .A2(n5016), .ZN(n6551) );
  NAND2_X1 U6472 ( .A1(n6552), .A2(n6551), .ZN(n6550) );
  OR2_X1 U6473 ( .A1(n5018), .A2(n5503), .ZN(n5019) );
  AND2_X1 U6474 ( .A1(n6550), .A2(n5019), .ZN(n6578) );
  NAND2_X1 U6475 ( .A1(n6577), .A2(n6578), .ZN(n5024) );
  INV_X1 U6476 ( .A(n5020), .ZN(n5021) );
  NAND2_X1 U6477 ( .A1(n5022), .A2(n5021), .ZN(n5023) );
  NAND2_X1 U6478 ( .A1(n5024), .A2(n5023), .ZN(n6597) );
  NAND2_X1 U6479 ( .A1(n5058), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5029) );
  INV_X1 U6480 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9034) );
  INV_X1 U6481 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7811) );
  OR2_X1 U6482 ( .A1(n5089), .A2(n7811), .ZN(n5027) );
  INV_X1 U6483 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7840) );
  NAND4_X4 U6484 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n5814)
         );
  NAND2_X1 U6485 ( .A1(n5814), .A2(n5173), .ZN(n5049) );
  NAND2_X1 U6486 ( .A1(n5031), .A2(n5030), .ZN(n5034) );
  NAND2_X1 U6487 ( .A1(n5032), .A2(SI_1_), .ZN(n5033) );
  NAND2_X1 U6488 ( .A1(n5034), .A2(n5033), .ZN(n5097) );
  OAI21_X1 U6489 ( .B1(n5063), .B2(n5036), .A(n5035), .ZN(n5068) );
  INV_X1 U6490 ( .A(SI_2_), .ZN(n5037) );
  XNOR2_X1 U6491 ( .A(n5068), .B(n5037), .ZN(n5095) );
  XNOR2_X1 U6492 ( .A(n5097), .B(n5095), .ZN(n6459) );
  INV_X1 U6493 ( .A(n6459), .ZN(n5038) );
  NAND2_X1 U6494 ( .A1(n5094), .A2(n5038), .ZN(n5047) );
  OR2_X1 U6495 ( .A1(n5041), .A2(n4945), .ZN(n5111) );
  INV_X1 U6496 ( .A(n5111), .ZN(n5042) );
  NAND2_X1 U6497 ( .A1(n5042), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5044) );
  INV_X1 U6498 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6499 ( .A1(n5111), .A2(n5043), .ZN(n5072) );
  AND2_X1 U6500 ( .A1(n5044), .A2(n5072), .ZN(n9037) );
  NAND2_X1 U6501 ( .A1(n6478), .A2(n9037), .ZN(n5045) );
  INV_X1 U6502 ( .A(n5813), .ZN(n6600) );
  NAND2_X1 U6503 ( .A1(n6600), .A2(n5077), .ZN(n5048) );
  NAND2_X1 U6504 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  XNOR2_X1 U6505 ( .A(n5050), .B(n5788), .ZN(n5055) );
  NAND2_X1 U6506 ( .A1(n5814), .A2(n5694), .ZN(n5052) );
  OR2_X1 U6507 ( .A1(n5813), .A2(n5310), .ZN(n5051) );
  NAND2_X1 U6508 ( .A1(n5052), .A2(n5051), .ZN(n5053) );
  XNOR2_X1 U6509 ( .A(n5055), .B(n5053), .ZN(n6598) );
  NAND2_X1 U6510 ( .A1(n6597), .A2(n6598), .ZN(n5057) );
  INV_X1 U6511 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6512 ( .A1(n5055), .A2(n5054), .ZN(n5056) );
  NAND2_X1 U6513 ( .A1(n5057), .A2(n5056), .ZN(n6657) );
  NAND2_X1 U6514 ( .A1(n5058), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5062) );
  OR2_X1 U6515 ( .A1(n5088), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5061) );
  INV_X1 U6516 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7815) );
  OR2_X1 U6517 ( .A1(n5089), .A2(n7815), .ZN(n5060) );
  INV_X1 U6518 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7844) );
  OR2_X1 U6519 ( .A1(n5025), .A2(n7844), .ZN(n5059) );
  NAND2_X1 U6520 ( .A1(n9012), .A2(n5173), .ZN(n5079) );
  INV_X1 U6521 ( .A(SI_3_), .ZN(n5067) );
  XNOR2_X1 U6522 ( .A(n5098), .B(n5067), .ZN(n5101) );
  NAND2_X1 U6523 ( .A1(n5097), .A2(n5095), .ZN(n5069) );
  NAND2_X1 U6524 ( .A1(n5068), .A2(SI_2_), .ZN(n5099) );
  NAND2_X1 U6525 ( .A1(n5069), .A2(n5099), .ZN(n5070) );
  XNOR2_X1 U6526 ( .A(n5101), .B(n5070), .ZN(n6465) );
  INV_X1 U6527 ( .A(n6465), .ZN(n5071) );
  NAND2_X1 U6528 ( .A1(n4352), .A2(n5071), .ZN(n5076) );
  NAND2_X1 U6529 ( .A1(n5039), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6530 ( .A1(n5072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6531 ( .A(n5073), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U6532 ( .A1(n6478), .A2(n9050), .ZN(n5074) );
  AND3_X2 U6533 ( .A1(n5076), .A2(n5075), .A3(n5074), .ZN(n6813) );
  INV_X1 U6534 ( .A(n6813), .ZN(n5816) );
  NAND2_X1 U6535 ( .A1(n5816), .A2(n5711), .ZN(n5078) );
  NAND2_X1 U6536 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  XNOR2_X1 U6537 ( .A(n5080), .B(n5788), .ZN(n5085) );
  NAND2_X1 U6538 ( .A1(n9012), .A2(n5694), .ZN(n5082) );
  OR2_X1 U6539 ( .A1(n6813), .A2(n5310), .ZN(n5081) );
  NAND2_X1 U6540 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  XNOR2_X1 U6541 ( .A(n5085), .B(n5083), .ZN(n6658) );
  INV_X1 U6542 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6543 ( .A1(n5085), .A2(n5084), .ZN(n5086) );
  NAND2_X1 U6544 ( .A1(n5518), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5093) );
  INV_X1 U6545 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5087) );
  OR2_X1 U6546 ( .A1(n5888), .A2(n5087), .ZN(n5092) );
  NAND2_X1 U6547 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5140) );
  OAI21_X1 U6548 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5140), .ZN(n6805) );
  OR2_X1 U6549 ( .A1(n5664), .A2(n6805), .ZN(n5091) );
  INV_X1 U6550 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6802) );
  OR2_X1 U6551 ( .A1(n5089), .A2(n6802), .ZN(n5090) );
  NAND2_X1 U6552 ( .A1(n9011), .A2(n5173), .ZN(n5120) );
  AND2_X1 U6553 ( .A1(n5101), .A2(n5095), .ZN(n5096) );
  NAND2_X1 U6554 ( .A1(n5097), .A2(n5096), .ZN(n5105) );
  NAND2_X1 U6555 ( .A1(n5098), .A2(SI_3_), .ZN(n5103) );
  INV_X1 U6556 ( .A(n5099), .ZN(n5100) );
  NAND2_X1 U6557 ( .A1(n5105), .A2(n5104), .ZN(n5129) );
  OAI21_X1 U6558 ( .B1(n5267), .B2(n5107), .A(n5106), .ZN(n5130) );
  INV_X1 U6559 ( .A(SI_4_), .ZN(n5108) );
  XNOR2_X1 U6560 ( .A(n5130), .B(n5108), .ZN(n5128) );
  XNOR2_X1 U6561 ( .A(n5129), .B(n5128), .ZN(n6461) );
  OR2_X1 U6562 ( .A1(n5212), .A2(n6461), .ZN(n5117) );
  OR2_X1 U6563 ( .A1(n5109), .A2(n4945), .ZN(n5110) );
  AND2_X1 U6564 ( .A1(n5111), .A2(n5110), .ZN(n5114) );
  INV_X1 U6565 ( .A(n5114), .ZN(n5112) );
  NAND2_X1 U6566 ( .A1(n5112), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5115) );
  INV_X1 U6567 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6568 ( .A1(n5114), .A2(n5113), .ZN(n5133) );
  AND2_X1 U6569 ( .A1(n5115), .A2(n5133), .ZN(n9587) );
  NAND2_X1 U6570 ( .A1(n9770), .A2(n4351), .ZN(n5119) );
  NAND2_X1 U6571 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  XNOR2_X1 U6572 ( .A(n5121), .B(n5503), .ZN(n5126) );
  NAND2_X1 U6573 ( .A1(n4349), .A2(n5694), .ZN(n5123) );
  NAND2_X1 U6574 ( .A1(n9770), .A2(n5173), .ZN(n5122) );
  NAND2_X1 U6575 ( .A1(n5123), .A2(n5122), .ZN(n5125) );
  XNOR2_X1 U6576 ( .A(n5126), .B(n5125), .ZN(n6693) );
  INV_X1 U6577 ( .A(n6693), .ZN(n5124) );
  NAND2_X1 U6578 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  NAND2_X1 U6579 ( .A1(n6694), .A2(n5127), .ZN(n5149) );
  NAND2_X1 U6580 ( .A1(n5129), .A2(n5128), .ZN(n5132) );
  NAND2_X1 U6581 ( .A1(n5130), .A2(SI_4_), .ZN(n5131) );
  NAND2_X1 U6582 ( .A1(n5132), .A2(n5131), .ZN(n5163) );
  MUX2_X1 U6583 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5267), .Z(n5164) );
  INV_X1 U6584 ( .A(SI_5_), .ZN(n10198) );
  XNOR2_X1 U6585 ( .A(n5163), .B(n5162), .ZN(n6463) );
  OR2_X1 U6586 ( .A1(n6463), .A2(n5212), .ZN(n5136) );
  NAND2_X1 U6587 ( .A1(n5133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5134) );
  XNOR2_X1 U6588 ( .A(n5134), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9602) );
  AOI22_X1 U6589 ( .A1(n7645), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6478), .B2(
        n9602), .ZN(n5135) );
  NAND2_X1 U6590 ( .A1(n5518), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5146) );
  INV_X1 U6591 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6592 ( .A1(n5888), .A2(n5137), .ZN(n5145) );
  INV_X1 U6593 ( .A(n5140), .ZN(n5138) );
  NAND2_X1 U6594 ( .A1(n5138), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5156) );
  INV_X1 U6595 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6596 ( .A1(n5140), .A2(n5139), .ZN(n5141) );
  NAND2_X1 U6597 ( .A1(n5156), .A2(n5141), .ZN(n6952) );
  OR2_X1 U6598 ( .A1(n5664), .A2(n6952), .ZN(n5144) );
  INV_X1 U6599 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5142) );
  OR2_X1 U6600 ( .A1(n5089), .A2(n5142), .ZN(n5143) );
  NAND4_X1 U6601 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n9010)
         );
  NAND2_X1 U6602 ( .A1(n9010), .A2(n5173), .ZN(n5147) );
  OAI21_X1 U6603 ( .B1(n7544), .B2(n5118), .A(n5147), .ZN(n5148) );
  XNOR2_X1 U6604 ( .A(n5148), .B(n5503), .ZN(n5150) );
  NAND2_X1 U6605 ( .A1(n5149), .A2(n5150), .ZN(n6942) );
  INV_X2 U6606 ( .A(n5310), .ZN(n5690) );
  AOI22_X1 U6607 ( .A1(n7541), .A2(n5690), .B1(n9010), .B2(n5694), .ZN(n6945)
         );
  NAND2_X1 U6608 ( .A1(n6942), .A2(n6945), .ZN(n5153) );
  INV_X1 U6609 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6610 ( .A1(n6495), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5161) );
  INV_X1 U6611 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7849) );
  OR2_X1 U6612 ( .A1(n6498), .A2(n7849), .ZN(n5160) );
  INV_X1 U6613 ( .A(n5156), .ZN(n5154) );
  NAND2_X1 U6614 ( .A1(n5154), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5189) );
  INV_X1 U6615 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6616 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6617 ( .A1(n5189), .A2(n5157), .ZN(n6891) );
  OR2_X1 U6618 ( .A1(n5664), .A2(n6891), .ZN(n5159) );
  INV_X1 U6619 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7820) );
  OR2_X1 U6620 ( .A1(n5089), .A2(n7820), .ZN(n5158) );
  NAND2_X1 U6621 ( .A1(n5164), .A2(SI_5_), .ZN(n5165) );
  INV_X1 U6622 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5166) );
  MUX2_X1 U6623 ( .A(n6501), .B(n5166), .S(n5267), .Z(n5179) );
  XNOR2_X1 U6624 ( .A(n5179), .B(SI_6_), .ZN(n5177) );
  XNOR2_X1 U6625 ( .A(n5178), .B(n5177), .ZN(n6467) );
  OR2_X1 U6626 ( .A1(n6467), .A2(n5212), .ZN(n5170) );
  NAND2_X1 U6627 ( .A1(n5167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5168) );
  XNOR2_X1 U6628 ( .A(n5168), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9063) );
  AOI22_X1 U6629 ( .A1(n7645), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6478), .B2(
        n9063), .ZN(n5169) );
  NAND2_X1 U6630 ( .A1(n5170), .A2(n5169), .ZN(n7537) );
  NAND2_X1 U6631 ( .A1(n7537), .A2(n5492), .ZN(n5171) );
  OAI21_X1 U6632 ( .B1(n7536), .B2(n5310), .A(n5171), .ZN(n5172) );
  XNOR2_X1 U6633 ( .A(n5172), .B(n5788), .ZN(n7006) );
  OR2_X1 U6634 ( .A1(n7536), .A2(n5790), .ZN(n5175) );
  NAND2_X1 U6635 ( .A1(n7537), .A2(n5173), .ZN(n5174) );
  AND2_X1 U6636 ( .A1(n5175), .A2(n5174), .ZN(n7005) );
  AND2_X1 U6637 ( .A1(n7006), .A2(n7005), .ZN(n5176) );
  INV_X1 U6638 ( .A(n5179), .ZN(n5180) );
  MUX2_X1 U6639 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5267), .Z(n5204) );
  INV_X1 U6640 ( .A(SI_7_), .ZN(n5181) );
  XNOR2_X1 U6641 ( .A(n5204), .B(n5181), .ZN(n5202) );
  XNOR2_X1 U6642 ( .A(n5203), .B(n5202), .ZN(n6471) );
  OR2_X1 U6643 ( .A1(n6471), .A2(n5212), .ZN(n5185) );
  NAND2_X1 U6644 ( .A1(n5182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U6645 ( .A(n5183), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U6646 ( .A1(n7645), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6478), .B2(
        n9508), .ZN(n5184) );
  NAND2_X1 U6647 ( .A1(n5185), .A2(n5184), .ZN(n6961) );
  NAND2_X1 U6648 ( .A1(n6961), .A2(n5492), .ZN(n5197) );
  NAND2_X1 U6649 ( .A1(n5518), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5195) );
  INV_X1 U6650 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6651 ( .A1(n5888), .A2(n5186), .ZN(n5194) );
  INV_X1 U6652 ( .A(n5189), .ZN(n5187) );
  NAND2_X1 U6653 ( .A1(n5187), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5221) );
  INV_X1 U6654 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6655 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  NAND2_X1 U6656 ( .A1(n5221), .A2(n5190), .ZN(n6972) );
  OR2_X1 U6657 ( .A1(n5664), .A2(n6972), .ZN(n5193) );
  INV_X1 U6658 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5191) );
  OR2_X1 U6659 ( .A1(n5089), .A2(n5191), .ZN(n5192) );
  OR2_X1 U6660 ( .A1(n9739), .A2(n5310), .ZN(n5196) );
  NAND2_X1 U6661 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  XNOR2_X1 U6662 ( .A(n5198), .B(n5788), .ZN(n5200) );
  INV_X1 U6663 ( .A(n9739), .ZN(n9009) );
  AOI22_X1 U6664 ( .A1(n6961), .A2(n5690), .B1(n9009), .B2(n5694), .ZN(n5199)
         );
  NAND2_X1 U6665 ( .A1(n5200), .A2(n5199), .ZN(n6967) );
  NAND2_X1 U6666 ( .A1(n6966), .A2(n6967), .ZN(n5201) );
  OR2_X1 U6667 ( .A1(n5200), .A2(n5199), .ZN(n6968) );
  NAND2_X1 U6668 ( .A1(n5201), .A2(n6968), .ZN(n5232) );
  NAND2_X1 U6669 ( .A1(n5203), .A2(n5202), .ZN(n5206) );
  NAND2_X1 U6670 ( .A1(n5204), .A2(SI_7_), .ZN(n5205) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5207) );
  MUX2_X1 U6672 ( .A(n6473), .B(n5207), .S(n5267), .Z(n5208) );
  NAND2_X1 U6673 ( .A1(n5208), .A2(n10116), .ZN(n5237) );
  INV_X1 U6674 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6675 ( .A1(n5209), .A2(SI_8_), .ZN(n5210) );
  NAND2_X1 U6676 ( .A1(n5237), .A2(n5210), .ZN(n5235) );
  INV_X1 U6677 ( .A(n5235), .ZN(n5211) );
  XNOR2_X1 U6678 ( .A(n5236), .B(n5211), .ZN(n6474) );
  OR2_X1 U6679 ( .A1(n6474), .A2(n5212), .ZN(n5218) );
  NOR2_X1 U6680 ( .A1(n5182), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5276) );
  OR2_X1 U6681 ( .A1(n5276), .A2(n4945), .ZN(n5215) );
  INV_X1 U6682 ( .A(n5215), .ZN(n5213) );
  NAND2_X1 U6683 ( .A1(n5213), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5216) );
  INV_X1 U6684 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6685 ( .A1(n5215), .A2(n5214), .ZN(n5243) );
  AOI22_X1 U6686 ( .A1(n7645), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6478), .B2(
        n9521), .ZN(n5217) );
  NAND2_X1 U6687 ( .A1(n5218), .A2(n5217), .ZN(n7138) );
  NAND2_X1 U6688 ( .A1(n7138), .A2(n5492), .ZN(n5229) );
  NAND2_X1 U6689 ( .A1(n5518), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5227) );
  INV_X1 U6690 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5219) );
  OR2_X1 U6691 ( .A1(n5888), .A2(n5219), .ZN(n5226) );
  NAND2_X1 U6692 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  NAND2_X1 U6693 ( .A1(n5249), .A2(n5222), .ZN(n9752) );
  OR2_X1 U6694 ( .A1(n5664), .A2(n9752), .ZN(n5225) );
  INV_X1 U6695 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5223) );
  OR2_X1 U6696 ( .A1(n5089), .A2(n5223), .ZN(n5224) );
  NAND4_X1 U6697 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n9008)
         );
  NAND2_X1 U6698 ( .A1(n9008), .A2(n5690), .ZN(n5228) );
  NAND2_X1 U6699 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  XNOR2_X1 U6700 ( .A(n5230), .B(n5788), .ZN(n5233) );
  AND2_X1 U6701 ( .A1(n9008), .A2(n5694), .ZN(n5231) );
  AOI21_X1 U6702 ( .B1(n7138), .B2(n5690), .A(n5231), .ZN(n7142) );
  INV_X1 U6703 ( .A(n5232), .ZN(n5234) );
  NAND2_X1 U6704 ( .A1(n5234), .A2(n5233), .ZN(n7161) );
  INV_X1 U6705 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5239) );
  MUX2_X1 U6706 ( .A(n6504), .B(n5239), .S(n5267), .Z(n5240) );
  NAND2_X1 U6707 ( .A1(n5240), .A2(n10088), .ZN(n5266) );
  INV_X1 U6708 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6709 ( .A1(n5241), .A2(SI_9_), .ZN(n5242) );
  XNOR2_X1 U6710 ( .A(n5265), .B(n4924), .ZN(n6475) );
  NAND2_X1 U6711 ( .A1(n6475), .A2(n4352), .ZN(n5246) );
  NAND2_X1 U6712 ( .A1(n5243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5244) );
  XNOR2_X1 U6713 ( .A(n5244), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9537) );
  AOI22_X1 U6714 ( .A1(n7645), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6478), .B2(
        n9537), .ZN(n5245) );
  NAND2_X1 U6715 ( .A1(n9788), .A2(n5492), .ZN(n5256) );
  NAND2_X1 U6716 ( .A1(n6495), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5254) );
  INV_X1 U6717 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7839) );
  OR2_X1 U6718 ( .A1(n6498), .A2(n7839), .ZN(n5253) );
  INV_X1 U6719 ( .A(n5249), .ZN(n5247) );
  NAND2_X1 U6720 ( .A1(n5247), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5301) );
  INV_X1 U6721 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6722 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  NAND2_X1 U6723 ( .A1(n5301), .A2(n5250), .ZN(n7164) );
  OR2_X1 U6724 ( .A1(n5664), .A2(n7164), .ZN(n5252) );
  INV_X1 U6725 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7099) );
  OR2_X1 U6726 ( .A1(n5089), .A2(n7099), .ZN(n5251) );
  OR2_X1 U6727 ( .A1(n9741), .A2(n5310), .ZN(n5255) );
  NAND2_X1 U6728 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  XNOR2_X1 U6729 ( .A(n5257), .B(n5503), .ZN(n5262) );
  INV_X1 U6730 ( .A(n5262), .ZN(n5259) );
  NOR2_X1 U6731 ( .A1(n9741), .A2(n5790), .ZN(n5258) );
  AOI21_X1 U6732 ( .B1(n9788), .B2(n5690), .A(n5258), .ZN(n5261) );
  NAND2_X1 U6733 ( .A1(n5259), .A2(n5261), .ZN(n5260) );
  INV_X1 U6734 ( .A(n5260), .ZN(n5263) );
  XNOR2_X1 U6735 ( .A(n5262), .B(n5261), .ZN(n7163) );
  MUX2_X1 U6736 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5267), .Z(n5269) );
  XNOR2_X1 U6737 ( .A(n5269), .B(n5268), .ZN(n5293) );
  NAND2_X1 U6738 ( .A1(n5269), .A2(SI_10_), .ZN(n5270) );
  INV_X1 U6739 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5271) );
  MUX2_X1 U6740 ( .A(n6508), .B(n5271), .S(n5267), .Z(n5272) );
  NAND2_X1 U6741 ( .A1(n5272), .A2(n10099), .ZN(n5323) );
  INV_X1 U6742 ( .A(n5272), .ZN(n5273) );
  NAND2_X1 U6743 ( .A1(n5273), .A2(SI_11_), .ZN(n5274) );
  NAND2_X1 U6744 ( .A1(n5323), .A2(n5274), .ZN(n5321) );
  XNOR2_X1 U6745 ( .A(n5322), .B(n5321), .ZN(n6506) );
  NAND2_X1 U6746 ( .A1(n6506), .A2(n4352), .ZN(n5279) );
  NOR2_X1 U6747 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5275) );
  NAND2_X1 U6748 ( .A1(n5276), .A2(n5275), .ZN(n5295) );
  NAND2_X1 U6749 ( .A1(n5326), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5277) );
  XNOR2_X1 U6750 ( .A(n5277), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9619) );
  AOI22_X1 U6751 ( .A1(n7645), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6478), .B2(
        n9619), .ZN(n5278) );
  NAND2_X1 U6752 ( .A1(n8961), .A2(n5492), .ZN(n5289) );
  NAND2_X1 U6753 ( .A1(n6495), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5287) );
  INV_X1 U6754 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5280) );
  OR2_X1 U6755 ( .A1(n6498), .A2(n5280), .ZN(n5286) );
  INV_X1 U6756 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6757 ( .A1(n5303), .A2(n5282), .ZN(n5283) );
  NAND2_X1 U6758 ( .A1(n5333), .A2(n5283), .ZN(n8959) );
  OR2_X1 U6759 ( .A1(n5664), .A2(n8959), .ZN(n5285) );
  INV_X1 U6760 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7211) );
  OR2_X1 U6761 ( .A1(n5089), .A2(n7211), .ZN(n5284) );
  OR2_X1 U6762 ( .A1(n7317), .A2(n5310), .ZN(n5288) );
  NAND2_X1 U6763 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  XNOR2_X1 U6764 ( .A(n5290), .B(n5503), .ZN(n5315) );
  NAND2_X1 U6765 ( .A1(n8961), .A2(n5690), .ZN(n5292) );
  OR2_X1 U6766 ( .A1(n7317), .A2(n5790), .ZN(n5291) );
  NAND2_X1 U6767 ( .A1(n5292), .A2(n5291), .ZN(n8952) );
  XNOR2_X1 U6768 ( .A(n5294), .B(n5293), .ZN(n6481) );
  NAND2_X1 U6769 ( .A1(n6481), .A2(n4352), .ZN(n5298) );
  NAND2_X1 U6770 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5296) );
  XNOR2_X1 U6771 ( .A(n5296), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9489) );
  AOI22_X1 U6772 ( .A1(n7645), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6478), .B2(
        n9489), .ZN(n5297) );
  NAND2_X1 U6773 ( .A1(n5298), .A2(n5297), .ZN(n9797) );
  NAND2_X1 U6774 ( .A1(n9797), .A2(n5690), .ZN(n5309) );
  NAND2_X1 U6775 ( .A1(n6495), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5307) );
  INV_X1 U6776 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5299) );
  OR2_X1 U6777 ( .A1(n5089), .A2(n5299), .ZN(n5306) );
  NAND2_X1 U6778 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  NAND2_X1 U6779 ( .A1(n5303), .A2(n5302), .ZN(n7052) );
  OR2_X1 U6780 ( .A1(n5664), .A2(n7052), .ZN(n5305) );
  OR2_X1 U6781 ( .A1(n6498), .A2(n9822), .ZN(n5304) );
  OR2_X1 U6782 ( .A1(n8956), .A2(n5790), .ZN(n5308) );
  NAND2_X1 U6783 ( .A1(n5309), .A2(n5308), .ZN(n7314) );
  NAND2_X1 U6784 ( .A1(n9797), .A2(n5492), .ZN(n5312) );
  OR2_X1 U6785 ( .A1(n8956), .A2(n5310), .ZN(n5311) );
  NAND2_X1 U6786 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  XNOR2_X1 U6787 ( .A(n5313), .B(n5673), .ZN(n5316) );
  AOI22_X1 U6788 ( .A1(n5315), .A2(n8952), .B1(n7314), .B2(n5316), .ZN(n5314)
         );
  NAND2_X1 U6789 ( .A1(n7313), .A2(n5314), .ZN(n5320) );
  INV_X1 U6790 ( .A(n5315), .ZN(n8953) );
  OAI21_X1 U6791 ( .B1(n5316), .B2(n7314), .A(n8952), .ZN(n5318) );
  NOR2_X1 U6792 ( .A1(n8952), .A2(n7314), .ZN(n5317) );
  INV_X1 U6793 ( .A(n5316), .ZN(n8951) );
  AOI22_X1 U6794 ( .A1(n8953), .A2(n5318), .B1(n5317), .B2(n8951), .ZN(n5319)
         );
  NAND2_X1 U6795 ( .A1(n5320), .A2(n5319), .ZN(n7294) );
  MUX2_X1 U6796 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5267), .Z(n5349) );
  XNOR2_X1 U6797 ( .A(n5349), .B(n5325), .ZN(n5348) );
  XNOR2_X1 U6798 ( .A(n5352), .B(n5348), .ZN(n6514) );
  NAND2_X1 U6799 ( .A1(n6514), .A2(n4352), .ZN(n5331) );
  NOR2_X1 U6800 ( .A1(n5326), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5379) );
  NOR2_X1 U6801 ( .A1(n5379), .A2(n4945), .ZN(n5327) );
  NAND2_X1 U6802 ( .A1(n5327), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5329) );
  INV_X1 U6803 ( .A(n5327), .ZN(n5328) );
  INV_X1 U6804 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6805 ( .A1(n5328), .A2(n5377), .ZN(n5354) );
  AOI22_X1 U6806 ( .A1(n7645), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6478), .B2(
        n9635), .ZN(n5330) );
  NAND2_X1 U6807 ( .A1(n9807), .A2(n5492), .ZN(n5341) );
  NAND2_X1 U6808 ( .A1(n6495), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5339) );
  INV_X1 U6809 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7855) );
  OR2_X1 U6810 ( .A1(n6498), .A2(n7855), .ZN(n5338) );
  NAND2_X1 U6811 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  NAND2_X1 U6812 ( .A1(n5359), .A2(n5334), .ZN(n7300) );
  OR2_X1 U6813 ( .A1(n5664), .A2(n7300), .ZN(n5337) );
  INV_X1 U6814 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6815 ( .A1(n5089), .A2(n5335), .ZN(n5336) );
  OR2_X1 U6816 ( .A1(n7400), .A2(n5310), .ZN(n5340) );
  NAND2_X1 U6817 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  XNOR2_X1 U6818 ( .A(n5342), .B(n5503), .ZN(n5344) );
  NOR2_X1 U6819 ( .A1(n7400), .A2(n5790), .ZN(n5343) );
  AOI21_X1 U6820 ( .B1(n9807), .B2(n5690), .A(n5343), .ZN(n5345) );
  XNOR2_X1 U6821 ( .A(n5344), .B(n5345), .ZN(n7295) );
  INV_X1 U6822 ( .A(n5344), .ZN(n5346) );
  NAND2_X1 U6823 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  INV_X1 U6824 ( .A(n5348), .ZN(n5351) );
  NAND2_X1 U6825 ( .A1(n5349), .A2(SI_12_), .ZN(n5350) );
  MUX2_X1 U6826 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7525), .Z(n5373) );
  XNOR2_X1 U6827 ( .A(n5373), .B(SI_13_), .ZN(n5353) );
  XNOR2_X1 U6828 ( .A(n5374), .B(n5353), .ZN(n6522) );
  NAND2_X1 U6829 ( .A1(n6522), .A2(n4352), .ZN(n5357) );
  NAND2_X1 U6830 ( .A1(n5354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5355) );
  XNOR2_X1 U6831 ( .A(n5355), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9652) );
  AOI22_X1 U6832 ( .A1(n7645), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6478), .B2(
        n9652), .ZN(n5356) );
  NAND2_X1 U6833 ( .A1(n7433), .A2(n5492), .ZN(n5367) );
  NAND2_X1 U6834 ( .A1(n6495), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5365) );
  INV_X1 U6835 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7287) );
  OR2_X1 U6836 ( .A1(n5089), .A2(n7287), .ZN(n5364) );
  NAND2_X1 U6837 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  NAND2_X1 U6838 ( .A1(n5387), .A2(n5360), .ZN(n7403) );
  OR2_X1 U6839 ( .A1(n5664), .A2(n7403), .ZN(n5363) );
  INV_X1 U6840 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5361) );
  OR2_X1 U6841 ( .A1(n6498), .A2(n5361), .ZN(n5362) );
  OR2_X1 U6842 ( .A1(n7296), .A2(n5310), .ZN(n5366) );
  NAND2_X1 U6843 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  XNOR2_X1 U6844 ( .A(n5368), .B(n5503), .ZN(n5370) );
  NOR2_X1 U6845 ( .A1(n7296), .A2(n5790), .ZN(n5369) );
  AOI21_X1 U6846 ( .B1(n7433), .B2(n5690), .A(n5369), .ZN(n5371) );
  INV_X1 U6847 ( .A(n5370), .ZN(n5372) );
  NAND2_X1 U6848 ( .A1(n5375), .A2(n10210), .ZN(n5376) );
  MUX2_X1 U6849 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7525), .Z(n5403) );
  XNOR2_X1 U6850 ( .A(n5403), .B(n10231), .ZN(n5401) );
  XNOR2_X1 U6851 ( .A(n5402), .B(n5401), .ZN(n6583) );
  NAND2_X1 U6852 ( .A1(n6583), .A2(n4352), .ZN(n5383) );
  INV_X1 U6853 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5378) );
  NAND3_X1 U6854 ( .A1(n5379), .A2(n5378), .A3(n5377), .ZN(n5380) );
  NAND2_X1 U6855 ( .A1(n5380), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5381) );
  XNOR2_X1 U6856 ( .A(n5381), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9669) );
  AOI22_X1 U6857 ( .A1(n7645), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6478), .B2(
        n9669), .ZN(n5382) );
  NAND2_X1 U6858 ( .A1(n7344), .A2(n5492), .ZN(n5394) );
  NAND2_X1 U6859 ( .A1(n6495), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5392) );
  INV_X1 U6860 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5384) );
  OR2_X1 U6861 ( .A1(n6498), .A2(n5384), .ZN(n5391) );
  INV_X1 U6862 ( .A(n5387), .ZN(n5385) );
  INV_X1 U6863 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6864 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  NAND2_X1 U6865 ( .A1(n5416), .A2(n5388), .ZN(n8862) );
  OR2_X1 U6866 ( .A1(n5664), .A2(n8862), .ZN(n5390) );
  INV_X1 U6867 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7340) );
  OR2_X1 U6868 ( .A1(n5089), .A2(n7340), .ZN(n5389) );
  NAND4_X1 U6869 ( .A1(n5392), .A2(n5391), .A3(n5390), .A4(n5389), .ZN(n9005)
         );
  NAND2_X1 U6870 ( .A1(n9005), .A2(n5690), .ZN(n5393) );
  NAND2_X1 U6871 ( .A1(n5394), .A2(n5393), .ZN(n5395) );
  XNOR2_X1 U6872 ( .A(n5395), .B(n5503), .ZN(n5398) );
  AND2_X1 U6873 ( .A1(n9005), .A2(n5694), .ZN(n5396) );
  AOI21_X1 U6874 ( .B1(n7344), .B2(n5690), .A(n5396), .ZN(n8860) );
  NAND2_X1 U6875 ( .A1(n8859), .A2(n8860), .ZN(n8858) );
  INV_X1 U6876 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6877 ( .A1(n5397), .A2(n5399), .ZN(n5400) );
  NAND2_X2 U6878 ( .A1(n8858), .A2(n5400), .ZN(n5428) );
  NAND2_X1 U6879 ( .A1(n5402), .A2(n5401), .ZN(n5406) );
  INV_X1 U6880 ( .A(n5403), .ZN(n5404) );
  NAND2_X1 U6881 ( .A1(n5404), .A2(n10231), .ZN(n5405) );
  MUX2_X1 U6882 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7525), .Z(n5434) );
  XNOR2_X1 U6883 ( .A(n5434), .B(n10188), .ZN(n5407) );
  XNOR2_X1 U6884 ( .A(n5430), .B(n5407), .ZN(n6606) );
  NAND2_X1 U6885 ( .A1(n6606), .A2(n4352), .ZN(n5413) );
  NAND2_X1 U6886 ( .A1(n5408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5409) );
  MUX2_X1 U6887 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5409), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5411) );
  NAND2_X1 U6888 ( .A1(n5411), .A2(n5410), .ZN(n7858) );
  INV_X1 U6889 ( .A(n7858), .ZN(n9688) );
  AOI22_X1 U6890 ( .A1(n7645), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6478), .B2(
        n9688), .ZN(n5412) );
  NAND2_X1 U6891 ( .A1(n7443), .A2(n5492), .ZN(n5423) );
  NAND2_X1 U6892 ( .A1(n6495), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5421) );
  INV_X1 U6893 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9682) );
  OR2_X1 U6894 ( .A1(n6498), .A2(n9682), .ZN(n5420) );
  INV_X1 U6895 ( .A(n5416), .ZN(n5414) );
  INV_X1 U6896 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6897 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  NAND2_X1 U6898 ( .A1(n5441), .A2(n5417), .ZN(n8995) );
  OR2_X1 U6899 ( .A1(n5664), .A2(n8995), .ZN(n5419) );
  INV_X1 U6900 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7444) );
  OR2_X1 U6901 ( .A1(n5089), .A2(n7444), .ZN(n5418) );
  NAND4_X1 U6902 ( .A1(n5421), .A2(n5420), .A3(n5419), .A4(n5418), .ZN(n9302)
         );
  NAND2_X1 U6903 ( .A1(n9302), .A2(n5690), .ZN(n5422) );
  NAND2_X1 U6904 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  XNOR2_X1 U6905 ( .A(n5424), .B(n5503), .ZN(n5426) );
  XNOR2_X2 U6906 ( .A(n5428), .B(n5426), .ZN(n8989) );
  AND2_X1 U6907 ( .A1(n9302), .A2(n5694), .ZN(n5425) );
  AOI21_X1 U6908 ( .B1(n7443), .B2(n5690), .A(n5425), .ZN(n8990) );
  INV_X1 U6909 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U6910 ( .A1(n5428), .A2(n5427), .ZN(n5429) );
  INV_X1 U6911 ( .A(n5430), .ZN(n5433) );
  INV_X1 U6912 ( .A(n5434), .ZN(n5431) );
  NAND2_X1 U6913 ( .A1(n5431), .A2(n10188), .ZN(n5432) );
  NAND2_X1 U6914 ( .A1(n5434), .A2(SI_15_), .ZN(n5435) );
  MUX2_X1 U6915 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7525), .Z(n5456) );
  XNOR2_X1 U6916 ( .A(n5456), .B(SI_16_), .ZN(n5436) );
  NAND2_X1 U6917 ( .A1(n5410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5437) );
  XNOR2_X1 U6918 ( .A(n5437), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7860) );
  AOI22_X1 U6919 ( .A1(n7645), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6478), .B2(
        n7860), .ZN(n5438) );
  NAND2_X1 U6920 ( .A1(n9398), .A2(n5492), .ZN(n5449) );
  INV_X1 U6921 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6922 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  AND2_X1 U6923 ( .A1(n5464), .A2(n5442), .ZN(n9294) );
  NAND2_X1 U6924 ( .A1(n9294), .A2(n5798), .ZN(n5447) );
  NAND2_X1 U6925 ( .A1(n6495), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5446) );
  INV_X1 U6926 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5443) );
  OR2_X1 U6927 ( .A1(n5089), .A2(n5443), .ZN(n5445) );
  INV_X1 U6928 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7861) );
  OR2_X1 U6929 ( .A1(n6498), .A2(n7861), .ZN(n5444) );
  OR2_X1 U6930 ( .A1(n8993), .A2(n5310), .ZN(n5448) );
  NAND2_X1 U6931 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XNOR2_X1 U6932 ( .A(n5450), .B(n5673), .ZN(n5452) );
  NOR2_X1 U6933 ( .A1(n8993), .A2(n5790), .ZN(n5451) );
  AOI21_X1 U6934 ( .B1(n9398), .B2(n5690), .A(n5451), .ZN(n5453) );
  XNOR2_X1 U6935 ( .A(n5452), .B(n5453), .ZN(n8905) );
  INV_X1 U6936 ( .A(n5452), .ZN(n5454) );
  NAND2_X1 U6937 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  NAND2_X1 U6938 ( .A1(n5457), .A2(n10213), .ZN(n5481) );
  NAND2_X1 U6939 ( .A1(n5486), .A2(n5481), .ZN(n5458) );
  MUX2_X1 U6940 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7525), .Z(n5479) );
  XNOR2_X1 U6941 ( .A(n5479), .B(n10182), .ZN(n5483) );
  XNOR2_X1 U6942 ( .A(n5458), .B(n5483), .ZN(n6705) );
  NAND2_X1 U6943 ( .A1(n6705), .A2(n4352), .ZN(n5461) );
  XNOR2_X1 U6944 ( .A(n5459), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9710) );
  AOI22_X1 U6945 ( .A1(n7645), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6478), .B2(
        n9710), .ZN(n5460) );
  NAND2_X1 U6946 ( .A1(n9285), .A2(n5492), .ZN(n5471) );
  INV_X1 U6947 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7828) );
  INV_X1 U6948 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6949 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6950 ( .A1(n5515), .A2(n5465), .ZN(n9276) );
  OR2_X1 U6951 ( .A1(n9276), .A2(n5664), .ZN(n5469) );
  INV_X1 U6952 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9459) );
  OR2_X1 U6953 ( .A1(n5888), .A2(n9459), .ZN(n5467) );
  INV_X1 U6954 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9395) );
  OR2_X1 U6955 ( .A1(n6498), .A2(n9395), .ZN(n5466) );
  AND2_X1 U6956 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  OAI211_X1 U6957 ( .C1(n5089), .C2(n7828), .A(n5469), .B(n5468), .ZN(n9301)
         );
  NAND2_X1 U6958 ( .A1(n9301), .A2(n5690), .ZN(n5470) );
  NAND2_X1 U6959 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  XNOR2_X1 U6960 ( .A(n5472), .B(n5503), .ZN(n5474) );
  AND2_X1 U6961 ( .A1(n9301), .A2(n5694), .ZN(n5473) );
  AOI21_X1 U6962 ( .B1(n9285), .B2(n5690), .A(n5473), .ZN(n5475) );
  XNOR2_X1 U6963 ( .A(n5474), .B(n5475), .ZN(n8914) );
  NAND2_X1 U6964 ( .A1(n8913), .A2(n8914), .ZN(n5478) );
  INV_X1 U6965 ( .A(n5474), .ZN(n5476) );
  NAND2_X1 U6966 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  NAND2_X2 U6967 ( .A1(n5478), .A2(n5477), .ZN(n8876) );
  INV_X1 U6968 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6969 ( .A1(n5480), .A2(n10182), .ZN(n5482) );
  AND2_X1 U6970 ( .A1(n5481), .A2(n5482), .ZN(n5485) );
  INV_X1 U6971 ( .A(n5482), .ZN(n5484) );
  MUX2_X1 U6972 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7525), .Z(n5487) );
  NAND2_X1 U6973 ( .A1(n5487), .A2(SI_18_), .ZN(n5488) );
  OAI21_X1 U6974 ( .B1(n5487), .B2(SI_18_), .A(n5488), .ZN(n5507) );
  NAND2_X2 U6975 ( .A1(n5510), .A2(n5488), .ZN(n5533) );
  MUX2_X1 U6976 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7525), .Z(n5535) );
  XNOR2_X1 U6977 ( .A(n5535), .B(SI_19_), .ZN(n5534) );
  XNOR2_X1 U6978 ( .A(n5533), .B(n5534), .ZN(n6879) );
  NAND2_X1 U6979 ( .A1(n6879), .A2(n4352), .ZN(n5491) );
  AOI22_X1 U6980 ( .A1(n7645), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7662), .B2(
        n6478), .ZN(n5490) );
  NAND2_X1 U6981 ( .A1(n9245), .A2(n5492), .ZN(n5502) );
  INV_X1 U6982 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5514) );
  INV_X1 U6983 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6984 ( .A1(n5517), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U6985 ( .A1(n5542), .A2(n5495), .ZN(n9246) );
  OR2_X1 U6986 ( .A1(n9246), .A2(n5664), .ZN(n5500) );
  INV_X1 U6987 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U6988 ( .A1(n5794), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6989 ( .A1(n6495), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5496) );
  OAI211_X1 U6990 ( .C1(n6498), .C2(n9383), .A(n5497), .B(n5496), .ZN(n5498)
         );
  INV_X1 U6991 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U6992 ( .A1(n5500), .A2(n5499), .ZN(n9265) );
  NAND2_X1 U6993 ( .A1(n9265), .A2(n5690), .ZN(n5501) );
  NAND2_X1 U6994 ( .A1(n5502), .A2(n5501), .ZN(n5504) );
  XNOR2_X1 U6995 ( .A(n5504), .B(n5503), .ZN(n8879) );
  NAND2_X1 U6996 ( .A1(n9245), .A2(n5690), .ZN(n5506) );
  NAND2_X1 U6997 ( .A1(n9265), .A2(n5694), .ZN(n5505) );
  NAND2_X1 U6998 ( .A1(n5506), .A2(n5505), .ZN(n5528) );
  NAND2_X1 U6999 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  AND2_X1 U7000 ( .A1(n5510), .A2(n5509), .ZN(n6729) );
  NAND2_X1 U7001 ( .A1(n6729), .A2(n4352), .ZN(n5513) );
  XNOR2_X1 U7002 ( .A(n5511), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U7003 ( .A1(n7645), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6478), .B2(
        n9725), .ZN(n5512) );
  NAND2_X1 U7004 ( .A1(n9386), .A2(n5690), .ZN(n5522) );
  NAND2_X1 U7005 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U7006 ( .A1(n5517), .A2(n5516), .ZN(n9258) );
  AOI22_X1 U7007 ( .A1(n5518), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6495), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7008 ( .A1(n5794), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U7009 ( .C1(n9258), .C2(n5664), .A(n5520), .B(n5519), .ZN(n9242)
         );
  NAND2_X1 U7010 ( .A1(n9242), .A2(n5694), .ZN(n5521) );
  NAND2_X1 U7011 ( .A1(n5522), .A2(n5521), .ZN(n8965) );
  NAND2_X1 U7012 ( .A1(n9386), .A2(n5492), .ZN(n5524) );
  NAND2_X1 U7013 ( .A1(n9242), .A2(n5690), .ZN(n5523) );
  NAND2_X1 U7014 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  XNOR2_X1 U7015 ( .A(n5525), .B(n5673), .ZN(n8875) );
  OAI22_X1 U7016 ( .A1(n8879), .A2(n5528), .B1(n8965), .B2(n8875), .ZN(n5526)
         );
  NAND2_X1 U7017 ( .A1(n8875), .A2(n8965), .ZN(n5527) );
  INV_X1 U7018 ( .A(n5528), .ZN(n8878) );
  NAND2_X1 U7019 ( .A1(n5527), .A2(n8878), .ZN(n5530) );
  INV_X1 U7020 ( .A(n5527), .ZN(n5529) );
  AOI22_X1 U7021 ( .A1(n8879), .A2(n5530), .B1(n5529), .B2(n5528), .ZN(n5531)
         );
  INV_X1 U7022 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U7023 ( .A1(n5536), .A2(n10223), .ZN(n5537) );
  MUX2_X1 U7024 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7525), .Z(n5557) );
  XNOR2_X1 U7025 ( .A(n5557), .B(n5559), .ZN(n5538) );
  XNOR2_X1 U7026 ( .A(n5560), .B(n5538), .ZN(n6991) );
  NAND2_X1 U7027 ( .A1(n6991), .A2(n4352), .ZN(n5540) );
  NAND2_X1 U7028 ( .A1(n5039), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7029 ( .A1(n9234), .A2(n5492), .ZN(n5550) );
  INV_X1 U7030 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7031 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  AND2_X1 U7032 ( .A1(n5567), .A2(n5543), .ZN(n9229) );
  NAND2_X1 U7033 ( .A1(n9229), .A2(n5798), .ZN(n5548) );
  INV_X1 U7034 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U7035 ( .A1(n6495), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7036 ( .A1(n5794), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7037 ( .C1(n9378), .C2(n6498), .A(n5545), .B(n5544), .ZN(n5546)
         );
  INV_X1 U7038 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7039 ( .A1(n5548), .A2(n5547), .ZN(n9364) );
  NAND2_X1 U7040 ( .A1(n9364), .A2(n5690), .ZN(n5549) );
  NAND2_X1 U7041 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  XNOR2_X1 U7042 ( .A(n5551), .B(n5788), .ZN(n8931) );
  AND2_X1 U7043 ( .A1(n9364), .A2(n5694), .ZN(n5552) );
  AOI21_X1 U7044 ( .B1(n9234), .B2(n5690), .A(n5552), .ZN(n5554) );
  NAND2_X1 U7045 ( .A1(n8931), .A2(n5554), .ZN(n5553) );
  INV_X1 U7046 ( .A(n8931), .ZN(n5555) );
  INV_X1 U7047 ( .A(n5554), .ZN(n8930) );
  NAND2_X1 U7048 ( .A1(n5555), .A2(n8930), .ZN(n5556) );
  NAND2_X1 U7049 ( .A1(n5558), .A2(n5557), .ZN(n5561) );
  NAND2_X1 U7050 ( .A1(n5561), .A2(n4912), .ZN(n5584) );
  MUX2_X1 U7051 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7525), .Z(n5580) );
  XNOR2_X1 U7052 ( .A(n5580), .B(SI_21_), .ZN(n5562) );
  XNOR2_X1 U7053 ( .A(n5584), .B(n5562), .ZN(n7088) );
  NAND2_X1 U7054 ( .A1(n7088), .A2(n4352), .ZN(n5564) );
  NAND2_X1 U7055 ( .A1(n5039), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7056 ( .A1(n9222), .A2(n5492), .ZN(n5575) );
  INV_X1 U7057 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7058 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND2_X1 U7059 ( .A1(n5610), .A2(n5568), .ZN(n9212) );
  OR2_X1 U7060 ( .A1(n9212), .A2(n5664), .ZN(n5573) );
  INV_X1 U7061 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U7062 ( .A1(n6495), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7063 ( .A1(n5794), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U7064 ( .C1(n9371), .C2(n6498), .A(n5570), .B(n5569), .ZN(n5571)
         );
  INV_X1 U7065 ( .A(n5571), .ZN(n5572) );
  NAND2_X1 U7066 ( .A1(n5573), .A2(n5572), .ZN(n9355) );
  NAND2_X1 U7067 ( .A1(n9355), .A2(n5690), .ZN(n5574) );
  NAND2_X1 U7068 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  XNOR2_X1 U7069 ( .A(n5576), .B(n5788), .ZN(n5579) );
  AND2_X1 U7070 ( .A1(n9355), .A2(n5694), .ZN(n5577) );
  AOI21_X1 U7071 ( .B1(n9222), .B2(n5690), .A(n5577), .ZN(n5578) );
  XNOR2_X1 U7072 ( .A(n5579), .B(n5578), .ZN(n8888) );
  NOR2_X1 U7073 ( .A1(n5581), .A2(n10199), .ZN(n5583) );
  NAND2_X1 U7074 ( .A1(n5581), .A2(n10199), .ZN(n5582) );
  MUX2_X1 U7075 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7525), .Z(n5601) );
  XNOR2_X1 U7076 ( .A(n5601), .B(n10123), .ZN(n5599) );
  XNOR2_X1 U7077 ( .A(n5600), .B(n5599), .ZN(n7172) );
  NAND2_X1 U7078 ( .A1(n7172), .A2(n4352), .ZN(n5586) );
  NAND2_X1 U7079 ( .A1(n5039), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7080 ( .A1(n9203), .A2(n5492), .ZN(n5593) );
  XNOR2_X1 U7081 ( .A(n5610), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U7082 ( .A1(n9196), .A2(n5798), .ZN(n5591) );
  INV_X1 U7083 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U7084 ( .A1(n5794), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7085 ( .A1(n6495), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7086 ( .C1(n6498), .C2(n9362), .A(n5588), .B(n5587), .ZN(n5589)
         );
  INV_X1 U7087 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7088 ( .A1(n5591), .A2(n5590), .ZN(n9365) );
  NAND2_X1 U7089 ( .A1(n9365), .A2(n5690), .ZN(n5592) );
  NAND2_X1 U7090 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  XNOR2_X1 U7091 ( .A(n5594), .B(n5788), .ZN(n5597) );
  NOR2_X1 U7092 ( .A1(n5598), .A2(n5597), .ZN(n8941) );
  NAND2_X1 U7093 ( .A1(n9203), .A2(n5690), .ZN(n5596) );
  NAND2_X1 U7094 ( .A1(n9365), .A2(n5694), .ZN(n5595) );
  NAND2_X1 U7095 ( .A1(n5596), .A2(n5595), .ZN(n8940) );
  AND2_X2 U7096 ( .A1(n5598), .A2(n5597), .ZN(n8943) );
  NAND2_X1 U7097 ( .A1(n5600), .A2(n5599), .ZN(n5604) );
  INV_X1 U7098 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7099 ( .A1(n5602), .A2(n10123), .ZN(n5603) );
  NAND2_X1 U7100 ( .A1(n5604), .A2(n5603), .ZN(n5627) );
  MUX2_X1 U7101 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7525), .Z(n5628) );
  XNOR2_X1 U7102 ( .A(n5628), .B(n10214), .ZN(n5626) );
  XNOR2_X1 U7103 ( .A(n5627), .B(n5626), .ZN(n6230) );
  NAND2_X1 U7104 ( .A1(n6230), .A2(n4352), .ZN(n5606) );
  NAND2_X1 U7105 ( .A1(n7645), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7106 ( .A1(n9187), .A2(n5492), .ZN(n5618) );
  INV_X1 U7107 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5608) );
  INV_X1 U7108 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5607) );
  OAI21_X1 U7109 ( .B1(n5610), .B2(n5608), .A(n5607), .ZN(n5611) );
  NAND2_X1 U7110 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5609) );
  NAND2_X1 U7111 ( .A1(n5611), .A2(n5635), .ZN(n9175) );
  OR2_X1 U7112 ( .A1(n9175), .A2(n5664), .ZN(n5616) );
  INV_X1 U7113 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U7114 ( .A1(n5794), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7115 ( .A1(n6495), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7116 ( .C1(n6498), .C2(n9353), .A(n5613), .B(n5612), .ZN(n5614)
         );
  INV_X1 U7117 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7118 ( .A1(n9356), .A2(n5690), .ZN(n5617) );
  NAND2_X1 U7119 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U7120 ( .A(n5619), .B(n5788), .ZN(n5621) );
  AND2_X1 U7121 ( .A1(n9356), .A2(n5694), .ZN(n5620) );
  AOI21_X1 U7122 ( .B1(n9187), .B2(n5690), .A(n5620), .ZN(n5622) );
  NAND2_X1 U7123 ( .A1(n5621), .A2(n5622), .ZN(n8921) );
  INV_X1 U7124 ( .A(n5621), .ZN(n5624) );
  INV_X1 U7125 ( .A(n5622), .ZN(n5623) );
  NAND2_X1 U7126 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  AND2_X1 U7127 ( .A1(n8921), .A2(n5625), .ZN(n8867) );
  NAND2_X1 U7128 ( .A1(n5627), .A2(n5626), .ZN(n5631) );
  INV_X1 U7129 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7130 ( .A1(n5629), .A2(n10214), .ZN(n5630) );
  MUX2_X1 U7131 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7525), .Z(n5655) );
  XNOR2_X1 U7132 ( .A(n5655), .B(n10184), .ZN(n5653) );
  NAND2_X1 U7133 ( .A1(n7645), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7134 ( .A1(n5882), .A2(n5492), .ZN(n5643) );
  INV_X1 U7135 ( .A(n5635), .ZN(n5633) );
  NAND2_X1 U7136 ( .A1(n5633), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5662) );
  INV_X1 U7137 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7138 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  NAND2_X1 U7139 ( .A1(n5662), .A2(n5636), .ZN(n9165) );
  OR2_X1 U7140 ( .A1(n9165), .A2(n5664), .ZN(n5641) );
  INV_X1 U7141 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U7142 ( .A1(n6495), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7143 ( .A1(n5794), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U7144 ( .C1(n6498), .C2(n9345), .A(n5638), .B(n5637), .ZN(n5639)
         );
  INV_X1 U7145 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7146 ( .A1(n9347), .A2(n5690), .ZN(n5642) );
  NAND2_X1 U7147 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  XNOR2_X1 U7148 ( .A(n5644), .B(n5788), .ZN(n5646) );
  AND2_X1 U7149 ( .A1(n9347), .A2(n5694), .ZN(n5645) );
  AOI21_X1 U7150 ( .B1(n5882), .B2(n5690), .A(n5645), .ZN(n5647) );
  NAND2_X1 U7151 ( .A1(n5646), .A2(n5647), .ZN(n5651) );
  INV_X1 U7152 ( .A(n5646), .ZN(n5649) );
  INV_X1 U7153 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U7154 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  NAND2_X1 U7155 ( .A1(n5651), .A2(n5650), .ZN(n8920) );
  INV_X1 U7156 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U7157 ( .A1(n5654), .A2(n5653), .ZN(n5658) );
  INV_X1 U7158 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7159 ( .A1(n5656), .A2(n10184), .ZN(n5657) );
  NAND2_X1 U7160 ( .A1(n5658), .A2(n5657), .ZN(n5675) );
  MUX2_X1 U7161 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7525), .Z(n5676) );
  XNOR2_X1 U7162 ( .A(n5676), .B(n10114), .ZN(n5674) );
  XNOR2_X1 U7163 ( .A(n5675), .B(n5674), .ZN(n7407) );
  NAND2_X1 U7164 ( .A1(n7407), .A2(n4352), .ZN(n5660) );
  NAND2_X1 U7165 ( .A1(n7645), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7166 ( .A1(n9148), .A2(n5492), .ZN(n5671) );
  INV_X1 U7167 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7168 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  NAND2_X1 U7169 ( .A1(n5683), .A2(n5663), .ZN(n9149) );
  INV_X1 U7170 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U7171 ( .A1(n5794), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7172 ( .A1(n6495), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U7173 ( .C1(n6498), .C2(n9340), .A(n5666), .B(n5665), .ZN(n5667)
         );
  INV_X1 U7174 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U7175 ( .A1(n9159), .A2(n5690), .ZN(n5670) );
  NAND2_X1 U7176 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  XNOR2_X1 U7177 ( .A(n5673), .B(n5672), .ZN(n5697) );
  OAI22_X1 U7178 ( .A1(n5883), .A2(n5310), .B1(n9326), .B2(n5790), .ZN(n5696)
         );
  XNOR2_X1 U7179 ( .A(n5697), .B(n5696), .ZN(n8896) );
  NAND2_X1 U7180 ( .A1(n5675), .A2(n5674), .ZN(n5679) );
  INV_X1 U7181 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7182 ( .A1(n5677), .A2(n10114), .ZN(n5678) );
  MUX2_X1 U7183 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7525), .Z(n5705) );
  XNOR2_X1 U7184 ( .A(n5705), .B(n10090), .ZN(n5703) );
  XNOR2_X1 U7185 ( .A(n5704), .B(n5703), .ZN(n7450) );
  NAND2_X1 U7186 ( .A1(n7450), .A2(n4352), .ZN(n5681) );
  NAND2_X1 U7187 ( .A1(n7645), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5680) );
  NAND2_X2 U7188 ( .A1(n5681), .A2(n5680), .ZN(n9127) );
  NAND2_X1 U7189 ( .A1(n9127), .A2(n5492), .ZN(n5692) );
  INV_X1 U7190 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7191 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  NAND2_X1 U7192 ( .A1(n9128), .A2(n5798), .ZN(n5689) );
  INV_X1 U7193 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U7194 ( .A1(n5794), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7195 ( .A1(n6495), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5685) );
  OAI211_X1 U7196 ( .C1(n6498), .C2(n9335), .A(n5686), .B(n5685), .ZN(n5687)
         );
  INV_X1 U7197 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7198 ( .A1(n9140), .A2(n5690), .ZN(n5691) );
  NAND2_X1 U7199 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  XNOR2_X1 U7200 ( .A(n5693), .B(n5788), .ZN(n5699) );
  AND2_X1 U7201 ( .A1(n9140), .A2(n5694), .ZN(n5695) );
  AOI21_X1 U7202 ( .B1(n9127), .B2(n5690), .A(n5695), .ZN(n5700) );
  XNOR2_X1 U7203 ( .A(n5699), .B(n5700), .ZN(n8976) );
  NOR2_X1 U7204 ( .A1(n5697), .A2(n5696), .ZN(n8977) );
  NOR2_X2 U7205 ( .A1(n8895), .A2(n5698), .ZN(n8975) );
  INV_X1 U7206 ( .A(n5699), .ZN(n5702) );
  INV_X1 U7207 ( .A(n5700), .ZN(n5701) );
  NAND2_X1 U7208 ( .A1(n5704), .A2(n5703), .ZN(n5708) );
  INV_X1 U7209 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7210 ( .A1(n5706), .A2(n10090), .ZN(n5707) );
  MUX2_X1 U7211 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7525), .Z(n5782) );
  XNOR2_X1 U7212 ( .A(n5782), .B(n10065), .ZN(n5780) );
  NAND2_X1 U7213 ( .A1(n7480), .A2(n4352), .ZN(n5710) );
  NAND2_X1 U7214 ( .A1(n5039), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5709) );
  NAND2_X2 U7215 ( .A1(n5710), .A2(n5709), .ZN(n9118) );
  NAND2_X1 U7216 ( .A1(n9118), .A2(n5492), .ZN(n5719) );
  XNOR2_X1 U7217 ( .A(n5763), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U7218 ( .A1(n9114), .A2(n5798), .ZN(n5717) );
  INV_X1 U7219 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7220 ( .A1(n6495), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7221 ( .A1(n5794), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5712) );
  OAI211_X1 U7222 ( .C1(n6498), .C2(n5714), .A(n5713), .B(n5712), .ZN(n5715)
         );
  INV_X1 U7223 ( .A(n5715), .ZN(n5716) );
  NAND2_X1 U7224 ( .A1(n9131), .A2(n5690), .ZN(n5718) );
  NAND2_X1 U7225 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  XNOR2_X1 U7226 ( .A(n5720), .B(n5788), .ZN(n5723) );
  NOR2_X1 U7227 ( .A1(n9327), .A2(n5790), .ZN(n5721) );
  AOI21_X1 U7228 ( .B1(n9118), .B2(n5690), .A(n5721), .ZN(n5722) );
  NAND2_X1 U7229 ( .A1(n5723), .A2(n5722), .ZN(n5804) );
  OAI21_X1 U7230 ( .B1(n5723), .B2(n5722), .A(n5804), .ZN(n5725) );
  NOR3_X2 U7231 ( .A1(n8975), .A2(n5724), .A3(n5725), .ZN(n5807) );
  INV_X1 U7232 ( .A(n5726), .ZN(n5750) );
  NAND2_X1 U7233 ( .A1(n7408), .A2(P1_B_REG_SCAN_IN), .ZN(n5728) );
  MUX2_X1 U7234 ( .A(n5728), .B(P1_B_REG_SCAN_IN), .S(n5727), .Z(n5729) );
  NOR4_X1 U7235 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5733) );
  NOR4_X1 U7236 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5732) );
  NOR4_X1 U7237 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5731) );
  NOR4_X1 U7238 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5730) );
  AND4_X1 U7239 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n5739)
         );
  NOR2_X1 U7240 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5737) );
  NOR4_X1 U7241 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5736) );
  NOR4_X1 U7242 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5735) );
  NOR4_X1 U7243 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5734) );
  AND4_X1 U7244 ( .A1(n5737), .A2(n5736), .A3(n5735), .A4(n5734), .ZN(n5738)
         );
  NAND2_X1 U7245 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  NAND2_X1 U7246 ( .A1(n6485), .A2(n5740), .ZN(n5751) );
  NAND2_X1 U7247 ( .A1(n5741), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7248 ( .A1(n5751), .A2(n6554), .ZN(n5906) );
  INV_X1 U7249 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U7250 ( .A1(n6485), .A2(n6489), .ZN(n5743) );
  NAND2_X1 U7251 ( .A1(n4972), .A2(n7408), .ZN(n6487) );
  NAND2_X1 U7252 ( .A1(n5743), .A2(n6487), .ZN(n5905) );
  NOR2_X1 U7253 ( .A1(n5906), .A2(n5905), .ZN(n6746) );
  INV_X1 U7254 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7255 ( .A1(n6485), .A2(n5744), .ZN(n5746) );
  INV_X1 U7256 ( .A(n5727), .ZN(n5745) );
  NAND2_X1 U7257 ( .A1(n5745), .A2(n4972), .ZN(n9470) );
  AND2_X1 U7258 ( .A1(n6746), .A2(n5910), .ZN(n5774) );
  NAND2_X1 U7259 ( .A1(n5747), .A2(n7669), .ZN(n6519) );
  INV_X1 U7260 ( .A(n6519), .ZN(n6749) );
  NOR2_X1 U7261 ( .A1(n9806), .A2(n7735), .ZN(n5749) );
  OAI21_X1 U7262 ( .B1(n5807), .B2(n5750), .A(n8991), .ZN(n5779) );
  INV_X1 U7263 ( .A(n5905), .ZN(n5752) );
  NAND3_X1 U7264 ( .A1(n5752), .A2(n5910), .A3(n5751), .ZN(n5757) );
  NAND2_X1 U7265 ( .A1(n9787), .A2(n7669), .ZN(n5904) );
  NAND2_X1 U7266 ( .A1(n5757), .A2(n5904), .ZN(n5753) );
  NAND2_X1 U7267 ( .A1(n7735), .A2(n5856), .ZN(n6744) );
  NAND2_X1 U7268 ( .A1(n5753), .A2(n6744), .ZN(n6553) );
  OAI21_X1 U7269 ( .B1(n6553), .B2(n5754), .A(P1_STATE_REG_SCAN_IN), .ZN(n5755) );
  OR2_X1 U7270 ( .A1(n6479), .A2(P1_U3086), .ZN(n7802) );
  INV_X1 U7271 ( .A(n5856), .ZN(n5756) );
  NAND2_X1 U7272 ( .A1(n7735), .A2(n5756), .ZN(n5859) );
  INV_X1 U7273 ( .A(n5859), .ZN(n6750) );
  NAND2_X1 U7274 ( .A1(n6554), .A2(n6750), .ZN(n7800) );
  NOR2_X1 U7275 ( .A1(n5757), .A2(n7800), .ZN(n5771) );
  NAND2_X1 U7276 ( .A1(n5771), .A2(n4355), .ZN(n8983) );
  INV_X1 U7277 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5762) );
  OAI22_X1 U7278 ( .A1(n9316), .A2(n8983), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5762), .ZN(n5773) );
  INV_X1 U7279 ( .A(n5763), .ZN(n5760) );
  AND2_X1 U7280 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5759) );
  NAND2_X1 U7281 ( .A1(n5760), .A2(n5759), .ZN(n5793) );
  INV_X1 U7282 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5761) );
  OAI21_X1 U7283 ( .B1(n5763), .B2(n5762), .A(n5761), .ZN(n5764) );
  NAND2_X1 U7284 ( .A1(n9100), .A2(n5798), .ZN(n5769) );
  INV_X1 U7285 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U7286 ( .A1(n5794), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7287 ( .A1(n6495), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5765) );
  OAI211_X1 U7288 ( .C1(n6498), .C2(n7511), .A(n5766), .B(n5765), .ZN(n5767)
         );
  INV_X1 U7289 ( .A(n5767), .ZN(n5768) );
  INV_X1 U7290 ( .A(n4355), .ZN(n5770) );
  NAND2_X1 U7291 ( .A1(n5771), .A2(n5770), .ZN(n8994) );
  NOR2_X1 U7292 ( .A1(n9317), .A2(n8994), .ZN(n5772) );
  AOI211_X1 U7293 ( .C1(n9114), .C2(n8980), .A(n5773), .B(n5772), .ZN(n5778)
         );
  INV_X1 U7294 ( .A(n5774), .ZN(n5775) );
  OR2_X1 U7295 ( .A1(n6519), .A2(n7740), .ZN(n6748) );
  OR2_X1 U7296 ( .A1(n5775), .A2(n6748), .ZN(n5777) );
  INV_X1 U7297 ( .A(n5904), .ZN(n5776) );
  NAND3_X1 U7298 ( .A1(n5779), .A2(n5778), .A3(n4917), .ZN(P1_U3214) );
  NAND2_X1 U7299 ( .A1(n5781), .A2(n5780), .ZN(n5785) );
  INV_X1 U7300 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U7301 ( .A1(n5783), .A2(n10065), .ZN(n5784) );
  MUX2_X1 U7302 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7525), .Z(n5848) );
  XNOR2_X1 U7303 ( .A(n5848), .B(n10201), .ZN(n5846) );
  XNOR2_X2 U7304 ( .A(n5847), .B(n5846), .ZN(n6277) );
  NAND2_X1 U7305 ( .A1(n7645), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5786) );
  OAI22_X1 U7306 ( .A1(n9098), .A2(n5118), .B1(n9317), .B2(n5310), .ZN(n5789)
         );
  XNOR2_X1 U7307 ( .A(n5789), .B(n5788), .ZN(n5792) );
  OAI22_X1 U7308 ( .A1(n9098), .A2(n5310), .B1(n9317), .B2(n5790), .ZN(n5791)
         );
  XNOR2_X1 U7309 ( .A(n5792), .B(n5791), .ZN(n5801) );
  NAND3_X1 U7310 ( .A1(n5807), .A2(n5801), .A3(n8991), .ZN(n5810) );
  INV_X1 U7311 ( .A(n5793), .ZN(n9087) );
  INV_X1 U7312 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7313 ( .A1(n5794), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7314 ( .A1(n6495), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5795) );
  OAI211_X1 U7315 ( .C1(n6498), .C2(n5908), .A(n5796), .B(n5795), .ZN(n5797)
         );
  AOI21_X1 U7316 ( .B1(n9087), .B2(n5798), .A(n5797), .ZN(n7502) );
  INV_X1 U7317 ( .A(n7502), .ZN(n9099) );
  AOI22_X1 U7318 ( .A1(n9099), .A2(n8985), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5800) );
  NAND2_X1 U7319 ( .A1(n9100), .A2(n8980), .ZN(n5799) );
  OAI211_X1 U7320 ( .C1(n9327), .C2(n8983), .A(n5800), .B(n5799), .ZN(n5803)
         );
  INV_X1 U7321 ( .A(n5801), .ZN(n5805) );
  NOR3_X1 U7322 ( .A1(n5805), .A2(n5804), .A3(n8973), .ZN(n5802) );
  AOI211_X1 U7323 ( .C1(n7504), .C2(n8971), .A(n5803), .B(n5802), .ZN(n5809)
         );
  NAND3_X1 U7324 ( .A1(n5805), .A2(n8991), .A3(n5804), .ZN(n5806) );
  OR2_X1 U7325 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  NAND2_X1 U7326 ( .A1(n5863), .A2(n6556), .ZN(n6527) );
  NAND2_X1 U7327 ( .A1(n6526), .A2(n5812), .ZN(n6588) );
  NAND2_X1 U7328 ( .A1(n6588), .A2(n6587), .ZN(n6586) );
  OR2_X1 U7329 ( .A1(n5814), .A2(n6600), .ZN(n5815) );
  NAND2_X1 U7330 ( .A1(n6586), .A2(n5815), .ZN(n6646) );
  OR2_X1 U7331 ( .A1(n9012), .A2(n5816), .ZN(n5817) );
  XNOR2_X1 U7332 ( .A(n4349), .B(n6806), .ZN(n6797) );
  OR2_X1 U7333 ( .A1(n4349), .A2(n9770), .ZN(n5818) );
  NAND2_X1 U7334 ( .A1(n6792), .A2(n5818), .ZN(n6821) );
  OR2_X1 U7335 ( .A1(n7544), .A2(n9010), .ZN(n7535) );
  NAND2_X1 U7336 ( .A1(n9010), .A2(n7544), .ZN(n7752) );
  NAND2_X1 U7337 ( .A1(n7535), .A2(n7752), .ZN(n7670) );
  NAND2_X1 U7338 ( .A1(n6821), .A2(n7670), .ZN(n6820) );
  OR2_X1 U7339 ( .A1(n9010), .A2(n7541), .ZN(n5819) );
  NAND2_X1 U7340 ( .A1(n6820), .A2(n5819), .ZN(n6888) );
  NAND2_X1 U7341 ( .A1(n7536), .A2(n7537), .ZN(n7674) );
  NAND2_X1 U7342 ( .A1(n7543), .A2(n7674), .ZN(n6887) );
  NAND2_X1 U7343 ( .A1(n6888), .A2(n6887), .ZN(n6886) );
  INV_X1 U7344 ( .A(n7536), .ZN(n6955) );
  OR2_X1 U7345 ( .A1(n7537), .A2(n6955), .ZN(n5820) );
  NAND2_X1 U7346 ( .A1(n6886), .A2(n5820), .ZN(n6897) );
  OR2_X1 U7347 ( .A1(n6961), .A2(n9739), .ZN(n7555) );
  NAND2_X1 U7348 ( .A1(n6961), .A2(n9739), .ZN(n7675) );
  NAND2_X1 U7349 ( .A1(n7555), .A2(n7675), .ZN(n7533) );
  OR2_X1 U7350 ( .A1(n6961), .A2(n9009), .ZN(n5821) );
  NOR2_X1 U7351 ( .A1(n7138), .A2(n9008), .ZN(n9735) );
  NAND2_X1 U7352 ( .A1(n7138), .A2(n9008), .ZN(n9733) );
  NAND2_X1 U7353 ( .A1(n9788), .A2(n9741), .ZN(n7573) );
  INV_X1 U7354 ( .A(n9741), .ZN(n9795) );
  OR2_X1 U7355 ( .A1(n9788), .A2(n9795), .ZN(n5822) );
  OR2_X1 U7356 ( .A1(n9797), .A2(n8956), .ZN(n7576) );
  NAND2_X1 U7357 ( .A1(n9797), .A2(n8956), .ZN(n7581) );
  NAND2_X1 U7358 ( .A1(n7576), .A2(n7581), .ZN(n7679) );
  INV_X1 U7359 ( .A(n8956), .ZN(n9007) );
  OR2_X1 U7360 ( .A1(n9797), .A2(n9007), .ZN(n5823) );
  NAND2_X1 U7361 ( .A1(n8961), .A2(n7317), .ZN(n7582) );
  NAND2_X1 U7362 ( .A1(n7574), .A2(n7582), .ZN(n7201) );
  INV_X1 U7363 ( .A(n7317), .ZN(n7298) );
  NAND2_X1 U7364 ( .A1(n9807), .A2(n7400), .ZN(n7583) );
  NAND2_X1 U7365 ( .A1(n7575), .A2(n7583), .ZN(n7222) );
  INV_X1 U7366 ( .A(n7400), .ZN(n9006) );
  OR2_X1 U7367 ( .A1(n9807), .A2(n9006), .ZN(n5824) );
  OR2_X1 U7368 ( .A1(n7433), .A2(n7296), .ZN(n7587) );
  NAND2_X1 U7369 ( .A1(n7433), .A2(n7296), .ZN(n7761) );
  NAND2_X1 U7370 ( .A1(n7587), .A2(n7761), .ZN(n7684) );
  OR2_X1 U7371 ( .A1(n7433), .A2(n9804), .ZN(n5825) );
  NAND2_X1 U7372 ( .A1(n7344), .A2(n9005), .ZN(n5826) );
  OR2_X1 U7373 ( .A1(n7344), .A2(n9005), .ZN(n5827) );
  NOR2_X1 U7374 ( .A1(n7443), .A2(n9302), .ZN(n5829) );
  NAND2_X1 U7375 ( .A1(n7443), .A2(n9302), .ZN(n5828) );
  OAI21_X1 U7376 ( .B1(n7442), .B2(n5829), .A(n5828), .ZN(n9289) );
  NAND2_X1 U7377 ( .A1(n7770), .A2(n7774), .ZN(n9290) );
  NAND2_X1 U7378 ( .A1(n9289), .A2(n9290), .ZN(n5831) );
  NAND2_X1 U7379 ( .A1(n9398), .A2(n9271), .ZN(n5830) );
  AND2_X1 U7380 ( .A1(n9285), .A2(n9301), .ZN(n5833) );
  OR2_X1 U7381 ( .A1(n9285), .A2(n9301), .ZN(n5832) );
  NOR2_X1 U7382 ( .A1(n9234), .A2(n9364), .ZN(n5834) );
  NAND2_X1 U7383 ( .A1(n9234), .A2(n9364), .ZN(n5835) );
  OR2_X1 U7384 ( .A1(n9203), .A2(n9365), .ZN(n5836) );
  OR2_X1 U7385 ( .A1(n9222), .A2(n9355), .ZN(n9193) );
  AND2_X1 U7386 ( .A1(n5836), .A2(n9193), .ZN(n5837) );
  NAND2_X1 U7387 ( .A1(n9203), .A2(n9365), .ZN(n5838) );
  OR2_X1 U7388 ( .A1(n9187), .A2(n9356), .ZN(n5840) );
  NOR2_X1 U7389 ( .A1(n5882), .A2(n9347), .ZN(n5841) );
  AND2_X1 U7390 ( .A1(n9148), .A2(n9159), .ZN(n5843) );
  OR2_X1 U7391 ( .A1(n9148), .A2(n9159), .ZN(n5842) );
  NOR2_X1 U7392 ( .A1(n9127), .A2(n9140), .ZN(n5844) );
  NAND2_X1 U7393 ( .A1(n9118), .A2(n9327), .ZN(n7636) );
  NOR2_X1 U7394 ( .A1(n9098), .A2(n9317), .ZN(n5845) );
  INV_X1 U7395 ( .A(n9317), .ZN(n9004) );
  OAI22_X1 U7396 ( .A1(n7499), .A2(n5845), .B1(n9004), .B2(n7504), .ZN(n5855)
         );
  NAND2_X1 U7397 ( .A1(n5847), .A2(n5846), .ZN(n5851) );
  INV_X1 U7398 ( .A(n5848), .ZN(n5849) );
  NAND2_X1 U7399 ( .A1(n5849), .A2(n10201), .ZN(n5850) );
  INV_X1 U7400 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8854) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5852) );
  MUX2_X1 U7402 ( .A(n8854), .B(n5852), .S(n7525), .Z(n7513) );
  NAND2_X1 U7403 ( .A1(n8852), .A2(n4352), .ZN(n5854) );
  NAND2_X1 U7404 ( .A1(n7645), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5853) );
  OR2_X2 U7405 ( .A1(n5897), .A2(n7502), .ZN(n7701) );
  NAND2_X1 U7406 ( .A1(n5897), .A2(n7502), .ZN(n7712) );
  XNOR2_X1 U7407 ( .A(n5855), .B(n7697), .ZN(n9094) );
  NAND2_X1 U7408 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  AND2_X1 U7409 ( .A1(n5858), .A2(n6519), .ZN(n5860) );
  NAND2_X1 U7410 ( .A1(n5860), .A2(n5859), .ZN(n9737) );
  INV_X1 U7411 ( .A(n9787), .ZN(n5861) );
  INV_X1 U7412 ( .A(n5862), .ZN(n7666) );
  INV_X1 U7413 ( .A(n6556), .ZN(n6755) );
  NAND2_X1 U7414 ( .A1(n7666), .A2(n6524), .ZN(n5865) );
  OR2_X1 U7415 ( .A1(n9013), .A2(n7745), .ZN(n5864) );
  NAND2_X1 U7416 ( .A1(n5865), .A2(n5864), .ZN(n6585) );
  INV_X1 U7417 ( .A(n6587), .ZN(n7667) );
  OR2_X1 U7418 ( .A1(n5814), .A2(n5813), .ZN(n5866) );
  NAND2_X1 U7419 ( .A1(n9012), .A2(n6813), .ZN(n7751) );
  OR2_X1 U7420 ( .A1(n9012), .A2(n6813), .ZN(n5867) );
  NAND2_X1 U7421 ( .A1(n4349), .A2(n6806), .ZN(n7750) );
  NAND2_X1 U7422 ( .A1(n6798), .A2(n7750), .ZN(n7550) );
  OR2_X1 U7423 ( .A1(n4349), .A2(n6806), .ZN(n7534) );
  NAND2_X1 U7424 ( .A1(n7550), .A2(n7534), .ZN(n7532) );
  INV_X1 U7425 ( .A(n7535), .ZN(n5868) );
  OAI21_X1 U7426 ( .B1(n7532), .B2(n5868), .A(n7752), .ZN(n6882) );
  INV_X1 U7427 ( .A(n9008), .ZN(n7165) );
  NAND2_X1 U7428 ( .A1(n7138), .A2(n7165), .ZN(n7554) );
  NAND2_X1 U7429 ( .A1(n7573), .A2(n7554), .ZN(n7678) );
  INV_X1 U7430 ( .A(n7675), .ZN(n5869) );
  OR2_X1 U7431 ( .A1(n7138), .A2(n7165), .ZN(n9742) );
  NAND2_X1 U7432 ( .A1(n7563), .A2(n9742), .ZN(n7559) );
  NAND2_X1 U7433 ( .A1(n7559), .A2(n7573), .ZN(n5870) );
  NAND2_X1 U7434 ( .A1(n5871), .A2(n5870), .ZN(n7757) );
  NAND2_X1 U7435 ( .A1(n7555), .A2(n7543), .ZN(n5872) );
  OR2_X1 U7436 ( .A1(n7559), .A2(n5872), .ZN(n7754) );
  NAND2_X1 U7437 ( .A1(n7757), .A2(n7754), .ZN(n5873) );
  INV_X1 U7438 ( .A(n7679), .ZN(n7049) );
  INV_X1 U7439 ( .A(n7581), .ZN(n5874) );
  NOR2_X1 U7440 ( .A1(n7201), .A2(n5874), .ZN(n5875) );
  NAND2_X1 U7441 ( .A1(n7203), .A2(n5875), .ZN(n5876) );
  NAND2_X1 U7442 ( .A1(n5876), .A2(n7574), .ZN(n7218) );
  INV_X1 U7443 ( .A(n7222), .ZN(n7682) );
  NAND2_X1 U7444 ( .A1(n7218), .A2(n7682), .ZN(n7279) );
  INV_X1 U7445 ( .A(n7575), .ZN(n5877) );
  NOR2_X1 U7446 ( .A1(n7684), .A2(n5877), .ZN(n5878) );
  NAND2_X1 U7447 ( .A1(n7279), .A2(n5878), .ZN(n7280) );
  INV_X1 U7448 ( .A(n9005), .ZN(n7284) );
  OR2_X1 U7449 ( .A1(n7344), .A2(n7284), .ZN(n7591) );
  NAND2_X1 U7450 ( .A1(n7344), .A2(n7284), .ZN(n7765) );
  NAND2_X1 U7451 ( .A1(n7591), .A2(n7765), .ZN(n7685) );
  INV_X1 U7452 ( .A(n7761), .ZN(n7567) );
  NOR2_X1 U7453 ( .A1(n7685), .A2(n7567), .ZN(n7590) );
  INV_X1 U7454 ( .A(n9302), .ZN(n8908) );
  OR2_X1 U7455 ( .A1(n7443), .A2(n8908), .ZN(n7769) );
  NAND2_X1 U7456 ( .A1(n7443), .A2(n8908), .ZN(n7764) );
  NAND2_X1 U7457 ( .A1(n7769), .A2(n7764), .ZN(n7686) );
  INV_X1 U7458 ( .A(n9290), .ZN(n9300) );
  NAND2_X1 U7459 ( .A1(n9299), .A2(n9300), .ZN(n9298) );
  INV_X1 U7460 ( .A(n9301), .ZN(n7600) );
  XNOR2_X1 U7461 ( .A(n9285), .B(n7600), .ZN(n7689) );
  OR2_X1 U7462 ( .A1(n9285), .A2(n7600), .ZN(n7602) );
  INV_X1 U7463 ( .A(n9242), .ZN(n9392) );
  OR2_X1 U7464 ( .A1(n9386), .A2(n9392), .ZN(n7776) );
  NAND2_X1 U7465 ( .A1(n9386), .A2(n9392), .ZN(n7599) );
  NAND2_X1 U7466 ( .A1(n9262), .A2(n7599), .ZN(n9239) );
  INV_X1 U7467 ( .A(n9265), .ZN(n8967) );
  OR2_X1 U7468 ( .A1(n9245), .A2(n8967), .ZN(n7777) );
  NAND2_X1 U7469 ( .A1(n9245), .A2(n8967), .ZN(n7782) );
  NAND2_X1 U7470 ( .A1(n9239), .A2(n9240), .ZN(n9238) );
  INV_X1 U7471 ( .A(n9364), .ZN(n9217) );
  XNOR2_X1 U7472 ( .A(n9234), .B(n9217), .ZN(n9227) );
  OR2_X1 U7473 ( .A1(n9234), .A2(n9217), .ZN(n7608) );
  XNOR2_X1 U7474 ( .A(n9222), .B(n9355), .ZN(n9209) );
  NAND2_X1 U7475 ( .A1(n9222), .A2(n9375), .ZN(n7610) );
  NAND2_X1 U7476 ( .A1(n9206), .A2(n7610), .ZN(n9191) );
  INV_X1 U7477 ( .A(n9365), .ZN(n9181) );
  OR2_X1 U7478 ( .A1(n9203), .A2(n9181), .ZN(n7615) );
  NAND2_X1 U7479 ( .A1(n9203), .A2(n9181), .ZN(n7614) );
  NAND2_X1 U7480 ( .A1(n9191), .A2(n9195), .ZN(n5879) );
  NAND2_X1 U7481 ( .A1(n5879), .A2(n7614), .ZN(n9172) );
  INV_X1 U7482 ( .A(n9356), .ZN(n5880) );
  OR2_X2 U7483 ( .A1(n9187), .A2(n5880), .ZN(n7620) );
  NAND2_X1 U7484 ( .A1(n9172), .A2(n9173), .ZN(n5881) );
  OR2_X2 U7485 ( .A1(n5882), .A2(n8900), .ZN(n7705) );
  NAND2_X1 U7486 ( .A1(n9148), .A2(n9326), .ZN(n7725) );
  NAND2_X1 U7487 ( .A1(n5884), .A2(n7725), .ZN(n9125) );
  XNOR2_X1 U7488 ( .A(n9127), .B(n9140), .ZN(n9124) );
  NAND2_X1 U7489 ( .A1(n9125), .A2(n9124), .ZN(n9123) );
  NAND2_X1 U7490 ( .A1(n9127), .A2(n9316), .ZN(n7711) );
  INV_X1 U7491 ( .A(n9111), .ZN(n7693) );
  NAND2_X1 U7492 ( .A1(n7504), .A2(n9317), .ZN(n7638) );
  XNOR2_X1 U7493 ( .A(n5885), .B(n7697), .ZN(n5895) );
  OR2_X1 U7494 ( .A1(n5747), .A2(n5886), .ZN(n7663) );
  NAND2_X1 U7495 ( .A1(n7746), .A2(n4909), .ZN(n7661) );
  INV_X1 U7496 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9313) );
  OR2_X1 U7497 ( .A1(n6498), .A2(n9313), .ZN(n5891) );
  INV_X1 U7498 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7499 ( .A1(n4361), .A2(n5887), .ZN(n5890) );
  INV_X1 U7500 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9419) );
  OR2_X1 U7501 ( .A1(n5888), .A2(n9419), .ZN(n5889) );
  INV_X1 U7502 ( .A(n7735), .ZN(n5892) );
  NOR2_X2 U7503 ( .A1(n5892), .A2(n4355), .ZN(n9805) );
  NAND2_X1 U7504 ( .A1(n4358), .A2(P1_B_REG_SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7505 ( .A1(n9805), .A2(n5894), .ZN(n9074) );
  OAI22_X1 U7506 ( .A1(n5895), .A2(n9746), .B1(n7664), .B2(n9074), .ZN(n5896)
         );
  INV_X1 U7507 ( .A(n5896), .ZN(n9096) );
  NAND2_X1 U7508 ( .A1(n7735), .A2(n4355), .ZN(n9738) );
  INV_X1 U7509 ( .A(n9187), .ZN(n9440) );
  INV_X1 U7510 ( .A(n9386), .ZN(n9261) );
  AND2_X1 U7511 ( .A1(n6589), .A2(n5813), .ZN(n6648) );
  NAND2_X1 U7512 ( .A1(n6648), .A2(n6813), .ZN(n6804) );
  INV_X1 U7513 ( .A(n7537), .ZN(n9778) );
  AND2_X1 U7514 ( .A1(n6890), .A2(n9778), .ZN(n6901) );
  INV_X1 U7515 ( .A(n6961), .ZN(n6970) );
  INV_X1 U7516 ( .A(n9797), .ZN(n7318) );
  NAND2_X1 U7517 ( .A1(n9440), .A2(n9182), .ZN(n9183) );
  AOI21_X1 U7518 ( .B1(n9090), .B2(n7503), .A(n9291), .ZN(n5900) );
  NAND2_X1 U7519 ( .A1(n5900), .A2(n9079), .ZN(n9092) );
  OAI21_X1 U7520 ( .B1(n9317), .B2(n9738), .A(n9092), .ZN(n5901) );
  INV_X1 U7521 ( .A(n5901), .ZN(n5902) );
  NAND2_X1 U7522 ( .A1(n9096), .A2(n5902), .ZN(n5903) );
  AOI21_X1 U7523 ( .B1(n9094), .B2(n9812), .A(n5903), .ZN(n5912) );
  NAND3_X1 U7524 ( .A1(n5905), .A2(n5904), .A3(n6744), .ZN(n5907) );
  MUX2_X1 U7525 ( .A(n5908), .B(n5912), .S(n9826), .Z(n5909) );
  NAND2_X1 U7526 ( .A1(n5909), .A2(n4915), .ZN(P1_U3551) );
  INV_X1 U7527 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5913) );
  MUX2_X1 U7528 ( .A(n5913), .B(n5912), .S(n9816), .Z(n5914) );
  NAND2_X1 U7529 ( .A1(n5914), .A2(n4914), .ZN(P1_U3519) );
  NOR2_X4 U7530 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5980) );
  INV_X2 U7531 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U7532 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5923) );
  NOR2_X1 U7533 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5922) );
  NAND3_X1 U7534 ( .A1(n6354), .A2(n6377), .A3(n6352), .ZN(n5926) );
  NAND2_X1 U7535 ( .A1(n6346), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7536 ( .A1(n5934), .A2(n5933), .ZN(n6303) );
  NAND2_X1 U7537 ( .A1(n7172), .A2(n8115), .ZN(n5936) );
  INV_X1 U7538 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7233) );
  OR2_X1 U7539 ( .A1(n4353), .A2(n7233), .ZN(n5935) );
  INV_X1 U7540 ( .A(n8050), .ZN(n8729) );
  NAND2_X1 U7541 ( .A1(n5940), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7542 ( .A1(n6270), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5945) );
  NAND2_X2 U7543 ( .A1(n5949), .A2(n5943), .ZN(n5989) );
  INV_X4 U7544 ( .A(n5989), .ZN(n6305) );
  NAND2_X1 U7545 ( .A1(n6305), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5944) );
  AND2_X1 U7546 ( .A1(n5945), .A2(n5944), .ZN(n5953) );
  NAND2_X1 U7547 ( .A1(n6013), .A2(n6014), .ZN(n6026) );
  NAND2_X1 U7548 ( .A1(n6122), .A2(n6121), .ZN(n6133) );
  NOR2_X1 U7549 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5946) );
  INV_X1 U7550 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7551 ( .A1(n6224), .A2(n5947), .ZN(n5948) );
  NAND2_X1 U7552 ( .A1(n6233), .A2(n5948), .ZN(n8578) );
  OR2_X2 U7553 ( .A1(n5949), .A2(n8856), .ZN(n5974) );
  NAND2_X1 U7554 ( .A1(n8578), .A2(n4357), .ZN(n5952) );
  INV_X1 U7555 ( .A(n5949), .ZN(n5950) );
  NAND2_X1 U7556 ( .A1(n6001), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7557 ( .A1(n5973), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5957) );
  INV_X1 U7558 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6402) );
  INV_X1 U7559 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6691) );
  OR2_X1 U7560 ( .A1(n5974), .A2(n6691), .ZN(n5955) );
  OR2_X1 U7561 ( .A1(n5961), .A2(n6847), .ZN(n5954) );
  INV_X1 U7562 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5959) );
  INV_X1 U7563 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U7564 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5958) );
  NAND2_X1 U7565 ( .A1(n9923), .A2(n6845), .ZN(n8169) );
  INV_X1 U7566 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5960) );
  INV_X1 U7567 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10098) );
  OR2_X1 U7568 ( .A1(n5974), .A2(n10098), .ZN(n5964) );
  INV_X1 U7569 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6791) );
  OR2_X1 U7570 ( .A1(n5961), .A2(n6791), .ZN(n5963) );
  NAND2_X1 U7571 ( .A1(n5973), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5962) );
  INV_X1 U7572 ( .A(n6317), .ZN(n6608) );
  NAND2_X1 U7573 ( .A1(n5064), .A2(SI_0_), .ZN(n5967) );
  INV_X1 U7574 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7575 ( .A1(n5967), .A2(n5966), .ZN(n5969) );
  AND2_X1 U7576 ( .A1(n5969), .A2(n5968), .ZN(n8857) );
  MUX2_X1 U7577 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8857), .S(n5970), .Z(n6788) );
  NAND2_X1 U7578 ( .A1(n6757), .A2(n6761), .ZN(n5972) );
  NAND2_X1 U7579 ( .A1(n9923), .A2(n6687), .ZN(n5971) );
  NAND2_X1 U7580 ( .A1(n5972), .A2(n5971), .ZN(n9915) );
  INV_X1 U7581 ( .A(n5961), .ZN(n6001) );
  NAND2_X1 U7582 ( .A1(n6001), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7583 ( .A1(n5973), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5978) );
  INV_X1 U7584 ( .A(n5974), .ZN(n5975) );
  NAND2_X1 U7585 ( .A1(n4356), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7586 ( .A1(n6305), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5976) );
  OR2_X1 U7587 ( .A1(n4353), .A2(n5036), .ZN(n5985) );
  OR2_X1 U7588 ( .A1(n5995), .A2(n6459), .ZN(n5984) );
  OR2_X1 U7589 ( .A1(n5970), .A2(n4350), .ZN(n5983) );
  NAND2_X1 U7590 ( .A1(n4354), .A2(n9930), .ZN(n8155) );
  NAND2_X1 U7591 ( .A1(n9915), .A2(n6319), .ZN(n5988) );
  INV_X1 U7592 ( .A(n9930), .ZN(n9938) );
  OR2_X1 U7593 ( .A1(n4354), .A2(n9938), .ZN(n5987) );
  NAND2_X1 U7594 ( .A1(n5988), .A2(n5987), .ZN(n6723) );
  NAND2_X1 U7595 ( .A1(n5973), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5993) );
  INV_X1 U7596 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6400) );
  OR2_X1 U7597 ( .A1(n5989), .A2(n6400), .ZN(n5992) );
  OR2_X1 U7598 ( .A1(n5974), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5991) );
  INV_X1 U7599 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6401) );
  OR2_X1 U7600 ( .A1(n5961), .A2(n6401), .ZN(n5990) );
  INV_X1 U7601 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6454) );
  OR2_X1 U7602 ( .A1(n4353), .A2(n6454), .ZN(n5997) );
  OR2_X1 U7603 ( .A1(n5995), .A2(n6465), .ZN(n5996) );
  OAI211_X1 U7604 ( .C1(n5970), .C2(n6536), .A(n5997), .B(n5996), .ZN(n7105)
         );
  NAND2_X1 U7605 ( .A1(n9921), .A2(n7105), .ZN(n8181) );
  NAND2_X1 U7606 ( .A1(n8181), .A2(n8174), .ZN(n8122) );
  NAND2_X1 U7607 ( .A1(n6723), .A2(n8122), .ZN(n5999) );
  NAND2_X1 U7608 ( .A1(n9921), .A2(n6994), .ZN(n5998) );
  NAND2_X1 U7609 ( .A1(n6305), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7610 ( .A1(n5973), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6004) );
  AND2_X1 U7611 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6000) );
  NOR2_X1 U7612 ( .A1(n6013), .A2(n6000), .ZN(n7020) );
  OR2_X1 U7613 ( .A1(n5974), .A2(n7020), .ZN(n6003) );
  NAND2_X1 U7614 ( .A1(n6001), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6002) );
  NAND4_X1 U7615 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n8335)
         );
  NAND2_X1 U7616 ( .A1(n6006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  INV_X1 U7617 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7618 ( .A(n6008), .B(n6007), .ZN(n6929) );
  OR2_X1 U7619 ( .A1(n5995), .A2(n6461), .ZN(n6010) );
  OR2_X1 U7620 ( .A1(n4353), .A2(n5107), .ZN(n6009) );
  OAI211_X1 U7621 ( .C1(n5970), .C2(n6929), .A(n6010), .B(n6009), .ZN(n6836)
         );
  NOR2_X1 U7622 ( .A1(n8335), .A2(n6836), .ZN(n6012) );
  NAND2_X1 U7623 ( .A1(n8335), .A2(n6836), .ZN(n6011) );
  NAND2_X1 U7624 ( .A1(n6305), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7625 ( .A1(n5973), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7626 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  AND2_X1 U7627 ( .A1(n6026), .A2(n6015), .ZN(n7029) );
  OR2_X1 U7628 ( .A1(n5974), .A2(n7029), .ZN(n6018) );
  INV_X1 U7629 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6016) );
  NAND4_X1 U7630 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n8334)
         );
  OR2_X1 U7631 ( .A1(n6021), .A2(n8847), .ZN(n6022) );
  XNOR2_X1 U7632 ( .A(n6022), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6930) );
  OR2_X1 U7633 ( .A1(n5995), .A2(n6463), .ZN(n6024) );
  INV_X1 U7634 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6457) );
  OR2_X1 U7635 ( .A1(n4353), .A2(n6457), .ZN(n6023) );
  OAI211_X1 U7636 ( .C1(n5970), .C2(n9870), .A(n6024), .B(n6023), .ZN(n6985)
         );
  INV_X1 U7637 ( .A(n6985), .ZN(n9948) );
  NAND2_X1 U7638 ( .A1(n6305), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6031) );
  INV_X1 U7639 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6025) );
  OR2_X1 U7640 ( .A1(n6040), .A2(n6025), .ZN(n6030) );
  NAND2_X1 U7641 ( .A1(n6026), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6027) );
  AND2_X1 U7642 ( .A1(n6038), .A2(n6027), .ZN(n7152) );
  OR2_X1 U7643 ( .A1(n6157), .A2(n7152), .ZN(n6029) );
  INV_X1 U7644 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6915) );
  OR2_X1 U7645 ( .A1(n6308), .A2(n6915), .ZN(n6028) );
  NAND2_X1 U7646 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  MUX2_X1 U7647 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6033), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n6034) );
  NAND2_X1 U7648 ( .A1(n6034), .A2(n4372), .ZN(n6933) );
  OR2_X1 U7649 ( .A1(n5995), .A2(n6467), .ZN(n6036) );
  OR2_X1 U7650 ( .A1(n4353), .A2(n6501), .ZN(n6035) );
  OAI211_X1 U7651 ( .C1(n5970), .C2(n6933), .A(n6036), .B(n6035), .ZN(n7046)
         );
  NAND2_X1 U7652 ( .A1(n7194), .A2(n7046), .ZN(n8179) );
  INV_X1 U7653 ( .A(n7046), .ZN(n9953) );
  NAND2_X1 U7654 ( .A1(n8333), .A2(n9953), .ZN(n8188) );
  NAND2_X1 U7655 ( .A1(n8179), .A2(n8188), .ZN(n7154) );
  NAND2_X1 U7656 ( .A1(n7155), .A2(n7154), .ZN(n7153) );
  NAND2_X1 U7657 ( .A1(n8333), .A2(n7046), .ZN(n6037) );
  NAND2_X1 U7658 ( .A1(n6305), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6044) );
  AND2_X1 U7659 ( .A1(n6038), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6039) );
  NOR2_X1 U7660 ( .A1(n6052), .A2(n6039), .ZN(n7199) );
  OR2_X1 U7661 ( .A1(n5974), .A2(n7199), .ZN(n6043) );
  INV_X1 U7662 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7184) );
  OR2_X1 U7663 ( .A1(n6308), .A2(n7184), .ZN(n6042) );
  INV_X2 U7664 ( .A(n6040), .ZN(n6270) );
  NAND2_X1 U7665 ( .A1(n6270), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6041) );
  NAND4_X1 U7666 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(n8332)
         );
  OR2_X1 U7667 ( .A1(n5995), .A2(n6471), .ZN(n6050) );
  INV_X1 U7668 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6470) );
  OR2_X1 U7669 ( .A1(n4353), .A2(n6470), .ZN(n6049) );
  NAND2_X1 U7670 ( .A1(n4372), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6045) );
  MUX2_X1 U7671 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6045), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6047) );
  AND2_X1 U7672 ( .A1(n6047), .A2(n6046), .ZN(n7074) );
  OR2_X1 U7673 ( .A1(n5970), .A2(n7060), .ZN(n6048) );
  XNOR2_X1 U7674 ( .A(n8332), .B(n9957), .ZN(n8193) );
  INV_X1 U7675 ( .A(n8332), .ZN(n7043) );
  NAND2_X1 U7676 ( .A1(n7043), .A2(n9957), .ZN(n6051) );
  NAND2_X1 U7677 ( .A1(n6305), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7678 ( .A1(n6270), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6056) );
  NOR2_X1 U7679 ( .A1(n6052), .A2(n7255), .ZN(n6053) );
  OR2_X1 U7680 ( .A1(n6069), .A2(n6053), .ZN(n7260) );
  NAND2_X1 U7681 ( .A1(n4357), .A2(n7260), .ZN(n6055) );
  NAND2_X1 U7682 ( .A1(n6001), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6054) );
  NAND4_X1 U7683 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n8331)
         );
  OR2_X1 U7684 ( .A1(n6474), .A2(n5995), .ZN(n6062) );
  NAND2_X1 U7685 ( .A1(n6046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6059) );
  INV_X1 U7686 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7687 ( .A(n6059), .B(n6058), .ZN(n9893) );
  OR2_X1 U7688 ( .A1(n4360), .A2(n9893), .ZN(n6061) );
  OR2_X1 U7689 ( .A1(n4353), .A2(n6473), .ZN(n6060) );
  NAND2_X1 U7690 ( .A1(n8331), .A2(n9962), .ZN(n8194) );
  NAND2_X1 U7691 ( .A1(n6064), .A2(n6063), .ZN(n7236) );
  INV_X1 U7692 ( .A(n9962), .ZN(n6065) );
  NAND2_X1 U7693 ( .A1(n8331), .A2(n6065), .ZN(n6066) );
  NAND2_X1 U7694 ( .A1(n6270), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6074) );
  INV_X1 U7695 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6067) );
  OR2_X1 U7696 ( .A1(n5989), .A2(n6067), .ZN(n6073) );
  OR2_X1 U7697 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  AND2_X1 U7698 ( .A1(n6087), .A2(n6070), .ZN(n7326) );
  OR2_X1 U7699 ( .A1(n6157), .A2(n7326), .ZN(n6072) );
  INV_X1 U7700 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7327) );
  OR2_X1 U7701 ( .A1(n6308), .A2(n7327), .ZN(n6071) );
  NAND2_X1 U7702 ( .A1(n6475), .A2(n8115), .ZN(n6077) );
  NOR2_X1 U7703 ( .A1(n6046), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6080) );
  INV_X1 U7704 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8847) );
  OR2_X1 U7705 ( .A1(n6080), .A2(n8847), .ZN(n6075) );
  XNOR2_X1 U7706 ( .A(n6075), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7125) );
  AOI22_X1 U7707 ( .A1(n6204), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6399), .B2(
        n7125), .ZN(n6076) );
  NAND2_X1 U7708 ( .A1(n6077), .A2(n6076), .ZN(n7265) );
  NAND2_X1 U7709 ( .A1(n7458), .A2(n7265), .ZN(n8200) );
  NAND2_X1 U7710 ( .A1(n8330), .A2(n7492), .ZN(n8195) );
  NAND2_X1 U7711 ( .A1(n8200), .A2(n8195), .ZN(n8127) );
  NAND2_X1 U7712 ( .A1(n7458), .A2(n7492), .ZN(n6078) );
  NAND2_X1 U7713 ( .A1(n6481), .A2(n8115), .ZN(n6086) );
  INV_X1 U7714 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6079) );
  NOR2_X1 U7715 ( .A1(n6083), .A2(n8847), .ZN(n6081) );
  MUX2_X1 U7716 ( .A(n8847), .B(n6081), .S(P2_IR_REG_10__SCAN_IN), .Z(n6084)
         );
  INV_X1 U7717 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6082) );
  AOI22_X1 U7718 ( .A1(n6204), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6399), .B2(
        n7382), .ZN(n6085) );
  NAND2_X1 U7719 ( .A1(n6086), .A2(n6085), .ZN(n7456) );
  NAND2_X1 U7720 ( .A1(n6305), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7721 ( .A1(n6270), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7722 ( .A1(n6087), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6088) );
  AND2_X1 U7723 ( .A1(n6097), .A2(n6088), .ZN(n7464) );
  OR2_X1 U7724 ( .A1(n5974), .A2(n7464), .ZN(n6090) );
  NAND2_X1 U7725 ( .A1(n6001), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6089) );
  NAND4_X1 U7726 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n8329)
         );
  NAND2_X1 U7727 ( .A1(n7456), .A2(n8329), .ZN(n7347) );
  OR2_X1 U7728 ( .A1(n8329), .A2(n7456), .ZN(n7348) );
  NAND2_X1 U7729 ( .A1(n6093), .A2(n7348), .ZN(n7475) );
  NAND2_X1 U7730 ( .A1(n6506), .A2(n8115), .ZN(n6096) );
  OR2_X1 U7731 ( .A1(n6104), .A2(n8847), .ZN(n6094) );
  XNOR2_X1 U7732 ( .A(n6094), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7386) );
  AOI22_X1 U7733 ( .A1(n6204), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6399), .B2(
        n7386), .ZN(n6095) );
  NAND2_X1 U7734 ( .A1(n6096), .A2(n6095), .ZN(n9978) );
  NAND2_X1 U7735 ( .A1(n6305), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7736 ( .A1(n6270), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7737 ( .A1(n6097), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6098) );
  AND2_X1 U7738 ( .A1(n6108), .A2(n6098), .ZN(n8055) );
  OR2_X1 U7739 ( .A1(n6157), .A2(n8055), .ZN(n6100) );
  NAND2_X1 U7740 ( .A1(n6001), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6099) );
  NAND4_X1 U7741 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n8686)
         );
  NAND2_X1 U7742 ( .A1(n6514), .A2(n8115), .ZN(n6107) );
  INV_X1 U7743 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7744 ( .A1(n6104), .A2(n6103), .ZN(n6117) );
  NAND2_X1 U7745 ( .A1(n6117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6105) );
  XNOR2_X1 U7746 ( .A(n6105), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7390) );
  AOI22_X1 U7747 ( .A1(n6204), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6399), .B2(
        n7390), .ZN(n6106) );
  NAND2_X1 U7748 ( .A1(n6107), .A2(n6106), .ZN(n9984) );
  NAND2_X1 U7749 ( .A1(n6270), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6113) );
  INV_X1 U7750 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7376) );
  OR2_X1 U7751 ( .A1(n5989), .A2(n7376), .ZN(n6112) );
  AND2_X1 U7752 ( .A1(n6108), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6109) );
  NOR2_X1 U7753 ( .A1(n6122), .A2(n6109), .ZN(n7977) );
  OR2_X1 U7754 ( .A1(n6157), .A2(n7977), .ZN(n6111) );
  INV_X1 U7755 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7388) );
  OR2_X1 U7756 ( .A1(n6308), .A2(n7388), .ZN(n6110) );
  OR2_X1 U7757 ( .A1(n9984), .A2(n9558), .ZN(n8219) );
  NAND2_X1 U7758 ( .A1(n9984), .A2(n9558), .ZN(n8218) );
  NAND2_X1 U7759 ( .A1(n8219), .A2(n8218), .ZN(n8222) );
  OAI21_X1 U7760 ( .B1(n9978), .B2(n8686), .A(n8222), .ZN(n6116) );
  AND2_X1 U7761 ( .A1(n9978), .A2(n8686), .ZN(n6114) );
  INV_X1 U7762 ( .A(n9558), .ZN(n8328) );
  AOI22_X1 U7763 ( .A1(n8222), .A2(n6114), .B1(n8328), .B2(n9984), .ZN(n6115)
         );
  NAND2_X1 U7764 ( .A1(n6522), .A2(n8115), .ZN(n6120) );
  NAND2_X1 U7765 ( .A1(n6118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7766 ( .A(n6129), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8376) );
  AOI22_X1 U7767 ( .A1(n6204), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6399), .B2(
        n8376), .ZN(n6119) );
  NAND2_X1 U7768 ( .A1(n6120), .A2(n6119), .ZN(n9550) );
  NAND2_X1 U7769 ( .A1(n6305), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7770 ( .A1(n6270), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6126) );
  OR2_X1 U7771 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  AND2_X1 U7772 ( .A1(n6123), .A2(n6133), .ZN(n9554) );
  OR2_X1 U7773 ( .A1(n6157), .A2(n9554), .ZN(n6125) );
  NAND2_X1 U7774 ( .A1(n6001), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6124) );
  NAND4_X1 U7775 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n8685)
         );
  OR2_X1 U7776 ( .A1(n9550), .A2(n8685), .ZN(n8133) );
  NAND2_X1 U7777 ( .A1(n9550), .A2(n8685), .ZN(n8132) );
  NAND2_X1 U7778 ( .A1(n6583), .A2(n8115), .ZN(n6132) );
  INV_X1 U7779 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7780 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  NAND2_X1 U7781 ( .A1(n6130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7782 ( .A(n6141), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8380) );
  AOI22_X1 U7783 ( .A1(n6204), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6399), .B2(
        n8380), .ZN(n6131) );
  INV_X1 U7784 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8379) );
  OR2_X1 U7785 ( .A1(n5989), .A2(n8379), .ZN(n6139) );
  NAND2_X1 U7786 ( .A1(n6133), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6134) );
  AND2_X1 U7787 ( .A1(n6146), .A2(n6134), .ZN(n7937) );
  OR2_X1 U7788 ( .A1(n5974), .A2(n7937), .ZN(n6138) );
  INV_X1 U7789 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7790 ( .A1(n6308), .A2(n6135), .ZN(n6137) );
  NAND2_X1 U7791 ( .A1(n6270), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6136) );
  NAND4_X1 U7792 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n8659)
         );
  NAND2_X1 U7793 ( .A1(n6606), .A2(n8115), .ZN(n6145) );
  INV_X1 U7794 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7795 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U7796 ( .A1(n6142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U7797 ( .A(n6143), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8421) );
  AOI22_X1 U7798 ( .A1(n6204), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8421), .B2(
        n6399), .ZN(n6144) );
  INV_X1 U7799 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8752) );
  OR2_X1 U7800 ( .A1(n5989), .A2(n8752), .ZN(n6151) );
  AND2_X1 U7801 ( .A1(n6146), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6147) );
  NOR2_X1 U7802 ( .A1(n6155), .A2(n6147), .ZN(n8090) );
  OR2_X1 U7803 ( .A1(n5974), .A2(n8090), .ZN(n6150) );
  INV_X1 U7804 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8662) );
  OR2_X1 U7805 ( .A1(n6308), .A2(n8662), .ZN(n6149) );
  NAND2_X1 U7806 ( .A1(n6270), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6148) );
  NAND4_X1 U7807 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n8669)
         );
  NAND2_X1 U7808 ( .A1(n8837), .A2(n8669), .ZN(n8643) );
  NAND2_X1 U7809 ( .A1(n6662), .A2(n8115), .ZN(n6154) );
  XNOR2_X1 U7810 ( .A(n6152), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8424) );
  AOI22_X1 U7811 ( .A1(n6204), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6399), .B2(
        n8424), .ZN(n6153) );
  NAND2_X1 U7812 ( .A1(n6270), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6161) );
  INV_X1 U7813 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8750) );
  OR2_X1 U7814 ( .A1(n5989), .A2(n8750), .ZN(n6160) );
  NOR2_X1 U7815 ( .A1(n6155), .A2(n10119), .ZN(n6156) );
  OR2_X1 U7816 ( .A1(n6174), .A2(n6156), .ZN(n8001) );
  INV_X1 U7817 ( .A(n8001), .ZN(n8651) );
  OR2_X1 U7818 ( .A1(n6157), .A2(n8651), .ZN(n6159) );
  INV_X1 U7819 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8652) );
  OR2_X1 U7820 ( .A1(n6308), .A2(n8652), .ZN(n6158) );
  NAND2_X1 U7821 ( .A1(n8749), .A2(n8660), .ZN(n6163) );
  AND2_X1 U7822 ( .A1(n8643), .A2(n6163), .ZN(n6162) );
  NAND2_X1 U7823 ( .A1(n8658), .A2(n6162), .ZN(n6168) );
  INV_X1 U7824 ( .A(n6163), .ZN(n6166) );
  OR2_X1 U7825 ( .A1(n8837), .A2(n8669), .ZN(n8644) );
  INV_X1 U7826 ( .A(n8644), .ZN(n6164) );
  NAND2_X1 U7827 ( .A1(n8749), .A2(n8094), .ZN(n8236) );
  NOR2_X1 U7828 ( .A1(n6164), .A2(n8646), .ZN(n6165) );
  OR2_X1 U7829 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  NAND2_X1 U7830 ( .A1(n6705), .A2(n8115), .ZN(n6172) );
  NAND2_X1 U7831 ( .A1(n6180), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7832 ( .A(n6170), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8460) );
  AOI22_X1 U7833 ( .A1(n6204), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6399), .B2(
        n8460), .ZN(n6171) );
  NAND2_X1 U7834 ( .A1(n6270), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6179) );
  INV_X1 U7835 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8638) );
  OR2_X1 U7836 ( .A1(n6308), .A2(n8638), .ZN(n6178) );
  OR2_X1 U7837 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  AND2_X1 U7838 ( .A1(n6190), .A2(n6175), .ZN(n8009) );
  OR2_X1 U7839 ( .A1(n5974), .A2(n8009), .ZN(n6177) );
  INV_X1 U7840 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8745) );
  OR2_X1 U7841 ( .A1(n5989), .A2(n8745), .ZN(n6176) );
  NAND2_X1 U7842 ( .A1(n8826), .A2(n8650), .ZN(n8241) );
  NAND2_X1 U7843 ( .A1(n8245), .A2(n8241), .ZN(n8635) );
  NAND2_X1 U7844 ( .A1(n6729), .A2(n8115), .ZN(n6189) );
  INV_X1 U7845 ( .A(n6180), .ZN(n6182) );
  NAND2_X1 U7846 ( .A1(n6183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6186) );
  INV_X1 U7847 ( .A(n6186), .ZN(n6184) );
  NAND2_X1 U7848 ( .A1(n6184), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7849 ( .A1(n6186), .A2(n6185), .ZN(n6201) );
  AND2_X1 U7850 ( .A1(n6187), .A2(n6201), .ZN(n8476) );
  AOI22_X1 U7851 ( .A1(n6204), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6399), .B2(
        n8476), .ZN(n6188) );
  NAND2_X1 U7852 ( .A1(n6270), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7853 ( .A1(n6305), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7854 ( .A1(n6190), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6191) );
  AND2_X1 U7855 ( .A1(n6207), .A2(n6191), .ZN(n8067) );
  OR2_X1 U7856 ( .A1(n5974), .A2(n8067), .ZN(n6193) );
  NAND2_X1 U7857 ( .A1(n6001), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6192) );
  NAND4_X1 U7858 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n8636)
         );
  OR2_X1 U7859 ( .A1(n8820), .A2(n8636), .ZN(n6196) );
  AND2_X1 U7860 ( .A1(n8635), .A2(n6196), .ZN(n6200) );
  INV_X1 U7861 ( .A(n6196), .ZN(n6199) );
  INV_X1 U7862 ( .A(n8650), .ZN(n8626) );
  NAND2_X1 U7863 ( .A1(n8826), .A2(n8626), .ZN(n8622) );
  NAND2_X1 U7864 ( .A1(n8820), .A2(n8636), .ZN(n6197) );
  AND2_X1 U7865 ( .A1(n8622), .A2(n6197), .ZN(n6198) );
  NAND2_X1 U7866 ( .A1(n6879), .A2(n8115), .ZN(n6206) );
  NAND2_X1 U7867 ( .A1(n6201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6203) );
  AOI22_X1 U7868 ( .A1(n6204), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8472), .B2(
        n6399), .ZN(n6205) );
  NAND2_X1 U7869 ( .A1(n6270), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7870 ( .A1(n6305), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6211) );
  INV_X1 U7871 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8617) );
  OR2_X1 U7872 ( .A1(n6308), .A2(n8617), .ZN(n6210) );
  AND2_X1 U7873 ( .A1(n6207), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6208) );
  OR2_X1 U7874 ( .A1(n6208), .A2(n6222), .ZN(n8618) );
  NAND2_X1 U7875 ( .A1(n4357), .A2(n8618), .ZN(n6209) );
  NAND4_X1 U7876 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n8627)
         );
  INV_X1 U7877 ( .A(n8814), .ZN(n6213) );
  NAND2_X1 U7878 ( .A1(n6991), .A2(n8115), .ZN(n6215) );
  INV_X1 U7879 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7034) );
  OR2_X1 U7880 ( .A1(n4353), .A2(n7034), .ZN(n6214) );
  INV_X1 U7881 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10208) );
  XNOR2_X1 U7882 ( .A(n6222), .B(n10208), .ZN(n8606) );
  NAND2_X1 U7883 ( .A1(n8606), .A2(n4357), .ZN(n6219) );
  NAND2_X1 U7884 ( .A1(n6305), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7885 ( .A1(n6270), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7886 ( .A1(n6001), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7887 ( .A1(n8735), .A2(n8614), .ZN(n8256) );
  OR2_X1 U7888 ( .A1(n8735), .A2(n8589), .ZN(n8585) );
  NAND2_X1 U7889 ( .A1(n8600), .A2(n8585), .ZN(n6229) );
  NAND2_X1 U7890 ( .A1(n7088), .A2(n8115), .ZN(n6221) );
  INV_X1 U7891 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7136) );
  OR2_X1 U7892 ( .A1(n4353), .A2(n7136), .ZN(n6220) );
  INV_X1 U7893 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10153) );
  AOI21_X1 U7894 ( .B1(n6222), .B2(n10208), .A(n10153), .ZN(n6223) );
  OR2_X1 U7895 ( .A1(n6224), .A2(n6223), .ZN(n8593) );
  NAND2_X1 U7896 ( .A1(n8593), .A2(n4357), .ZN(n6228) );
  NAND2_X1 U7897 ( .A1(n6305), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7898 ( .A1(n6270), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7899 ( .A1(n6001), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7900 ( .A1(n8802), .A2(n8570), .ZN(n8253) );
  NAND2_X1 U7901 ( .A1(n8259), .A2(n8253), .ZN(n8584) );
  NAND2_X1 U7902 ( .A1(n6229), .A2(n8584), .ZN(n8588) );
  INV_X1 U7903 ( .A(n8570), .ZN(n8602) );
  OR2_X1 U7904 ( .A1(n8802), .A2(n8602), .ZN(n8567) );
  NAND2_X1 U7905 ( .A1(n8050), .A2(n7947), .ZN(n8264) );
  NAND2_X1 U7906 ( .A1(n6230), .A2(n8115), .ZN(n6232) );
  INV_X1 U7907 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7232) );
  OR2_X1 U7908 ( .A1(n4353), .A2(n7232), .ZN(n6231) );
  NAND2_X1 U7909 ( .A1(n6233), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7910 ( .A1(n6241), .A2(n6234), .ZN(n8564) );
  NAND2_X1 U7911 ( .A1(n8564), .A2(n4357), .ZN(n6237) );
  AOI22_X1 U7912 ( .A1(n6305), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n6270), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7913 ( .A1(n6001), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6235) );
  NOR2_X1 U7914 ( .A1(n7910), .A2(n8571), .ZN(n6238) );
  NAND2_X1 U7915 ( .A1(n7304), .A2(n8115), .ZN(n6240) );
  INV_X1 U7916 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7335) );
  OR2_X1 U7917 ( .A1(n4353), .A2(n7335), .ZN(n6239) );
  NAND2_X1 U7918 ( .A1(n6241), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7919 ( .A1(n6249), .A2(n6242), .ZN(n8551) );
  NAND2_X1 U7920 ( .A1(n8551), .A2(n4357), .ZN(n6245) );
  AOI22_X1 U7921 ( .A1(n6305), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n6270), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7922 ( .A1(n6001), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7923 ( .A1(n7407), .A2(n8115), .ZN(n6248) );
  INV_X1 U7924 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7804) );
  OR2_X1 U7925 ( .A1(n4353), .A2(n7804), .ZN(n6247) );
  AND2_X1 U7926 ( .A1(n6249), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6250) );
  OR2_X1 U7927 ( .A1(n6250), .A2(n6258), .ZN(n8540) );
  INV_X1 U7928 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U7929 ( .A1(n6305), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7930 ( .A1(n6270), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6251) );
  OAI211_X1 U7931 ( .C1(n8544), .C2(n6308), .A(n6252), .B(n6251), .ZN(n6253)
         );
  NAND2_X1 U7932 ( .A1(n8784), .A2(n8549), .ZN(n8280) );
  NAND2_X1 U7933 ( .A1(n8279), .A2(n8280), .ZN(n8543) );
  NAND2_X1 U7934 ( .A1(n8537), .A2(n8543), .ZN(n8536) );
  INV_X1 U7935 ( .A(n8549), .ZN(n8326) );
  NAND2_X1 U7936 ( .A1(n7450), .A2(n8115), .ZN(n6256) );
  INV_X1 U7937 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7453) );
  OR2_X1 U7938 ( .A1(n4353), .A2(n7453), .ZN(n6255) );
  INV_X1 U7939 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7940 ( .A1(n6258), .A2(n6257), .ZN(n6268) );
  OR2_X1 U7941 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  NAND2_X1 U7942 ( .A1(n6268), .A2(n6259), .ZN(n8529) );
  NAND2_X1 U7943 ( .A1(n8529), .A2(n4357), .ZN(n6264) );
  INV_X1 U7944 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U7945 ( .A1(n6305), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7946 ( .A1(n6270), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6260) );
  OAI211_X1 U7947 ( .C1(n8530), .C2(n6308), .A(n6261), .B(n6260), .ZN(n6262)
         );
  INV_X1 U7948 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U7949 ( .A1(n8712), .A2(n8538), .ZN(n8143) );
  NOR2_X1 U7950 ( .A1(n8712), .A2(n8538), .ZN(n8145) );
  NAND2_X1 U7951 ( .A1(n7480), .A2(n8115), .ZN(n6267) );
  INV_X1 U7952 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6265) );
  OR2_X1 U7953 ( .A1(n4353), .A2(n6265), .ZN(n6266) );
  NAND2_X1 U7954 ( .A1(n6268), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7955 ( .A1(n6280), .A2(n6269), .ZN(n8520) );
  NAND2_X1 U7956 ( .A1(n8520), .A2(n4357), .ZN(n6275) );
  INV_X1 U7957 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U7958 ( .A1(n6305), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7959 ( .A1(n6270), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U7960 ( .C1(n8519), .C2(n6308), .A(n6272), .B(n6271), .ZN(n6273)
         );
  INV_X1 U7961 ( .A(n6273), .ZN(n6274) );
  NAND2_X1 U7962 ( .A1(n6277), .A2(n8115), .ZN(n6279) );
  INV_X1 U7963 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7498) );
  OR2_X1 U7964 ( .A1(n4353), .A2(n7498), .ZN(n6278) );
  AND2_X1 U7965 ( .A1(n6280), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6281) );
  INV_X1 U7966 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U7967 ( .A1(n6305), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7968 ( .A1(n6270), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6282) );
  OAI211_X1 U7969 ( .C1(n8510), .C2(n6308), .A(n6283), .B(n6282), .ZN(n6284)
         );
  AOI21_X1 U7970 ( .B1(n8511), .B2(n4357), .A(n6284), .ZN(n8153) );
  NAND2_X1 U7971 ( .A1(n8852), .A2(n8115), .ZN(n6286) );
  OR2_X1 U7972 ( .A1(n4353), .A2(n8854), .ZN(n6285) );
  NAND2_X1 U7973 ( .A1(n8492), .A2(n4357), .ZN(n8113) );
  INV_X1 U7974 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7975 ( .A1(n6270), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7976 ( .A1(n6305), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6287) );
  OAI211_X1 U7977 ( .C1(n6308), .C2(n6289), .A(n6288), .B(n6287), .ZN(n6290)
         );
  INV_X1 U7978 ( .A(n6290), .ZN(n6291) );
  NAND2_X1 U7979 ( .A1(n8291), .A2(n8503), .ZN(n8105) );
  NAND2_X1 U7980 ( .A1(n8293), .A2(n8105), .ZN(n6337) );
  XNOR2_X1 U7981 ( .A(n6292), .B(n6337), .ZN(n6316) );
  NAND2_X1 U7982 ( .A1(n6294), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6295) );
  MUX2_X1 U7983 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6295), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6297) );
  NAND2_X1 U7984 ( .A1(n6673), .A2(n8299), .ZN(n8118) );
  INV_X1 U7985 ( .A(n6298), .ZN(n6299) );
  NAND2_X1 U7986 ( .A1(n6299), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7987 ( .A1(n8472), .A2(n8319), .ZN(n6301) );
  INV_X1 U7988 ( .A(n6302), .ZN(n6410) );
  INV_X1 U7989 ( .A(n8473), .ZN(n8317) );
  NAND2_X1 U7990 ( .A1(n6410), .A2(n8317), .ZN(n6304) );
  NAND2_X1 U7991 ( .A1(n5970), .A2(n6304), .ZN(n6312) );
  INV_X1 U7992 ( .A(n6312), .ZN(n6685) );
  INV_X1 U7993 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7994 ( .A1(n6305), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7995 ( .A1(n6270), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6306) );
  OAI211_X1 U7996 ( .C1(n6309), .C2(n6308), .A(n6307), .B(n6306), .ZN(n6310)
         );
  INV_X1 U7997 ( .A(n6310), .ZN(n6311) );
  NAND2_X1 U7998 ( .A1(n8113), .A2(n6311), .ZN(n8324) );
  AND2_X1 U7999 ( .A1(n5970), .A2(P2_B_REG_SCAN_IN), .ZN(n6313) );
  NOR2_X1 U8000 ( .A1(n9920), .A2(n6313), .ZN(n8493) );
  AOI22_X1 U8001 ( .A1(n8517), .A2(n8687), .B1(n8324), .B2(n8493), .ZN(n6314)
         );
  INV_X1 U8002 ( .A(n6757), .ZN(n6318) );
  NAND2_X1 U8003 ( .A1(n6318), .A2(n6759), .ZN(n6758) );
  NAND2_X1 U8004 ( .A1(n6758), .A2(n8169), .ZN(n9918) );
  NAND2_X1 U8005 ( .A1(n9916), .A2(n8154), .ZN(n6722) );
  INV_X1 U8006 ( .A(n8122), .ZN(n6724) );
  NAND2_X1 U8007 ( .A1(n6722), .A2(n6724), .ZN(n6721) );
  NAND2_X1 U8008 ( .A1(n6721), .A2(n8181), .ZN(n7018) );
  INV_X1 U8009 ( .A(n8335), .ZN(n6831) );
  NAND2_X1 U8010 ( .A1(n6831), .A2(n6836), .ZN(n8175) );
  INV_X1 U8011 ( .A(n6836), .ZN(n9944) );
  NAND2_X1 U8012 ( .A1(n8335), .A2(n9944), .ZN(n8183) );
  NAND2_X1 U8013 ( .A1(n7018), .A2(n8172), .ZN(n6320) );
  NAND2_X1 U8014 ( .A1(n6320), .A2(n8175), .ZN(n7028) );
  NAND2_X1 U8015 ( .A1(n7044), .A2(n6985), .ZN(n8176) );
  NAND2_X1 U8016 ( .A1(n8334), .A2(n9948), .ZN(n8182) );
  AND2_X1 U8017 ( .A1(n8176), .A2(n8179), .ZN(n8186) );
  NAND2_X1 U8018 ( .A1(n7150), .A2(n8186), .ZN(n7175) );
  NAND2_X1 U8019 ( .A1(n7175), .A2(n8188), .ZN(n6322) );
  INV_X1 U8020 ( .A(n8193), .ZN(n6321) );
  NAND2_X1 U8021 ( .A1(n6322), .A2(n6321), .ZN(n7174) );
  NAND2_X1 U8022 ( .A1(n8332), .A2(n9957), .ZN(n7242) );
  AND2_X1 U8023 ( .A1(n8194), .A2(n7242), .ZN(n8192) );
  INV_X1 U8024 ( .A(n8127), .ZN(n6323) );
  INV_X1 U8025 ( .A(n7456), .ZN(n9968) );
  NAND2_X1 U8026 ( .A1(n9968), .A2(n8329), .ZN(n8210) );
  AND2_X1 U8027 ( .A1(n8210), .A2(n8195), .ZN(n8206) );
  NAND2_X1 U8028 ( .A1(n7330), .A2(n8206), .ZN(n7473) );
  NAND2_X1 U8029 ( .A1(n9978), .A2(n8680), .ZN(n8212) );
  INV_X1 U8030 ( .A(n8329), .ZN(n7879) );
  NAND2_X1 U8031 ( .A1(n7456), .A2(n7879), .ZN(n8201) );
  AND2_X1 U8032 ( .A1(n8212), .A2(n8201), .ZN(n8209) );
  NAND2_X1 U8033 ( .A1(n7473), .A2(n8209), .ZN(n6324) );
  NAND2_X1 U8034 ( .A1(n6324), .A2(n8211), .ZN(n8692) );
  NAND2_X1 U8035 ( .A1(n8692), .A2(n8691), .ZN(n8694) );
  NAND2_X1 U8036 ( .A1(n9550), .A2(n7981), .ZN(n8224) );
  OR2_X1 U8037 ( .A1(n9550), .A2(n7981), .ZN(n8225) );
  INV_X1 U8038 ( .A(n8225), .ZN(n6325) );
  XNOR2_X1 U8039 ( .A(n8757), .B(n9559), .ZN(n8226) );
  NAND2_X1 U8040 ( .A1(n8677), .A2(n8676), .ZN(n8675) );
  NAND2_X1 U8041 ( .A1(n8757), .A2(n9559), .ZN(n6326) );
  NAND2_X1 U8042 ( .A1(n8675), .A2(n6326), .ZN(n8656) );
  INV_X1 U8043 ( .A(n8669), .ZN(n8649) );
  OR2_X1 U8044 ( .A1(n8837), .A2(n8649), .ZN(n8232) );
  NAND2_X1 U8045 ( .A1(n8656), .A2(n8232), .ZN(n6327) );
  NAND2_X1 U8046 ( .A1(n8837), .A2(n8649), .ZN(n8231) );
  INV_X1 U8047 ( .A(n8236), .ZN(n6328) );
  NAND2_X1 U8048 ( .A1(n8633), .A2(n8241), .ZN(n6329) );
  INV_X1 U8049 ( .A(n8820), .ZN(n6330) );
  AND2_X1 U8050 ( .A1(n6330), .A2(n8636), .ZN(n8242) );
  NAND2_X1 U8051 ( .A1(n8820), .A2(n7955), .ZN(n8247) );
  NAND2_X1 U8052 ( .A1(n6331), .A2(n8251), .ZN(n8596) );
  INV_X1 U8053 ( .A(n8253), .ZN(n8260) );
  NOR2_X1 U8054 ( .A1(n8795), .A2(n8571), .ZN(n8271) );
  INV_X1 U8055 ( .A(n8271), .ZN(n6332) );
  NAND2_X1 U8056 ( .A1(n6333), .A2(n7911), .ZN(n8140) );
  NAND2_X1 U8057 ( .A1(n8795), .A2(n8571), .ZN(n8552) );
  NAND2_X1 U8058 ( .A1(n6334), .A2(n8274), .ZN(n8542) );
  NAND2_X1 U8059 ( .A1(n8542), .A2(n8280), .ZN(n6335) );
  NAND2_X1 U8060 ( .A1(n6335), .A2(n8279), .ZN(n8523) );
  INV_X1 U8061 ( .A(n8538), .ZN(n7991) );
  NOR2_X1 U8062 ( .A1(n8712), .A2(n7991), .ZN(n8283) );
  NAND2_X1 U8063 ( .A1(n8712), .A2(n7991), .ZN(n8282) );
  NAND2_X1 U8064 ( .A1(n8774), .A2(n8504), .ZN(n8288) );
  NOR2_X1 U8065 ( .A1(n8512), .A2(n8153), .ZN(n6336) );
  INV_X1 U8066 ( .A(n6337), .ZN(n6338) );
  AOI21_X1 U8067 ( .B1(n8299), .B2(n7235), .A(n8472), .ZN(n6339) );
  AND2_X1 U8068 ( .A1(n6339), .A2(n9967), .ZN(n6341) );
  NAND2_X1 U8069 ( .A1(n8310), .A2(n8482), .ZN(n6384) );
  INV_X1 U8070 ( .A(n6384), .ZN(n6340) );
  NAND2_X1 U8071 ( .A1(n8290), .A2(n6340), .ZN(n6623) );
  NAND2_X1 U8072 ( .A1(n7875), .A2(n9919), .ZN(n6342) );
  NAND2_X1 U8073 ( .A1(n4481), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U8074 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6348), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6349) );
  NAND2_X1 U8075 ( .A1(n6376), .A2(n6377), .ZN(n6351) );
  XNOR2_X1 U8076 ( .A(n6362), .B(P2_B_REG_SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8077 ( .A1(n7806), .A2(n7455), .ZN(n6360) );
  NAND2_X1 U8078 ( .A1(n7455), .A2(n6362), .ZN(n6511) );
  NOR2_X1 U8079 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6366) );
  NOR4_X1 U8080 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6365) );
  NOR4_X1 U8081 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6364) );
  NOR4_X1 U8082 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6363) );
  NAND4_X1 U8083 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n6372)
         );
  NOR4_X1 U8084 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6370) );
  NOR4_X1 U8085 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6369) );
  NOR4_X1 U8086 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6368) );
  NOR4_X1 U8087 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6367) );
  NAND4_X1 U8088 ( .A1(n6370), .A2(n6369), .A3(n6368), .A4(n6367), .ZN(n6371)
         );
  NOR2_X1 U8089 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  NAND2_X1 U8090 ( .A1(n6772), .A2(n6614), .ZN(n6625) );
  INV_X1 U8091 ( .A(n7806), .ZN(n6375) );
  NOR2_X1 U8092 ( .A1(n6362), .A2(n7455), .ZN(n6374) );
  XNOR2_X1 U8093 ( .A(n6376), .B(n6377), .ZN(n6731) );
  INV_X1 U8094 ( .A(n6637), .ZN(n8843) );
  NOR2_X1 U8095 ( .A1(n9985), .A2(n8290), .ZN(n6378) );
  NOR2_X1 U8096 ( .A1(n6673), .A2(n8482), .ZN(n6676) );
  NOR2_X1 U8097 ( .A1(n8310), .A2(n7235), .ZN(n6385) );
  NAND2_X1 U8098 ( .A1(n6676), .A2(n6385), .ZN(n6613) );
  NAND2_X1 U8099 ( .A1(n6378), .A2(n6613), .ZN(n6632) );
  INV_X1 U8100 ( .A(n6844), .ZN(n9551) );
  NAND2_X1 U8101 ( .A1(n9985), .A2(n9551), .ZN(n9929) );
  NAND2_X1 U8102 ( .A1(n6632), .A2(n9929), .ZN(n6615) );
  NAND2_X1 U8103 ( .A1(n6631), .A2(n6615), .ZN(n6382) );
  NAND2_X1 U8104 ( .A1(n6614), .A2(n6637), .ZN(n6379) );
  NAND2_X1 U8105 ( .A1(n6613), .A2(n6623), .ZN(n6380) );
  NAND2_X1 U8106 ( .A1(n6636), .A2(n6380), .ZN(n6381) );
  NAND2_X1 U8107 ( .A1(n6383), .A2(n4910), .ZN(P2_U3456) );
  NAND2_X1 U8108 ( .A1(n8290), .A2(n6384), .ZN(n6618) );
  NAND3_X1 U8109 ( .A1(n6614), .A2(n6637), .A3(n6618), .ZN(n6773) );
  NOR2_X1 U8110 ( .A1(n6773), .A2(n6638), .ZN(n6391) );
  NAND2_X1 U8111 ( .A1(n6385), .A2(n8482), .ZN(n6386) );
  NAND2_X1 U8112 ( .A1(n6387), .A2(n6774), .ZN(n6389) );
  INV_X1 U8113 ( .A(n6774), .ZN(n6775) );
  NAND2_X1 U8114 ( .A1(n6672), .A2(n6775), .ZN(n6388) );
  OR2_X1 U8115 ( .A1(n10003), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8116 ( .A1(n4415), .A2(n6393), .ZN(n6394) );
  NAND2_X1 U8117 ( .A1(n6394), .A2(n4913), .ZN(P2_U3488) );
  NOR2_X1 U8118 ( .A1(n6395), .A2(P1_U3086), .ZN(n6396) );
  INV_X1 U8119 ( .A(n6513), .ZN(n6628) );
  INV_X1 U8120 ( .A(n6731), .ZN(n6397) );
  OR2_X1 U8121 ( .A1(n6619), .A2(n6397), .ZN(n6414) );
  NAND2_X1 U8122 ( .A1(n8290), .A2(n6731), .ZN(n6398) );
  NAND2_X1 U8123 ( .A1(n6414), .A2(n6398), .ZN(n6426) );
  OAI21_X1 U8124 ( .B1(n6426), .B2(n6399), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  MUX2_X1 U8125 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8473), .Z(n6918) );
  XNOR2_X1 U8126 ( .A(n6918), .B(n6929), .ZN(n6413) );
  MUX2_X1 U8127 ( .A(n6401), .B(n6400), .S(n8473), .Z(n6408) );
  INV_X1 U8128 ( .A(n6408), .ZN(n6409) );
  MUX2_X1 U8129 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8473), .Z(n6407) );
  MUX2_X1 U8130 ( .A(n6847), .B(n6402), .S(n8473), .Z(n6403) );
  XNOR2_X1 U8131 ( .A(n6403), .B(n6568), .ZN(n6574) );
  MUX2_X1 U8132 ( .A(n6791), .B(n5960), .S(n8473), .Z(n9828) );
  NAND2_X1 U8133 ( .A1(n9828), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6573) );
  INV_X1 U8134 ( .A(n6403), .ZN(n6404) );
  NAND2_X1 U8135 ( .A1(n6404), .A2(n6568), .ZN(n6405) );
  INV_X1 U8136 ( .A(n4350), .ZN(n6406) );
  XNOR2_X1 U8137 ( .A(n6407), .B(n6406), .ZN(n9844) );
  XNOR2_X1 U8138 ( .A(n6408), .B(n6536), .ZN(n6533) );
  NAND2_X1 U8139 ( .A1(n6534), .A2(n6533), .ZN(n6532) );
  OAI21_X1 U8140 ( .B1(n6409), .B2(n6536), .A(n6532), .ZN(n6412) );
  NOR2_X1 U8141 ( .A1(n6412), .A2(n6413), .ZN(n6917) );
  AOI211_X1 U8142 ( .C1(n6413), .C2(n6412), .A(n9857), .B(n6917), .ZN(n6452)
         );
  INV_X1 U8143 ( .A(n6414), .ZN(n6429) );
  INV_X1 U8144 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6415) );
  NOR2_X1 U8145 ( .A1(n9841), .A2(n6415), .ZN(n6451) );
  AND2_X1 U8146 ( .A1(n9833), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8147 ( .A1(n6420), .A2(n6419), .ZN(n6418) );
  OAI21_X1 U8148 ( .B1(n6420), .B2(n6419), .A(n6418), .ZN(n9852) );
  NAND2_X1 U8149 ( .A1(n9851), .A2(n9852), .ZN(n9850) );
  NAND2_X1 U8150 ( .A1(n4350), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6421) );
  INV_X1 U8151 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9991) );
  MUX2_X1 U8152 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9991), .S(n6929), .Z(n6422)
         );
  INV_X1 U8153 ( .A(n6422), .ZN(n6424) );
  NAND3_X1 U8154 ( .A1(n6544), .A2(n6424), .A3(n6423), .ZN(n6425) );
  OR2_X1 U8155 ( .A1(n6302), .A2(n9827), .ZN(n7496) );
  NOR2_X1 U8156 ( .A1(n6426), .A2(n7496), .ZN(n9830) );
  NAND2_X1 U8157 ( .A1(n9830), .A2(n8473), .ZN(n9909) );
  AOI21_X1 U8158 ( .B1(n6909), .B2(n6425), .A(n9909), .ZN(n6450) );
  INV_X1 U8159 ( .A(n6426), .ZN(n6433) );
  NOR2_X1 U8160 ( .A1(n8473), .A2(P2_U3151), .ZN(n7481) );
  AND2_X1 U8161 ( .A1(n7481), .A2(n6302), .ZN(n6427) );
  NAND2_X1 U8162 ( .A1(n6433), .A2(n6427), .ZN(n6431) );
  INV_X1 U8163 ( .A(n7496), .ZN(n6428) );
  NAND2_X1 U8164 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  INV_X1 U8165 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10185) );
  NOR2_X1 U8166 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10185), .ZN(n6835) );
  INV_X1 U8167 ( .A(n6835), .ZN(n6448) );
  NOR2_X1 U8168 ( .A1(n7496), .A2(n8473), .ZN(n6432) );
  INV_X1 U8169 ( .A(n9905), .ZN(n9838) );
  AND2_X1 U8170 ( .A1(n9833), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6436) );
  OAI21_X1 U8171 ( .B1(n6437), .B2(n6436), .A(n6438), .ZN(n6562) );
  INV_X1 U8172 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6847) );
  OR2_X1 U8173 ( .A1(n6562), .A2(n6847), .ZN(n6564) );
  NAND2_X1 U8174 ( .A1(n6564), .A2(n6438), .ZN(n9835) );
  NAND2_X1 U8175 ( .A1(n4350), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6439) );
  OAI21_X1 U8176 ( .B1(n6440), .B2(n6536), .A(n6443), .ZN(n6539) );
  NAND2_X1 U8177 ( .A1(n6537), .A2(n6443), .ZN(n6441) );
  INV_X1 U8178 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7019) );
  MUX2_X1 U8179 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7019), .S(n6929), .Z(n6442)
         );
  NAND2_X1 U8180 ( .A1(n6441), .A2(n6442), .ZN(n6928) );
  INV_X1 U8181 ( .A(n6442), .ZN(n6444) );
  NAND3_X1 U8182 ( .A1(n6537), .A2(n6444), .A3(n6443), .ZN(n6445) );
  NAND2_X1 U8183 ( .A1(n6928), .A2(n6445), .ZN(n6446) );
  NAND2_X1 U8184 ( .A1(n9838), .A2(n6446), .ZN(n6447) );
  OAI211_X1 U8185 ( .C1(n9871), .C2(n6929), .A(n6448), .B(n6447), .ZN(n6449)
         );
  OR4_X1 U8186 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(P2_U3186)
         );
  AOI22_X1 U8187 ( .A1(n9479), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9018), .ZN(n6453) );
  OAI21_X1 U8188 ( .B1(n6455), .B2(n6469), .A(n6453), .ZN(P1_U3354) );
  AND2_X1 U8189 ( .A1(n7525), .A2(P2_U3151), .ZN(n8850) );
  INV_X2 U8190 ( .A(n8850), .ZN(n8853) );
  INV_X2 U8191 ( .A(n7495), .ZN(n8855) );
  OAI222_X1 U8192 ( .A1(n8853), .A2(n6454), .B1(n8855), .B2(n6465), .C1(n6536), 
        .C2(n9827), .ZN(P2_U3292) );
  INV_X1 U8193 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6456) );
  OAI222_X1 U8194 ( .A1(n8853), .A2(n6456), .B1(n8855), .B2(n6455), .C1(n6568), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  OAI222_X1 U8195 ( .A1(n8853), .A2(n5036), .B1(n8855), .B2(n6459), .C1(n4350), 
        .C2(n9827), .ZN(P2_U3293) );
  OAI222_X1 U8196 ( .A1(n6929), .A2(P2_U3151), .B1(n8855), .B2(n6461), .C1(
        n5107), .C2(n8853), .ZN(P2_U3291) );
  OAI222_X1 U8197 ( .A1(n9870), .A2(n9827), .B1(n8855), .B2(n6463), .C1(n6457), 
        .C2(n8853), .ZN(P2_U3290) );
  OAI222_X1 U8198 ( .A1(n6933), .A2(P2_U3151), .B1(n8855), .B2(n6467), .C1(
        n6501), .C2(n8853), .ZN(P2_U3289) );
  CLKBUF_X1 U8199 ( .A(n9479), .Z(n9475) );
  AOI22_X1 U8200 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n9475), .B1(n9037), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6458) );
  OAI21_X1 U8201 ( .B1(n6459), .B2(n6469), .A(n6458), .ZN(P1_U3353) );
  AOI22_X1 U8202 ( .A1(n9587), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9475), .ZN(n6460) );
  OAI21_X1 U8203 ( .B1(n6461), .B2(n6469), .A(n6460), .ZN(P1_U3351) );
  AOI22_X1 U8204 ( .A1(n9602), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9475), .ZN(n6462) );
  OAI21_X1 U8205 ( .B1(n6463), .B2(n6469), .A(n6462), .ZN(P1_U3350) );
  AOI22_X1 U8206 ( .A1(n9050), .A2(P1_STATE_REG_SCAN_IN), .B1(n9475), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6464) );
  OAI21_X1 U8207 ( .B1(n6465), .B2(n6469), .A(n6464), .ZN(P1_U3352) );
  AOI22_X1 U8208 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9063), .B1(n9475), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6466) );
  OAI21_X1 U8209 ( .B1(n6467), .B2(n6469), .A(n6466), .ZN(P1_U3349) );
  AOI22_X1 U8210 ( .A1(n9508), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9475), .ZN(n6468) );
  OAI21_X1 U8211 ( .B1(n6471), .B2(n6469), .A(n6468), .ZN(P1_U3348) );
  OAI222_X1 U8212 ( .A1(n7060), .A2(n9827), .B1(n8855), .B2(n6471), .C1(n6470), 
        .C2(n8853), .ZN(P2_U3288) );
  AOI22_X1 U8213 ( .A1(n9521), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9475), .ZN(n6472) );
  OAI21_X1 U8214 ( .B1(n6474), .B2(n6469), .A(n6472), .ZN(P1_U3347) );
  OAI222_X1 U8215 ( .A1(n9893), .A2(P2_U3151), .B1(n8855), .B2(n6474), .C1(
        n6473), .C2(n8853), .ZN(P2_U3287) );
  INV_X1 U8216 ( .A(n6475), .ZN(n6491) );
  AOI22_X1 U8217 ( .A1(n9537), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9475), .ZN(n6476) );
  OAI21_X1 U8218 ( .B1(n6491), .B2(n6469), .A(n6476), .ZN(P1_U3346) );
  AND2_X1 U8219 ( .A1(n6510), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8220 ( .A1(n6510), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8221 ( .A1(n6510), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8222 ( .A1(n6510), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8223 ( .A1(n6510), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8224 ( .A1(n6510), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8225 ( .A1(n6510), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8226 ( .A1(n6510), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8227 ( .A1(n6510), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8228 ( .A1(n6510), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8229 ( .A1(n6510), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AOI21_X1 U8230 ( .B1(n6479), .B2(n7735), .A(n6478), .ZN(n7833) );
  INV_X1 U8231 ( .A(n7833), .ZN(n6480) );
  INV_X1 U8232 ( .A(n7802), .ZN(n7798) );
  OR2_X1 U8233 ( .A1(n6554), .A2(n7798), .ZN(n7834) );
  AND2_X1 U8234 ( .A1(n6480), .A2(n7834), .ZN(n9593) );
  NOR2_X1 U8235 ( .A1(n9593), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8236 ( .A(n6481), .ZN(n6484) );
  AOI22_X1 U8237 ( .A1(n9489), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9479), .ZN(n6482) );
  OAI21_X1 U8238 ( .B1(n6484), .B2(n6469), .A(n6482), .ZN(P1_U3345) );
  AOI22_X1 U8239 ( .A1(n7382), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8850), .ZN(n6483) );
  OAI21_X1 U8240 ( .B1(n6484), .B2(n8855), .A(n6483), .ZN(P2_U3285) );
  INV_X1 U8241 ( .A(n6485), .ZN(n6486) );
  INV_X1 U8242 ( .A(n9768), .ZN(n6490) );
  NAND2_X1 U8243 ( .A1(n6490), .A2(n6487), .ZN(n6488) );
  OAI21_X1 U8244 ( .B1(n6490), .B2(n6489), .A(n6488), .ZN(P1_U3440) );
  OAI222_X1 U8245 ( .A1(n9827), .A2(n7078), .B1(n8855), .B2(n6491), .C1(n6504), 
        .C2(n8853), .ZN(P2_U3286) );
  INV_X1 U8246 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8247 ( .A1(n6608), .A2(P2_U3893), .ZN(n6492) );
  OAI21_X1 U8248 ( .B1(P2_U3893), .B2(n6493), .A(n6492), .ZN(P2_U3491) );
  INV_X1 U8249 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6500) );
  INV_X1 U8250 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9309) );
  INV_X1 U8251 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6494) );
  OR2_X1 U8252 ( .A1(n5089), .A2(n6494), .ZN(n6497) );
  NAND2_X1 U8253 ( .A1(n6495), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6496) );
  OAI211_X1 U8254 ( .C1(n6498), .C2(n9309), .A(n6497), .B(n6496), .ZN(n9076)
         );
  NAND2_X1 U8255 ( .A1(n9076), .A2(P1_U3973), .ZN(n6499) );
  OAI21_X1 U8256 ( .B1(P1_U3973), .B2(n6500), .A(n6499), .ZN(P1_U3585) );
  MUX2_X1 U8257 ( .A(n6501), .B(n7536), .S(P1_U3973), .Z(n6502) );
  INV_X1 U8258 ( .A(n6502), .ZN(P1_U3560) );
  MUX2_X1 U8259 ( .A(n6508), .B(n7317), .S(P1_U3973), .Z(n6503) );
  INV_X1 U8260 ( .A(n6503), .ZN(P1_U3565) );
  MUX2_X1 U8261 ( .A(n6504), .B(n9741), .S(P1_U3973), .Z(n6505) );
  INV_X1 U8262 ( .A(n6505), .ZN(P1_U3563) );
  INV_X1 U8263 ( .A(n6506), .ZN(n6509) );
  AOI22_X1 U8264 ( .A1(n9619), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9479), .ZN(n6507) );
  OAI21_X1 U8265 ( .B1(n6509), .B2(n6469), .A(n6507), .ZN(P1_U3344) );
  INV_X1 U8266 ( .A(n7386), .ZN(n7417) );
  OAI222_X1 U8267 ( .A1(n7417), .A2(n9827), .B1(n8855), .B2(n6509), .C1(n6508), 
        .C2(n8853), .ZN(P2_U3284) );
  INV_X1 U8268 ( .A(n6511), .ZN(n6512) );
  AOI22_X1 U8269 ( .A1(n6510), .A2(n4728), .B1(n6513), .B2(n6512), .ZN(
        P2_U3376) );
  INV_X1 U8270 ( .A(n6514), .ZN(n6517) );
  AOI22_X1 U8271 ( .A1(n7390), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8850), .ZN(n6515) );
  OAI21_X1 U8272 ( .B1(n6517), .B2(n8855), .A(n6515), .ZN(P2_U3283) );
  AOI22_X1 U8273 ( .A1(n9635), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9479), .ZN(n6516) );
  OAI21_X1 U8274 ( .B1(n6517), .B2(n6469), .A(n6516), .ZN(P1_U3343) );
  INV_X1 U8275 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6521) );
  AND2_X1 U8276 ( .A1(n9014), .A2(n6755), .ZN(n7744) );
  NOR2_X1 U8277 ( .A1(n6524), .A2(n7744), .ZN(n7668) );
  NOR2_X1 U8278 ( .A1(n9812), .A2(n9331), .ZN(n6518) );
  INV_X1 U8279 ( .A(n9013), .ZN(n6591) );
  OAI222_X1 U8280 ( .A1(n6755), .A2(n6519), .B1(n7668), .B2(n6518), .C1(n9740), 
        .C2(n6591), .ZN(n9413) );
  NAND2_X1 U8281 ( .A1(n9413), .A2(n9816), .ZN(n6520) );
  OAI21_X1 U8282 ( .B1(n9816), .B2(n6521), .A(n6520), .ZN(P1_U3453) );
  AND2_X1 U8283 ( .A1(n6510), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8284 ( .A1(n6510), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8285 ( .A1(n6510), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8286 ( .A1(n6510), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8287 ( .A1(n6510), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8288 ( .A1(n6510), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8289 ( .A1(n6510), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8290 ( .A1(n6510), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8291 ( .A1(n6510), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8292 ( .A1(n6510), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8293 ( .A1(n6510), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8294 ( .A1(n6510), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8295 ( .A1(n6510), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8296 ( .A1(n6510), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8297 ( .A1(n6510), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8298 ( .A1(n6510), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8299 ( .A1(n6510), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8300 ( .A1(n6510), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8301 ( .A1(n6510), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  INV_X1 U8302 ( .A(n6522), .ZN(n6560) );
  AOI22_X1 U8303 ( .A1(n9652), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9479), .ZN(n6523) );
  OAI21_X1 U8304 ( .B1(n6560), .B2(n6469), .A(n6523), .ZN(P1_U3342) );
  XNOR2_X1 U8305 ( .A(n7666), .B(n6524), .ZN(n6525) );
  NAND2_X1 U8306 ( .A1(n6525), .A2(n9331), .ZN(n6878) );
  AOI22_X1 U8307 ( .A1(n9796), .A2(n9014), .B1(n5814), .B2(n9805), .ZN(n6530)
         );
  OAI21_X1 U8308 ( .B1(n5862), .B2(n6527), .A(n6526), .ZN(n6873) );
  NAND2_X1 U8309 ( .A1(n6873), .A2(n9812), .ZN(n6529) );
  OAI21_X1 U8310 ( .B1(n7745), .B2(n6755), .A(n9761), .ZN(n6528) );
  OR2_X1 U8311 ( .A1(n6528), .A2(n6589), .ZN(n6870) );
  AND4_X1 U8312 ( .A1(n6878), .A2(n6530), .A3(n6529), .A4(n6870), .ZN(n6671)
         );
  INV_X1 U8313 ( .A(n9406), .ZN(n7430) );
  AOI22_X1 U8314 ( .A1(n7430), .A2(n6579), .B1(P1_REG1_REG_1__SCAN_IN), .B2(
        n9824), .ZN(n6531) );
  OAI21_X1 U8315 ( .B1(n6671), .B2(n9824), .A(n6531), .ZN(P1_U3523) );
  INV_X1 U8316 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6549) );
  OAI21_X1 U8317 ( .B1(n6534), .B2(n6533), .A(n6532), .ZN(n6535) );
  NAND2_X1 U8318 ( .A1(n6535), .A2(n6411), .ZN(n6548) );
  INV_X1 U8319 ( .A(n6537), .ZN(n6538) );
  AOI21_X1 U8320 ( .B1(n6401), .B2(n6539), .A(n6538), .ZN(n6541) );
  INV_X1 U8321 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U8322 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10211), .ZN(n6739) );
  INV_X1 U8323 ( .A(n6739), .ZN(n6540) );
  OAI21_X1 U8324 ( .B1(n9905), .B2(n6541), .A(n6540), .ZN(n6546) );
  NAND2_X1 U8325 ( .A1(n6542), .A2(n6400), .ZN(n6543) );
  AOI21_X1 U8326 ( .B1(n6544), .B2(n6543), .A(n9909), .ZN(n6545) );
  AOI211_X1 U8327 ( .C1(n4783), .C2(n9896), .A(n6546), .B(n6545), .ZN(n6547)
         );
  OAI211_X1 U8328 ( .C1(n9841), .C2(n6549), .A(n6548), .B(n6547), .ZN(P2_U3185) );
  OAI21_X1 U8329 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(n9026) );
  INV_X1 U8330 ( .A(n6553), .ZN(n6555) );
  NAND2_X1 U8331 ( .A1(n6555), .A2(n6554), .ZN(n6599) );
  AOI22_X1 U8332 ( .A1(n8971), .A2(n6556), .B1(n6599), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U8333 ( .A1(n8985), .A2(n9013), .ZN(n6557) );
  OAI211_X1 U8334 ( .C1(n9026), .C2(n8973), .A(n6558), .B(n6557), .ZN(P1_U3232) );
  INV_X1 U8335 ( .A(n8376), .ZN(n8364) );
  INV_X1 U8336 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6559) );
  OAI222_X1 U8337 ( .A1(n8364), .A2(P2_U3151), .B1(n8855), .B2(n6560), .C1(
        n6559), .C2(n8853), .ZN(P2_U3282) );
  XNOR2_X1 U8338 ( .A(n6561), .B(n6402), .ZN(n6571) );
  INV_X1 U8339 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U8340 ( .A1(n9841), .A2(n10009), .ZN(n6570) );
  NAND2_X1 U8341 ( .A1(P2_U3151), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8342 ( .A1(n6562), .A2(n6847), .ZN(n6563) );
  NAND2_X1 U8343 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  NAND2_X1 U8344 ( .A1(n9838), .A2(n6565), .ZN(n6566) );
  OAI211_X1 U8345 ( .C1(n9871), .C2(n6568), .A(n6567), .B(n6566), .ZN(n6569)
         );
  AOI211_X1 U8346 ( .C1(n8489), .C2(n6571), .A(n6570), .B(n6569), .ZN(n6576)
         );
  OAI211_X1 U8347 ( .C1(n6574), .C2(n6573), .A(n6572), .B(n6411), .ZN(n6575)
         );
  NAND2_X1 U8348 ( .A1(n6576), .A2(n6575), .ZN(P2_U3183) );
  XOR2_X1 U8349 ( .A(n6577), .B(n6578), .Z(n6582) );
  INV_X1 U8350 ( .A(n8983), .ZN(n8999) );
  AOI22_X1 U8351 ( .A1(n8999), .A2(n9014), .B1(n8985), .B2(n5814), .ZN(n6581)
         );
  AOI22_X1 U8352 ( .A1(n8971), .A2(n6579), .B1(n6599), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U8353 ( .C1(n6582), .C2(n8973), .A(n6581), .B(n6580), .ZN(P1_U3222) );
  INV_X1 U8354 ( .A(n6583), .ZN(n6605) );
  AOI22_X1 U8355 ( .A1(n9669), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9479), .ZN(n6584) );
  OAI21_X1 U8356 ( .B1(n6605), .B2(n6469), .A(n6584), .ZN(P1_U3341) );
  XNOR2_X1 U8357 ( .A(n6587), .B(n6585), .ZN(n6869) );
  OAI21_X1 U8358 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(n6867) );
  OAI21_X1 U8359 ( .B1(n6589), .B2(n5813), .A(n9761), .ZN(n6590) );
  OR2_X1 U8360 ( .A1(n6590), .A2(n6648), .ZN(n6860) );
  INV_X1 U8361 ( .A(n6860), .ZN(n6593) );
  INV_X1 U8362 ( .A(n9012), .ZN(n6861) );
  OAI22_X1 U8363 ( .A1(n6861), .A2(n9740), .B1(n6591), .B2(n9738), .ZN(n6592)
         );
  AOI211_X1 U8364 ( .C1(n6867), .C2(n9812), .A(n6593), .B(n6592), .ZN(n6594)
         );
  OAI21_X1 U8365 ( .B1(n9746), .B2(n6869), .A(n6594), .ZN(n6701) );
  OAI22_X1 U8366 ( .A1(n9406), .A2(n5813), .B1(n9826), .B2(n7840), .ZN(n6595)
         );
  AOI21_X1 U8367 ( .B1(n6701), .B2(n9826), .A(n6595), .ZN(n6596) );
  INV_X1 U8368 ( .A(n6596), .ZN(P1_U3524) );
  XOR2_X1 U8369 ( .A(n6598), .B(n6597), .Z(n6603) );
  AOI22_X1 U8370 ( .A1(n8985), .A2(n9012), .B1(n8999), .B2(n9013), .ZN(n6602)
         );
  AOI22_X1 U8371 ( .A1(n8971), .A2(n6600), .B1(n6599), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6601) );
  OAI211_X1 U8372 ( .C1(n6603), .C2(n8973), .A(n6602), .B(n6601), .ZN(P1_U3237) );
  INV_X1 U8373 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6604) );
  OAI222_X1 U8374 ( .A1(P2_U3151), .A2(n8397), .B1(n8855), .B2(n6605), .C1(
        n6604), .C2(n8853), .ZN(P2_U3281) );
  INV_X1 U8375 ( .A(n6606), .ZN(n6654) );
  AOI22_X1 U8376 ( .A1(n9688), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9479), .ZN(n6607) );
  OAI21_X1 U8377 ( .B1(n6654), .B2(n6469), .A(n6607), .ZN(P1_U3340) );
  INV_X1 U8378 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6612) );
  INV_X1 U8379 ( .A(n6788), .ZN(n6640) );
  AND2_X1 U8380 ( .A1(n6608), .A2(n6640), .ZN(n8160) );
  INV_X1 U8381 ( .A(n8160), .ZN(n8164) );
  NAND2_X1 U8382 ( .A1(n8159), .A2(n8164), .ZN(n8121) );
  OAI21_X1 U8383 ( .B1(n8671), .B2(n9980), .A(n8121), .ZN(n6610) );
  NAND2_X1 U8384 ( .A1(n6609), .A2(n8684), .ZN(n6783) );
  OAI211_X1 U8385 ( .C1(n6640), .C2(n9967), .A(n6610), .B(n6783), .ZN(n6842)
         );
  NAND2_X1 U8386 ( .A1(n6842), .A2(n9986), .ZN(n6611) );
  OAI21_X1 U8387 ( .B1(n6612), .B2(n9986), .A(n6611), .ZN(P2_U3390) );
  INV_X1 U8388 ( .A(n6613), .ZN(n6630) );
  NAND2_X1 U8389 ( .A1(n6625), .A2(n6630), .ZN(n6621) );
  INV_X1 U8390 ( .A(n6614), .ZN(n6616) );
  OAI21_X1 U8391 ( .B1(n6617), .B2(n6616), .A(n6615), .ZN(n6620) );
  NAND4_X1 U8392 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6622)
         );
  NAND2_X1 U8393 ( .A1(n6622), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6627) );
  INV_X1 U8394 ( .A(n6623), .ZN(n6781) );
  NAND2_X1 U8395 ( .A1(n6637), .A2(n6781), .ZN(n8318) );
  INV_X1 U8396 ( .A(n8318), .ZN(n6624) );
  NAND2_X1 U8397 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  NAND2_X1 U8398 ( .A1(n6627), .A2(n6626), .ZN(n6733) );
  NOR2_X1 U8399 ( .A1(n6733), .A2(n6628), .ZN(n6720) );
  AND2_X1 U8400 ( .A1(n6631), .A2(n6781), .ZN(n6686) );
  INV_X1 U8401 ( .A(n6686), .ZN(n6629) );
  INV_X1 U8402 ( .A(n8121), .ZN(n6782) );
  NAND2_X1 U8403 ( .A1(n6631), .A2(n6630), .ZN(n6635) );
  INV_X1 U8404 ( .A(n6632), .ZN(n6633) );
  NAND2_X1 U8405 ( .A1(n6636), .A2(n6633), .ZN(n6634) );
  NAND2_X1 U8406 ( .A1(n6636), .A2(n9985), .ZN(n6639) );
  OAI22_X1 U8407 ( .A1(n6782), .A2(n8082), .B1(n8099), .B2(n6640), .ZN(n6641)
         );
  AOI21_X1 U8408 ( .B1(n8066), .B2(n6609), .A(n6641), .ZN(n6642) );
  OAI21_X1 U8409 ( .B1(n6720), .B2(n10098), .A(n6642), .ZN(P2_U3172) );
  INV_X1 U8410 ( .A(n7671), .ZN(n6643) );
  XNOR2_X1 U8411 ( .A(n6644), .B(n6643), .ZN(n6816) );
  OAI21_X1 U8412 ( .B1(n6646), .B2(n7671), .A(n6645), .ZN(n6647) );
  INV_X1 U8413 ( .A(n6647), .ZN(n6819) );
  INV_X1 U8414 ( .A(n9812), .ZN(n9773) );
  AOI22_X1 U8415 ( .A1(n9805), .A2(n4349), .B1(n5814), .B2(n9796), .ZN(n6649)
         );
  OAI211_X1 U8416 ( .C1(n6648), .C2(n6813), .A(n9761), .B(n6804), .ZN(n6812)
         );
  OAI211_X1 U8417 ( .C1(n6819), .C2(n9773), .A(n6649), .B(n6812), .ZN(n6650)
         );
  AOI21_X1 U8418 ( .B1(n9331), .B2(n6816), .A(n6650), .ZN(n6667) );
  OAI22_X1 U8419 ( .A1(n9406), .A2(n6813), .B1(n9826), .B2(n7844), .ZN(n6651)
         );
  INV_X1 U8420 ( .A(n6651), .ZN(n6652) );
  OAI21_X1 U8421 ( .B1(n6667), .B2(n9824), .A(n6652), .ZN(P1_U3525) );
  INV_X1 U8422 ( .A(n8421), .ZN(n8412) );
  INV_X1 U8423 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6653) );
  OAI222_X1 U8424 ( .A1(n9827), .A2(n8412), .B1(n8855), .B2(n6654), .C1(n6653), 
        .C2(n8853), .ZN(P2_U3280) );
  NAND2_X1 U8425 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9047) );
  INV_X1 U8426 ( .A(n9047), .ZN(n6656) );
  INV_X1 U8427 ( .A(n5814), .ZN(n6871) );
  OAI22_X1 U8428 ( .A1(n6813), .A2(n9002), .B1(n8983), .B2(n6871), .ZN(n6655)
         );
  AOI211_X1 U8429 ( .C1(n8985), .C2(n4349), .A(n6656), .B(n6655), .ZN(n6661)
         );
  XNOR2_X1 U8430 ( .A(n6658), .B(n6657), .ZN(n6659) );
  NAND2_X1 U8431 ( .A1(n6659), .A2(n8991), .ZN(n6660) );
  OAI211_X1 U8432 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8996), .A(n6661), .B(
        n6660), .ZN(P1_U3218) );
  INV_X1 U8433 ( .A(n6662), .ZN(n6704) );
  AOI22_X1 U8434 ( .A1(n7860), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9479), .ZN(n6663) );
  OAI21_X1 U8435 ( .B1(n6704), .B2(n6469), .A(n6663), .ZN(P1_U3339) );
  INV_X1 U8436 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6664) );
  OAI22_X1 U8437 ( .A1(n9466), .A2(n6813), .B1(n9816), .B2(n6664), .ZN(n6665)
         );
  INV_X1 U8438 ( .A(n6665), .ZN(n6666) );
  OAI21_X1 U8439 ( .B1(n6667), .B2(n9814), .A(n6666), .ZN(P1_U3462) );
  INV_X1 U8440 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6668) );
  OAI22_X1 U8441 ( .A1(n9466), .A2(n7745), .B1(n9816), .B2(n6668), .ZN(n6669)
         );
  INV_X1 U8442 ( .A(n6669), .ZN(n6670) );
  OAI21_X1 U8443 ( .B1(n6671), .B2(n9814), .A(n6670), .ZN(P1_U3456) );
  INV_X1 U8444 ( .A(n6676), .ZN(n6677) );
  XNOR2_X1 U8445 ( .A(n6712), .B(n6687), .ZN(n6680) );
  NOR2_X1 U8446 ( .A1(n6680), .A2(n6609), .ZN(n6709) );
  AND2_X1 U8447 ( .A1(n6680), .A2(n6609), .ZN(n6681) );
  NOR2_X1 U8448 ( .A1(n6709), .A2(n6681), .ZN(n6683) );
  OAI21_X1 U8449 ( .B1(n6788), .B2(n7922), .A(n8159), .ZN(n6682) );
  NAND2_X1 U8450 ( .A1(n6683), .A2(n6682), .ZN(n6711) );
  OAI21_X1 U8451 ( .B1(n6683), .B2(n6682), .A(n6711), .ZN(n6684) );
  NAND2_X1 U8452 ( .A1(n6684), .A2(n8088), .ZN(n6690) );
  OAI22_X1 U8453 ( .A1(n8070), .A2(n6317), .B1(n6687), .B2(n8099), .ZN(n6688)
         );
  AOI21_X1 U8454 ( .B1(n8066), .B2(n4354), .A(n6688), .ZN(n6689) );
  OAI211_X1 U8455 ( .C1(n6720), .C2(n6691), .A(n6690), .B(n6689), .ZN(P2_U3162) );
  AOI21_X1 U8456 ( .B1(n6692), .B2(n6693), .A(n8973), .ZN(n6695) );
  NAND2_X1 U8457 ( .A1(n6695), .A2(n6694), .ZN(n6698) );
  AND2_X1 U8458 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9592) );
  OAI22_X1 U8459 ( .A1(n6806), .A2(n9002), .B1(n8983), .B2(n6861), .ZN(n6696)
         );
  AOI211_X1 U8460 ( .C1(n8985), .C2(n9010), .A(n9592), .B(n6696), .ZN(n6697)
         );
  OAI211_X1 U8461 ( .C1(n8996), .C2(n6805), .A(n6698), .B(n6697), .ZN(P1_U3230) );
  INV_X1 U8462 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6699) );
  OAI22_X1 U8463 ( .A1(n9466), .A2(n5813), .B1(n9816), .B2(n6699), .ZN(n6700)
         );
  AOI21_X1 U8464 ( .B1(n6701), .B2(n9816), .A(n6700), .ZN(n6702) );
  INV_X1 U8465 ( .A(n6702), .ZN(P1_U3459) );
  INV_X1 U8466 ( .A(n8424), .ZN(n8437) );
  INV_X1 U8467 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6703) );
  OAI222_X1 U8468 ( .A1(n8437), .A2(n9827), .B1(n8855), .B2(n6704), .C1(n6703), 
        .C2(n8853), .ZN(P2_U3279) );
  INV_X1 U8469 ( .A(n6705), .ZN(n6708) );
  AOI22_X1 U8470 ( .A1(n9710), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9475), .ZN(n6706) );
  OAI21_X1 U8471 ( .B1(n6708), .B2(n6469), .A(n6706), .ZN(P1_U3338) );
  INV_X1 U8472 ( .A(n8460), .ZN(n8440) );
  INV_X1 U8473 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6707) );
  OAI222_X1 U8474 ( .A1(P2_U3151), .A2(n8440), .B1(n8855), .B2(n6708), .C1(
        n6707), .C2(n8853), .ZN(P2_U3278) );
  INV_X1 U8475 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6719) );
  INV_X1 U8476 ( .A(n6709), .ZN(n6710) );
  NAND2_X1 U8477 ( .A1(n6711), .A2(n6710), .ZN(n6714) );
  XNOR2_X1 U8478 ( .A(n6734), .B(n4354), .ZN(n6713) );
  NAND2_X1 U8479 ( .A1(n6714), .A2(n6713), .ZN(n6736) );
  OAI21_X1 U8480 ( .B1(n6714), .B2(n6713), .A(n6736), .ZN(n6715) );
  NAND2_X1 U8481 ( .A1(n6715), .A2(n8088), .ZN(n6718) );
  OAI22_X1 U8482 ( .A1(n8070), .A2(n9923), .B1(n9930), .B2(n8099), .ZN(n6716)
         );
  AOI21_X1 U8483 ( .B1(n8066), .B2(n8336), .A(n6716), .ZN(n6717) );
  OAI211_X1 U8484 ( .C1(n6720), .C2(n6719), .A(n6718), .B(n6717), .ZN(P2_U3177) );
  OAI21_X1 U8485 ( .B1(n6722), .B2(n6724), .A(n6721), .ZN(n6998) );
  INV_X1 U8486 ( .A(n4354), .ZN(n6760) );
  XNOR2_X1 U8487 ( .A(n6724), .B(n6723), .ZN(n6725) );
  OAI222_X1 U8488 ( .A1(n9920), .A2(n6831), .B1(n9922), .B2(n6760), .C1(n9928), 
        .C2(n6725), .ZN(n6995) );
  AOI21_X1 U8489 ( .B1(n9980), .B2(n6998), .A(n6995), .ZN(n7107) );
  INV_X1 U8490 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6726) );
  OAI22_X1 U8491 ( .A1(n6994), .A2(n8807), .B1(n9986), .B2(n6726), .ZN(n6727)
         );
  INV_X1 U8492 ( .A(n6727), .ZN(n6728) );
  OAI21_X1 U8493 ( .B1(n7107), .B2(n9988), .A(n6728), .ZN(P2_U3399) );
  INV_X1 U8494 ( .A(n6729), .ZN(n6770) );
  AOI22_X1 U8495 ( .A1(n9725), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9475), .ZN(n6730) );
  OAI21_X1 U8496 ( .B1(n6770), .B2(n6469), .A(n6730), .ZN(P1_U3337) );
  OR2_X1 U8497 ( .A1(n6731), .A2(n9827), .ZN(n8322) );
  INV_X1 U8498 ( .A(n8322), .ZN(n6732) );
  NAND2_X1 U8499 ( .A1(n6734), .A2(n6760), .ZN(n6735) );
  AND2_X1 U8500 ( .A1(n6736), .A2(n6735), .ZN(n6738) );
  XNOR2_X1 U8501 ( .A(n7922), .B(n6994), .ZN(n6828) );
  XNOR2_X1 U8502 ( .A(n6828), .B(n9921), .ZN(n6737) );
  NAND3_X1 U8503 ( .A1(n6736), .A2(n6735), .A3(n6737), .ZN(n6829) );
  OAI211_X1 U8504 ( .C1(n6738), .C2(n6737), .A(n8088), .B(n6829), .ZN(n6743)
         );
  AOI21_X1 U8505 ( .B1(n8080), .B2(n7105), .A(n6739), .ZN(n6740) );
  OAI21_X1 U8506 ( .B1(n8070), .B2(n6760), .A(n6740), .ZN(n6741) );
  AOI21_X1 U8507 ( .B1(n8066), .B2(n8335), .A(n6741), .ZN(n6742) );
  OAI211_X1 U8508 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8040), .A(n6743), .B(
        n6742), .ZN(P2_U3158) );
  NAND3_X1 U8509 ( .A1(n6746), .A2(n6745), .A3(n6744), .ZN(n6747) );
  AOI21_X1 U8510 ( .B1(n9764), .B2(n9761), .A(n9286), .ZN(n6756) );
  OR2_X1 U8511 ( .A1(n9295), .A2(n9740), .ZN(n9279) );
  INV_X1 U8512 ( .A(n9279), .ZN(n9211) );
  NOR4_X1 U8513 ( .A1(n9295), .A2(n7668), .A3(n6750), .A4(n6749), .ZN(n6753)
         );
  OAI22_X1 U8514 ( .A1(n9251), .A2(n9029), .B1(n6751), .B2(n9753), .ZN(n6752)
         );
  AOI211_X1 U8515 ( .C1(n9211), .C2(n9013), .A(n6753), .B(n6752), .ZN(n6754)
         );
  OAI21_X1 U8516 ( .B1(n6756), .B2(n6755), .A(n6754), .ZN(P1_U3293) );
  INV_X1 U8517 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6767) );
  INV_X1 U8518 ( .A(n8159), .ZN(n6759) );
  OAI21_X1 U8519 ( .B1(n6318), .B2(n6759), .A(n6758), .ZN(n6849) );
  OAI22_X1 U8520 ( .A1(n6317), .A2(n9922), .B1(n6760), .B2(n9920), .ZN(n6764)
         );
  XNOR2_X1 U8521 ( .A(n6318), .B(n6761), .ZN(n6762) );
  NOR2_X1 U8522 ( .A1(n6762), .A2(n9928), .ZN(n6763) );
  AOI211_X1 U8523 ( .C1(n9919), .C2(n6849), .A(n6764), .B(n6763), .ZN(n6851)
         );
  AOI22_X1 U8524 ( .A1(n6849), .A2(n6344), .B1(n9985), .B2(n6845), .ZN(n6765)
         );
  NAND2_X1 U8525 ( .A1(n6851), .A2(n6765), .ZN(n6768) );
  NAND2_X1 U8526 ( .A1(n6768), .A2(n9986), .ZN(n6766) );
  OAI21_X1 U8527 ( .B1(n6767), .B2(n9986), .A(n6766), .ZN(P2_U3393) );
  NAND2_X1 U8528 ( .A1(n6768), .A2(n10003), .ZN(n6769) );
  OAI21_X1 U8529 ( .B1(n10003), .B2(n6402), .A(n6769), .ZN(P2_U3460) );
  INV_X1 U8530 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6771) );
  INV_X1 U8531 ( .A(n8476), .ZN(n8462) );
  OAI222_X1 U8532 ( .A1(n8853), .A2(n6771), .B1(n8855), .B2(n6770), .C1(
        P2_U3151), .C2(n8462), .ZN(P2_U3277) );
  INV_X1 U8533 ( .A(n6772), .ZN(n6780) );
  INV_X1 U8534 ( .A(n6773), .ZN(n6779) );
  NAND2_X1 U8535 ( .A1(n8844), .A2(n6774), .ZN(n6778) );
  NAND2_X1 U8536 ( .A1(n6776), .A2(n6775), .ZN(n6777) );
  NAND4_X1 U8537 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6786)
         );
  NOR3_X1 U8538 ( .A1(n6782), .A2(n9985), .A3(n6781), .ZN(n6785) );
  INV_X1 U8539 ( .A(n6783), .ZN(n6784) );
  OAI21_X1 U8540 ( .B1(n6785), .B2(n6784), .A(n9562), .ZN(n6790) );
  INV_X1 U8541 ( .A(n6786), .ZN(n6787) );
  INV_X1 U8542 ( .A(n9929), .ZN(n8673) );
  AOI22_X1 U8543 ( .A1(n8664), .A2(n6788), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9934), .ZN(n6789) );
  OAI211_X1 U8544 ( .C1(n6791), .C2(n9562), .A(n6790), .B(n6789), .ZN(P2_U3233) );
  OAI21_X1 U8545 ( .B1(n6793), .B2(n6797), .A(n6792), .ZN(n6794) );
  INV_X1 U8546 ( .A(n6794), .ZN(n9774) );
  NAND2_X1 U8547 ( .A1(n6795), .A2(n7662), .ZN(n7202) );
  AND2_X1 U8548 ( .A1(n9737), .A2(n7202), .ZN(n6796) );
  INV_X1 U8549 ( .A(n6797), .ZN(n7673) );
  XNOR2_X1 U8550 ( .A(n6798), .B(n7673), .ZN(n6799) );
  NAND2_X1 U8551 ( .A1(n6799), .A2(n9331), .ZN(n6801) );
  AOI22_X1 U8552 ( .A1(n9796), .A2(n9012), .B1(n9010), .B2(n9805), .ZN(n6800)
         );
  AND2_X1 U8553 ( .A1(n6801), .A2(n6800), .ZN(n9772) );
  MUX2_X1 U8554 ( .A(n9772), .B(n6802), .S(n9295), .Z(n6809) );
  INV_X1 U8555 ( .A(n6822), .ZN(n6803) );
  AOI211_X1 U8556 ( .C1(n9770), .C2(n6804), .A(n9291), .B(n6803), .ZN(n9769)
         );
  OAI22_X1 U8557 ( .A1(n9756), .A2(n6806), .B1(n6805), .B2(n9753), .ZN(n6807)
         );
  AOI21_X1 U8558 ( .B1(n9769), .B2(n9764), .A(n6807), .ZN(n6808) );
  OAI211_X1 U8559 ( .C1(n9774), .C2(n9307), .A(n6809), .B(n6808), .ZN(P1_U3289) );
  OR2_X1 U8560 ( .A1(n9295), .A2(n9738), .ZN(n9216) );
  INV_X1 U8561 ( .A(n9216), .ZN(n9113) );
  INV_X2 U8562 ( .A(n9251), .ZN(n9295) );
  INV_X1 U8563 ( .A(n9753), .ZN(n9293) );
  INV_X1 U8564 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U8565 ( .A1(n9295), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9293), .B2(
        n6810), .ZN(n6811) );
  OAI21_X1 U8566 ( .B1(n9282), .B2(n6812), .A(n6811), .ZN(n6815) );
  INV_X1 U8567 ( .A(n4349), .ZN(n6947) );
  OAI22_X1 U8568 ( .A1(n6947), .A2(n9279), .B1(n9756), .B2(n6813), .ZN(n6814)
         );
  AOI211_X1 U8569 ( .C1(n9113), .C2(n5814), .A(n6815), .B(n6814), .ZN(n6818)
         );
  NOR2_X1 U8570 ( .A1(n9295), .A2(n9746), .ZN(n9135) );
  NAND2_X1 U8571 ( .A1(n6816), .A2(n9135), .ZN(n6817) );
  OAI211_X1 U8572 ( .C1(n6819), .C2(n9307), .A(n6818), .B(n6817), .ZN(P1_U3290) );
  OAI21_X1 U8573 ( .B1(n6821), .B2(n7670), .A(n6820), .ZN(n6852) );
  AOI211_X1 U8574 ( .C1(n7541), .C2(n6822), .A(n9291), .B(n6890), .ZN(n6856)
         );
  XNOR2_X1 U8575 ( .A(n7532), .B(n7670), .ZN(n6823) );
  OAI222_X1 U8576 ( .A1(n9740), .A2(n7536), .B1(n9738), .B2(n6947), .C1(n6823), 
        .C2(n9746), .ZN(n6853) );
  AOI211_X1 U8577 ( .C1(n9812), .C2(n6852), .A(n6856), .B(n6853), .ZN(n6827)
         );
  OAI22_X1 U8578 ( .A1(n9466), .A2(n7544), .B1(n9816), .B2(n5137), .ZN(n6824)
         );
  INV_X1 U8579 ( .A(n6824), .ZN(n6825) );
  OAI21_X1 U8580 ( .B1(n6827), .B2(n9814), .A(n6825), .ZN(P1_U3468) );
  INV_X1 U8581 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7847) );
  AOI22_X1 U8582 ( .A1(n7430), .A2(n7541), .B1(n9824), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6826) );
  OAI21_X1 U8583 ( .B1(n6827), .B2(n9824), .A(n6826), .ZN(P1_U3527) );
  INV_X1 U8584 ( .A(n6828), .ZN(n6830) );
  OAI21_X1 U8585 ( .B1(n9921), .B2(n6830), .A(n6829), .ZN(n6834) );
  XNOR2_X1 U8586 ( .A(n7922), .B(n6836), .ZN(n6832) );
  NAND2_X1 U8587 ( .A1(n6832), .A2(n6831), .ZN(n6980) );
  OAI21_X1 U8588 ( .B1(n6832), .B2(n6831), .A(n6980), .ZN(n6833) );
  AOI21_X1 U8589 ( .B1(n6834), .B2(n6833), .A(n6982), .ZN(n6841) );
  AOI21_X1 U8590 ( .B1(n8080), .B2(n6836), .A(n6835), .ZN(n6837) );
  OAI21_X1 U8591 ( .B1(n8093), .B2(n7044), .A(n6837), .ZN(n6839) );
  NOR2_X1 U8592 ( .A1(n8040), .A2(n7020), .ZN(n6838) );
  AOI211_X1 U8593 ( .C1(n8091), .C2(n8336), .A(n6839), .B(n6838), .ZN(n6840)
         );
  OAI21_X1 U8594 ( .B1(n6841), .B2(n8082), .A(n6840), .ZN(P2_U3170) );
  NAND2_X1 U8595 ( .A1(n6842), .A2(n10003), .ZN(n6843) );
  OAI21_X1 U8596 ( .B1(n10003), .B2(n5960), .A(n6843), .ZN(P2_U3459) );
  NAND2_X1 U8597 ( .A1(n6844), .A2(n6673), .ZN(n9931) );
  NOR2_X1 U8598 ( .A1(n9936), .A2(n9931), .ZN(n7874) );
  AOI22_X1 U8599 ( .A1(n8664), .A2(n6845), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9934), .ZN(n6846) );
  OAI21_X1 U8600 ( .B1(n6847), .B2(n9562), .A(n6846), .ZN(n6848) );
  AOI21_X1 U8601 ( .B1(n7874), .B2(n6849), .A(n6848), .ZN(n6850) );
  OAI21_X1 U8602 ( .B1(n6851), .B2(n9936), .A(n6850), .ZN(P2_U3232) );
  INV_X1 U8603 ( .A(n6852), .ZN(n6859) );
  NAND2_X1 U8604 ( .A1(n6853), .A2(n9251), .ZN(n6858) );
  NOR2_X1 U8605 ( .A1(n9756), .A2(n7544), .ZN(n6855) );
  OAI22_X1 U8606 ( .A1(n9251), .A2(n5142), .B1(n6952), .B2(n9753), .ZN(n6854)
         );
  AOI211_X1 U8607 ( .C1(n6856), .C2(n9764), .A(n6855), .B(n6854), .ZN(n6857)
         );
  OAI211_X1 U8608 ( .C1(n6859), .C2(n9307), .A(n6858), .B(n6857), .ZN(P1_U3288) );
  INV_X1 U8609 ( .A(n9135), .ZN(n9225) );
  OAI22_X1 U8610 ( .A1(n6861), .A2(n9279), .B1(n9282), .B2(n6860), .ZN(n6866)
         );
  NAND2_X1 U8611 ( .A1(n9113), .A2(n9013), .ZN(n6864) );
  OR2_X1 U8612 ( .A1(n9753), .A2(n9034), .ZN(n6862) );
  MUX2_X1 U8613 ( .A(n6862), .B(n7811), .S(n9295), .Z(n6863) );
  OAI211_X1 U8614 ( .C1(n5813), .C2(n9756), .A(n6864), .B(n6863), .ZN(n6865)
         );
  AOI211_X1 U8615 ( .C1(n9275), .C2(n6867), .A(n6866), .B(n6865), .ZN(n6868)
         );
  OAI21_X1 U8616 ( .B1(n6869), .B2(n9225), .A(n6868), .ZN(P1_U3291) );
  OAI22_X1 U8617 ( .A1(n6871), .A2(n9279), .B1(n9282), .B2(n6870), .ZN(n6872)
         );
  AOI21_X1 U8618 ( .B1(n9275), .B2(n6873), .A(n6872), .ZN(n6877) );
  AOI22_X1 U8619 ( .A1(n9295), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9293), .ZN(n6874) );
  OAI21_X1 U8620 ( .B1(n9756), .B2(n7745), .A(n6874), .ZN(n6875) );
  AOI21_X1 U8621 ( .B1(n9113), .B2(n9014), .A(n6875), .ZN(n6876) );
  OAI211_X1 U8622 ( .C1(n9295), .C2(n6878), .A(n6877), .B(n6876), .ZN(P1_U3292) );
  INV_X1 U8623 ( .A(n6879), .ZN(n6954) );
  AOI22_X1 U8624 ( .A1(n7662), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n9475), .ZN(n6880) );
  OAI21_X1 U8625 ( .B1(n6954), .B2(n6469), .A(n6880), .ZN(P1_U3336) );
  INV_X1 U8626 ( .A(n6898), .ZN(n7756) );
  INV_X1 U8627 ( .A(n6887), .ZN(n6881) );
  OAI21_X1 U8628 ( .B1(n6882), .B2(n6881), .A(n9331), .ZN(n6883) );
  AOI21_X1 U8629 ( .B1(n7756), .B2(n7543), .A(n6883), .ZN(n6885) );
  INV_X1 U8630 ( .A(n9010), .ZN(n7003) );
  OAI22_X1 U8631 ( .A1(n7003), .A2(n9738), .B1(n9739), .B2(n9740), .ZN(n6884)
         );
  NOR2_X1 U8632 ( .A1(n6885), .A2(n6884), .ZN(n9777) );
  OAI21_X1 U8633 ( .B1(n6888), .B2(n6887), .A(n6886), .ZN(n9780) );
  INV_X1 U8634 ( .A(n6901), .ZN(n6889) );
  OAI211_X1 U8635 ( .C1(n9778), .C2(n6890), .A(n6889), .B(n9761), .ZN(n9776)
         );
  INV_X1 U8636 ( .A(n6891), .ZN(n7011) );
  AOI22_X1 U8637 ( .A1(n9295), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7011), .B2(
        n9293), .ZN(n6893) );
  NAND2_X1 U8638 ( .A1(n9286), .A2(n7537), .ZN(n6892) );
  OAI211_X1 U8639 ( .C1(n9776), .C2(n9282), .A(n6893), .B(n6892), .ZN(n6894)
         );
  AOI21_X1 U8640 ( .B1(n9780), .B2(n9275), .A(n6894), .ZN(n6895) );
  OAI21_X1 U8641 ( .B1(n9777), .B2(n9295), .A(n6895), .ZN(P1_U3287) );
  OAI21_X1 U8642 ( .B1(n6897), .B2(n7533), .A(n6896), .ZN(n6960) );
  INV_X1 U8643 ( .A(n6960), .ZN(n6908) );
  NAND2_X1 U8644 ( .A1(n6898), .A2(n7543), .ZN(n6899) );
  OR2_X1 U8645 ( .A1(n6899), .A2(n7533), .ZN(n7090) );
  NAND2_X1 U8646 ( .A1(n6899), .A2(n7533), .ZN(n6900) );
  AOI21_X1 U8647 ( .B1(n7090), .B2(n6900), .A(n9746), .ZN(n6958) );
  OAI211_X1 U8648 ( .C1(n6901), .C2(n6970), .A(n9761), .B(n9759), .ZN(n6957)
         );
  OAI22_X1 U8649 ( .A1(n9251), .A2(n5191), .B1(n6972), .B2(n9753), .ZN(n6902)
         );
  AOI21_X1 U8650 ( .B1(n9211), .B2(n9008), .A(n6902), .ZN(n6903) );
  OAI21_X1 U8651 ( .B1(n7536), .B2(n9216), .A(n6903), .ZN(n6904) );
  AOI21_X1 U8652 ( .B1(n9286), .B2(n6961), .A(n6904), .ZN(n6905) );
  OAI21_X1 U8653 ( .B1(n9282), .B2(n6957), .A(n6905), .ZN(n6906) );
  AOI21_X1 U8654 ( .B1(n6958), .B2(n9251), .A(n6906), .ZN(n6907) );
  OAI21_X1 U8655 ( .B1(n6908), .B2(n9307), .A(n6907), .ZN(P1_U3286) );
  INV_X1 U8656 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U8657 ( .A1(n6930), .A2(n6910), .ZN(n6911) );
  INV_X1 U8658 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9993) );
  XNOR2_X1 U8659 ( .A(n6933), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U8660 ( .A1(n6933), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6912) );
  AOI21_X1 U8661 ( .B1(n9996), .B2(n6913), .A(n7076), .ZN(n6941) );
  INV_X1 U8662 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6914) );
  MUX2_X1 U8663 ( .A(n6915), .B(n6914), .S(n8473), .Z(n6916) );
  INV_X1 U8664 ( .A(n6933), .ZN(n9873) );
  NAND2_X1 U8665 ( .A1(n6916), .A2(n9873), .ZN(n6922) );
  XNOR2_X1 U8666 ( .A(n6916), .B(n6933), .ZN(n9876) );
  MUX2_X1 U8667 ( .A(n6016), .B(n9993), .S(n8473), .Z(n6919) );
  NOR2_X1 U8668 ( .A1(n6919), .A2(n6930), .ZN(n6921) );
  AOI21_X1 U8669 ( .B1(n6918), .B2(n6929), .A(n6917), .ZN(n9859) );
  AOI21_X1 U8670 ( .B1(n6930), .B2(n6919), .A(n6921), .ZN(n6920) );
  INV_X1 U8671 ( .A(n6920), .ZN(n9858) );
  NOR2_X1 U8672 ( .A1(n9859), .A2(n9858), .ZN(n9856) );
  MUX2_X1 U8673 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8473), .Z(n7061) );
  XNOR2_X1 U8674 ( .A(n7061), .B(n7074), .ZN(n6923) );
  OAI21_X1 U8675 ( .B1(n6924), .B2(n6923), .A(n7062), .ZN(n6939) );
  INV_X1 U8676 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8677 ( .A1(n9896), .A2(n7074), .ZN(n6926) );
  INV_X1 U8678 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10127) );
  NOR2_X1 U8679 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10127), .ZN(n7192) );
  INV_X1 U8680 ( .A(n7192), .ZN(n6925) );
  OAI211_X1 U8681 ( .C1(n6927), .C2(n9841), .A(n6926), .B(n6925), .ZN(n6938)
         );
  NOR2_X1 U8682 ( .A1(n6930), .A2(n6931), .ZN(n6932) );
  NOR2_X1 U8683 ( .A1(n6932), .A2(n9862), .ZN(n9880) );
  XNOR2_X1 U8684 ( .A(n6933), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U8685 ( .A1(n6933), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6934) );
  AOI21_X1 U8686 ( .B1(n7184), .B2(n6935), .A(n7069), .ZN(n6936) );
  NOR2_X1 U8687 ( .A1(n6936), .A2(n9905), .ZN(n6937) );
  AOI211_X1 U8688 ( .C1(n6411), .C2(n6939), .A(n6938), .B(n6937), .ZN(n6940)
         );
  OAI21_X1 U8689 ( .B1(n6941), .B2(n9909), .A(n6940), .ZN(P2_U3189) );
  NAND2_X1 U8690 ( .A1(n6943), .A2(n6942), .ZN(n6944) );
  XOR2_X1 U8691 ( .A(n6945), .B(n6944), .Z(n6946) );
  NAND2_X1 U8692 ( .A1(n6946), .A2(n8991), .ZN(n6951) );
  NAND2_X1 U8693 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9611) );
  INV_X1 U8694 ( .A(n9611), .ZN(n6949) );
  OAI22_X1 U8695 ( .A1(n7544), .A2(n9002), .B1(n8983), .B2(n6947), .ZN(n6948)
         );
  AOI211_X1 U8696 ( .C1(n8985), .C2(n6955), .A(n6949), .B(n6948), .ZN(n6950)
         );
  OAI211_X1 U8697 ( .C1(n8996), .C2(n6952), .A(n6951), .B(n6950), .ZN(P1_U3227) );
  INV_X1 U8698 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6953) );
  OAI222_X1 U8699 ( .A1(n9827), .A2(n8482), .B1(n8855), .B2(n6954), .C1(n6953), 
        .C2(n8853), .ZN(P2_U3276) );
  AOI22_X1 U8700 ( .A1(n6955), .A2(n9796), .B1(n9805), .B2(n9008), .ZN(n6956)
         );
  NAND2_X1 U8701 ( .A1(n6957), .A2(n6956), .ZN(n6959) );
  AOI211_X1 U8702 ( .C1(n9812), .C2(n6960), .A(n6959), .B(n6958), .ZN(n6965)
         );
  AOI22_X1 U8703 ( .A1(n7430), .A2(n6961), .B1(n9824), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6962) );
  OAI21_X1 U8704 ( .B1(n6965), .B2(n9824), .A(n6962), .ZN(P1_U3529) );
  OAI22_X1 U8705 ( .A1(n9466), .A2(n6970), .B1(n9816), .B2(n5186), .ZN(n6963)
         );
  INV_X1 U8706 ( .A(n6963), .ZN(n6964) );
  OAI21_X1 U8707 ( .B1(n6965), .B2(n9814), .A(n6964), .ZN(P1_U3474) );
  NAND2_X1 U8708 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  XNOR2_X1 U8709 ( .A(n6966), .B(n6969), .ZN(n6978) );
  NOR2_X1 U8710 ( .A1(n9002), .A2(n6970), .ZN(n6977) );
  NAND2_X1 U8711 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9513) );
  INV_X1 U8712 ( .A(n9513), .ZN(n6971) );
  AOI21_X1 U8713 ( .B1(n8985), .B2(n9008), .A(n6971), .ZN(n6975) );
  INV_X1 U8714 ( .A(n6972), .ZN(n6973) );
  NAND2_X1 U8715 ( .A1(n8980), .A2(n6973), .ZN(n6974) );
  OAI211_X1 U8716 ( .C1(n7536), .C2(n8983), .A(n6975), .B(n6974), .ZN(n6976)
         );
  AOI211_X1 U8717 ( .C1(n6978), .C2(n8991), .A(n6977), .B(n6976), .ZN(n6979)
         );
  INV_X1 U8718 ( .A(n6979), .ZN(P1_U3213) );
  INV_X1 U8719 ( .A(n6980), .ZN(n6981) );
  XNOR2_X1 U8720 ( .A(n7961), .B(n6985), .ZN(n7036) );
  XNOR2_X1 U8721 ( .A(n7036), .B(n8334), .ZN(n6983) );
  AOI21_X1 U8722 ( .B1(n4456), .B2(n6983), .A(n4377), .ZN(n6990) );
  NAND2_X1 U8723 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9868) );
  INV_X1 U8724 ( .A(n9868), .ZN(n6984) );
  AOI21_X1 U8725 ( .B1(n8080), .B2(n6985), .A(n6984), .ZN(n6986) );
  OAI21_X1 U8726 ( .B1(n8093), .B2(n7194), .A(n6986), .ZN(n6988) );
  NOR2_X1 U8727 ( .A1(n8040), .A2(n7029), .ZN(n6987) );
  AOI211_X1 U8728 ( .C1(n8091), .C2(n8335), .A(n6988), .B(n6987), .ZN(n6989)
         );
  OAI21_X1 U8729 ( .B1(n6990), .B2(n8082), .A(n6989), .ZN(P2_U3167) );
  INV_X1 U8730 ( .A(n6991), .ZN(n7035) );
  AOI22_X1 U8731 ( .A1(n4909), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n9475), .ZN(n6992) );
  OAI21_X1 U8732 ( .B1(n7035), .B2(n6469), .A(n6992), .ZN(P1_U3335) );
  INV_X1 U8733 ( .A(n9931), .ZN(n6993) );
  OR2_X1 U8734 ( .A1(n9919), .A2(n6993), .ZN(n9561) );
  OAI22_X1 U8735 ( .A1(n8695), .A2(n6994), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9553), .ZN(n6997) );
  MUX2_X1 U8736 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6995), .S(n9562), .Z(n6996)
         );
  AOI211_X1 U8737 ( .C1(n8698), .C2(n6998), .A(n6997), .B(n6996), .ZN(n6999)
         );
  INV_X1 U8738 ( .A(n6999), .ZN(P2_U3230) );
  NAND2_X1 U8739 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9060) );
  INV_X1 U8740 ( .A(n9060), .ZN(n7000) );
  AOI21_X1 U8741 ( .B1(n8985), .B2(n9009), .A(n7000), .ZN(n7002) );
  NAND2_X1 U8742 ( .A1(n8971), .A2(n7537), .ZN(n7001) );
  OAI211_X1 U8743 ( .C1(n7003), .C2(n8983), .A(n7002), .B(n7001), .ZN(n7010)
         );
  XNOR2_X1 U8744 ( .A(n7006), .B(n7005), .ZN(n7007) );
  XNOR2_X1 U8745 ( .A(n7004), .B(n7007), .ZN(n7008) );
  NOR2_X1 U8746 ( .A1(n7008), .A2(n8973), .ZN(n7009) );
  AOI211_X1 U8747 ( .C1(n7011), .C2(n8980), .A(n7010), .B(n7009), .ZN(n7012)
         );
  INV_X1 U8748 ( .A(n7012), .ZN(P1_U3239) );
  INV_X1 U8749 ( .A(n8172), .ZN(n7013) );
  XNOR2_X1 U8750 ( .A(n7014), .B(n7013), .ZN(n7017) );
  NAND2_X1 U8751 ( .A1(n8334), .A2(n8684), .ZN(n7015) );
  OAI21_X1 U8752 ( .B1(n9921), .B2(n9922), .A(n7015), .ZN(n7016) );
  AOI21_X1 U8753 ( .B1(n7017), .B2(n8671), .A(n7016), .ZN(n9943) );
  XNOR2_X1 U8754 ( .A(n7018), .B(n8172), .ZN(n9946) );
  NOR2_X1 U8755 ( .A1(n9562), .A2(n7019), .ZN(n7022) );
  OAI22_X1 U8756 ( .A1(n8695), .A2(n9944), .B1(n7020), .B2(n9553), .ZN(n7021)
         );
  AOI211_X1 U8757 ( .C1(n9946), .C2(n8698), .A(n7022), .B(n7021), .ZN(n7023)
         );
  OAI21_X1 U8758 ( .B1(n9936), .B2(n9943), .A(n7023), .ZN(P2_U3229) );
  XNOR2_X1 U8759 ( .A(n7024), .B(n8124), .ZN(n7025) );
  NAND2_X1 U8760 ( .A1(n7025), .A2(n8671), .ZN(n7027) );
  AOI22_X1 U8761 ( .A1(n8333), .A2(n8684), .B1(n8687), .B2(n8335), .ZN(n7026)
         );
  NAND2_X1 U8762 ( .A1(n7027), .A2(n7026), .ZN(n9949) );
  INV_X1 U8763 ( .A(n9949), .ZN(n7033) );
  OAI21_X1 U8764 ( .B1(n7028), .B2(n8124), .A(n7150), .ZN(n9951) );
  NOR2_X1 U8765 ( .A1(n9562), .A2(n6016), .ZN(n7031) );
  OAI22_X1 U8766 ( .A1(n8695), .A2(n9948), .B1(n7029), .B2(n9553), .ZN(n7030)
         );
  AOI211_X1 U8767 ( .C1(n9951), .C2(n8698), .A(n7031), .B(n7030), .ZN(n7032)
         );
  OAI21_X1 U8768 ( .B1(n9936), .B2(n7033), .A(n7032), .ZN(P2_U3228) );
  OAI222_X1 U8769 ( .A1(n8310), .A2(P2_U3151), .B1(n8855), .B2(n7035), .C1(
        n7034), .C2(n8853), .ZN(P2_U3275) );
  NOR2_X1 U8770 ( .A1(n7036), .A2(n8334), .ZN(n7040) );
  INV_X1 U8771 ( .A(n7040), .ZN(n7038) );
  XNOR2_X1 U8772 ( .A(n7922), .B(n9953), .ZN(n7186) );
  XNOR2_X1 U8773 ( .A(n7186), .B(n8333), .ZN(n7039) );
  INV_X1 U8774 ( .A(n7187), .ZN(n7042) );
  OAI21_X1 U8775 ( .B1(n4377), .B2(n7040), .A(n7039), .ZN(n7041) );
  NAND3_X1 U8776 ( .A1(n7042), .A2(n8088), .A3(n7041), .ZN(n7048) );
  INV_X1 U8777 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U8778 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10130), .ZN(n9872) );
  OAI22_X1 U8779 ( .A1(n8070), .A2(n7044), .B1(n7043), .B2(n8093), .ZN(n7045)
         );
  AOI211_X1 U8780 ( .C1(n7046), .C2(n8080), .A(n9872), .B(n7045), .ZN(n7047)
         );
  OAI211_X1 U8781 ( .C1(n7152), .C2(n8040), .A(n7048), .B(n7047), .ZN(P2_U3179) );
  OAI21_X1 U8782 ( .B1(n7049), .B2(n4461), .A(n7203), .ZN(n7050) );
  AOI22_X1 U8783 ( .A1(n7050), .A2(n9331), .B1(n9805), .B2(n7298), .ZN(n9800)
         );
  XNOR2_X1 U8784 ( .A(n7051), .B(n7679), .ZN(n9802) );
  NAND2_X1 U8785 ( .A1(n9802), .A2(n9275), .ZN(n7057) );
  INV_X1 U8786 ( .A(n7052), .ZN(n7321) );
  AOI22_X1 U8787 ( .A1(n9295), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7321), .B2(
        n9293), .ZN(n7053) );
  OAI21_X1 U8788 ( .B1(n9216), .B2(n9741), .A(n7053), .ZN(n7055) );
  OAI211_X1 U8789 ( .C1(n4455), .C2(n7318), .A(n9761), .B(n7209), .ZN(n9798)
         );
  NOR2_X1 U8790 ( .A1(n9798), .A2(n9282), .ZN(n7054) );
  AOI211_X1 U8791 ( .C1(n9286), .C2(n9797), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OAI211_X1 U8792 ( .C1(n9295), .C2(n9800), .A(n7057), .B(n7056), .ZN(P1_U3283) );
  MUX2_X1 U8793 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8473), .Z(n7058) );
  NOR2_X1 U8794 ( .A1(n7058), .A2(n7078), .ZN(n7109) );
  AND2_X1 U8795 ( .A1(n7058), .A2(n7078), .ZN(n7108) );
  NOR2_X1 U8796 ( .A1(n7109), .A2(n7108), .ZN(n7065) );
  MUX2_X1 U8797 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8473), .Z(n7059) );
  OR2_X1 U8798 ( .A1(n7059), .A2(n9893), .ZN(n7064) );
  XOR2_X1 U8799 ( .A(n9893), .B(n7059), .Z(n9899) );
  OR2_X1 U8800 ( .A1(n7061), .A2(n7060), .ZN(n7063) );
  NAND2_X1 U8801 ( .A1(n7063), .A2(n7062), .ZN(n9898) );
  NAND2_X1 U8802 ( .A1(n9899), .A2(n9898), .ZN(n9897) );
  NAND2_X1 U8803 ( .A1(n7064), .A2(n9897), .ZN(n7110) );
  XNOR2_X1 U8804 ( .A(n7065), .B(n7110), .ZN(n7086) );
  NOR2_X1 U8805 ( .A1(n7074), .A2(n7067), .ZN(n7068) );
  XNOR2_X1 U8806 ( .A(n9893), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n9904) );
  AOI21_X1 U8807 ( .B1(n7071), .B2(n7327), .A(n7118), .ZN(n7072) );
  NOR2_X1 U8808 ( .A1(n7072), .A2(n9905), .ZN(n7085) );
  INV_X1 U8809 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7083) );
  NOR2_X1 U8810 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  XNOR2_X1 U8811 ( .A(n9893), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U8812 ( .A1(n9893), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7077) );
  AOI21_X1 U8813 ( .B1(n6067), .B2(n7079), .A(n7126), .ZN(n7080) );
  OR2_X1 U8814 ( .A1(n7080), .A2(n9909), .ZN(n7082) );
  NOR2_X1 U8815 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6068), .ZN(n7270) );
  AOI21_X1 U8816 ( .B1(n9896), .B2(n7125), .A(n7270), .ZN(n7081) );
  OAI211_X1 U8817 ( .C1(n7083), .C2(n9841), .A(n7082), .B(n7081), .ZN(n7084)
         );
  AOI211_X1 U8818 ( .C1(n7086), .C2(n6411), .A(n7085), .B(n7084), .ZN(n7087)
         );
  INV_X1 U8819 ( .A(n7087), .ZN(P2_U3191) );
  INV_X1 U8820 ( .A(n7088), .ZN(n7137) );
  AOI22_X1 U8821 ( .A1(n7746), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n9475), .ZN(n7089) );
  OAI21_X1 U8822 ( .B1(n7137), .B2(n6469), .A(n7089), .ZN(P1_U3334) );
  NAND2_X1 U8823 ( .A1(n7090), .A2(n7675), .ZN(n9747) );
  INV_X1 U8824 ( .A(n7554), .ZN(n7091) );
  OR2_X1 U8825 ( .A1(n9747), .A2(n7091), .ZN(n9744) );
  NAND2_X1 U8826 ( .A1(n9744), .A2(n9742), .ZN(n7092) );
  XNOR2_X1 U8827 ( .A(n7092), .B(n4382), .ZN(n7093) );
  NAND2_X1 U8828 ( .A1(n7093), .A2(n9331), .ZN(n7095) );
  NAND2_X1 U8829 ( .A1(n9008), .A2(n9796), .ZN(n7094) );
  NAND2_X1 U8830 ( .A1(n7095), .A2(n7094), .ZN(n9791) );
  INV_X1 U8831 ( .A(n9791), .ZN(n7104) );
  OAI21_X1 U8832 ( .B1(n7097), .B2(n4382), .A(n7096), .ZN(n9793) );
  XOR2_X1 U8833 ( .A(n9788), .B(n9760), .Z(n7098) );
  AOI22_X1 U8834 ( .A1(n7098), .A2(n9761), .B1(n9805), .B2(n9007), .ZN(n9789)
         );
  OAI22_X1 U8835 ( .A1(n9251), .A2(n7099), .B1(n7164), .B2(n9753), .ZN(n7100)
         );
  AOI21_X1 U8836 ( .B1(n9286), .B2(n9788), .A(n7100), .ZN(n7101) );
  OAI21_X1 U8837 ( .B1(n9789), .B2(n9282), .A(n7101), .ZN(n7102) );
  AOI21_X1 U8838 ( .B1(n9793), .B2(n9275), .A(n7102), .ZN(n7103) );
  OAI21_X1 U8839 ( .B1(n9295), .B2(n7104), .A(n7103), .ZN(P1_U3284) );
  AOI22_X1 U8840 ( .A1(n8753), .A2(n7105), .B1(n10004), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7106) );
  OAI21_X1 U8841 ( .B1(n7107), .B2(n10004), .A(n7106), .ZN(P2_U3462) );
  INV_X1 U8842 ( .A(n7108), .ZN(n7111) );
  AOI21_X1 U8843 ( .B1(n7111), .B2(n7110), .A(n7109), .ZN(n7115) );
  INV_X1 U8844 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7381) );
  INV_X1 U8845 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7359) );
  MUX2_X1 U8846 ( .A(n7381), .B(n7359), .S(n8473), .Z(n7113) );
  AND2_X1 U8847 ( .A1(n7113), .A2(n7382), .ZN(n7370) );
  INV_X1 U8848 ( .A(n7370), .ZN(n7112) );
  OAI21_X1 U8849 ( .B1(n7382), .B2(n7113), .A(n7112), .ZN(n7114) );
  AOI21_X1 U8850 ( .B1(n7115), .B2(n7114), .A(n7369), .ZN(n7135) );
  INV_X1 U8851 ( .A(n7116), .ZN(n7117) );
  NOR2_X1 U8852 ( .A1(n7125), .A2(n7117), .ZN(n7119) );
  MUX2_X1 U8853 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7381), .S(n7382), .Z(n7120)
         );
  OAI21_X1 U8854 ( .B1(n4579), .B2(n4578), .A(n7384), .ZN(n7133) );
  INV_X1 U8855 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7123) );
  INV_X1 U8856 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7121) );
  NOR2_X1 U8857 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7121), .ZN(n7465) );
  AOI21_X1 U8858 ( .B1(n9896), .B2(n7382), .A(n7465), .ZN(n7122) );
  OAI21_X1 U8859 ( .B1(n7123), .B2(n9841), .A(n7122), .ZN(n7132) );
  NOR2_X1 U8860 ( .A1(n7125), .A2(n7124), .ZN(n7127) );
  MUX2_X1 U8861 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7359), .S(n7382), .Z(n7128)
         );
  NAND2_X1 U8862 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  AOI21_X1 U8863 ( .B1(n7361), .B2(n7130), .A(n9909), .ZN(n7131) );
  AOI211_X1 U8864 ( .C1(n9838), .C2(n7133), .A(n7132), .B(n7131), .ZN(n7134)
         );
  OAI21_X1 U8865 ( .B1(n7135), .B2(n9857), .A(n7134), .ZN(P2_U3192) );
  OAI222_X1 U8866 ( .A1(P2_U3151), .A2(n6674), .B1(n8855), .B2(n7137), .C1(
        n7136), .C2(n8853), .ZN(P2_U3274) );
  OAI21_X1 U8867 ( .B1(n7139), .B2(n7142), .A(n7141), .ZN(n7143) );
  NAND2_X1 U8868 ( .A1(n7143), .A2(n8991), .ZN(n7149) );
  INV_X1 U8869 ( .A(n9752), .ZN(n7147) );
  NAND2_X1 U8870 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9530) );
  INV_X1 U8871 ( .A(n9530), .ZN(n7144) );
  AOI21_X1 U8872 ( .B1(n8985), .B2(n9795), .A(n7144), .ZN(n7145) );
  OAI21_X1 U8873 ( .B1(n9739), .B2(n8983), .A(n7145), .ZN(n7146) );
  AOI21_X1 U8874 ( .B1(n7147), .B2(n8980), .A(n7146), .ZN(n7148) );
  OAI211_X1 U8875 ( .C1(n4642), .C2(n9002), .A(n7149), .B(n7148), .ZN(P1_U3221) );
  NAND2_X1 U8876 ( .A1(n7150), .A2(n8176), .ZN(n7151) );
  INV_X1 U8877 ( .A(n7154), .ZN(n8125) );
  XNOR2_X1 U8878 ( .A(n7151), .B(n8125), .ZN(n9956) );
  OAI22_X1 U8879 ( .A1(n8695), .A2(n9953), .B1(n7152), .B2(n9553), .ZN(n7159)
         );
  OAI211_X1 U8880 ( .C1(n7155), .C2(n7154), .A(n7153), .B(n8671), .ZN(n7157)
         );
  AOI22_X1 U8881 ( .A1(n8687), .A2(n8334), .B1(n8332), .B2(n8684), .ZN(n7156)
         );
  NAND2_X1 U8882 ( .A1(n7157), .A2(n7156), .ZN(n9954) );
  MUX2_X1 U8883 ( .A(n9954), .B(P2_REG2_REG_6__SCAN_IN), .S(n9936), .Z(n7158)
         );
  AOI211_X1 U8884 ( .C1(n8698), .C2(n9956), .A(n7159), .B(n7158), .ZN(n7160)
         );
  INV_X1 U8885 ( .A(n7160), .ZN(P2_U3227) );
  NAND2_X1 U8886 ( .A1(n7141), .A2(n7161), .ZN(n7162) );
  XOR2_X1 U8887 ( .A(n7163), .B(n7162), .Z(n7171) );
  INV_X1 U8888 ( .A(n7164), .ZN(n7168) );
  OR2_X1 U8889 ( .A1(n8983), .A2(n7165), .ZN(n7166) );
  NAND2_X1 U8890 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9546) );
  OAI211_X1 U8891 ( .C1(n8994), .C2(n8956), .A(n7166), .B(n9546), .ZN(n7167)
         );
  AOI21_X1 U8892 ( .B1(n7168), .B2(n8980), .A(n7167), .ZN(n7170) );
  NAND2_X1 U8893 ( .A1(n8971), .A2(n9788), .ZN(n7169) );
  OAI211_X1 U8894 ( .C1(n7171), .C2(n8973), .A(n7170), .B(n7169), .ZN(P1_U3231) );
  INV_X1 U8895 ( .A(n7172), .ZN(n7234) );
  AOI22_X1 U8896 ( .A1(n4959), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n9475), .ZN(n7173) );
  OAI21_X1 U8897 ( .B1(n7234), .B2(n6469), .A(n7173), .ZN(P1_U3333) );
  INV_X1 U8898 ( .A(n9919), .ZN(n7181) );
  NAND3_X1 U8899 ( .A1(n7175), .A2(n8193), .A3(n8188), .ZN(n7176) );
  NAND2_X1 U8900 ( .A1(n7174), .A2(n7176), .ZN(n9958) );
  OAI21_X1 U8901 ( .B1(n8193), .B2(n4460), .A(n7177), .ZN(n7179) );
  INV_X1 U8902 ( .A(n8331), .ZN(n7263) );
  OAI22_X1 U8903 ( .A1(n7263), .A2(n9920), .B1(n7194), .B2(n9922), .ZN(n7178)
         );
  AOI21_X1 U8904 ( .B1(n7179), .B2(n8671), .A(n7178), .ZN(n7180) );
  OAI21_X1 U8905 ( .B1(n7181), .B2(n9958), .A(n7180), .ZN(n9960) );
  OAI22_X1 U8906 ( .A1(n9958), .A2(n9931), .B1(n7199), .B2(n9553), .ZN(n7182)
         );
  NOR2_X1 U8907 ( .A1(n9960), .A2(n7182), .ZN(n7183) );
  MUX2_X1 U8908 ( .A(n7184), .B(n7183), .S(n9562), .Z(n7185) );
  OAI21_X1 U8909 ( .B1(n9957), .B2(n8695), .A(n7185), .ZN(P2_U3226) );
  XNOR2_X1 U8910 ( .A(n7922), .B(n9957), .ZN(n7188) );
  NOR2_X1 U8911 ( .A1(n7188), .A2(n8332), .ZN(n7249) );
  AOI21_X1 U8912 ( .B1(n7188), .B2(n8332), .A(n7249), .ZN(n7189) );
  NAND2_X1 U8913 ( .A1(n7190), .A2(n7189), .ZN(n7251) );
  OAI21_X1 U8914 ( .B1(n7190), .B2(n7189), .A(n7251), .ZN(n7191) );
  NAND2_X1 U8915 ( .A1(n7191), .A2(n8088), .ZN(n7198) );
  INV_X1 U8916 ( .A(n9957), .ZN(n7196) );
  AOI21_X1 U8917 ( .B1(n8066), .B2(n8331), .A(n7192), .ZN(n7193) );
  OAI21_X1 U8918 ( .B1(n8070), .B2(n7194), .A(n7193), .ZN(n7195) );
  AOI21_X1 U8919 ( .B1(n7196), .B2(n8080), .A(n7195), .ZN(n7197) );
  OAI211_X1 U8920 ( .C1(n7199), .C2(n8040), .A(n7198), .B(n7197), .ZN(P2_U3153) );
  INV_X1 U8921 ( .A(n7201), .ZN(n7681) );
  XNOR2_X1 U8922 ( .A(n7200), .B(n7681), .ZN(n7306) );
  OR2_X1 U8923 ( .A1(n9295), .A2(n7202), .ZN(n9758) );
  NAND2_X1 U8924 ( .A1(n7203), .A2(n7581), .ZN(n7204) );
  XNOR2_X1 U8925 ( .A(n7204), .B(n7681), .ZN(n7206) );
  OAI22_X1 U8926 ( .A1(n8956), .A2(n9738), .B1(n7400), .B2(n9740), .ZN(n7205)
         );
  AOI21_X1 U8927 ( .B1(n7206), .B2(n9331), .A(n7205), .ZN(n7207) );
  OAI21_X1 U8928 ( .B1(n7306), .B2(n9737), .A(n7207), .ZN(n7307) );
  NAND2_X1 U8929 ( .A1(n7307), .A2(n9251), .ZN(n7215) );
  INV_X1 U8930 ( .A(n7208), .ZN(n7226) );
  AOI211_X1 U8931 ( .C1(n8961), .C2(n7209), .A(n9291), .B(n7226), .ZN(n7308)
         );
  INV_X1 U8932 ( .A(n8961), .ZN(n7210) );
  NOR2_X1 U8933 ( .A1(n7210), .A2(n9756), .ZN(n7213) );
  OAI22_X1 U8934 ( .A1(n9251), .A2(n7211), .B1(n8959), .B2(n9753), .ZN(n7212)
         );
  AOI211_X1 U8935 ( .C1(n7308), .C2(n9764), .A(n7213), .B(n7212), .ZN(n7214)
         );
  OAI211_X1 U8936 ( .C1(n7306), .C2(n9758), .A(n7215), .B(n7214), .ZN(P1_U3282) );
  INV_X1 U8937 ( .A(n6230), .ZN(n7217) );
  AOI21_X1 U8938 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9479), .A(n7798), .ZN(
        n7216) );
  OAI21_X1 U8939 ( .B1(n7217), .B2(n6469), .A(n7216), .ZN(P1_U3332) );
  XNOR2_X1 U8940 ( .A(n7218), .B(n7222), .ZN(n7220) );
  NOR2_X1 U8941 ( .A1(n7317), .A2(n9738), .ZN(n7219) );
  AOI21_X1 U8942 ( .B1(n7220), .B2(n9331), .A(n7219), .ZN(n9810) );
  XNOR2_X1 U8943 ( .A(n7221), .B(n7222), .ZN(n9813) );
  NAND2_X1 U8944 ( .A1(n9813), .A2(n9275), .ZN(n7230) );
  INV_X1 U8945 ( .A(n7300), .ZN(n7223) );
  AOI22_X1 U8946 ( .A1(n9295), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7223), .B2(
        n9293), .ZN(n7224) );
  OAI21_X1 U8947 ( .B1(n9279), .B2(n7296), .A(n7224), .ZN(n7228) );
  INV_X1 U8948 ( .A(n9807), .ZN(n7225) );
  OAI211_X1 U8949 ( .C1(n7226), .C2(n7225), .A(n9761), .B(n7285), .ZN(n9808)
         );
  NOR2_X1 U8950 ( .A1(n9808), .A2(n9282), .ZN(n7227) );
  AOI211_X1 U8951 ( .C1(n9286), .C2(n9807), .A(n7228), .B(n7227), .ZN(n7229)
         );
  OAI211_X1 U8952 ( .C1(n9295), .C2(n9810), .A(n7230), .B(n7229), .ZN(P1_U3281) );
  NAND2_X1 U8953 ( .A1(n6230), .A2(n7495), .ZN(n7231) );
  OAI211_X1 U8954 ( .C1(n7232), .C2(n8853), .A(n7231), .B(n8322), .ZN(P2_U3272) );
  OAI222_X1 U8955 ( .A1(n7235), .A2(n9827), .B1(n8855), .B2(n7234), .C1(n7233), 
        .C2(n8853), .ZN(P2_U3273) );
  NAND2_X1 U8956 ( .A1(n7237), .A2(n7243), .ZN(n7238) );
  NAND3_X1 U8957 ( .A1(n7236), .A2(n8671), .A3(n7238), .ZN(n7240) );
  AOI22_X1 U8958 ( .A1(n8330), .A2(n8684), .B1(n8687), .B2(n8332), .ZN(n7239)
         );
  NAND2_X1 U8959 ( .A1(n7240), .A2(n7239), .ZN(n9963) );
  MUX2_X1 U8960 ( .A(n9963), .B(P2_REG2_REG_8__SCAN_IN), .S(n9936), .Z(n7241)
         );
  INV_X1 U8961 ( .A(n7241), .ZN(n7248) );
  NAND2_X1 U8962 ( .A1(n7174), .A2(n7242), .ZN(n7244) );
  XNOR2_X1 U8963 ( .A(n7244), .B(n6063), .ZN(n9965) );
  INV_X1 U8964 ( .A(n7260), .ZN(n7245) );
  OAI22_X1 U8965 ( .A1(n8695), .A2(n9962), .B1(n7245), .B2(n9553), .ZN(n7246)
         );
  AOI21_X1 U8966 ( .B1(n9965), .B2(n8698), .A(n7246), .ZN(n7247) );
  NAND2_X1 U8967 ( .A1(n7248), .A2(n7247), .ZN(P2_U3225) );
  INV_X1 U8968 ( .A(n7249), .ZN(n7250) );
  NAND2_X1 U8969 ( .A1(n7251), .A2(n7250), .ZN(n7253) );
  XNOR2_X1 U8970 ( .A(n7961), .B(n9962), .ZN(n7264) );
  XNOR2_X1 U8971 ( .A(n7264), .B(n8331), .ZN(n7252) );
  NAND2_X1 U8972 ( .A1(n7253), .A2(n7252), .ZN(n7269) );
  OAI21_X1 U8973 ( .B1(n7253), .B2(n7252), .A(n7269), .ZN(n7254) );
  NAND2_X1 U8974 ( .A1(n7254), .A2(n8088), .ZN(n7262) );
  NOR2_X1 U8975 ( .A1(n8099), .A2(n9962), .ZN(n7259) );
  NAND2_X1 U8976 ( .A1(n8091), .A2(n8332), .ZN(n7257) );
  NOR2_X1 U8977 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7255), .ZN(n9894) );
  INV_X1 U8978 ( .A(n9894), .ZN(n7256) );
  OAI211_X1 U8979 ( .C1(n7458), .C2(n8093), .A(n7257), .B(n7256), .ZN(n7258)
         );
  AOI211_X1 U8980 ( .C1(n7260), .C2(n8096), .A(n7259), .B(n7258), .ZN(n7261)
         );
  NAND2_X1 U8981 ( .A1(n7262), .A2(n7261), .ZN(P2_U3161) );
  NAND2_X1 U8982 ( .A1(n7264), .A2(n7263), .ZN(n7268) );
  XNOR2_X1 U8983 ( .A(n7922), .B(n7265), .ZN(n7457) );
  XNOR2_X1 U8984 ( .A(n7457), .B(n8330), .ZN(n7267) );
  NAND2_X1 U8985 ( .A1(n7269), .A2(n7266), .ZN(n7461) );
  NAND2_X1 U8986 ( .A1(n7461), .A2(n8088), .ZN(n7278) );
  AOI21_X1 U8987 ( .B1(n7269), .B2(n7268), .A(n7267), .ZN(n7277) );
  INV_X1 U8988 ( .A(n7326), .ZN(n7275) );
  NOR2_X1 U8989 ( .A1(n8099), .A2(n7492), .ZN(n7274) );
  NAND2_X1 U8990 ( .A1(n8091), .A2(n8331), .ZN(n7272) );
  INV_X1 U8991 ( .A(n7270), .ZN(n7271) );
  OAI211_X1 U8992 ( .C1(n7879), .C2(n8093), .A(n7272), .B(n7271), .ZN(n7273)
         );
  AOI211_X1 U8993 ( .C1(n7275), .C2(n8096), .A(n7274), .B(n7273), .ZN(n7276)
         );
  OAI21_X1 U8994 ( .B1(n7278), .B2(n7277), .A(n7276), .ZN(P2_U3171) );
  NAND2_X1 U8995 ( .A1(n7279), .A2(n7575), .ZN(n7282) );
  INV_X1 U8996 ( .A(n7280), .ZN(n7281) );
  AOI21_X1 U8997 ( .B1(n7684), .B2(n7282), .A(n7281), .ZN(n7283) );
  OAI222_X1 U8998 ( .A1(n9738), .A2(n7400), .B1(n9740), .B2(n7284), .C1(n9746), 
        .C2(n7283), .ZN(n7427) );
  INV_X1 U8999 ( .A(n7427), .ZN(n7293) );
  AOI211_X1 U9000 ( .C1(n7433), .C2(n7285), .A(n9291), .B(n7341), .ZN(n7428)
         );
  INV_X1 U9001 ( .A(n7433), .ZN(n7286) );
  NOR2_X1 U9002 ( .A1(n7286), .A2(n9756), .ZN(n7289) );
  OAI22_X1 U9003 ( .A1(n9251), .A2(n7287), .B1(n7403), .B2(n9753), .ZN(n7288)
         );
  AOI211_X1 U9004 ( .C1(n7428), .C2(n9764), .A(n7289), .B(n7288), .ZN(n7292)
         );
  XNOR2_X1 U9005 ( .A(n7290), .B(n7684), .ZN(n7429) );
  NAND2_X1 U9006 ( .A1(n7429), .A2(n9275), .ZN(n7291) );
  OAI211_X1 U9007 ( .C1(n7293), .C2(n9295), .A(n7292), .B(n7291), .ZN(P1_U3280) );
  XOR2_X1 U9008 ( .A(n7294), .B(n7295), .Z(n7303) );
  NAND2_X1 U9009 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9644) );
  OAI21_X1 U9010 ( .B1(n8994), .B2(n7296), .A(n9644), .ZN(n7297) );
  AOI21_X1 U9011 ( .B1(n8999), .B2(n7298), .A(n7297), .ZN(n7299) );
  OAI21_X1 U9012 ( .B1(n8996), .B2(n7300), .A(n7299), .ZN(n7301) );
  AOI21_X1 U9013 ( .B1(n9807), .B2(n8971), .A(n7301), .ZN(n7302) );
  OAI21_X1 U9014 ( .B1(n7303), .B2(n8973), .A(n7302), .ZN(P1_U3224) );
  INV_X1 U9015 ( .A(n7304), .ZN(n7336) );
  AOI22_X1 U9016 ( .A1(n5727), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n9475), .ZN(n7305) );
  OAI21_X1 U9017 ( .B1(n7336), .B2(n6469), .A(n7305), .ZN(P1_U3331) );
  INV_X1 U9018 ( .A(n7306), .ZN(n7309) );
  AOI211_X1 U9019 ( .C1(n9787), .C2(n7309), .A(n7308), .B(n7307), .ZN(n7312)
         );
  INV_X1 U9020 ( .A(n9466), .ZN(n7432) );
  AOI22_X1 U9021 ( .A1(n8961), .A2(n7432), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9814), .ZN(n7310) );
  OAI21_X1 U9022 ( .B1(n7312), .B2(n9814), .A(n7310), .ZN(P1_U3486) );
  AOI22_X1 U9023 ( .A1(n8961), .A2(n7430), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9824), .ZN(n7311) );
  OAI21_X1 U9024 ( .B1(n7312), .B2(n9824), .A(n7311), .ZN(P1_U3533) );
  XNOR2_X1 U9025 ( .A(n7313), .B(n8951), .ZN(n7315) );
  NOR2_X1 U9026 ( .A1(n7315), .A2(n7314), .ZN(n8950) );
  AOI21_X1 U9027 ( .B1(n7315), .B2(n7314), .A(n8950), .ZN(n7323) );
  OR2_X1 U9028 ( .A1(n8983), .A2(n9741), .ZN(n7316) );
  NAND2_X1 U9029 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9498) );
  OAI211_X1 U9030 ( .C1(n8994), .C2(n7317), .A(n7316), .B(n9498), .ZN(n7320)
         );
  NOR2_X1 U9031 ( .A1(n7318), .A2(n9002), .ZN(n7319) );
  AOI211_X1 U9032 ( .C1(n7321), .C2(n8980), .A(n7320), .B(n7319), .ZN(n7322)
         );
  OAI21_X1 U9033 ( .B1(n7323), .B2(n8973), .A(n7322), .ZN(P1_U3217) );
  OAI21_X1 U9034 ( .B1(n4453), .B2(n8127), .A(n7324), .ZN(n7325) );
  AOI222_X1 U9035 ( .A1(n8671), .A2(n7325), .B1(n8329), .B2(n8684), .C1(n8331), 
        .C2(n8687), .ZN(n7485) );
  NOR2_X1 U9036 ( .A1(n8695), .A2(n7492), .ZN(n7329) );
  OAI22_X1 U9037 ( .A1(n9562), .A2(n7327), .B1(n7326), .B2(n9553), .ZN(n7328)
         );
  NOR2_X1 U9038 ( .A1(n7329), .A2(n7328), .ZN(n7334) );
  NAND2_X1 U9039 ( .A1(n7331), .A2(n8127), .ZN(n7332) );
  AND2_X1 U9040 ( .A1(n7330), .A2(n7332), .ZN(n7487) );
  NAND2_X1 U9041 ( .A1(n7487), .A2(n8698), .ZN(n7333) );
  OAI211_X1 U9042 ( .C1(n7485), .C2(n9936), .A(n7334), .B(n7333), .ZN(P2_U3224) );
  OAI222_X1 U9043 ( .A1(n6362), .A2(P2_U3151), .B1(n8855), .B2(n7336), .C1(
        n7335), .C2(n8853), .ZN(P2_U3271) );
  NAND2_X1 U9044 ( .A1(n7280), .A2(n7761), .ZN(n7337) );
  XOR2_X1 U9045 ( .A(n7685), .B(n7337), .Z(n7338) );
  AOI222_X1 U9046 ( .A1(n9331), .A2(n7338), .B1(n9302), .B2(n9805), .C1(n9804), 
        .C2(n9796), .ZN(n9408) );
  XNOR2_X1 U9047 ( .A(n7339), .B(n7685), .ZN(n9411) );
  NAND2_X1 U9048 ( .A1(n9411), .A2(n9275), .ZN(n7346) );
  OAI22_X1 U9049 ( .A1(n9251), .A2(n7340), .B1(n8862), .B2(n9753), .ZN(n7343)
         );
  OAI211_X1 U9050 ( .C1(n9409), .C2(n7341), .A(n4378), .B(n9761), .ZN(n9407)
         );
  NOR2_X1 U9051 ( .A1(n9407), .A2(n9282), .ZN(n7342) );
  AOI211_X1 U9052 ( .C1(n9286), .C2(n7344), .A(n7343), .B(n7342), .ZN(n7345)
         );
  OAI211_X1 U9053 ( .C1(n9295), .C2(n9408), .A(n7346), .B(n7345), .ZN(P1_U3279) );
  NAND2_X1 U9054 ( .A1(n7348), .A2(n7347), .ZN(n8129) );
  NAND2_X1 U9055 ( .A1(n7330), .A2(n8195), .ZN(n7349) );
  XOR2_X1 U9056 ( .A(n8129), .B(n7349), .Z(n7352) );
  INV_X1 U9057 ( .A(n7352), .ZN(n9970) );
  INV_X1 U9058 ( .A(n7874), .ZN(n7358) );
  XNOR2_X1 U9059 ( .A(n7350), .B(n8129), .ZN(n7354) );
  OAI22_X1 U9060 ( .A1(n8680), .A2(n9920), .B1(n7458), .B2(n9922), .ZN(n7351)
         );
  AOI21_X1 U9061 ( .B1(n7352), .B2(n9919), .A(n7351), .ZN(n7353) );
  OAI21_X1 U9062 ( .B1(n7354), .B2(n9928), .A(n7353), .ZN(n9972) );
  NAND2_X1 U9063 ( .A1(n9972), .A2(n9562), .ZN(n7357) );
  OAI22_X1 U9064 ( .A1(n9562), .A2(n7381), .B1(n7464), .B2(n9553), .ZN(n7355)
         );
  AOI21_X1 U9065 ( .B1(n8664), .B2(n7456), .A(n7355), .ZN(n7356) );
  OAI211_X1 U9066 ( .C1(n9970), .C2(n7358), .A(n7357), .B(n7356), .ZN(P2_U3223) );
  OR2_X1 U9067 ( .A1(n7382), .A2(n7359), .ZN(n7360) );
  NOR2_X1 U9068 ( .A1(n7386), .A2(n7362), .ZN(n7363) );
  INV_X1 U9069 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10001) );
  OR2_X1 U9070 ( .A1(n7390), .A2(n7376), .ZN(n8342) );
  NAND2_X1 U9071 ( .A1(n7390), .A2(n7376), .ZN(n7364) );
  NAND2_X1 U9072 ( .A1(n8342), .A2(n7364), .ZN(n7366) );
  INV_X1 U9073 ( .A(n8343), .ZN(n7365) );
  AOI21_X1 U9074 ( .B1(n7367), .B2(n7366), .A(n7365), .ZN(n7397) );
  INV_X1 U9075 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7368) );
  MUX2_X1 U9076 ( .A(n7368), .B(n10001), .S(n8473), .Z(n7372) );
  AND2_X1 U9077 ( .A1(n7372), .A2(n7386), .ZN(n7373) );
  INV_X1 U9078 ( .A(n7373), .ZN(n7371) );
  OAI21_X1 U9079 ( .B1(n7386), .B2(n7372), .A(n7371), .ZN(n7420) );
  MUX2_X1 U9080 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8473), .Z(n7375) );
  INV_X1 U9081 ( .A(n7390), .ZN(n7374) );
  AND2_X1 U9082 ( .A1(n7375), .A2(n7374), .ZN(n8337) );
  INV_X1 U9083 ( .A(n8337), .ZN(n7378) );
  MUX2_X1 U9084 ( .A(n7388), .B(n7376), .S(n8473), .Z(n7377) );
  NAND2_X1 U9085 ( .A1(n7377), .A2(n7390), .ZN(n8338) );
  NAND2_X1 U9086 ( .A1(n7378), .A2(n8338), .ZN(n7379) );
  XNOR2_X1 U9087 ( .A(n8339), .B(n7379), .ZN(n7380) );
  NAND2_X1 U9088 ( .A1(n7380), .A2(n6411), .ZN(n7396) );
  OR2_X1 U9089 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  XNOR2_X1 U9090 ( .A(n7386), .B(n7385), .ZN(n7414) );
  NOR2_X1 U9091 ( .A1(n7386), .A2(n7385), .ZN(n7387) );
  OR2_X1 U9092 ( .A1(n7390), .A2(n7388), .ZN(n8346) );
  NAND2_X1 U9093 ( .A1(n7390), .A2(n7388), .ZN(n7389) );
  OAI21_X1 U9094 ( .B1(n4450), .B2(n4462), .A(n8347), .ZN(n7394) );
  INV_X1 U9095 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7392) );
  INV_X1 U9096 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U9097 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10222), .ZN(n7978) );
  AOI21_X1 U9098 ( .B1(n9896), .B2(n7390), .A(n7978), .ZN(n7391) );
  OAI21_X1 U9099 ( .B1(n7392), .B2(n9841), .A(n7391), .ZN(n7393) );
  AOI21_X1 U9100 ( .B1(n7394), .B2(n9838), .A(n7393), .ZN(n7395) );
  OAI211_X1 U9101 ( .C1(n7397), .C2(n9909), .A(n7396), .B(n7395), .ZN(P2_U3194) );
  XOR2_X1 U9102 ( .A(n7398), .B(n7399), .Z(n7406) );
  NAND2_X1 U9103 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9661) );
  OAI21_X1 U9104 ( .B1(n8983), .B2(n7400), .A(n9661), .ZN(n7401) );
  AOI21_X1 U9105 ( .B1(n8985), .B2(n9005), .A(n7401), .ZN(n7402) );
  OAI21_X1 U9106 ( .B1(n8996), .B2(n7403), .A(n7402), .ZN(n7404) );
  AOI21_X1 U9107 ( .B1(n7433), .B2(n8971), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9108 ( .B1(n7406), .B2(n8973), .A(n7405), .ZN(P1_U3234) );
  INV_X1 U9109 ( .A(n7407), .ZN(n7805) );
  INV_X1 U9110 ( .A(n7408), .ZN(n7409) );
  AOI22_X1 U9111 ( .A1(n7409), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9475), .ZN(n7410) );
  OAI21_X1 U9112 ( .B1(n7805), .B2(n6469), .A(n7410), .ZN(P1_U3330) );
  AOI21_X1 U9113 ( .B1(n10001), .B2(n7412), .A(n7411), .ZN(n7426) );
  AOI21_X1 U9114 ( .B1(n7368), .B2(n7414), .A(n7413), .ZN(n7415) );
  NOR2_X1 U9115 ( .A1(n7415), .A2(n9905), .ZN(n7424) );
  INV_X1 U9116 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7416) );
  OAI22_X1 U9117 ( .A1(n9871), .A2(n7417), .B1(n9841), .B2(n7416), .ZN(n7423)
         );
  AOI21_X1 U9118 ( .B1(n7420), .B2(n7419), .A(n7418), .ZN(n7421) );
  NAND2_X1 U9119 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8057) );
  OAI21_X1 U9120 ( .B1(n7421), .B2(n9857), .A(n8057), .ZN(n7422) );
  NOR3_X1 U9121 ( .A1(n7424), .A2(n7423), .A3(n7422), .ZN(n7425) );
  OAI21_X1 U9122 ( .B1(n7426), .B2(n9909), .A(n7425), .ZN(P2_U3193) );
  AOI211_X1 U9123 ( .C1(n9812), .C2(n7429), .A(n7428), .B(n7427), .ZN(n7435)
         );
  AOI22_X1 U9124 ( .A1(n7433), .A2(n7430), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9824), .ZN(n7431) );
  OAI21_X1 U9125 ( .B1(n7435), .B2(n9824), .A(n7431), .ZN(P1_U3535) );
  AOI22_X1 U9126 ( .A1(n7433), .A2(n7432), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9814), .ZN(n7434) );
  OAI21_X1 U9127 ( .B1(n7435), .B2(n9814), .A(n7434), .ZN(P1_U3492) );
  NAND2_X1 U9128 ( .A1(n7436), .A2(n7686), .ZN(n7437) );
  NAND2_X1 U9129 ( .A1(n7438), .A2(n7437), .ZN(n7439) );
  NAND2_X1 U9130 ( .A1(n7439), .A2(n9331), .ZN(n7441) );
  AOI22_X1 U9131 ( .A1(n9271), .A2(n9805), .B1(n9796), .B2(n9005), .ZN(n7440)
         );
  NAND2_X1 U9132 ( .A1(n7441), .A2(n7440), .ZN(n9402) );
  INV_X1 U9133 ( .A(n9402), .ZN(n7449) );
  XNOR2_X1 U9134 ( .A(n7442), .B(n7686), .ZN(n9404) );
  NAND2_X1 U9135 ( .A1(n9404), .A2(n9275), .ZN(n7448) );
  AOI211_X1 U9136 ( .C1(n7443), .C2(n4378), .A(n9291), .B(n4653), .ZN(n9403)
         );
  NOR2_X1 U9137 ( .A1(n9467), .A2(n9756), .ZN(n7446) );
  OAI22_X1 U9138 ( .A1(n9251), .A2(n7444), .B1(n8995), .B2(n9753), .ZN(n7445)
         );
  AOI211_X1 U9139 ( .C1(n9403), .C2(n9764), .A(n7446), .B(n7445), .ZN(n7447)
         );
  OAI211_X1 U9140 ( .C1(n9295), .C2(n7449), .A(n7448), .B(n7447), .ZN(P1_U3278) );
  INV_X1 U9141 ( .A(n7450), .ZN(n7454) );
  AOI22_X1 U9142 ( .A1(n7451), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9475), .ZN(n7452) );
  OAI21_X1 U9143 ( .B1(n7454), .B2(n6469), .A(n7452), .ZN(P1_U3329) );
  OAI222_X1 U9144 ( .A1(n7455), .A2(n9827), .B1(n8855), .B2(n7454), .C1(n7453), 
        .C2(n8853), .ZN(P2_U3269) );
  XNOR2_X1 U9145 ( .A(n7456), .B(n7961), .ZN(n7463) );
  INV_X1 U9146 ( .A(n7457), .ZN(n7459) );
  NAND2_X1 U9147 ( .A1(n7459), .A2(n8330), .ZN(n7460) );
  AOI21_X1 U9148 ( .B1(n7463), .B2(n7462), .A(n7882), .ZN(n7472) );
  INV_X1 U9149 ( .A(n7464), .ZN(n7470) );
  NOR2_X1 U9150 ( .A1(n8099), .A2(n9968), .ZN(n7469) );
  NAND2_X1 U9151 ( .A1(n8091), .A2(n8330), .ZN(n7467) );
  INV_X1 U9152 ( .A(n7465), .ZN(n7466) );
  OAI211_X1 U9153 ( .C1(n8680), .C2(n8093), .A(n7467), .B(n7466), .ZN(n7468)
         );
  AOI211_X1 U9154 ( .C1(n7470), .C2(n8096), .A(n7469), .B(n7468), .ZN(n7471)
         );
  OAI21_X1 U9155 ( .B1(n7472), .B2(n8082), .A(n7471), .ZN(P2_U3157) );
  NAND2_X1 U9156 ( .A1(n7473), .A2(n8201), .ZN(n7474) );
  XOR2_X1 U9157 ( .A(n8130), .B(n7474), .Z(n9975) );
  XNOR2_X1 U9158 ( .A(n7475), .B(n8130), .ZN(n7476) );
  OAI222_X1 U9159 ( .A1(n9920), .A2(n9558), .B1(n9922), .B2(n7879), .C1(n9928), 
        .C2(n7476), .ZN(n9976) );
  NAND2_X1 U9160 ( .A1(n9976), .A2(n9562), .ZN(n7479) );
  OAI22_X1 U9161 ( .A1(n9562), .A2(n7368), .B1(n8055), .B2(n9553), .ZN(n7477)
         );
  AOI21_X1 U9162 ( .B1(n8664), .B2(n9978), .A(n7477), .ZN(n7478) );
  OAI211_X1 U9163 ( .C1(n8667), .C2(n9975), .A(n7479), .B(n7478), .ZN(P2_U3222) );
  INV_X1 U9164 ( .A(n7480), .ZN(n7484) );
  AOI21_X1 U9165 ( .B1(n8850), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7481), .ZN(
        n7482) );
  OAI21_X1 U9166 ( .B1(n7484), .B2(n8855), .A(n7482), .ZN(P2_U3268) );
  AOI22_X1 U9167 ( .A1(n4358), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9475), .ZN(n7483) );
  OAI21_X1 U9168 ( .B1(n7484), .B2(n6469), .A(n7483), .ZN(P1_U3328) );
  INV_X1 U9169 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7488) );
  INV_X1 U9170 ( .A(n7485), .ZN(n7486) );
  AOI21_X1 U9171 ( .B1(n7487), .B2(n9980), .A(n7486), .ZN(n7490) );
  MUX2_X1 U9172 ( .A(n7488), .B(n7490), .S(n9986), .Z(n7489) );
  OAI21_X1 U9173 ( .B1(n7492), .B2(n8807), .A(n7489), .ZN(P2_U3417) );
  MUX2_X1 U9174 ( .A(n6067), .B(n7490), .S(n10003), .Z(n7491) );
  OAI21_X1 U9175 ( .B1(n7492), .B2(n8736), .A(n7491), .ZN(P2_U3468) );
  INV_X1 U9176 ( .A(n6277), .ZN(n7494) );
  AOI22_X1 U9177 ( .A1(n4355), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9475), .ZN(n7493) );
  OAI21_X1 U9178 ( .B1(n7494), .B2(n6469), .A(n7493), .ZN(P1_U3327) );
  NAND2_X1 U9179 ( .A1(n6277), .A2(n7495), .ZN(n7497) );
  OAI211_X1 U9180 ( .C1(n8853), .C2(n7498), .A(n7497), .B(n7496), .ZN(P2_U3267) );
  INV_X1 U9181 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7508) );
  XNOR2_X1 U9182 ( .A(n7499), .B(n7694), .ZN(n9097) );
  OAI21_X1 U9183 ( .B1(n7501), .B2(n7694), .A(n7500), .ZN(n9106) );
  OAI22_X1 U9184 ( .A1(n9327), .A2(n9738), .B1(n7502), .B2(n9740), .ZN(n7505)
         );
  AOI211_X1 U9185 ( .C1(n7504), .C2(n9112), .A(n9291), .B(n5899), .ZN(n9105)
         );
  AOI211_X1 U9186 ( .C1(n9331), .C2(n9106), .A(n7505), .B(n9105), .ZN(n7506)
         );
  INV_X1 U9187 ( .A(n7506), .ZN(n7507) );
  AOI21_X1 U9188 ( .B1(n9097), .B2(n9812), .A(n7507), .ZN(n7510) );
  MUX2_X1 U9189 ( .A(n7508), .B(n7510), .S(n9816), .Z(n7509) );
  OAI21_X1 U9190 ( .B1(n9098), .B2(n9466), .A(n7509), .ZN(P1_U3518) );
  MUX2_X1 U9191 ( .A(n7511), .B(n7510), .S(n9826), .Z(n7512) );
  OAI21_X1 U9192 ( .B1(n9098), .B2(n9406), .A(n7512), .ZN(P1_U3550) );
  INV_X1 U9193 ( .A(SI_29_), .ZN(n7516) );
  INV_X1 U9194 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8102) );
  INV_X1 U9195 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7518) );
  MUX2_X1 U9196 ( .A(n8102), .B(n7518), .S(n7525), .Z(n7519) );
  INV_X1 U9197 ( .A(SI_30_), .ZN(n10226) );
  NAND2_X1 U9198 ( .A1(n7519), .A2(n10226), .ZN(n7522) );
  INV_X1 U9199 ( .A(n7519), .ZN(n7520) );
  NAND2_X1 U9200 ( .A1(n7520), .A2(SI_30_), .ZN(n7521) );
  NAND2_X1 U9201 ( .A1(n7522), .A2(n7521), .ZN(n7523) );
  INV_X1 U9202 ( .A(n8101), .ZN(n9478) );
  OAI222_X1 U9203 ( .A1(n5949), .A2(P2_U3151), .B1(n8855), .B2(n9478), .C1(
        n8102), .C2(n8853), .ZN(P2_U3265) );
  MUX2_X1 U9204 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7525), .Z(n7527) );
  INV_X1 U9205 ( .A(SI_31_), .ZN(n7526) );
  XNOR2_X1 U9206 ( .A(n7527), .B(n7526), .ZN(n7528) );
  XNOR2_X1 U9207 ( .A(n7529), .B(n7528), .ZN(n8845) );
  NAND2_X1 U9208 ( .A1(n8845), .A2(n4352), .ZN(n7531) );
  NAND2_X1 U9209 ( .A1(n7645), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7530) );
  NOR2_X1 U9210 ( .A1(n9417), .A2(n9076), .ZN(n7786) );
  NAND2_X1 U9211 ( .A1(n7608), .A2(n7777), .ZN(n7607) );
  INV_X1 U9212 ( .A(n7769), .ZN(n7569) );
  NAND4_X1 U9213 ( .A1(n7532), .A2(n7654), .A3(n7543), .A4(n7752), .ZN(n7553)
         );
  INV_X1 U9214 ( .A(n7533), .ZN(n7552) );
  AND4_X1 U9215 ( .A1(n7535), .A2(n7674), .A3(n7534), .A4(n7660), .ZN(n7549)
         );
  OAI21_X1 U9216 ( .B1(n7536), .B2(n7654), .A(n9778), .ZN(n7540) );
  NAND2_X1 U9217 ( .A1(n7536), .A2(n7654), .ZN(n7538) );
  NAND2_X1 U9218 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  NAND2_X1 U9219 ( .A1(n7540), .A2(n7539), .ZN(n7547) );
  NOR2_X1 U9220 ( .A1(n9010), .A2(n7660), .ZN(n7542) );
  NAND3_X1 U9221 ( .A1(n7543), .A2(n7542), .A3(n7541), .ZN(n7546) );
  NAND4_X1 U9222 ( .A1(n7674), .A2(n7544), .A3(n9010), .A4(n7660), .ZN(n7545)
         );
  NAND3_X1 U9223 ( .A1(n7547), .A2(n7546), .A3(n7545), .ZN(n7548) );
  AOI21_X1 U9224 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7551) );
  NAND3_X1 U9225 ( .A1(n7553), .A2(n7552), .A3(n7551), .ZN(n7562) );
  NAND2_X1 U9226 ( .A1(n7554), .A2(n7675), .ZN(n7557) );
  NAND2_X1 U9227 ( .A1(n9742), .A2(n7555), .ZN(n7556) );
  MUX2_X1 U9228 ( .A(n7557), .B(n7556), .S(n7654), .Z(n7558) );
  INV_X1 U9229 ( .A(n7558), .ZN(n7561) );
  MUX2_X1 U9230 ( .A(n7678), .B(n7559), .S(n7660), .Z(n7560) );
  INV_X1 U9231 ( .A(n7563), .ZN(n7564) );
  OAI21_X1 U9232 ( .B1(n7578), .B2(n7564), .A(n7581), .ZN(n7565) );
  NAND3_X1 U9233 ( .A1(n7565), .A2(n7574), .A3(n7576), .ZN(n7566) );
  NAND2_X1 U9234 ( .A1(n7591), .A2(n7587), .ZN(n7766) );
  AOI21_X1 U9235 ( .B1(n7569), .B2(n7774), .A(n7568), .ZN(n7570) );
  INV_X1 U9236 ( .A(n7571), .ZN(n7572) );
  INV_X1 U9237 ( .A(n7573), .ZN(n7579) );
  NAND2_X1 U9238 ( .A1(n7575), .A2(n7574), .ZN(n7580) );
  INV_X1 U9239 ( .A(n7576), .ZN(n7577) );
  NOR2_X1 U9240 ( .A1(n7580), .A2(n7577), .ZN(n7758) );
  OAI21_X1 U9241 ( .B1(n7579), .B2(n7578), .A(n7758), .ZN(n7586) );
  INV_X1 U9242 ( .A(n7580), .ZN(n7585) );
  NAND2_X1 U9243 ( .A1(n7582), .A2(n7581), .ZN(n7584) );
  AOI21_X1 U9244 ( .B1(n7585), .B2(n7584), .A(n4514), .ZN(n7762) );
  NAND2_X1 U9245 ( .A1(n7586), .A2(n7762), .ZN(n7588) );
  NAND2_X1 U9246 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  NAND2_X1 U9247 ( .A1(n7590), .A2(n7589), .ZN(n7592) );
  NAND4_X1 U9248 ( .A1(n7770), .A2(n7592), .A3(n7769), .A4(n7591), .ZN(n7593)
         );
  INV_X1 U9249 ( .A(n7689), .ZN(n9273) );
  INV_X1 U9250 ( .A(n7599), .ZN(n7603) );
  AOI21_X1 U9251 ( .B1(n7600), .B2(n9285), .A(n7603), .ZN(n7775) );
  NAND3_X1 U9252 ( .A1(n7777), .A2(n7776), .A3(n7660), .ZN(n7601) );
  AOI21_X1 U9253 ( .B1(n7604), .B2(n7775), .A(n7601), .ZN(n7606) );
  NAND2_X1 U9254 ( .A1(n9234), .A2(n9217), .ZN(n7609) );
  NAND2_X1 U9255 ( .A1(n7609), .A2(n7782), .ZN(n7605) );
  AND2_X1 U9256 ( .A1(n7776), .A2(n7602), .ZN(n7771) );
  OR2_X1 U9257 ( .A1(n9222), .A2(n9375), .ZN(n7715) );
  NAND2_X1 U9258 ( .A1(n7715), .A2(n7608), .ZN(n7709) );
  NAND2_X1 U9259 ( .A1(n7610), .A2(n7609), .ZN(n7716) );
  MUX2_X1 U9260 ( .A(n7709), .B(n7716), .S(n7654), .Z(n7612) );
  MUX2_X1 U9261 ( .A(n7610), .B(n7715), .S(n7654), .Z(n7611) );
  OAI21_X1 U9262 ( .B1(n7613), .B2(n7612), .A(n7611), .ZN(n7619) );
  NAND2_X1 U9263 ( .A1(n7704), .A2(n7614), .ZN(n7717) );
  AOI21_X1 U9264 ( .B1(n7619), .B2(n9195), .A(n7618), .ZN(n7625) );
  INV_X1 U9265 ( .A(n9163), .ZN(n7622) );
  MUX2_X1 U9266 ( .A(n7620), .B(n7704), .S(n7654), .Z(n7621) );
  NAND2_X1 U9267 ( .A1(n7622), .A2(n7621), .ZN(n7624) );
  OAI21_X1 U9268 ( .B1(n7625), .B2(n7624), .A(n7623), .ZN(n7628) );
  INV_X1 U9269 ( .A(n7725), .ZN(n7665) );
  INV_X1 U9270 ( .A(n7708), .ZN(n7626) );
  OAI21_X1 U9271 ( .B1(n7628), .B2(n7665), .A(n7626), .ZN(n7627) );
  AOI21_X1 U9272 ( .B1(n7627), .B2(n7711), .A(n7724), .ZN(n7632) );
  OAI21_X1 U9273 ( .B1(n7628), .B2(n7708), .A(n7725), .ZN(n7630) );
  INV_X1 U9274 ( .A(n7724), .ZN(n7629) );
  INV_X1 U9275 ( .A(n7711), .ZN(n7785) );
  AOI21_X1 U9276 ( .B1(n7630), .B2(n7629), .A(n7785), .ZN(n7631) );
  MUX2_X2 U9277 ( .A(n7632), .B(n7631), .S(n7654), .Z(n7637) );
  NAND2_X1 U9278 ( .A1(n7638), .A2(n7636), .ZN(n7727) );
  AOI21_X1 U9279 ( .B1(n7637), .B2(n7728), .A(n7727), .ZN(n7634) );
  INV_X1 U9280 ( .A(n7633), .ZN(n7635) );
  NOR2_X1 U9281 ( .A1(n7634), .A2(n7635), .ZN(n7642) );
  INV_X1 U9282 ( .A(n7728), .ZN(n7702) );
  INV_X1 U9283 ( .A(n7638), .ZN(n7639) );
  NOR2_X1 U9284 ( .A1(n7640), .A2(n7639), .ZN(n7641) );
  MUX2_X1 U9285 ( .A(n7701), .B(n7712), .S(n7654), .Z(n7643) );
  OAI21_X2 U9286 ( .B1(n7644), .B2(n7697), .A(n7643), .ZN(n7653) );
  NAND2_X1 U9287 ( .A1(n8101), .A2(n4352), .ZN(n7647) );
  NAND2_X1 U9288 ( .A1(n7645), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7646) );
  INV_X1 U9289 ( .A(n7664), .ZN(n9003) );
  OAI21_X1 U9290 ( .B1(n9417), .B2(n9003), .A(n9076), .ZN(n7649) );
  OAI21_X1 U9291 ( .B1(n7660), .B2(n7652), .A(n4401), .ZN(n7797) );
  AOI211_X1 U9292 ( .C1(n7790), .C2(n7662), .A(n4959), .B(n7661), .ZN(n7796)
         );
  NAND2_X1 U9293 ( .A1(n9084), .A2(n7664), .ZN(n7713) );
  INV_X1 U9294 ( .A(n7713), .ZN(n7698) );
  NOR2_X1 U9295 ( .A1(n9084), .A2(n7664), .ZN(n7787) );
  INV_X1 U9296 ( .A(n9240), .ZN(n7690) );
  NAND4_X1 U9297 ( .A1(n7669), .A2(n7668), .A3(n7667), .A4(n7666), .ZN(n7672)
         );
  NOR3_X1 U9298 ( .A1(n7672), .A2(n7671), .A3(n7670), .ZN(n7676) );
  NAND4_X1 U9299 ( .A1(n7676), .A2(n7675), .A3(n7674), .A4(n7673), .ZN(n7677)
         );
  NOR4_X1 U9300 ( .A1(n7679), .A2(n7754), .A3(n7678), .A4(n7677), .ZN(n7680)
         );
  NAND3_X1 U9301 ( .A1(n7682), .A2(n7681), .A3(n7680), .ZN(n7683) );
  NOR4_X1 U9302 ( .A1(n7686), .A2(n7685), .A3(n7684), .A4(n7683), .ZN(n7687)
         );
  NAND3_X1 U9303 ( .A1(n9263), .A2(n9300), .A3(n7687), .ZN(n7688) );
  NOR4_X1 U9304 ( .A1(n9227), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n7691)
         );
  NAND4_X1 U9305 ( .A1(n9195), .A2(n9173), .A3(n7691), .A4(n9209), .ZN(n7692)
         );
  NOR4_X1 U9306 ( .A1(n7693), .A2(n9143), .A3(n9163), .A4(n7692), .ZN(n7695)
         );
  NAND3_X1 U9307 ( .A1(n7695), .A2(n7694), .A3(n9124), .ZN(n7696) );
  NOR4_X1 U9308 ( .A1(n7698), .A2(n7787), .A3(n7697), .A4(n7696), .ZN(n7700)
         );
  INV_X1 U9309 ( .A(n7790), .ZN(n7699) );
  NAND3_X1 U9310 ( .A1(n7700), .A2(n7699), .A3(n7652), .ZN(n7737) );
  NAND2_X1 U9311 ( .A1(n7701), .A2(n7633), .ZN(n7731) );
  NOR3_X2 U9312 ( .A1(n7731), .A2(n7702), .A3(n7724), .ZN(n7783) );
  NAND3_X1 U9313 ( .A1(n7719), .A2(n7704), .A3(n7703), .ZN(n7706) );
  NAND2_X1 U9314 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  NOR2_X1 U9315 ( .A1(n7708), .A2(n7707), .ZN(n7723) );
  INV_X1 U9316 ( .A(n7709), .ZN(n7710) );
  NAND2_X1 U9317 ( .A1(n7723), .A2(n7710), .ZN(n7780) );
  OAI21_X1 U9318 ( .B1(n7780), .B2(n4383), .A(n7711), .ZN(n7714) );
  NAND2_X1 U9319 ( .A1(n7713), .A2(n7712), .ZN(n7742) );
  AOI21_X1 U9320 ( .B1(n7783), .B2(n7714), .A(n7742), .ZN(n7734) );
  INV_X1 U9321 ( .A(n9076), .ZN(n7732) );
  INV_X1 U9322 ( .A(n7715), .ZN(n7721) );
  INV_X1 U9323 ( .A(n7716), .ZN(n7720) );
  INV_X1 U9324 ( .A(n7717), .ZN(n7718) );
  OAI211_X1 U9325 ( .C1(n7721), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7722)
         );
  NAND2_X1 U9326 ( .A1(n7723), .A2(n7722), .ZN(n7726) );
  AOI21_X1 U9327 ( .B1(n7726), .B2(n7725), .A(n7724), .ZN(n7729) );
  AOI21_X1 U9328 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(n7730) );
  NOR2_X1 U9329 ( .A1(n7731), .A2(n7730), .ZN(n7743) );
  AOI21_X1 U9330 ( .B1(n7732), .B2(n9084), .A(n7743), .ZN(n7733) );
  AOI22_X1 U9331 ( .A1(n7734), .A2(n7733), .B1(n7787), .B2(n9076), .ZN(n7736)
         );
  OAI211_X1 U9332 ( .C1(n7736), .C2(n7790), .A(n7735), .B(n7652), .ZN(n7738)
         );
  AOI21_X1 U9333 ( .B1(n7738), .B2(n7737), .A(n7662), .ZN(n7739) );
  NOR2_X1 U9334 ( .A1(n7743), .A2(n7742), .ZN(n7789) );
  INV_X1 U9335 ( .A(n7744), .ZN(n7749) );
  NAND2_X1 U9336 ( .A1(n5814), .A2(n5813), .ZN(n7748) );
  NAND2_X1 U9337 ( .A1(n9013), .A2(n7745), .ZN(n7747) );
  AND4_X1 U9338 ( .A1(n7749), .A2(n7748), .A3(n7747), .A4(n7746), .ZN(n7753)
         );
  NAND4_X1 U9339 ( .A1(n7753), .A2(n7752), .A3(n7751), .A4(n7750), .ZN(n7755)
         );
  AOI21_X1 U9340 ( .B1(n7756), .B2(n7755), .A(n7754), .ZN(n7760) );
  INV_X1 U9341 ( .A(n7757), .ZN(n7759) );
  OAI21_X1 U9342 ( .B1(n7760), .B2(n7759), .A(n7758), .ZN(n7763) );
  AND3_X1 U9343 ( .A1(n7763), .A2(n7762), .A3(n7761), .ZN(n7767) );
  OAI211_X1 U9344 ( .C1(n7767), .C2(n7766), .A(n7765), .B(n7764), .ZN(n7768)
         );
  NAND3_X1 U9345 ( .A1(n7770), .A2(n7769), .A3(n7768), .ZN(n7773) );
  INV_X1 U9346 ( .A(n7771), .ZN(n7772) );
  AOI21_X1 U9347 ( .B1(n7774), .B2(n7773), .A(n7772), .ZN(n7779) );
  INV_X1 U9348 ( .A(n7775), .ZN(n7778) );
  OAI211_X1 U9349 ( .C1(n7779), .C2(n7778), .A(n7777), .B(n7776), .ZN(n7781)
         );
  AOI21_X1 U9350 ( .B1(n7782), .B2(n7781), .A(n7780), .ZN(n7784) );
  OAI21_X1 U9351 ( .B1(n7785), .B2(n7784), .A(n7783), .ZN(n7788) );
  AOI211_X1 U9352 ( .C1(n7789), .C2(n7788), .A(n7787), .B(n7786), .ZN(n7791)
         );
  NOR2_X1 U9353 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  XNOR2_X1 U9354 ( .A(n5886), .B(n7792), .ZN(n7793) );
  NOR2_X1 U9355 ( .A1(n7793), .A2(n4909), .ZN(n7794) );
  AOI211_X1 U9356 ( .C1(n7797), .C2(n7796), .A(n7795), .B(n7794), .ZN(n7803)
         );
  NAND2_X1 U9357 ( .A1(n4355), .A2(n4358), .ZN(n7835) );
  NAND2_X1 U9358 ( .A1(n7798), .A2(n5747), .ZN(n7799) );
  OAI211_X1 U9359 ( .C1(n7800), .C2(n7835), .A(P1_B_REG_SCAN_IN), .B(n7799), 
        .ZN(n7801) );
  OAI21_X1 U9360 ( .B1(n7803), .B2(n7802), .A(n7801), .ZN(P1_U3242) );
  OAI222_X1 U9361 ( .A1(n7806), .A2(n9827), .B1(n8855), .B2(n7805), .C1(n7804), 
        .C2(n8853), .ZN(P2_U3270) );
  NAND2_X1 U9362 ( .A1(n9652), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7807) );
  OAI21_X1 U9363 ( .B1(n9652), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7807), .ZN(
        n9655) );
  INV_X1 U9364 ( .A(n9635), .ZN(n7808) );
  AOI22_X1 U9365 ( .A1(n9635), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n5335), .B2(
        n7808), .ZN(n9638) );
  NAND2_X1 U9366 ( .A1(n9489), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7809) );
  OAI21_X1 U9367 ( .B1(n9489), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7809), .ZN(
        n9492) );
  INV_X1 U9368 ( .A(n9537), .ZN(n7810) );
  AOI22_X1 U9369 ( .A1(n9537), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7099), .B2(
        n7810), .ZN(n9540) );
  NAND2_X1 U9370 ( .A1(n9602), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7819) );
  XNOR2_X1 U9371 ( .A(n9037), .B(n7811), .ZN(n9043) );
  XNOR2_X1 U9372 ( .A(n9018), .B(n7812), .ZN(n9020) );
  AND2_X1 U9373 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9027) );
  NAND2_X1 U9374 ( .A1(n9020), .A2(n9027), .ZN(n9019) );
  NAND2_X1 U9375 ( .A1(n9018), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U9376 ( .A1(n9019), .A2(n7813), .ZN(n9042) );
  NAND2_X1 U9377 ( .A1(n9043), .A2(n9042), .ZN(n9041) );
  NAND2_X1 U9378 ( .A1(n9037), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U9379 ( .A1(n9041), .A2(n7814), .ZN(n9052) );
  XNOR2_X1 U9380 ( .A(n9050), .B(n7815), .ZN(n9053) );
  NAND2_X1 U9381 ( .A1(n9052), .A2(n9053), .ZN(n9051) );
  NAND2_X1 U9382 ( .A1(n9050), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U9383 ( .A1(n9051), .A2(n7816), .ZN(n9585) );
  MUX2_X1 U9384 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6802), .S(n9587), .Z(n9586)
         );
  AND2_X1 U9385 ( .A1(n9585), .A2(n9586), .ZN(n9583) );
  AOI21_X1 U9386 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9587), .A(n9583), .ZN(
        n9605) );
  INV_X1 U9387 ( .A(n9602), .ZN(n7817) );
  AOI22_X1 U9388 ( .A1(n9602), .A2(n5142), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n7817), .ZN(n9604) );
  NOR2_X1 U9389 ( .A1(n9605), .A2(n9604), .ZN(n9603) );
  INV_X1 U9390 ( .A(n9603), .ZN(n7818) );
  NAND2_X1 U9391 ( .A1(n7819), .A2(n7818), .ZN(n9065) );
  XNOR2_X1 U9392 ( .A(n9063), .B(n7820), .ZN(n9066) );
  NAND2_X1 U9393 ( .A1(n9065), .A2(n9066), .ZN(n9064) );
  NAND2_X1 U9394 ( .A1(n9063), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U9395 ( .A1(n9064), .A2(n7821), .ZN(n9506) );
  MUX2_X1 U9396 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n5191), .S(n9508), .Z(n9507)
         );
  AND2_X1 U9397 ( .A1(n9506), .A2(n9507), .ZN(n9504) );
  AOI21_X1 U9398 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9508), .A(n9504), .ZN(
        n9523) );
  INV_X1 U9399 ( .A(n9521), .ZN(n7822) );
  AOI22_X1 U9400 ( .A1(n9521), .A2(n5223), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n7822), .ZN(n9524) );
  NOR2_X1 U9401 ( .A1(n9523), .A2(n9524), .ZN(n9522) );
  AOI21_X1 U9402 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9521), .A(n9522), .ZN(
        n9539) );
  NAND2_X1 U9403 ( .A1(n9540), .A2(n9539), .ZN(n9538) );
  OAI21_X1 U9404 ( .B1(n9537), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9538), .ZN(
        n9491) );
  NOR2_X1 U9405 ( .A1(n9492), .A2(n9491), .ZN(n9490) );
  AOI21_X1 U9406 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9489), .A(n9490), .ZN(
        n9621) );
  NAND2_X1 U9407 ( .A1(n9619), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7823) );
  OAI21_X1 U9408 ( .B1(n9619), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7823), .ZN(
        n9622) );
  NOR2_X1 U9409 ( .A1(n9621), .A2(n9622), .ZN(n9620) );
  AOI21_X1 U9410 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9619), .A(n9620), .ZN(
        n9637) );
  NAND2_X1 U9411 ( .A1(n9638), .A2(n9637), .ZN(n9636) );
  OAI21_X1 U9412 ( .B1(n9635), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9636), .ZN(
        n9654) );
  NOR2_X1 U9413 ( .A1(n9655), .A2(n9654), .ZN(n9653) );
  AOI21_X1 U9414 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9652), .A(n9653), .ZN(
        n9671) );
  NAND2_X1 U9415 ( .A1(n9669), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7824) );
  OAI21_X1 U9416 ( .B1(n9669), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7824), .ZN(
        n9672) );
  NOR2_X1 U9417 ( .A1(n9671), .A2(n9672), .ZN(n9670) );
  AOI21_X1 U9418 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9669), .A(n9670), .ZN(
        n7825) );
  NOR2_X1 U9419 ( .A1(n7825), .A2(n7858), .ZN(n7826) );
  XNOR2_X1 U9420 ( .A(n7825), .B(n7858), .ZN(n9685) );
  NOR2_X1 U9421 ( .A1(n7444), .A2(n9685), .ZN(n9684) );
  NOR2_X1 U9422 ( .A1(n7826), .A2(n9684), .ZN(n9694) );
  XNOR2_X1 U9423 ( .A(n7860), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9693) );
  OR2_X1 U9424 ( .A1(n9694), .A2(n9693), .ZN(n9701) );
  NAND2_X1 U9425 ( .A1(n7860), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7827) );
  XNOR2_X1 U9426 ( .A(n9710), .B(n7828), .ZN(n9707) );
  NAND2_X1 U9427 ( .A1(n9706), .A2(n9707), .ZN(n9705) );
  OR2_X1 U9428 ( .A1(n9710), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U9429 ( .A1(n9725), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7831) );
  OR2_X1 U9430 ( .A1(n9725), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7830) );
  AND2_X1 U9431 ( .A1(n7831), .A2(n7830), .ZN(n9719) );
  NAND2_X1 U9432 ( .A1(n9720), .A2(n9719), .ZN(n9718) );
  NAND2_X1 U9433 ( .A1(n9718), .A2(n7831), .ZN(n7832) );
  XNOR2_X1 U9434 ( .A(n7832), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n7867) );
  INV_X1 U9435 ( .A(n7867), .ZN(n7864) );
  NAND2_X1 U9436 ( .A1(n7834), .A2(n7833), .ZN(n9579) );
  NOR2_X2 U9437 ( .A1(n9579), .A2(n7835), .ZN(n9717) );
  INV_X1 U9438 ( .A(n9579), .ZN(n7836) );
  INV_X1 U9439 ( .A(n4358), .ZN(n9025) );
  XNOR2_X1 U9440 ( .A(n9652), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9648) );
  OR2_X1 U9441 ( .A1(n9635), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7856) );
  OR2_X1 U9442 ( .A1(n9489), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U9443 ( .A1(n9489), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U9444 ( .A1(n7838), .A2(n7837), .ZN(n9484) );
  OR2_X1 U9445 ( .A1(n9537), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7854) );
  MUX2_X1 U9446 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7839), .S(n9537), .Z(n9535)
         );
  NAND2_X1 U9447 ( .A1(n9602), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7848) );
  XNOR2_X1 U9448 ( .A(n9037), .B(n7840), .ZN(n9040) );
  XNOR2_X1 U9449 ( .A(n9018), .B(n7841), .ZN(n9017) );
  AND2_X1 U9450 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9016) );
  NAND2_X1 U9451 ( .A1(n9017), .A2(n9016), .ZN(n9015) );
  NAND2_X1 U9452 ( .A1(n9018), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U9453 ( .A1(n9015), .A2(n7842), .ZN(n9039) );
  NAND2_X1 U9454 ( .A1(n9040), .A2(n9039), .ZN(n9038) );
  NAND2_X1 U9455 ( .A1(n9037), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U9456 ( .A1(n9038), .A2(n7843), .ZN(n9055) );
  XNOR2_X1 U9457 ( .A(n9050), .B(n7844), .ZN(n9056) );
  NAND2_X1 U9458 ( .A1(n9055), .A2(n9056), .ZN(n9054) );
  NAND2_X1 U9459 ( .A1(n9050), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U9460 ( .A1(n9054), .A2(n7845), .ZN(n9581) );
  INV_X1 U9461 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9817) );
  MUX2_X1 U9462 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9817), .S(n9587), .Z(n9582)
         );
  NAND2_X1 U9463 ( .A1(n9581), .A2(n9582), .ZN(n9580) );
  NAND2_X1 U9464 ( .A1(n9587), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7846) );
  AND2_X1 U9465 ( .A1(n9580), .A2(n7846), .ZN(n9599) );
  MUX2_X1 U9466 ( .A(n7847), .B(P1_REG1_REG_5__SCAN_IN), .S(n9602), .Z(n9598)
         );
  OR2_X1 U9467 ( .A1(n9599), .A2(n9598), .ZN(n9600) );
  NAND2_X1 U9468 ( .A1(n7848), .A2(n9600), .ZN(n9068) );
  XNOR2_X1 U9469 ( .A(n9063), .B(n7849), .ZN(n9069) );
  NAND2_X1 U9470 ( .A1(n9068), .A2(n9069), .ZN(n9067) );
  NAND2_X1 U9471 ( .A1(n9063), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U9472 ( .A1(n9067), .A2(n7850), .ZN(n9502) );
  INV_X1 U9473 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7851) );
  MUX2_X1 U9474 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7851), .S(n9508), .Z(n9503)
         );
  NAND2_X1 U9475 ( .A1(n9502), .A2(n9503), .ZN(n9501) );
  NAND2_X1 U9476 ( .A1(n9508), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7852) );
  AND2_X1 U9477 ( .A1(n9501), .A2(n7852), .ZN(n9517) );
  INV_X1 U9478 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7853) );
  MUX2_X1 U9479 ( .A(n7853), .B(P1_REG1_REG_8__SCAN_IN), .S(n9521), .Z(n9516)
         );
  NOR2_X1 U9480 ( .A1(n9517), .A2(n9516), .ZN(n9518) );
  AOI21_X1 U9481 ( .B1(n9521), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9518), .ZN(
        n9534) );
  NAND2_X1 U9482 ( .A1(n9535), .A2(n9534), .ZN(n9533) );
  NAND2_X1 U9483 ( .A1(n7854), .A2(n9533), .ZN(n9485) );
  NOR2_X1 U9484 ( .A1(n9484), .A2(n9485), .ZN(n9486) );
  AOI21_X1 U9485 ( .B1(n9489), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9486), .ZN(
        n9614) );
  XNOR2_X1 U9486 ( .A(n9619), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n9615) );
  NOR2_X1 U9487 ( .A1(n9614), .A2(n9615), .ZN(n9616) );
  AOI21_X1 U9488 ( .B1(n9619), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9616), .ZN(
        n9632) );
  MUX2_X1 U9489 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7855), .S(n9635), .Z(n9633)
         );
  NAND2_X1 U9490 ( .A1(n9632), .A2(n9633), .ZN(n9631) );
  NAND2_X1 U9491 ( .A1(n7856), .A2(n9631), .ZN(n9647) );
  NOR2_X1 U9492 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  AOI21_X1 U9493 ( .B1(n9652), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9649), .ZN(
        n9665) );
  XNOR2_X1 U9494 ( .A(n9669), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9664) );
  NOR2_X1 U9495 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  AOI21_X1 U9496 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9669), .A(n9666), .ZN(
        n7857) );
  NOR2_X1 U9497 ( .A1(n7857), .A2(n7858), .ZN(n7859) );
  XNOR2_X1 U9498 ( .A(n7858), .B(n7857), .ZN(n9683) );
  NOR2_X1 U9499 ( .A1(n9682), .A2(n9683), .ZN(n9681) );
  NOR2_X1 U9500 ( .A1(n7859), .A2(n9681), .ZN(n9695) );
  XNOR2_X1 U9501 ( .A(n7860), .B(n7861), .ZN(n9696) );
  INV_X1 U9502 ( .A(n7860), .ZN(n9698) );
  AOI22_X1 U9503 ( .A1(n9695), .A2(n9696), .B1(n9698), .B2(n7861), .ZN(n9709)
         );
  XNOR2_X1 U9504 ( .A(n9710), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9708) );
  OAI22_X1 U9505 ( .A1(n9709), .A2(n9708), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n9710), .ZN(n9723) );
  NAND2_X1 U9506 ( .A1(n9725), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7862) );
  OAI21_X1 U9507 ( .B1(n9725), .B2(P1_REG1_REG_18__SCAN_IN), .A(n7862), .ZN(
        n9722) );
  OR2_X1 U9508 ( .A1(n9723), .A2(n9722), .ZN(n9726) );
  NAND2_X1 U9509 ( .A1(n9726), .A2(n7862), .ZN(n7863) );
  XNOR2_X1 U9510 ( .A(n7863), .B(n9383), .ZN(n7865) );
  AOI22_X1 U9511 ( .A1(n7864), .A2(n9717), .B1(n9712), .B2(n7865), .ZN(n7869)
         );
  NOR2_X2 U9512 ( .A1(n9579), .A2(n4355), .ZN(n9724) );
  NOR2_X1 U9513 ( .A1(n7865), .A2(n9721), .ZN(n7866) );
  AOI211_X1 U9514 ( .C1(n7867), .C2(n9717), .A(n9724), .B(n7866), .ZN(n7868)
         );
  MUX2_X1 U9515 ( .A(n7869), .B(n7868), .S(n7662), .Z(n7870) );
  NAND2_X1 U9516 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8882) );
  OAI211_X1 U9517 ( .C1(n4822), .C2(n9732), .A(n7870), .B(n8882), .ZN(P1_U3262) );
  AOI22_X1 U9518 ( .A1(n8492), .A2(n9934), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9936), .ZN(n7871) );
  OAI21_X1 U9519 ( .B1(n7872), .B2(n8695), .A(n7871), .ZN(n7873) );
  AOI21_X1 U9520 ( .B1(n7875), .B2(n7874), .A(n7873), .ZN(n7876) );
  OAI21_X1 U9521 ( .B1(n7877), .B2(n9936), .A(n7876), .ZN(P2_U3204) );
  INV_X1 U9522 ( .A(n8774), .ZN(n7930) );
  XOR2_X1 U9523 ( .A(n7961), .B(n8130), .Z(n8054) );
  INV_X1 U9524 ( .A(n7878), .ZN(n7880) );
  OAI21_X1 U9525 ( .B1(n8680), .B2(n8054), .A(n8053), .ZN(n7976) );
  XNOR2_X1 U9526 ( .A(n9984), .B(n7961), .ZN(n7883) );
  XNOR2_X1 U9527 ( .A(n7883), .B(n9558), .ZN(n7975) );
  NAND2_X1 U9528 ( .A1(n7976), .A2(n7975), .ZN(n7885) );
  INV_X1 U9529 ( .A(n7883), .ZN(n7884) );
  NAND2_X1 U9530 ( .A1(n7885), .A2(n4930), .ZN(n7931) );
  XNOR2_X1 U9531 ( .A(n9550), .B(n7922), .ZN(n7886) );
  NAND2_X1 U9532 ( .A1(n7886), .A2(n7981), .ZN(n7932) );
  OAI21_X1 U9533 ( .B1(n7886), .B2(n7981), .A(n7932), .ZN(n8037) );
  XNOR2_X1 U9534 ( .A(n8757), .B(n7961), .ZN(n7888) );
  XNOR2_X1 U9535 ( .A(n7888), .B(n9559), .ZN(n7934) );
  INV_X1 U9536 ( .A(n7934), .ZN(n7887) );
  XNOR2_X1 U9537 ( .A(n8837), .B(n7961), .ZN(n7889) );
  XNOR2_X1 U9538 ( .A(n7889), .B(n8669), .ZN(n8084) );
  NOR2_X1 U9539 ( .A1(n7888), .A2(n8659), .ZN(n8085) );
  XNOR2_X1 U9540 ( .A(n8749), .B(n7922), .ZN(n7890) );
  NAND2_X1 U9541 ( .A1(n7890), .A2(n8094), .ZN(n7996) );
  NAND2_X1 U9542 ( .A1(n7997), .A2(n7996), .ZN(n8006) );
  XNOR2_X1 U9543 ( .A(n8826), .B(n7961), .ZN(n7894) );
  XNOR2_X1 U9544 ( .A(n7894), .B(n8626), .ZN(n8008) );
  INV_X1 U9545 ( .A(n8008), .ZN(n7892) );
  INV_X1 U9546 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U9547 ( .A1(n7891), .A2(n8660), .ZN(n8005) );
  AND2_X1 U9548 ( .A1(n7892), .A2(n8005), .ZN(n7893) );
  NAND2_X1 U9549 ( .A1(n8006), .A2(n7893), .ZN(n7897) );
  INV_X1 U9550 ( .A(n7894), .ZN(n7895) );
  NAND2_X1 U9551 ( .A1(n7895), .A2(n8650), .ZN(n7896) );
  NAND2_X1 U9552 ( .A1(n7897), .A2(n7896), .ZN(n8064) );
  XNOR2_X1 U9553 ( .A(n8820), .B(n7961), .ZN(n7898) );
  XNOR2_X1 U9554 ( .A(n7898), .B(n7955), .ZN(n8065) );
  INV_X1 U9555 ( .A(n7898), .ZN(n7899) );
  NAND2_X1 U9556 ( .A1(n7899), .A2(n7955), .ZN(n7900) );
  XNOR2_X1 U9557 ( .A(n8814), .B(n7961), .ZN(n7901) );
  XNOR2_X1 U9558 ( .A(n7901), .B(n8031), .ZN(n7952) );
  XNOR2_X1 U9559 ( .A(n8735), .B(n7961), .ZN(n7902) );
  XNOR2_X1 U9560 ( .A(n7902), .B(n8589), .ZN(n8028) );
  INV_X1 U9561 ( .A(n7902), .ZN(n7903) );
  XNOR2_X1 U9562 ( .A(n8802), .B(n7961), .ZN(n7904) );
  XNOR2_X1 U9563 ( .A(n7904), .B(n8570), .ZN(n7969) );
  NAND2_X1 U9564 ( .A1(n7968), .A2(n7969), .ZN(n7907) );
  INV_X1 U9565 ( .A(n7904), .ZN(n7905) );
  NAND2_X1 U9566 ( .A1(n7905), .A2(n8570), .ZN(n7906) );
  NAND2_X1 U9567 ( .A1(n7907), .A2(n7906), .ZN(n8044) );
  INV_X1 U9568 ( .A(n8044), .ZN(n7908) );
  XNOR2_X1 U9569 ( .A(n8050), .B(n7961), .ZN(n8045) );
  NAND2_X1 U9570 ( .A1(n8045), .A2(n8590), .ZN(n7909) );
  XNOR2_X1 U9571 ( .A(n7910), .B(n7961), .ZN(n7943) );
  INV_X1 U9572 ( .A(n7943), .ZN(n7913) );
  XNOR2_X1 U9573 ( .A(n8789), .B(n7961), .ZN(n7912) );
  NAND2_X1 U9574 ( .A1(n7912), .A2(n7911), .ZN(n7915) );
  OAI21_X1 U9575 ( .B1(n7912), .B2(n7911), .A(n7915), .ZN(n8015) );
  AOI21_X1 U9576 ( .B1(n7913), .B2(n8327), .A(n8015), .ZN(n7914) );
  NAND2_X1 U9577 ( .A1(n8020), .A2(n7915), .ZN(n7988) );
  XNOR2_X1 U9578 ( .A(n8784), .B(n7961), .ZN(n7916) );
  XNOR2_X1 U9579 ( .A(n7916), .B(n8549), .ZN(n7987) );
  NAND2_X1 U9580 ( .A1(n7988), .A2(n7987), .ZN(n7986) );
  INV_X1 U9581 ( .A(n7916), .ZN(n7917) );
  NAND2_X1 U9582 ( .A1(n7917), .A2(n8549), .ZN(n7918) );
  NAND2_X1 U9583 ( .A1(n7986), .A2(n7918), .ZN(n8074) );
  INV_X1 U9584 ( .A(n8074), .ZN(n7919) );
  XNOR2_X1 U9585 ( .A(n8712), .B(n7961), .ZN(n7920) );
  NAND2_X1 U9586 ( .A1(n7919), .A2(n4931), .ZN(n7921) );
  NAND2_X1 U9587 ( .A1(n7920), .A2(n8538), .ZN(n8075) );
  XNOR2_X1 U9588 ( .A(n8774), .B(n7922), .ZN(n7923) );
  NOR2_X1 U9589 ( .A1(n7923), .A2(n8504), .ZN(n7959) );
  AOI21_X1 U9590 ( .B1(n8504), .B2(n7923), .A(n7959), .ZN(n7924) );
  OAI211_X1 U9591 ( .C1(n7925), .C2(n7924), .A(n7960), .B(n8088), .ZN(n7929)
         );
  AOI22_X1 U9592 ( .A1(n8538), .A2(n8091), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7926) );
  OAI21_X1 U9593 ( .B1(n8153), .B2(n8093), .A(n7926), .ZN(n7927) );
  AOI21_X1 U9594 ( .B1(n8520), .B2(n8096), .A(n7927), .ZN(n7928) );
  OAI211_X1 U9595 ( .C1(n7930), .C2(n8099), .A(n7929), .B(n7928), .ZN(P2_U3154) );
  INV_X1 U9596 ( .A(n8757), .ZN(n7942) );
  OR2_X1 U9597 ( .A1(n7931), .A2(n8037), .ZN(n8035) );
  NAND2_X1 U9598 ( .A1(n8035), .A2(n7932), .ZN(n7935) );
  OAI21_X1 U9599 ( .B1(n7935), .B2(n7934), .A(n7933), .ZN(n7936) );
  NAND2_X1 U9600 ( .A1(n7936), .A2(n8088), .ZN(n7941) );
  INV_X1 U9601 ( .A(n7937), .ZN(n8672) );
  INV_X1 U9602 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U9603 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10129), .ZN(n8370) );
  AOI21_X1 U9604 ( .B1(n8066), .B2(n8669), .A(n8370), .ZN(n7938) );
  OAI21_X1 U9605 ( .B1(n8070), .B2(n7981), .A(n7938), .ZN(n7939) );
  AOI21_X1 U9606 ( .B1(n8672), .B2(n8096), .A(n7939), .ZN(n7940) );
  OAI211_X1 U9607 ( .C1(n7942), .C2(n8099), .A(n7941), .B(n7940), .ZN(P2_U3155) );
  NAND2_X1 U9608 ( .A1(n4384), .A2(n7943), .ZN(n8016) );
  OAI21_X1 U9609 ( .B1(n4384), .B2(n7943), .A(n8016), .ZN(n7944) );
  NOR2_X1 U9610 ( .A1(n7944), .A2(n8327), .ZN(n8019) );
  AOI21_X1 U9611 ( .B1(n8327), .B2(n7944), .A(n8019), .ZN(n7950) );
  AOI22_X1 U9612 ( .A1(n8561), .A2(n8066), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        n9827), .ZN(n7946) );
  NAND2_X1 U9613 ( .A1(n8096), .A2(n8564), .ZN(n7945) );
  OAI211_X1 U9614 ( .C1(n7947), .C2(n8070), .A(n7946), .B(n7945), .ZN(n7948)
         );
  AOI21_X1 U9615 ( .B1(n8795), .B2(n8080), .A(n7948), .ZN(n7949) );
  OAI21_X1 U9616 ( .B1(n7950), .B2(n8082), .A(n7949), .ZN(P2_U3156) );
  XOR2_X1 U9617 ( .A(n7952), .B(n7951), .Z(n7958) );
  AOI22_X1 U9618 ( .A1(n8066), .A2(n8589), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n7954) );
  NAND2_X1 U9619 ( .A1(n8096), .A2(n8618), .ZN(n7953) );
  OAI211_X1 U9620 ( .C1(n7955), .C2(n8070), .A(n7954), .B(n7953), .ZN(n7956)
         );
  AOI21_X1 U9621 ( .B1(n8814), .B2(n8080), .A(n7956), .ZN(n7957) );
  OAI21_X1 U9622 ( .B1(n7958), .B2(n8082), .A(n7957), .ZN(P2_U3159) );
  XNOR2_X1 U9623 ( .A(n8501), .B(n7961), .ZN(n7962) );
  AOI22_X1 U9624 ( .A1(n8528), .A2(n8091), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        n9827), .ZN(n7964) );
  NAND2_X1 U9625 ( .A1(n8511), .A2(n8096), .ZN(n7963) );
  OAI211_X1 U9626 ( .C1(n8503), .C2(n8093), .A(n7964), .B(n7963), .ZN(n7965)
         );
  AOI21_X1 U9627 ( .B1(n8512), .B2(n8080), .A(n7965), .ZN(n7966) );
  OAI21_X1 U9628 ( .B1(n7967), .B2(n8082), .A(n7966), .ZN(P2_U3160) );
  XOR2_X1 U9629 ( .A(n7969), .B(n7968), .Z(n7974) );
  AOI22_X1 U9630 ( .A1(n8066), .A2(n8590), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        n9827), .ZN(n7971) );
  NAND2_X1 U9631 ( .A1(n8096), .A2(n8593), .ZN(n7970) );
  OAI211_X1 U9632 ( .C1(n8614), .C2(n8070), .A(n7971), .B(n7970), .ZN(n7972)
         );
  AOI21_X1 U9633 ( .B1(n8802), .B2(n8080), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9634 ( .B1(n7974), .B2(n8082), .A(n7973), .ZN(P2_U3163) );
  XNOR2_X1 U9635 ( .A(n7976), .B(n7975), .ZN(n7985) );
  INV_X1 U9636 ( .A(n7977), .ZN(n8690) );
  NAND2_X1 U9637 ( .A1(n8091), .A2(n8686), .ZN(n7980) );
  INV_X1 U9638 ( .A(n7978), .ZN(n7979) );
  OAI211_X1 U9639 ( .C1(n7981), .C2(n8093), .A(n7980), .B(n7979), .ZN(n7983)
         );
  INV_X1 U9640 ( .A(n9984), .ZN(n8696) );
  NOR2_X1 U9641 ( .A1(n8696), .A2(n8099), .ZN(n7982) );
  AOI211_X1 U9642 ( .C1(n8690), .C2(n8096), .A(n7983), .B(n7982), .ZN(n7984)
         );
  OAI21_X1 U9643 ( .B1(n7985), .B2(n8082), .A(n7984), .ZN(P2_U3164) );
  INV_X1 U9644 ( .A(n8784), .ZN(n7995) );
  OAI21_X1 U9645 ( .B1(n7988), .B2(n7987), .A(n7986), .ZN(n7989) );
  NAND2_X1 U9646 ( .A1(n7989), .A2(n8088), .ZN(n7994) );
  AOI22_X1 U9647 ( .A1(n8561), .A2(n8091), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        n9827), .ZN(n7990) );
  OAI21_X1 U9648 ( .B1(n7991), .B2(n8093), .A(n7990), .ZN(n7992) );
  AOI21_X1 U9649 ( .B1(n8540), .B2(n8096), .A(n7992), .ZN(n7993) );
  OAI211_X1 U9650 ( .C1(n7995), .C2(n8099), .A(n7994), .B(n7993), .ZN(P2_U3165) );
  NAND2_X1 U9651 ( .A1(n8005), .A2(n7996), .ZN(n7998) );
  XOR2_X1 U9652 ( .A(n7998), .B(n7997), .Z(n8004) );
  NAND2_X1 U9653 ( .A1(n8091), .A2(n8669), .ZN(n7999) );
  NAND2_X1 U9654 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8418) );
  OAI211_X1 U9655 ( .C1(n8650), .C2(n8093), .A(n7999), .B(n8418), .ZN(n8000)
         );
  AOI21_X1 U9656 ( .B1(n8001), .B2(n8096), .A(n8000), .ZN(n8003) );
  NAND2_X1 U9657 ( .A1(n8749), .A2(n8080), .ZN(n8002) );
  OAI211_X1 U9658 ( .C1(n8004), .C2(n8082), .A(n8003), .B(n8002), .ZN(P2_U3166) );
  NAND2_X1 U9659 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  XOR2_X1 U9660 ( .A(n8008), .B(n8007), .Z(n8014) );
  AOI22_X1 U9661 ( .A1(n8066), .A2(n8636), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8011) );
  INV_X1 U9662 ( .A(n8009), .ZN(n8639) );
  NAND2_X1 U9663 ( .A1(n8096), .A2(n8639), .ZN(n8010) );
  OAI211_X1 U9664 ( .C1(n8094), .C2(n8070), .A(n8011), .B(n8010), .ZN(n8012)
         );
  AOI21_X1 U9665 ( .B1(n8826), .B2(n8080), .A(n8012), .ZN(n8013) );
  OAI21_X1 U9666 ( .B1(n8014), .B2(n8082), .A(n8013), .ZN(P2_U3168) );
  INV_X1 U9667 ( .A(n8015), .ZN(n8018) );
  INV_X1 U9668 ( .A(n8016), .ZN(n8017) );
  NOR3_X1 U9669 ( .A1(n8019), .A2(n8018), .A3(n8017), .ZN(n8022) );
  INV_X1 U9670 ( .A(n8020), .ZN(n8021) );
  OAI21_X1 U9671 ( .B1(n8022), .B2(n8021), .A(n8088), .ZN(n8026) );
  AOI22_X1 U9672 ( .A1(n8326), .A2(n8066), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        n9827), .ZN(n8023) );
  OAI21_X1 U9673 ( .B1(n8571), .B2(n8070), .A(n8023), .ZN(n8024) );
  AOI21_X1 U9674 ( .B1(n8551), .B2(n8096), .A(n8024), .ZN(n8025) );
  OAI211_X1 U9675 ( .C1(n8789), .C2(n8099), .A(n8026), .B(n8025), .ZN(P2_U3169) );
  XOR2_X1 U9676 ( .A(n8028), .B(n8027), .Z(n8034) );
  AOI22_X1 U9677 ( .A1(n8066), .A2(n8602), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8030) );
  NAND2_X1 U9678 ( .A1(n8096), .A2(n8606), .ZN(n8029) );
  OAI211_X1 U9679 ( .C1(n8031), .C2(n8070), .A(n8030), .B(n8029), .ZN(n8032)
         );
  AOI21_X1 U9680 ( .B1(n8735), .B2(n8080), .A(n8032), .ZN(n8033) );
  OAI21_X1 U9681 ( .B1(n8034), .B2(n8082), .A(n8033), .ZN(P2_U3173) );
  INV_X1 U9682 ( .A(n8035), .ZN(n8036) );
  AOI21_X1 U9683 ( .B1(n7931), .B2(n8037), .A(n8036), .ZN(n8043) );
  NOR2_X1 U9684 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6121), .ZN(n8350) );
  NOR2_X1 U9685 ( .A1(n8093), .A2(n9559), .ZN(n8038) );
  AOI211_X1 U9686 ( .C1(n8091), .C2(n8328), .A(n8350), .B(n8038), .ZN(n8039)
         );
  OAI21_X1 U9687 ( .B1(n9554), .B2(n8040), .A(n8039), .ZN(n8041) );
  AOI21_X1 U9688 ( .B1(n9550), .B2(n8080), .A(n8041), .ZN(n8042) );
  OAI21_X1 U9689 ( .B1(n8043), .B2(n8082), .A(n8042), .ZN(P2_U3174) );
  XNOR2_X1 U9690 ( .A(n8045), .B(n8590), .ZN(n8046) );
  XNOR2_X1 U9691 ( .A(n8044), .B(n8046), .ZN(n8052) );
  AOI22_X1 U9692 ( .A1(n8091), .A2(n8602), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8048) );
  NAND2_X1 U9693 ( .A1(n8096), .A2(n8578), .ZN(n8047) );
  OAI211_X1 U9694 ( .C1(n8571), .C2(n8093), .A(n8048), .B(n8047), .ZN(n8049)
         );
  AOI21_X1 U9695 ( .B1(n8050), .B2(n8080), .A(n8049), .ZN(n8051) );
  OAI21_X1 U9696 ( .B1(n8052), .B2(n8082), .A(n8051), .ZN(P2_U3175) );
  OAI211_X1 U9697 ( .C1(n4454), .C2(n8054), .A(n8053), .B(n8088), .ZN(n8063)
         );
  INV_X1 U9698 ( .A(n8055), .ZN(n8061) );
  INV_X1 U9699 ( .A(n9978), .ZN(n8056) );
  NOR2_X1 U9700 ( .A1(n8056), .A2(n8099), .ZN(n8060) );
  NAND2_X1 U9701 ( .A1(n8091), .A2(n8329), .ZN(n8058) );
  OAI211_X1 U9702 ( .C1(n9558), .C2(n8093), .A(n8058), .B(n8057), .ZN(n8059)
         );
  AOI211_X1 U9703 ( .C1(n8061), .C2(n8096), .A(n8060), .B(n8059), .ZN(n8062)
         );
  NAND2_X1 U9704 ( .A1(n8063), .A2(n8062), .ZN(P2_U3176) );
  XOR2_X1 U9705 ( .A(n8064), .B(n8065), .Z(n8073) );
  AND2_X1 U9706 ( .A1(n9827), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8458) );
  AOI21_X1 U9707 ( .B1(n8066), .B2(n8627), .A(n8458), .ZN(n8069) );
  INV_X1 U9708 ( .A(n8067), .ZN(n8630) );
  NAND2_X1 U9709 ( .A1(n8096), .A2(n8630), .ZN(n8068) );
  OAI211_X1 U9710 ( .C1(n8070), .C2(n8650), .A(n8069), .B(n8068), .ZN(n8071)
         );
  AOI21_X1 U9711 ( .B1(n8820), .B2(n8080), .A(n8071), .ZN(n8072) );
  OAI21_X1 U9712 ( .B1(n8073), .B2(n8082), .A(n8072), .ZN(P2_U3178) );
  NAND2_X1 U9713 ( .A1(n4931), .A2(n8075), .ZN(n8076) );
  XNOR2_X1 U9714 ( .A(n8074), .B(n8076), .ZN(n8083) );
  AOI22_X1 U9715 ( .A1(n8326), .A2(n8091), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        n9827), .ZN(n8078) );
  NAND2_X1 U9716 ( .A1(n8529), .A2(n8096), .ZN(n8077) );
  OAI211_X1 U9717 ( .C1(n8504), .C2(n8093), .A(n8078), .B(n8077), .ZN(n8079)
         );
  AOI21_X1 U9718 ( .B1(n8712), .B2(n8080), .A(n8079), .ZN(n8081) );
  OAI21_X1 U9719 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(P2_U3180) );
  INV_X1 U9720 ( .A(n8837), .ZN(n8100) );
  INV_X1 U9721 ( .A(n7933), .ZN(n8086) );
  OAI21_X1 U9722 ( .B1(n8086), .B2(n8085), .A(n8084), .ZN(n8089) );
  NAND3_X1 U9723 ( .A1(n8089), .A2(n8088), .A3(n8087), .ZN(n8098) );
  INV_X1 U9724 ( .A(n8090), .ZN(n8663) );
  INV_X1 U9725 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U9726 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10125), .ZN(n8401) );
  AOI21_X1 U9727 ( .B1(n8091), .B2(n8659), .A(n8401), .ZN(n8092) );
  OAI21_X1 U9728 ( .B1(n8094), .B2(n8093), .A(n8092), .ZN(n8095) );
  AOI21_X1 U9729 ( .B1(n8663), .B2(n8096), .A(n8095), .ZN(n8097) );
  OAI211_X1 U9730 ( .C1(n8100), .C2(n8099), .A(n8098), .B(n8097), .ZN(P2_U3181) );
  NAND2_X1 U9731 ( .A1(n8101), .A2(n8115), .ZN(n8104) );
  OR2_X1 U9732 ( .A1(n4353), .A2(n8102), .ZN(n8103) );
  NAND2_X1 U9733 ( .A1(n8104), .A2(n8103), .ZN(n8703) );
  INV_X1 U9734 ( .A(n8324), .ZN(n8117) );
  NAND2_X1 U9735 ( .A1(n8703), .A2(n8117), .ZN(n8300) );
  NAND2_X1 U9736 ( .A1(n8300), .A2(n8105), .ZN(n8302) );
  AOI21_X1 U9737 ( .B1(n8106), .B2(n8293), .A(n8302), .ZN(n8116) );
  INV_X1 U9738 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U9739 ( .A1(n6270), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8109) );
  INV_X1 U9740 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8107) );
  OR2_X1 U9741 ( .A1(n5989), .A2(n8107), .ZN(n8108) );
  OAI211_X1 U9742 ( .C1(n8110), .C2(n6308), .A(n8109), .B(n8108), .ZN(n8111)
         );
  INV_X1 U9743 ( .A(n8111), .ZN(n8112) );
  INV_X1 U9744 ( .A(n8703), .ZN(n8766) );
  NOR2_X1 U9745 ( .A1(n4353), .A2(n6500), .ZN(n8114) );
  NAND2_X1 U9746 ( .A1(n8763), .A2(n8494), .ZN(n8151) );
  AND2_X1 U9747 ( .A1(n8298), .A2(n8293), .ZN(n8311) );
  INV_X1 U9748 ( .A(n8247), .ZN(n8119) );
  NOR2_X1 U9749 ( .A1(n6673), .A2(n8310), .ZN(n8120) );
  AND4_X1 U9750 ( .A1(n6318), .A2(n8172), .A3(n9917), .A4(n8120), .ZN(n8126)
         );
  NOR2_X1 U9751 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  NAND4_X1 U9752 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n8128)
         );
  NOR4_X1 U9753 ( .A1(n8128), .A2(n8193), .A3(n8127), .A4(n6063), .ZN(n8131)
         );
  NAND4_X1 U9754 ( .A1(n8131), .A2(n8691), .A3(n8130), .A4(n8129), .ZN(n8134)
         );
  NAND2_X1 U9755 ( .A1(n8133), .A2(n8132), .ZN(n8221) );
  INV_X1 U9756 ( .A(n8221), .ZN(n9555) );
  NOR2_X1 U9757 ( .A1(n8134), .A2(n9555), .ZN(n8135) );
  INV_X1 U9758 ( .A(n8226), .ZN(n8676) );
  NAND4_X1 U9759 ( .A1(n8646), .A2(n8135), .A3(n8676), .A4(n4559), .ZN(n8136)
         );
  NOR3_X1 U9760 ( .A1(n8625), .A2(n8635), .A3(n8136), .ZN(n8137) );
  NAND3_X1 U9761 ( .A1(n8597), .A2(n8610), .A3(n8137), .ZN(n8138) );
  NOR2_X1 U9762 ( .A1(n8584), .A2(n8138), .ZN(n8139) );
  NAND2_X1 U9763 ( .A1(n8575), .A2(n8139), .ZN(n8142) );
  NAND2_X1 U9764 ( .A1(n8274), .A2(n8140), .ZN(n8555) );
  INV_X1 U9765 ( .A(n8552), .ZN(n8141) );
  OR4_X1 U9766 ( .A1(n8142), .A2(n8543), .A3(n8555), .A4(n8560), .ZN(n8146) );
  INV_X1 U9767 ( .A(n8143), .ZN(n8144) );
  INV_X1 U9768 ( .A(n8525), .ZN(n8524) );
  NAND2_X1 U9769 ( .A1(n8287), .A2(n8288), .ZN(n8515) );
  OR3_X1 U9770 ( .A1(n8146), .A2(n8524), .A3(n8515), .ZN(n8147) );
  NOR2_X1 U9771 ( .A1(n8501), .A2(n8147), .ZN(n8149) );
  INV_X1 U9772 ( .A(n8302), .ZN(n8148) );
  NAND4_X1 U9773 ( .A1(n8151), .A2(n8311), .A3(n8149), .A4(n8148), .ZN(n8150)
         );
  OAI21_X1 U9774 ( .B1(n8299), .B2(n8151), .A(n8150), .ZN(n8152) );
  INV_X1 U9775 ( .A(n8512), .ZN(n8768) );
  MUX2_X1 U9776 ( .A(n8153), .B(n8768), .S(n8297), .Z(n8305) );
  NAND2_X1 U9777 ( .A1(n8181), .A2(n8154), .ZN(n8157) );
  NAND2_X1 U9778 ( .A1(n8174), .A2(n8155), .ZN(n8156) );
  MUX2_X1 U9779 ( .A(n8157), .B(n8156), .S(n8290), .Z(n8158) );
  INV_X1 U9780 ( .A(n8158), .ZN(n8171) );
  NAND3_X1 U9781 ( .A1(n8159), .A2(n8169), .A3(n6674), .ZN(n8163) );
  NAND2_X1 U9782 ( .A1(n8169), .A2(n8160), .ZN(n8162) );
  NAND4_X1 U9783 ( .A1(n8163), .A2(n8162), .A3(n8297), .A4(n8161), .ZN(n8167)
         );
  NAND2_X1 U9784 ( .A1(n8164), .A2(n8161), .ZN(n8165) );
  NAND2_X1 U9785 ( .A1(n8165), .A2(n8290), .ZN(n8166) );
  NAND2_X1 U9786 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  OAI211_X1 U9787 ( .C1(n8169), .C2(n8297), .A(n8168), .B(n9917), .ZN(n8170)
         );
  NAND2_X1 U9788 ( .A1(n8171), .A2(n8170), .ZN(n8173) );
  NAND2_X1 U9789 ( .A1(n8173), .A2(n8172), .ZN(n8185) );
  INV_X1 U9790 ( .A(n8174), .ZN(n8177) );
  OAI211_X1 U9791 ( .C1(n8185), .C2(n8177), .A(n8176), .B(n8175), .ZN(n8178)
         );
  NAND3_X1 U9792 ( .A1(n8178), .A2(n8182), .A3(n8188), .ZN(n8180) );
  NAND2_X1 U9793 ( .A1(n8180), .A2(n8179), .ZN(n8191) );
  INV_X1 U9794 ( .A(n8181), .ZN(n8184) );
  OAI211_X1 U9795 ( .C1(n8185), .C2(n8184), .A(n8183), .B(n8182), .ZN(n8187)
         );
  NAND2_X1 U9796 ( .A1(n8187), .A2(n8186), .ZN(n8189) );
  NAND2_X1 U9797 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  NAND3_X1 U9798 ( .A1(n8195), .A2(n8194), .A3(n8290), .ZN(n8198) );
  NAND3_X1 U9799 ( .A1(n8200), .A2(n8297), .A3(n8199), .ZN(n8196) );
  NAND2_X1 U9800 ( .A1(n8198), .A2(n8196), .ZN(n8197) );
  INV_X1 U9801 ( .A(n8198), .ZN(n8204) );
  OAI21_X1 U9802 ( .B1(n9957), .B2(n8332), .A(n8199), .ZN(n8203) );
  NAND2_X1 U9803 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  AOI21_X1 U9804 ( .B1(n8204), .B2(n8203), .A(n8202), .ZN(n8205) );
  MUX2_X1 U9805 ( .A(n8206), .B(n8205), .S(n8290), .Z(n8207) );
  INV_X1 U9806 ( .A(n8211), .ZN(n8208) );
  AOI21_X1 U9807 ( .B1(n8215), .B2(n8209), .A(n8208), .ZN(n8217) );
  AND2_X1 U9808 ( .A1(n8211), .A2(n8210), .ZN(n8214) );
  INV_X1 U9809 ( .A(n8212), .ZN(n8213) );
  AOI21_X1 U9810 ( .B1(n8215), .B2(n8214), .A(n8213), .ZN(n8216) );
  MUX2_X1 U9811 ( .A(n8217), .B(n8216), .S(n8290), .Z(n8223) );
  MUX2_X1 U9812 ( .A(n8219), .B(n8218), .S(n8290), .Z(n8220) );
  MUX2_X1 U9813 ( .A(n8225), .B(n8224), .S(n8297), .Z(n8227) );
  AND2_X1 U9814 ( .A1(n8757), .A2(n8297), .ZN(n8229) );
  NOR2_X1 U9815 ( .A1(n8757), .A2(n8297), .ZN(n8228) );
  MUX2_X1 U9816 ( .A(n8229), .B(n8228), .S(n8659), .Z(n8230) );
  MUX2_X1 U9817 ( .A(n8232), .B(n8231), .S(n8290), .Z(n8233) );
  AND2_X1 U9818 ( .A1(n8646), .A2(n8233), .ZN(n8234) );
  MUX2_X1 U9819 ( .A(n8236), .B(n8235), .S(n8290), .Z(n8237) );
  INV_X1 U9820 ( .A(n8237), .ZN(n8238) );
  NOR2_X1 U9821 ( .A1(n8635), .A2(n8238), .ZN(n8239) );
  NAND2_X1 U9822 ( .A1(n8240), .A2(n8239), .ZN(n8246) );
  NAND3_X1 U9823 ( .A1(n8246), .A2(n8247), .A3(n8241), .ZN(n8243) );
  INV_X1 U9824 ( .A(n8242), .ZN(n8244) );
  NAND3_X1 U9825 ( .A1(n8243), .A2(n8244), .A3(n8251), .ZN(n8250) );
  NAND3_X1 U9826 ( .A1(n8246), .A2(n8245), .A3(n8244), .ZN(n8248) );
  NAND2_X1 U9827 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  AND2_X1 U9828 ( .A1(n8253), .A2(n8256), .ZN(n8255) );
  INV_X1 U9829 ( .A(n8259), .ZN(n8254) );
  NAND3_X1 U9830 ( .A1(n8257), .A2(n4869), .A3(n8256), .ZN(n8262) );
  AND2_X1 U9831 ( .A1(n8259), .A2(n8258), .ZN(n8261) );
  AOI21_X1 U9832 ( .B1(n8262), .B2(n8261), .A(n8260), .ZN(n8263) );
  INV_X1 U9833 ( .A(n8575), .ZN(n8269) );
  NAND3_X1 U9834 ( .A1(n8272), .A2(n8290), .A3(n8264), .ZN(n8267) );
  NAND2_X1 U9835 ( .A1(n8265), .A2(n8297), .ZN(n8266) );
  NAND2_X1 U9836 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  OAI21_X1 U9837 ( .B1(n8270), .B2(n8269), .A(n8268), .ZN(n8278) );
  NAND2_X1 U9838 ( .A1(n8272), .A2(n8271), .ZN(n8275) );
  OAI211_X1 U9839 ( .C1(n8290), .C2(n8272), .A(n8275), .B(n8274), .ZN(n8273)
         );
  INV_X1 U9840 ( .A(n8273), .ZN(n8277) );
  AOI21_X1 U9841 ( .B1(n8275), .B2(n8274), .A(n8290), .ZN(n8276) );
  MUX2_X1 U9842 ( .A(n8280), .B(n8279), .S(n8297), .Z(n8281) );
  INV_X1 U9843 ( .A(n8282), .ZN(n8284) );
  MUX2_X1 U9844 ( .A(n8284), .B(n8283), .S(n8290), .Z(n8285) );
  NOR2_X1 U9845 ( .A1(n8515), .A2(n8285), .ZN(n8286) );
  MUX2_X1 U9846 ( .A(n8288), .B(n8287), .S(n8297), .Z(n8289) );
  OR2_X1 U9847 ( .A1(n8503), .A2(n8297), .ZN(n8294) );
  AND2_X1 U9848 ( .A1(n8295), .A2(n8294), .ZN(n8304) );
  INV_X1 U9849 ( .A(n8314), .ZN(n8296) );
  NOR2_X1 U9850 ( .A1(n8296), .A2(n8517), .ZN(n8303) );
  NAND2_X1 U9851 ( .A1(n8298), .A2(n8297), .ZN(n8301) );
  AOI21_X1 U9852 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8307) );
  NAND4_X1 U9853 ( .A1(n8311), .A2(n8319), .A3(n6673), .A4(n8310), .ZN(n8312)
         );
  XNOR2_X1 U9854 ( .A(n8316), .B(n8482), .ZN(n8323) );
  NOR3_X1 U9855 ( .A1(n8318), .A2(n8317), .A3(n6302), .ZN(n8321) );
  OAI21_X1 U9856 ( .B1(n8322), .B2(n8319), .A(P2_B_REG_SCAN_IN), .ZN(n8320) );
  OAI22_X1 U9857 ( .A1(n8323), .A2(n8322), .B1(n8321), .B2(n8320), .ZN(
        P2_U3296) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8494), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8324), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U9860 ( .A(n8503), .ZN(n8325) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8325), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9862 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8517), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9863 ( .A(n8528), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8456), .Z(
        P2_U3518) );
  MUX2_X1 U9864 ( .A(n8538), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8456), .Z(
        P2_U3517) );
  MUX2_X1 U9865 ( .A(n8326), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8456), .Z(
        P2_U3516) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8561), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8327), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9868 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8590), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9869 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8602), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9870 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8589), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9871 ( .A(n8627), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8456), .Z(
        P2_U3510) );
  MUX2_X1 U9872 ( .A(n8636), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8456), .Z(
        P2_U3509) );
  MUX2_X1 U9873 ( .A(n8626), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8456), .Z(
        P2_U3508) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8660), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9875 ( .A(n8669), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8456), .Z(
        P2_U3506) );
  MUX2_X1 U9876 ( .A(n8659), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8456), .Z(
        P2_U3505) );
  MUX2_X1 U9877 ( .A(n8685), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8456), .Z(
        P2_U3504) );
  MUX2_X1 U9878 ( .A(n8328), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8456), .Z(
        P2_U3503) );
  MUX2_X1 U9879 ( .A(n8686), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8456), .Z(
        P2_U3502) );
  MUX2_X1 U9880 ( .A(n8329), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8456), .Z(
        P2_U3501) );
  MUX2_X1 U9881 ( .A(n8330), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8456), .Z(
        P2_U3500) );
  MUX2_X1 U9882 ( .A(n8331), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8456), .Z(
        P2_U3499) );
  MUX2_X1 U9883 ( .A(n8332), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8456), .Z(
        P2_U3498) );
  MUX2_X1 U9884 ( .A(n8333), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8456), .Z(
        P2_U3497) );
  MUX2_X1 U9885 ( .A(n8334), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8456), .Z(
        P2_U3496) );
  MUX2_X1 U9886 ( .A(n8335), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8456), .Z(
        P2_U3495) );
  MUX2_X1 U9887 ( .A(n8336), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8456), .Z(
        P2_U3494) );
  MUX2_X1 U9888 ( .A(n4354), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8456), .Z(
        P2_U3493) );
  MUX2_X1 U9889 ( .A(n6609), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8456), .Z(
        P2_U3492) );
  AOI21_X1 U9890 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8341) );
  MUX2_X1 U9891 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8473), .Z(n8365) );
  XNOR2_X1 U9892 ( .A(n8365), .B(n8376), .ZN(n8340) );
  NAND2_X1 U9893 ( .A1(n8341), .A2(n8340), .ZN(n8366) );
  OAI21_X1 U9894 ( .B1(n8341), .B2(n8340), .A(n8366), .ZN(n8356) );
  XNOR2_X1 U9895 ( .A(n8374), .B(n8364), .ZN(n8344) );
  INV_X1 U9896 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9568) );
  NOR2_X1 U9897 ( .A1(n9568), .A2(n8344), .ZN(n8377) );
  AOI21_X1 U9898 ( .B1(n8344), .B2(n9568), .A(n8377), .ZN(n8345) );
  NOR2_X1 U9899 ( .A1(n8345), .A2(n9909), .ZN(n8355) );
  INV_X1 U9900 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8353) );
  INV_X1 U9901 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9564) );
  NOR2_X1 U9902 ( .A1(n9564), .A2(n8348), .ZN(n8360) );
  AOI21_X1 U9903 ( .B1(n9564), .B2(n8348), .A(n8360), .ZN(n8349) );
  OR2_X1 U9904 ( .A1(n8349), .A2(n9905), .ZN(n8352) );
  AOI21_X1 U9905 ( .B1(n9896), .B2(n8376), .A(n8350), .ZN(n8351) );
  OAI211_X1 U9906 ( .C1(n8353), .C2(n9841), .A(n8352), .B(n8351), .ZN(n8354)
         );
  AOI211_X1 U9907 ( .C1(n8356), .C2(n6411), .A(n8355), .B(n8354), .ZN(n8357)
         );
  INV_X1 U9908 ( .A(n8357), .ZN(P2_U3195) );
  NOR2_X1 U9909 ( .A1(n8376), .A2(n8359), .ZN(n8361) );
  AOI22_X1 U9910 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8380), .B1(n8397), .B2(
        n6135), .ZN(n8362) );
  AOI21_X1 U9911 ( .B1(n8363), .B2(n8362), .A(n8389), .ZN(n8388) );
  MUX2_X1 U9912 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8473), .Z(n8391) );
  XNOR2_X1 U9913 ( .A(n8391), .B(n8380), .ZN(n8369) );
  OR2_X1 U9914 ( .A1(n8365), .A2(n8364), .ZN(n8367) );
  NAND2_X1 U9915 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND2_X1 U9916 ( .A1(n8369), .A2(n8368), .ZN(n8392) );
  OAI21_X1 U9917 ( .B1(n8369), .B2(n8368), .A(n8392), .ZN(n8386) );
  INV_X1 U9918 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U9919 ( .A1(n9896), .A2(n8380), .ZN(n8372) );
  INV_X1 U9920 ( .A(n8370), .ZN(n8371) );
  OAI211_X1 U9921 ( .C1(n8373), .C2(n9841), .A(n8372), .B(n8371), .ZN(n8385)
         );
  INV_X1 U9922 ( .A(n8374), .ZN(n8375) );
  NOR2_X1 U9923 ( .A1(n8376), .A2(n8375), .ZN(n8378) );
  XNOR2_X1 U9924 ( .A(n8380), .B(n8379), .ZN(n8381) );
  NOR2_X1 U9925 ( .A1(n8382), .A2(n8381), .ZN(n8396) );
  AOI21_X1 U9926 ( .B1(n8382), .B2(n8381), .A(n8396), .ZN(n8383) );
  NOR2_X1 U9927 ( .A1(n8383), .A2(n9909), .ZN(n8384) );
  AOI211_X1 U9928 ( .C1(n6411), .C2(n8386), .A(n8385), .B(n8384), .ZN(n8387)
         );
  OAI21_X1 U9929 ( .B1(n8388), .B2(n9905), .A(n8387), .ZN(P2_U3196) );
  AOI21_X1 U9930 ( .B1(n8662), .B2(n8390), .A(n8408), .ZN(n8407) );
  MUX2_X1 U9931 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8473), .Z(n8413) );
  XNOR2_X1 U9932 ( .A(n8413), .B(n8421), .ZN(n8395) );
  OR2_X1 U9933 ( .A1(n8391), .A2(n8397), .ZN(n8393) );
  NAND2_X1 U9934 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  NAND2_X1 U9935 ( .A1(n8395), .A2(n8394), .ZN(n8414) );
  OAI21_X1 U9936 ( .B1(n8395), .B2(n8394), .A(n8414), .ZN(n8405) );
  AOI21_X1 U9937 ( .B1(n8398), .B2(n8752), .A(n8422), .ZN(n8403) );
  INV_X1 U9938 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8399) );
  NOR2_X1 U9939 ( .A1(n9841), .A2(n8399), .ZN(n8400) );
  AOI211_X1 U9940 ( .C1(n8421), .C2(n9896), .A(n8401), .B(n8400), .ZN(n8402)
         );
  OAI21_X1 U9941 ( .B1(n8403), .B2(n9909), .A(n8402), .ZN(n8404) );
  AOI21_X1 U9942 ( .B1(n6411), .B2(n8405), .A(n8404), .ZN(n8406) );
  OAI21_X1 U9943 ( .B1(n8407), .B2(n9905), .A(n8406), .ZN(P2_U3197) );
  NOR2_X1 U9944 ( .A1(n8421), .A2(n4432), .ZN(n8409) );
  AOI22_X1 U9945 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8424), .B1(n8437), .B2(
        n8652), .ZN(n8410) );
  AOI21_X1 U9946 ( .B1(n8411), .B2(n8410), .A(n8432), .ZN(n8431) );
  MUX2_X1 U9947 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8473), .Z(n8435) );
  XNOR2_X1 U9948 ( .A(n8435), .B(n8424), .ZN(n8417) );
  OR2_X1 U9949 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  OAI21_X1 U9950 ( .B1(n8417), .B2(n8416), .A(n8434), .ZN(n8429) );
  INV_X1 U9951 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10011) );
  OR2_X1 U9952 ( .A1(n9871), .A2(n8437), .ZN(n8419) );
  OAI211_X1 U9953 ( .C1(n10011), .C2(n9841), .A(n8419), .B(n8418), .ZN(n8428)
         );
  NOR2_X1 U9954 ( .A1(n8421), .A2(n8420), .ZN(n8423) );
  XNOR2_X1 U9955 ( .A(n8424), .B(n8750), .ZN(n8425) );
  AOI21_X1 U9956 ( .B1(n4402), .B2(n8425), .A(n8436), .ZN(n8426) );
  NOR2_X1 U9957 ( .A1(n8426), .A2(n9909), .ZN(n8427) );
  AOI211_X1 U9958 ( .C1(n6411), .C2(n8429), .A(n8428), .B(n8427), .ZN(n8430)
         );
  OAI21_X1 U9959 ( .B1(n8431), .B2(n9905), .A(n8430), .ZN(P2_U3198) );
  AOI21_X1 U9960 ( .B1(n8638), .B2(n8433), .A(n8446), .ZN(n8444) );
  MUX2_X1 U9961 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8473), .Z(n8449) );
  XNOR2_X1 U9962 ( .A(n8449), .B(n8460), .ZN(n8452) );
  XNOR2_X1 U9963 ( .A(n8452), .B(n8451), .ZN(n8442) );
  INV_X1 U9964 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8439) );
  XNOR2_X1 U9965 ( .A(n8460), .B(n8459), .ZN(n8438) );
  OAI22_X1 U9966 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6173), .B1(n9871), .B2(
        n8440), .ZN(n8441) );
  OAI21_X1 U9967 ( .B1(n8444), .B2(n9905), .A(n8443), .ZN(P2_U3199) );
  NOR2_X1 U9968 ( .A1(n8460), .A2(n8445), .ZN(n8447) );
  NAND2_X1 U9969 ( .A1(n8462), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8468) );
  OAI21_X1 U9970 ( .B1(n8462), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8468), .ZN(
        n8448) );
  AOI21_X1 U9971 ( .B1(n4397), .B2(n8448), .A(n8470), .ZN(n8467) );
  INV_X1 U9972 ( .A(n9841), .ZN(n9900) );
  INV_X1 U9973 ( .A(n8449), .ZN(n8450) );
  MUX2_X1 U9974 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8473), .Z(n8453) );
  NOR2_X1 U9975 ( .A1(n8454), .A2(n8453), .ZN(n8477) );
  NAND2_X1 U9976 ( .A1(n8454), .A2(n8453), .ZN(n8475) );
  INV_X1 U9977 ( .A(n8475), .ZN(n8455) );
  NOR2_X1 U9978 ( .A1(n8477), .A2(n8455), .ZN(n8457) );
  NOR2_X1 U9979 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  NAND2_X1 U9980 ( .A1(n8462), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8484) );
  OAI21_X1 U9981 ( .B1(n8462), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8484), .ZN(
        n8463) );
  AOI21_X1 U9982 ( .B1(n4440), .B2(n8463), .A(n8485), .ZN(n8464) );
  OR2_X1 U9983 ( .A1(n8464), .A2(n9909), .ZN(n8465) );
  OAI211_X1 U9984 ( .C1(n8467), .C2(n9905), .A(n8466), .B(n8465), .ZN(P2_U3200) );
  INV_X1 U9985 ( .A(n8468), .ZN(n8469) );
  NOR2_X1 U9986 ( .A1(n8470), .A2(n8469), .ZN(n8471) );
  MUX2_X1 U9987 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8617), .S(n8482), .Z(n8474)
         );
  XNOR2_X1 U9988 ( .A(n8472), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8486) );
  MUX2_X1 U9989 ( .A(n8474), .B(n8486), .S(n8473), .Z(n8479) );
  OAI21_X1 U9990 ( .B1(n8477), .B2(n8476), .A(n8475), .ZN(n8478) );
  NAND2_X1 U9991 ( .A1(n9900), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U9992 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(n9827), .ZN(n8480) );
  OAI211_X1 U9993 ( .C1(n9871), .C2(n8482), .A(n8481), .B(n8480), .ZN(n8483)
         );
  INV_X1 U9994 ( .A(n8483), .ZN(n8491) );
  INV_X1 U9995 ( .A(n8486), .ZN(n8487) );
  XNOR2_X1 U9996 ( .A(n8488), .B(n8487), .ZN(n8490) );
  NAND2_X1 U9997 ( .A1(n8492), .A2(n9934), .ZN(n8495) );
  NAND2_X1 U9998 ( .A1(n8494), .A2(n8493), .ZN(n8761) );
  AOI21_X1 U9999 ( .B1(n8495), .B2(n8761), .A(n9936), .ZN(n8497) );
  AOI21_X1 U10000 ( .B1(n9936), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8497), .ZN(
        n8496) );
  OAI21_X1 U10001 ( .B1(n8763), .B2(n8695), .A(n8496), .ZN(P2_U3202) );
  AOI21_X1 U10002 ( .B1(n9936), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8497), .ZN(
        n8498) );
  OAI21_X1 U10003 ( .B1(n8766), .B2(n8695), .A(n8498), .ZN(P2_U3203) );
  XNOR2_X1 U10004 ( .A(n8499), .B(n8500), .ZN(n8769) );
  XNOR2_X1 U10005 ( .A(n8502), .B(n8501), .ZN(n8508) );
  NOR2_X1 U10006 ( .A1(n8503), .A2(n9920), .ZN(n8506) );
  INV_X1 U10007 ( .A(n8767), .ZN(n8509) );
  MUX2_X1 U10008 ( .A(n8510), .B(n8509), .S(n9562), .Z(n8514) );
  AOI22_X1 U10009 ( .A1(n8512), .A2(n8664), .B1(n9934), .B2(n8511), .ZN(n8513)
         );
  OAI211_X1 U10010 ( .C1(n8769), .C2(n8667), .A(n8514), .B(n8513), .ZN(
        P2_U3205) );
  XOR2_X1 U10011 ( .A(n8516), .B(n8515), .Z(n8518) );
  AOI222_X1 U10012 ( .A1(n8671), .A2(n8518), .B1(n8538), .B2(n8687), .C1(n8517), .C2(n8684), .ZN(n8772) );
  MUX2_X1 U10013 ( .A(n8519), .B(n8772), .S(n9562), .Z(n8522) );
  AOI22_X1 U10014 ( .A1(n8774), .A2(n8664), .B1(n9934), .B2(n8520), .ZN(n8521)
         );
  OAI211_X1 U10015 ( .C1(n8777), .C2(n8667), .A(n8522), .B(n8521), .ZN(
        P2_U3206) );
  XNOR2_X1 U10016 ( .A(n8523), .B(n8524), .ZN(n8715) );
  INV_X1 U10017 ( .A(n8715), .ZN(n8535) );
  XNOR2_X1 U10018 ( .A(n8526), .B(n8525), .ZN(n8527) );
  OAI22_X1 U10019 ( .A1(n8527), .A2(n9928), .B1(n8549), .B2(n9922), .ZN(n8713)
         );
  AND2_X1 U10020 ( .A1(n8528), .A2(n8684), .ZN(n8714) );
  OAI21_X1 U10021 ( .B1(n8713), .B2(n8714), .A(n9562), .ZN(n8534) );
  INV_X1 U10022 ( .A(n8529), .ZN(n8531) );
  OAI22_X1 U10023 ( .A1(n8531), .A2(n9553), .B1(n9562), .B2(n8530), .ZN(n8532)
         );
  AOI21_X1 U10024 ( .B1(n8712), .B2(n8664), .A(n8532), .ZN(n8533) );
  OAI211_X1 U10025 ( .C1(n8535), .C2(n8667), .A(n8534), .B(n8533), .ZN(
        P2_U3207) );
  OAI21_X1 U10026 ( .B1(n8537), .B2(n8543), .A(n8536), .ZN(n8539) );
  AOI222_X1 U10027 ( .A1(n8671), .A2(n8539), .B1(n8538), .B2(n8684), .C1(n8561), .C2(n8687), .ZN(n8782) );
  AOI22_X1 U10028 ( .A1(n8784), .A2(n8673), .B1(n9934), .B2(n8540), .ZN(n8541)
         );
  AOI21_X1 U10029 ( .B1(n8782), .B2(n8541), .A(n9936), .ZN(n8546) );
  XOR2_X1 U10030 ( .A(n8542), .B(n8543), .Z(n8787) );
  OAI22_X1 U10031 ( .A1(n8787), .A2(n8667), .B1(n8544), .B2(n9562), .ZN(n8545)
         );
  OR2_X1 U10032 ( .A1(n8546), .A2(n8545), .ZN(P2_U3208) );
  NOR2_X1 U10033 ( .A1(n8789), .A2(n9929), .ZN(n8550) );
  XOR2_X1 U10034 ( .A(n8547), .B(n8555), .Z(n8548) );
  OAI222_X1 U10035 ( .A1(n9920), .A2(n8549), .B1(n9922), .B2(n8571), .C1(n9928), .C2(n8548), .ZN(n8788) );
  AOI211_X1 U10036 ( .C1(n9934), .C2(n8551), .A(n8550), .B(n8788), .ZN(n8557)
         );
  NAND2_X1 U10037 ( .A1(n8553), .A2(n8552), .ZN(n8554) );
  XOR2_X1 U10038 ( .A(n8555), .B(n8554), .Z(n8721) );
  AOI22_X1 U10039 ( .A1(n8721), .A2(n8698), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9936), .ZN(n8556) );
  OAI21_X1 U10040 ( .B1(n8557), .B2(n9936), .A(n8556), .ZN(P2_U3209) );
  XOR2_X1 U10041 ( .A(n8558), .B(n8560), .Z(n8798) );
  INV_X1 U10042 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8563) );
  XOR2_X1 U10043 ( .A(n8560), .B(n8559), .Z(n8562) );
  AOI222_X1 U10044 ( .A1(n8671), .A2(n8562), .B1(n8561), .B2(n8684), .C1(n8590), .C2(n8687), .ZN(n8793) );
  MUX2_X1 U10045 ( .A(n8563), .B(n8793), .S(n9562), .Z(n8566) );
  AOI22_X1 U10046 ( .A1(n8795), .A2(n8664), .B1(n9934), .B2(n8564), .ZN(n8565)
         );
  OAI211_X1 U10047 ( .C1(n8798), .C2(n8667), .A(n8566), .B(n8565), .ZN(
        P2_U3210) );
  AND3_X1 U10048 ( .A1(n8588), .A2(n8575), .A3(n8567), .ZN(n8568) );
  OAI21_X1 U10049 ( .B1(n8569), .B2(n8568), .A(n8671), .ZN(n8574) );
  OAI22_X1 U10050 ( .A1(n8571), .A2(n9920), .B1(n8570), .B2(n9922), .ZN(n8572)
         );
  INV_X1 U10051 ( .A(n8572), .ZN(n8573) );
  NAND2_X1 U10052 ( .A1(n8574), .A2(n8573), .ZN(n8731) );
  OR2_X1 U10053 ( .A1(n8576), .A2(n8575), .ZN(n8727) );
  NAND3_X1 U10054 ( .A1(n8727), .A2(n8577), .A3(n8698), .ZN(n8580) );
  AOI22_X1 U10055 ( .A1(n9936), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9934), .B2(
        n8578), .ZN(n8579) );
  OAI211_X1 U10056 ( .C1(n8729), .C2(n8695), .A(n8580), .B(n8579), .ZN(n8581)
         );
  AOI21_X1 U10057 ( .B1(n8731), .B2(n9562), .A(n8581), .ZN(n8582) );
  INV_X1 U10058 ( .A(n8582), .ZN(P2_U3211) );
  XNOR2_X1 U10059 ( .A(n8583), .B(n8584), .ZN(n8805) );
  INV_X1 U10060 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8592) );
  INV_X1 U10061 ( .A(n8584), .ZN(n8586) );
  NAND3_X1 U10062 ( .A1(n8600), .A2(n8586), .A3(n8585), .ZN(n8587) );
  NAND2_X1 U10063 ( .A1(n8588), .A2(n8587), .ZN(n8591) );
  AOI222_X1 U10064 ( .A1(n8671), .A2(n8591), .B1(n8590), .B2(n8684), .C1(n8589), .C2(n8687), .ZN(n8800) );
  MUX2_X1 U10065 ( .A(n8592), .B(n8800), .S(n9562), .Z(n8595) );
  AOI22_X1 U10066 ( .A1(n8802), .A2(n8664), .B1(n9934), .B2(n8593), .ZN(n8594)
         );
  OAI211_X1 U10067 ( .C1(n8805), .C2(n8667), .A(n8595), .B(n8594), .ZN(
        P2_U3212) );
  XNOR2_X1 U10068 ( .A(n8596), .B(n8597), .ZN(n8809) );
  NAND2_X1 U10069 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10070 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  NAND2_X1 U10071 ( .A1(n8601), .A2(n8671), .ZN(n8604) );
  AOI22_X1 U10072 ( .A1(n8602), .A2(n8684), .B1(n8687), .B2(n8627), .ZN(n8603)
         );
  NAND2_X1 U10073 ( .A1(n8604), .A2(n8603), .ZN(n8806) );
  MUX2_X1 U10074 ( .A(n8806), .B(P2_REG2_REG_20__SCAN_IN), .S(n9936), .Z(n8605) );
  INV_X1 U10075 ( .A(n8605), .ZN(n8608) );
  AOI22_X1 U10076 ( .A1(n8735), .A2(n8664), .B1(n8606), .B2(n9934), .ZN(n8607)
         );
  OAI211_X1 U10077 ( .C1(n8809), .C2(n8667), .A(n8608), .B(n8607), .ZN(
        P2_U3213) );
  XOR2_X1 U10078 ( .A(n8609), .B(n8610), .Z(n8817) );
  INV_X1 U10079 ( .A(n8610), .ZN(n8611) );
  XNOR2_X1 U10080 ( .A(n8612), .B(n8611), .ZN(n8616) );
  NAND2_X1 U10081 ( .A1(n8636), .A2(n8687), .ZN(n8613) );
  OAI21_X1 U10082 ( .B1(n8614), .B2(n9920), .A(n8613), .ZN(n8615) );
  AOI21_X1 U10083 ( .B1(n8616), .B2(n8671), .A(n8615), .ZN(n8812) );
  MUX2_X1 U10084 ( .A(n8812), .B(n8617), .S(n9936), .Z(n8620) );
  AOI22_X1 U10085 ( .A1(n8814), .A2(n8664), .B1(n9934), .B2(n8618), .ZN(n8619)
         );
  OAI211_X1 U10086 ( .C1(n8817), .C2(n8667), .A(n8620), .B(n8619), .ZN(
        P2_U3214) );
  XOR2_X1 U10087 ( .A(n8621), .B(n8625), .Z(n8823) );
  INV_X1 U10088 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U10089 ( .A1(n8634), .A2(n8635), .ZN(n8623) );
  NAND2_X1 U10090 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  XOR2_X1 U10091 ( .A(n8625), .B(n8624), .Z(n8628) );
  AOI222_X1 U10092 ( .A1(n8671), .A2(n8628), .B1(n8627), .B2(n8684), .C1(n8626), .C2(n8687), .ZN(n8818) );
  MUX2_X1 U10093 ( .A(n8629), .B(n8818), .S(n9562), .Z(n8632) );
  AOI22_X1 U10094 ( .A1(n8820), .A2(n8664), .B1(n9934), .B2(n8630), .ZN(n8631)
         );
  OAI211_X1 U10095 ( .C1(n8823), .C2(n8667), .A(n8632), .B(n8631), .ZN(
        P2_U3215) );
  XOR2_X1 U10096 ( .A(n8633), .B(n8635), .Z(n8829) );
  XOR2_X1 U10097 ( .A(n8635), .B(n8634), .Z(n8637) );
  AOI222_X1 U10098 ( .A1(n8671), .A2(n8637), .B1(n8636), .B2(n8684), .C1(n8660), .C2(n8687), .ZN(n8824) );
  MUX2_X1 U10099 ( .A(n8638), .B(n8824), .S(n9562), .Z(n8641) );
  AOI22_X1 U10100 ( .A1(n8826), .A2(n8664), .B1(n9934), .B2(n8639), .ZN(n8640)
         );
  OAI211_X1 U10101 ( .C1(n8829), .C2(n8667), .A(n8641), .B(n8640), .ZN(
        P2_U3216) );
  XOR2_X1 U10102 ( .A(n8642), .B(n8646), .Z(n8833) );
  NAND2_X1 U10103 ( .A1(n8658), .A2(n8643), .ZN(n8645) );
  NAND2_X1 U10104 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  XNOR2_X1 U10105 ( .A(n8647), .B(n8646), .ZN(n8648) );
  OAI222_X1 U10106 ( .A1(n9920), .A2(n8650), .B1(n9922), .B2(n8649), .C1(n9928), .C2(n8648), .ZN(n8748) );
  NAND2_X1 U10107 ( .A1(n8748), .A2(n9562), .ZN(n8655) );
  OAI22_X1 U10108 ( .A1(n9562), .A2(n8652), .B1(n8651), .B2(n9553), .ZN(n8653)
         );
  AOI21_X1 U10109 ( .B1(n8749), .B2(n8664), .A(n8653), .ZN(n8654) );
  OAI211_X1 U10110 ( .C1(n8833), .C2(n8667), .A(n8655), .B(n8654), .ZN(
        P2_U3217) );
  XNOR2_X1 U10111 ( .A(n8656), .B(n8657), .ZN(n8841) );
  XNOR2_X1 U10112 ( .A(n8658), .B(n8657), .ZN(n8661) );
  AOI222_X1 U10113 ( .A1(n8671), .A2(n8661), .B1(n8660), .B2(n8684), .C1(n8659), .C2(n8687), .ZN(n8834) );
  MUX2_X1 U10114 ( .A(n8662), .B(n8834), .S(n9562), .Z(n8666) );
  AOI22_X1 U10115 ( .A1(n8837), .A2(n8664), .B1(n9934), .B2(n8663), .ZN(n8665)
         );
  OAI211_X1 U10116 ( .C1(n8841), .C2(n8667), .A(n8666), .B(n8665), .ZN(
        P2_U3218) );
  XNOR2_X1 U10117 ( .A(n8668), .B(n8676), .ZN(n8670) );
  AOI222_X1 U10118 ( .A1(n8671), .A2(n8670), .B1(n8685), .B2(n8687), .C1(n8669), .C2(n8684), .ZN(n8760) );
  AOI22_X1 U10119 ( .A1(n8757), .A2(n8673), .B1(n9934), .B2(n8672), .ZN(n8674)
         );
  AND2_X1 U10120 ( .A1(n8760), .A2(n8674), .ZN(n8679) );
  OAI21_X1 U10121 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8758) );
  AOI22_X1 U10122 ( .A1(n8758), .A2(n8698), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9936), .ZN(n8678) );
  OAI21_X1 U10123 ( .B1(n8679), .B2(n9936), .A(n8678), .ZN(P2_U3219) );
  NOR2_X1 U10124 ( .A1(n7475), .A2(n8680), .ZN(n8682) );
  INV_X1 U10125 ( .A(n7475), .ZN(n8681) );
  OAI22_X1 U10126 ( .A1(n8682), .A2(n9978), .B1(n8681), .B2(n8686), .ZN(n8683)
         );
  XNOR2_X1 U10127 ( .A(n8683), .B(n8691), .ZN(n8689) );
  AOI22_X1 U10128 ( .A1(n8687), .A2(n8686), .B1(n8685), .B2(n8684), .ZN(n8688)
         );
  OAI21_X1 U10129 ( .B1(n8689), .B2(n9928), .A(n8688), .ZN(n9982) );
  AOI21_X1 U10130 ( .B1(n9934), .B2(n8690), .A(n9982), .ZN(n8700) );
  OR2_X1 U10131 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  AND2_X1 U10132 ( .A1(n8694), .A2(n8693), .ZN(n9981) );
  OAI22_X1 U10133 ( .A1(n8696), .A2(n8695), .B1(n7388), .B2(n9562), .ZN(n8697)
         );
  AOI21_X1 U10134 ( .B1(n9981), .B2(n8698), .A(n8697), .ZN(n8699) );
  OAI21_X1 U10135 ( .B1(n8700), .B2(n9936), .A(n8699), .ZN(P2_U3221) );
  NAND2_X1 U10136 ( .A1(n4849), .A2(n8753), .ZN(n8702) );
  INV_X1 U10137 ( .A(n8761), .ZN(n8701) );
  NAND2_X1 U10138 ( .A1(n8701), .A2(n10003), .ZN(n8704) );
  OAI211_X1 U10139 ( .C1(n10003), .C2(n8107), .A(n8702), .B(n8704), .ZN(
        P2_U3490) );
  INV_X1 U10140 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U10141 ( .A1(n8703), .A2(n8753), .ZN(n8705) );
  OAI211_X1 U10142 ( .C1(n10003), .C2(n8706), .A(n8705), .B(n8704), .ZN(
        P2_U3489) );
  MUX2_X1 U10143 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8767), .S(n10003), .Z(
        n8708) );
  OAI22_X1 U10144 ( .A1(n8769), .A2(n8756), .B1(n8768), .B2(n8736), .ZN(n8707)
         );
  OR2_X1 U10145 ( .A1(n8708), .A2(n8707), .ZN(P2_U3487) );
  INV_X1 U10146 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8709) );
  MUX2_X1 U10147 ( .A(n8709), .B(n8772), .S(n10003), .Z(n8711) );
  NAND2_X1 U10148 ( .A1(n8774), .A2(n8753), .ZN(n8710) );
  OAI211_X1 U10149 ( .C1(n8756), .C2(n8777), .A(n8711), .B(n8710), .ZN(
        P2_U3486) );
  INV_X1 U10150 ( .A(n8712), .ZN(n8781) );
  INV_X1 U10151 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8716) );
  AOI211_X1 U10152 ( .C1(n8715), .C2(n9980), .A(n8714), .B(n8713), .ZN(n8778)
         );
  MUX2_X1 U10153 ( .A(n8716), .B(n8778), .S(n10003), .Z(n8717) );
  OAI21_X1 U10154 ( .B1(n8781), .B2(n8736), .A(n8717), .ZN(P2_U3485) );
  INV_X1 U10155 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8718) );
  MUX2_X1 U10156 ( .A(n8718), .B(n8782), .S(n10003), .Z(n8720) );
  NAND2_X1 U10157 ( .A1(n8784), .A2(n8753), .ZN(n8719) );
  OAI211_X1 U10158 ( .C1(n8787), .C2(n8756), .A(n8720), .B(n8719), .ZN(
        P2_U3484) );
  MUX2_X1 U10159 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8788), .S(n10003), .Z(
        n8723) );
  INV_X1 U10160 ( .A(n8721), .ZN(n8790) );
  OAI22_X1 U10161 ( .A1(n8790), .A2(n8756), .B1(n8789), .B2(n8736), .ZN(n8722)
         );
  OR2_X1 U10162 ( .A1(n8723), .A2(n8722), .ZN(P2_U3483) );
  INV_X1 U10163 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U10164 ( .A(n8724), .B(n8793), .S(n10003), .Z(n8726) );
  NAND2_X1 U10165 ( .A1(n8795), .A2(n8753), .ZN(n8725) );
  OAI211_X1 U10166 ( .C1(n8798), .C2(n8756), .A(n8726), .B(n8725), .ZN(
        P2_U3482) );
  NAND3_X1 U10167 ( .A1(n8577), .A2(n8727), .A3(n9980), .ZN(n8728) );
  OAI21_X1 U10168 ( .B1(n8729), .B2(n9967), .A(n8728), .ZN(n8730) );
  MUX2_X1 U10169 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8799), .S(n10003), .Z(
        P2_U3481) );
  INV_X1 U10170 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8732) );
  MUX2_X1 U10171 ( .A(n8732), .B(n8800), .S(n10003), .Z(n8734) );
  NAND2_X1 U10172 ( .A1(n8802), .A2(n8753), .ZN(n8733) );
  OAI211_X1 U10173 ( .C1(n8756), .C2(n8805), .A(n8734), .B(n8733), .ZN(
        P2_U3480) );
  MUX2_X1 U10174 ( .A(n8806), .B(P2_REG1_REG_20__SCAN_IN), .S(n10004), .Z(
        n8738) );
  INV_X1 U10175 ( .A(n8735), .ZN(n8808) );
  OAI22_X1 U10176 ( .A1(n8809), .A2(n8756), .B1(n8808), .B2(n8736), .ZN(n8737)
         );
  OR2_X1 U10177 ( .A1(n8738), .A2(n8737), .ZN(P2_U3479) );
  INV_X1 U10178 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8739) );
  MUX2_X1 U10179 ( .A(n8739), .B(n8812), .S(n10003), .Z(n8741) );
  NAND2_X1 U10180 ( .A1(n8814), .A2(n8753), .ZN(n8740) );
  OAI211_X1 U10181 ( .C1(n8756), .C2(n8817), .A(n8741), .B(n8740), .ZN(
        P2_U3478) );
  INV_X1 U10182 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8742) );
  MUX2_X1 U10183 ( .A(n8742), .B(n8818), .S(n10003), .Z(n8744) );
  NAND2_X1 U10184 ( .A1(n8820), .A2(n8753), .ZN(n8743) );
  OAI211_X1 U10185 ( .C1(n8823), .C2(n8756), .A(n8744), .B(n8743), .ZN(
        P2_U3477) );
  MUX2_X1 U10186 ( .A(n8745), .B(n8824), .S(n10003), .Z(n8747) );
  NAND2_X1 U10187 ( .A1(n8826), .A2(n8753), .ZN(n8746) );
  OAI211_X1 U10188 ( .C1(n8829), .C2(n8756), .A(n8747), .B(n8746), .ZN(
        P2_U3476) );
  AOI21_X1 U10189 ( .B1(n9985), .B2(n8749), .A(n8748), .ZN(n8830) );
  MUX2_X1 U10190 ( .A(n8750), .B(n8830), .S(n10003), .Z(n8751) );
  OAI21_X1 U10191 ( .B1(n8756), .B2(n8833), .A(n8751), .ZN(P2_U3475) );
  MUX2_X1 U10192 ( .A(n8752), .B(n8834), .S(n10003), .Z(n8755) );
  NAND2_X1 U10193 ( .A1(n8837), .A2(n8753), .ZN(n8754) );
  OAI211_X1 U10194 ( .C1(n8841), .C2(n8756), .A(n8755), .B(n8754), .ZN(
        P2_U3474) );
  AOI22_X1 U10195 ( .A1(n8758), .A2(n9980), .B1(n9985), .B2(n8757), .ZN(n8759)
         );
  NAND2_X1 U10196 ( .A1(n8760), .A2(n8759), .ZN(n8842) );
  MUX2_X1 U10197 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8842), .S(n10003), .Z(
        P2_U3473) );
  NOR2_X1 U10198 ( .A1(n8761), .A2(n9988), .ZN(n8764) );
  AOI21_X1 U10199 ( .B1(n9988), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8764), .ZN(
        n8762) );
  OAI21_X1 U10200 ( .B1(n8763), .B2(n8807), .A(n8762), .ZN(P2_U3458) );
  AOI21_X1 U10201 ( .B1(n9988), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8764), .ZN(
        n8765) );
  OAI21_X1 U10202 ( .B1(n8766), .B2(n8807), .A(n8765), .ZN(P2_U3457) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8767), .S(n9986), .Z(n8771) );
  INV_X1 U10204 ( .A(n9980), .ZN(n9974) );
  OAI22_X1 U10205 ( .A1(n8769), .A2(n8840), .B1(n8768), .B2(n8807), .ZN(n8770)
         );
  OR2_X1 U10206 ( .A1(n8771), .A2(n8770), .ZN(P2_U3455) );
  INV_X1 U10207 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8773) );
  MUX2_X1 U10208 ( .A(n8773), .B(n8772), .S(n9986), .Z(n8776) );
  NAND2_X1 U10209 ( .A1(n8774), .A2(n8836), .ZN(n8775) );
  OAI211_X1 U10210 ( .C1(n8777), .C2(n8840), .A(n8776), .B(n8775), .ZN(
        P2_U3454) );
  INV_X1 U10211 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8779) );
  MUX2_X1 U10212 ( .A(n8779), .B(n8778), .S(n9986), .Z(n8780) );
  OAI21_X1 U10213 ( .B1(n8781), .B2(n8807), .A(n8780), .ZN(P2_U3453) );
  INV_X1 U10214 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8783) );
  MUX2_X1 U10215 ( .A(n8783), .B(n8782), .S(n9986), .Z(n8786) );
  NAND2_X1 U10216 ( .A1(n8784), .A2(n8836), .ZN(n8785) );
  OAI211_X1 U10217 ( .C1(n8787), .C2(n8840), .A(n8786), .B(n8785), .ZN(
        P2_U3452) );
  MUX2_X1 U10218 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8788), .S(n9986), .Z(n8792) );
  OAI22_X1 U10219 ( .A1(n8790), .A2(n8840), .B1(n8789), .B2(n8807), .ZN(n8791)
         );
  OR2_X1 U10220 ( .A1(n8792), .A2(n8791), .ZN(P2_U3451) );
  INV_X1 U10221 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8794) );
  MUX2_X1 U10222 ( .A(n8794), .B(n8793), .S(n9986), .Z(n8797) );
  NAND2_X1 U10223 ( .A1(n8795), .A2(n8836), .ZN(n8796) );
  OAI211_X1 U10224 ( .C1(n8798), .C2(n8840), .A(n8797), .B(n8796), .ZN(
        P2_U3450) );
  MUX2_X1 U10225 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8799), .S(n9986), .Z(
        P2_U3449) );
  INV_X1 U10226 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8801) );
  MUX2_X1 U10227 ( .A(n8801), .B(n8800), .S(n9986), .Z(n8804) );
  NAND2_X1 U10228 ( .A1(n8802), .A2(n8836), .ZN(n8803) );
  OAI211_X1 U10229 ( .C1(n8805), .C2(n8840), .A(n8804), .B(n8803), .ZN(
        P2_U3448) );
  MUX2_X1 U10230 ( .A(n8806), .B(P2_REG0_REG_20__SCAN_IN), .S(n9988), .Z(n8811) );
  OAI22_X1 U10231 ( .A1(n8809), .A2(n8840), .B1(n8808), .B2(n8807), .ZN(n8810)
         );
  OR2_X1 U10232 ( .A1(n8811), .A2(n8810), .ZN(P2_U3447) );
  INV_X1 U10233 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8813) );
  MUX2_X1 U10234 ( .A(n8813), .B(n8812), .S(n9986), .Z(n8816) );
  NAND2_X1 U10235 ( .A1(n8814), .A2(n8836), .ZN(n8815) );
  OAI211_X1 U10236 ( .C1(n8817), .C2(n8840), .A(n8816), .B(n8815), .ZN(
        P2_U3446) );
  INV_X1 U10237 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8819) );
  MUX2_X1 U10238 ( .A(n8819), .B(n8818), .S(n9986), .Z(n8822) );
  NAND2_X1 U10239 ( .A1(n8820), .A2(n8836), .ZN(n8821) );
  OAI211_X1 U10240 ( .C1(n8823), .C2(n8840), .A(n8822), .B(n8821), .ZN(
        P2_U3444) );
  INV_X1 U10241 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8825) );
  MUX2_X1 U10242 ( .A(n8825), .B(n8824), .S(n9986), .Z(n8828) );
  NAND2_X1 U10243 ( .A1(n8826), .A2(n8836), .ZN(n8827) );
  OAI211_X1 U10244 ( .C1(n8829), .C2(n8840), .A(n8828), .B(n8827), .ZN(
        P2_U3441) );
  INV_X1 U10245 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8831) );
  MUX2_X1 U10246 ( .A(n8831), .B(n8830), .S(n9986), .Z(n8832) );
  OAI21_X1 U10247 ( .B1(n8833), .B2(n8840), .A(n8832), .ZN(P2_U3438) );
  INV_X1 U10248 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U10249 ( .A(n8835), .B(n8834), .S(n9986), .Z(n8839) );
  NAND2_X1 U10250 ( .A1(n8837), .A2(n8836), .ZN(n8838) );
  OAI211_X1 U10251 ( .C1(n8841), .C2(n8840), .A(n8839), .B(n8838), .ZN(
        P2_U3435) );
  MUX2_X1 U10252 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8842), .S(n9986), .Z(
        P2_U3432) );
  MUX2_X1 U10253 ( .A(n8844), .B(P2_D_REG_1__SCAN_IN), .S(n8843), .Z(P2_U3377)
         );
  INV_X1 U10254 ( .A(n8845), .ZN(n9474) );
  INV_X1 U10255 ( .A(n8846), .ZN(n8848) );
  NOR4_X1 U10256 ( .A1(n8848), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9827), .A4(
        n8847), .ZN(n8849) );
  AOI21_X1 U10257 ( .B1(n8850), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8849), .ZN(
        n8851) );
  OAI21_X1 U10258 ( .B1(n9474), .B2(n8855), .A(n8851), .ZN(P2_U3264) );
  INV_X1 U10259 ( .A(n8852), .ZN(n9482) );
  OAI222_X1 U10260 ( .A1(n9827), .A2(n8856), .B1(n8855), .B2(n9482), .C1(n8854), .C2(n8853), .ZN(P2_U3266) );
  MUX2_X1 U10261 ( .A(n8857), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10262 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n8861) );
  NAND2_X1 U10263 ( .A1(n8861), .A2(n8991), .ZN(n8866) );
  NAND2_X1 U10264 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9678) );
  OAI21_X1 U10265 ( .B1(n8994), .B2(n8908), .A(n9678), .ZN(n8864) );
  NOR2_X1 U10266 ( .A1(n8996), .A2(n8862), .ZN(n8863) );
  AOI211_X1 U10267 ( .C1(n8999), .C2(n9804), .A(n8864), .B(n8863), .ZN(n8865)
         );
  OAI211_X1 U10268 ( .C1(n9409), .C2(n9002), .A(n8866), .B(n8865), .ZN(
        P1_U3215) );
  INV_X1 U10269 ( .A(n8922), .ZN(n8869) );
  NOR3_X1 U10270 ( .A1(n8939), .A2(n8943), .A3(n8867), .ZN(n8868) );
  OAI21_X1 U10271 ( .B1(n8869), .B2(n8868), .A(n8991), .ZN(n8874) );
  AOI22_X1 U10272 ( .A1(n9347), .A2(n8985), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8871) );
  NAND2_X1 U10273 ( .A1(n9365), .A2(n8999), .ZN(n8870) );
  OAI211_X1 U10274 ( .C1(n8996), .C2(n9175), .A(n8871), .B(n8870), .ZN(n8872)
         );
  AOI21_X1 U10275 ( .B1(n9187), .B2(n8971), .A(n8872), .ZN(n8873) );
  NAND2_X1 U10276 ( .A1(n8874), .A2(n8873), .ZN(P1_U3216) );
  INV_X1 U10277 ( .A(n8875), .ZN(n8877) );
  XOR2_X1 U10278 ( .A(n8876), .B(n8875), .Z(n8966) );
  NOR2_X1 U10279 ( .A1(n8966), .A2(n8965), .ZN(n8964) );
  AOI21_X1 U10280 ( .B1(n8877), .B2(n8876), .A(n8964), .ZN(n8881) );
  XNOR2_X1 U10281 ( .A(n8879), .B(n8878), .ZN(n8880) );
  XNOR2_X1 U10282 ( .A(n8881), .B(n8880), .ZN(n8887) );
  OAI21_X1 U10283 ( .B1(n8994), .B2(n9217), .A(n8882), .ZN(n8883) );
  AOI21_X1 U10284 ( .B1(n8999), .B2(n9242), .A(n8883), .ZN(n8884) );
  OAI21_X1 U10285 ( .B1(n8996), .B2(n9246), .A(n8884), .ZN(n8885) );
  AOI21_X1 U10286 ( .B1(n9245), .B2(n8971), .A(n8885), .ZN(n8886) );
  OAI21_X1 U10287 ( .B1(n8887), .B2(n8973), .A(n8886), .ZN(P1_U3219) );
  XOR2_X1 U10288 ( .A(n8889), .B(n8888), .Z(n8894) );
  AOI22_X1 U10289 ( .A1(n9365), .A2(n8985), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8891) );
  NAND2_X1 U10290 ( .A1(n8999), .A2(n9364), .ZN(n8890) );
  OAI211_X1 U10291 ( .C1(n8996), .C2(n9212), .A(n8891), .B(n8890), .ZN(n8892)
         );
  AOI21_X1 U10292 ( .B1(n9222), .B2(n8971), .A(n8892), .ZN(n8893) );
  OAI21_X1 U10293 ( .B1(n8894), .B2(n8973), .A(n8893), .ZN(P1_U3223) );
  AOI21_X1 U10294 ( .B1(n8897), .B2(n8896), .A(n8895), .ZN(n8904) );
  NOR2_X1 U10295 ( .A1(n8996), .A2(n9149), .ZN(n8902) );
  NAND2_X1 U10296 ( .A1(n9140), .A2(n8985), .ZN(n8899) );
  NAND2_X1 U10297 ( .A1(P1_U3086), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8898) );
  OAI211_X1 U10298 ( .C1(n8900), .C2(n8983), .A(n8899), .B(n8898), .ZN(n8901)
         );
  AOI211_X1 U10299 ( .C1(n9148), .C2(n8971), .A(n8902), .B(n8901), .ZN(n8903)
         );
  OAI21_X1 U10300 ( .B1(n8904), .B2(n8973), .A(n8903), .ZN(P1_U3225) );
  XOR2_X1 U10301 ( .A(n8906), .B(n8905), .Z(n8912) );
  NAND2_X1 U10302 ( .A1(n8985), .A2(n9301), .ZN(n8907) );
  NAND2_X1 U10303 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9703) );
  OAI211_X1 U10304 ( .C1(n8908), .C2(n8983), .A(n8907), .B(n9703), .ZN(n8909)
         );
  AOI21_X1 U10305 ( .B1(n9294), .B2(n8980), .A(n8909), .ZN(n8911) );
  NAND2_X1 U10306 ( .A1(n9398), .A2(n8971), .ZN(n8910) );
  OAI211_X1 U10307 ( .C1(n8912), .C2(n8973), .A(n8911), .B(n8910), .ZN(
        P1_U3226) );
  XOR2_X1 U10308 ( .A(n8913), .B(n8914), .Z(n8919) );
  NAND2_X1 U10309 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9714) );
  OAI21_X1 U10310 ( .B1(n8994), .B2(n9392), .A(n9714), .ZN(n8915) );
  AOI21_X1 U10311 ( .B1(n8999), .B2(n9271), .A(n8915), .ZN(n8916) );
  OAI21_X1 U10312 ( .B1(n8996), .B2(n9276), .A(n8916), .ZN(n8917) );
  AOI21_X1 U10313 ( .B1(n9285), .B2(n8971), .A(n8917), .ZN(n8918) );
  OAI21_X1 U10314 ( .B1(n8919), .B2(n8973), .A(n8918), .ZN(P1_U3228) );
  AND3_X1 U10315 ( .A1(n8922), .A2(n8921), .A3(n8920), .ZN(n8923) );
  OAI21_X1 U10316 ( .B1(n8924), .B2(n8923), .A(n8991), .ZN(n8929) );
  AOI22_X1 U10317 ( .A1(n9159), .A2(n8985), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8926) );
  NAND2_X1 U10318 ( .A1(n9356), .A2(n8999), .ZN(n8925) );
  OAI211_X1 U10319 ( .C1(n8996), .C2(n9165), .A(n8926), .B(n8925), .ZN(n8927)
         );
  AOI21_X1 U10320 ( .B1(n5882), .B2(n8971), .A(n8927), .ZN(n8928) );
  NAND2_X1 U10321 ( .A1(n8929), .A2(n8928), .ZN(P1_U3229) );
  XNOR2_X1 U10322 ( .A(n8931), .B(n8930), .ZN(n8932) );
  XNOR2_X1 U10323 ( .A(n8933), .B(n8932), .ZN(n8938) );
  AOI22_X1 U10324 ( .A1(n8985), .A2(n9355), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8935) );
  NAND2_X1 U10325 ( .A1(n8980), .A2(n9229), .ZN(n8934) );
  OAI211_X1 U10326 ( .C1(n8967), .C2(n8983), .A(n8935), .B(n8934), .ZN(n8936)
         );
  AOI21_X1 U10327 ( .B1(n9234), .B2(n8971), .A(n8936), .ZN(n8937) );
  OAI21_X1 U10328 ( .B1(n8938), .B2(n8973), .A(n8937), .ZN(P1_U3233) );
  INV_X1 U10329 ( .A(n8939), .ZN(n8944) );
  OAI21_X1 U10330 ( .B1(n8941), .B2(n8943), .A(n8940), .ZN(n8942) );
  OAI21_X1 U10331 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(n8945) );
  NAND2_X1 U10332 ( .A1(n8945), .A2(n8991), .ZN(n8949) );
  AOI22_X1 U10333 ( .A1(n9356), .A2(n8985), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8946) );
  OAI21_X1 U10334 ( .B1(n9375), .B2(n8983), .A(n8946), .ZN(n8947) );
  AOI21_X1 U10335 ( .B1(n9196), .B2(n8980), .A(n8947), .ZN(n8948) );
  OAI211_X1 U10336 ( .C1(n9444), .C2(n9002), .A(n8949), .B(n8948), .ZN(
        P1_U3235) );
  AOI21_X1 U10337 ( .B1(n8951), .B2(n7313), .A(n8950), .ZN(n8955) );
  XNOR2_X1 U10338 ( .A(n8953), .B(n8952), .ZN(n8954) );
  XNOR2_X1 U10339 ( .A(n8955), .B(n8954), .ZN(n8963) );
  NAND2_X1 U10340 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9628) );
  OAI21_X1 U10341 ( .B1(n8983), .B2(n8956), .A(n9628), .ZN(n8957) );
  AOI21_X1 U10342 ( .B1(n8985), .B2(n9006), .A(n8957), .ZN(n8958) );
  OAI21_X1 U10343 ( .B1(n8996), .B2(n8959), .A(n8958), .ZN(n8960) );
  AOI21_X1 U10344 ( .B1(n8961), .B2(n8971), .A(n8960), .ZN(n8962) );
  OAI21_X1 U10345 ( .B1(n8963), .B2(n8973), .A(n8962), .ZN(P1_U3236) );
  AOI21_X1 U10346 ( .B1(n8966), .B2(n8965), .A(n8964), .ZN(n8974) );
  NAND2_X1 U10347 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9730) );
  OAI21_X1 U10348 ( .B1(n8994), .B2(n8967), .A(n9730), .ZN(n8968) );
  AOI21_X1 U10349 ( .B1(n8999), .B2(n9301), .A(n8968), .ZN(n8969) );
  OAI21_X1 U10350 ( .B1(n8996), .B2(n9258), .A(n8969), .ZN(n8970) );
  AOI21_X1 U10351 ( .B1(n9386), .B2(n8971), .A(n8970), .ZN(n8972) );
  OAI21_X1 U10352 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(P1_U3238) );
  OAI21_X1 U10353 ( .B1(n8895), .B2(n8977), .A(n8976), .ZN(n8978) );
  NAND3_X1 U10354 ( .A1(n8979), .A2(n8991), .A3(n8978), .ZN(n8987) );
  NAND2_X1 U10355 ( .A1(P1_U3086), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U10356 ( .A1(n9128), .A2(n8980), .ZN(n8981) );
  OAI211_X1 U10357 ( .C1(n9326), .C2(n8983), .A(n8982), .B(n8981), .ZN(n8984)
         );
  AOI21_X1 U10358 ( .B1(n9131), .B2(n8985), .A(n8984), .ZN(n8986) );
  OAI211_X1 U10359 ( .C1(n9429), .C2(n9002), .A(n8987), .B(n8986), .ZN(
        P1_U3240) );
  OAI21_X1 U10360 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8992) );
  NAND2_X1 U10361 ( .A1(n8992), .A2(n8991), .ZN(n9001) );
  NAND2_X1 U10362 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9689) );
  OAI21_X1 U10363 ( .B1(n8994), .B2(n8993), .A(n9689), .ZN(n8998) );
  NOR2_X1 U10364 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  AOI211_X1 U10365 ( .C1(n8999), .C2(n9005), .A(n8998), .B(n8997), .ZN(n9000)
         );
  OAI211_X1 U10366 ( .C1(n9467), .C2(n9002), .A(n9001), .B(n9000), .ZN(
        P1_U3241) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9003), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9099), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9004), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9131), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9159), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9347), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9356), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9365), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9355), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9364), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9265), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9242), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9301), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9271), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9302), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9005), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9804), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9006), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9007), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9008), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9009), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9010), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n4349), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9012), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5814), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9013), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9014), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10395 ( .C1(n9017), .C2(n9016), .A(n9712), .B(n9015), .ZN(n9024)
         );
  AOI22_X1 U10396 ( .A1(n9593), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9023) );
  NAND2_X1 U10397 ( .A1(n9724), .A2(n9018), .ZN(n9022) );
  OAI211_X1 U10398 ( .C1(n9020), .C2(n9027), .A(n9717), .B(n9019), .ZN(n9021)
         );
  NAND4_X1 U10399 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(
        P1_U3244) );
  MUX2_X1 U10400 ( .A(n9027), .B(n9026), .S(n9025), .Z(n9028) );
  NAND2_X1 U10401 ( .A1(n9028), .A2(n4355), .ZN(n9033) );
  NAND2_X1 U10402 ( .A1(n4358), .A2(n9029), .ZN(n9030) );
  NAND2_X1 U10403 ( .A1(n9030), .A2(n4355), .ZN(n9572) );
  INV_X1 U10404 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U10405 ( .A1(n9572), .A2(n9031), .ZN(n9575) );
  AND2_X1 U10406 ( .A1(P1_U3973), .A2(n9575), .ZN(n9032) );
  NAND2_X1 U10407 ( .A1(n9033), .A2(n9032), .ZN(n9595) );
  INV_X1 U10408 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9035) );
  OAI22_X1 U10409 ( .A1(n9732), .A2(n9035), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9034), .ZN(n9036) );
  AOI21_X1 U10410 ( .B1(n9037), .B2(n9724), .A(n9036), .ZN(n9046) );
  OAI211_X1 U10411 ( .C1(n9040), .C2(n9039), .A(n9712), .B(n9038), .ZN(n9045)
         );
  OAI211_X1 U10412 ( .C1(n9043), .C2(n9042), .A(n9717), .B(n9041), .ZN(n9044)
         );
  NAND4_X1 U10413 ( .A1(n9595), .A2(n9046), .A3(n9045), .A4(n9044), .ZN(
        P1_U3245) );
  INV_X1 U10414 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9048) );
  OAI21_X1 U10415 ( .B1(n9732), .B2(n9048), .A(n9047), .ZN(n9049) );
  AOI21_X1 U10416 ( .B1(n9050), .B2(n9724), .A(n9049), .ZN(n9059) );
  OAI211_X1 U10417 ( .C1(n9053), .C2(n9052), .A(n9717), .B(n9051), .ZN(n9058)
         );
  OAI211_X1 U10418 ( .C1(n9056), .C2(n9055), .A(n9712), .B(n9054), .ZN(n9057)
         );
  NAND3_X1 U10419 ( .A1(n9059), .A2(n9058), .A3(n9057), .ZN(P1_U3246) );
  INV_X1 U10420 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9061) );
  OAI21_X1 U10421 ( .B1(n9732), .B2(n9061), .A(n9060), .ZN(n9062) );
  AOI21_X1 U10422 ( .B1(n9063), .B2(n9724), .A(n9062), .ZN(n9072) );
  OAI211_X1 U10423 ( .C1(n9066), .C2(n9065), .A(n9717), .B(n9064), .ZN(n9071)
         );
  OAI211_X1 U10424 ( .C1(n9069), .C2(n9068), .A(n9712), .B(n9067), .ZN(n9070)
         );
  NAND3_X1 U10425 ( .A1(n9072), .A2(n9071), .A3(n9070), .ZN(P1_U3249) );
  XNOR2_X1 U10426 ( .A(n9417), .B(n9080), .ZN(n9073) );
  NAND2_X1 U10427 ( .A1(n9073), .A2(n9761), .ZN(n9308) );
  INV_X1 U10428 ( .A(n9074), .ZN(n9075) );
  NAND2_X1 U10429 ( .A1(n9076), .A2(n9075), .ZN(n9311) );
  NOR2_X1 U10430 ( .A1(n9295), .A2(n9311), .ZN(n9083) );
  NOR2_X1 U10431 ( .A1(n9417), .A2(n9756), .ZN(n9077) );
  AOI211_X1 U10432 ( .C1(n9295), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9083), .B(
        n9077), .ZN(n9078) );
  OAI21_X1 U10433 ( .B1(n9308), .B2(n9282), .A(n9078), .ZN(P1_U3263) );
  AOI21_X1 U10434 ( .B1(n9084), .B2(n9079), .A(n9291), .ZN(n9081) );
  NAND2_X1 U10435 ( .A1(n9081), .A2(n9080), .ZN(n9312) );
  AND2_X1 U10436 ( .A1(n9295), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9082) );
  NOR2_X1 U10437 ( .A1(n9083), .A2(n9082), .ZN(n9086) );
  NAND2_X1 U10438 ( .A1(n9084), .A2(n9286), .ZN(n9085) );
  OAI211_X1 U10439 ( .C1(n9312), .C2(n9282), .A(n9086), .B(n9085), .ZN(
        P1_U3264) );
  AOI22_X1 U10440 ( .A1(n9087), .A2(n9293), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9295), .ZN(n9088) );
  OAI21_X1 U10441 ( .B1(n9317), .B2(n9216), .A(n9088), .ZN(n9089) );
  AOI21_X1 U10442 ( .B1(n9090), .B2(n9286), .A(n9089), .ZN(n9091) );
  OAI21_X1 U10443 ( .B1(n9092), .B2(n9282), .A(n9091), .ZN(n9093) );
  AOI21_X1 U10444 ( .B1(n9094), .B2(n9275), .A(n9093), .ZN(n9095) );
  OAI21_X1 U10445 ( .B1(n9096), .B2(n9295), .A(n9095), .ZN(P1_U3356) );
  INV_X1 U10446 ( .A(n9097), .ZN(n9109) );
  NOR2_X1 U10447 ( .A1(n9098), .A2(n9756), .ZN(n9104) );
  NAND2_X1 U10448 ( .A1(n9099), .A2(n9211), .ZN(n9102) );
  AOI22_X1 U10449 ( .A1(n9100), .A2(n9293), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9295), .ZN(n9101) );
  OAI211_X1 U10450 ( .C1(n9327), .C2(n9216), .A(n9102), .B(n9101), .ZN(n9103)
         );
  AOI211_X1 U10451 ( .C1(n9105), .C2(n9764), .A(n9104), .B(n9103), .ZN(n9108)
         );
  NAND2_X1 U10452 ( .A1(n9106), .A2(n9135), .ZN(n9107) );
  OAI211_X1 U10453 ( .C1(n9109), .C2(n9307), .A(n9108), .B(n9107), .ZN(
        P1_U3265) );
  XNOR2_X1 U10454 ( .A(n9110), .B(n9111), .ZN(n9323) );
  OAI211_X1 U10455 ( .C1(n9425), .C2(n9126), .A(n9761), .B(n9112), .ZN(n9320)
         );
  AOI22_X1 U10456 ( .A1(n9140), .A2(n9113), .B1(n9295), .B2(
        P1_REG2_REG_27__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10457 ( .A1(n9114), .A2(n9293), .ZN(n9115) );
  OAI211_X1 U10458 ( .C1(n9317), .C2(n9279), .A(n9116), .B(n9115), .ZN(n9117)
         );
  AOI21_X1 U10459 ( .B1(n9118), .B2(n9286), .A(n9117), .ZN(n9119) );
  OAI21_X1 U10460 ( .B1(n9320), .B2(n9282), .A(n9119), .ZN(n9120) );
  AOI21_X1 U10461 ( .B1(n9315), .B2(n9275), .A(n9120), .ZN(n9121) );
  OAI21_X1 U10462 ( .B1(n9323), .B2(n9225), .A(n9121), .ZN(P1_U3266) );
  XOR2_X1 U10463 ( .A(n9124), .B(n9122), .Z(n9334) );
  INV_X1 U10464 ( .A(n9334), .ZN(n9137) );
  OAI21_X1 U10465 ( .B1(n9125), .B2(n9124), .A(n9123), .ZN(n9330) );
  AOI211_X1 U10466 ( .C1(n9127), .C2(n9146), .A(n9291), .B(n9126), .ZN(n9328)
         );
  NAND2_X1 U10467 ( .A1(n9328), .A2(n9764), .ZN(n9133) );
  AOI22_X1 U10468 ( .A1(n9128), .A2(n9293), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9295), .ZN(n9129) );
  OAI21_X1 U10469 ( .B1(n9326), .B2(n9216), .A(n9129), .ZN(n9130) );
  AOI21_X1 U10470 ( .B1(n9131), .B2(n9211), .A(n9130), .ZN(n9132) );
  OAI211_X1 U10471 ( .C1(n9429), .C2(n9756), .A(n9133), .B(n9132), .ZN(n9134)
         );
  AOI21_X1 U10472 ( .B1(n9135), .B2(n9330), .A(n9134), .ZN(n9136) );
  OAI21_X1 U10473 ( .B1(n9137), .B2(n9307), .A(n9136), .ZN(P1_U3267) );
  XNOR2_X1 U10474 ( .A(n9138), .B(n9143), .ZN(n9139) );
  NAND2_X1 U10475 ( .A1(n9139), .A2(n9331), .ZN(n9142) );
  AOI22_X1 U10476 ( .A1(n9140), .A2(n9805), .B1(n9796), .B2(n9347), .ZN(n9141)
         );
  NAND2_X1 U10477 ( .A1(n9142), .A2(n9141), .ZN(n9337) );
  INV_X1 U10478 ( .A(n9337), .ZN(n9155) );
  XOR2_X1 U10479 ( .A(n9144), .B(n9143), .Z(n9339) );
  NAND2_X1 U10480 ( .A1(n9339), .A2(n9275), .ZN(n9154) );
  INV_X1 U10481 ( .A(n9146), .ZN(n9147) );
  AOI211_X1 U10482 ( .C1(n9148), .C2(n9164), .A(n9291), .B(n9147), .ZN(n9338)
         );
  INV_X1 U10483 ( .A(n9149), .ZN(n9150) );
  AOI22_X1 U10484 ( .A1(n9150), .A2(n9293), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9295), .ZN(n9151) );
  OAI21_X1 U10485 ( .B1(n5883), .B2(n9756), .A(n9151), .ZN(n9152) );
  AOI21_X1 U10486 ( .B1(n9338), .B2(n9764), .A(n9152), .ZN(n9153) );
  OAI211_X1 U10487 ( .C1(n9295), .C2(n9155), .A(n9154), .B(n9153), .ZN(
        P1_U3268) );
  NAND2_X1 U10488 ( .A1(n9156), .A2(n9163), .ZN(n9157) );
  NAND3_X1 U10489 ( .A1(n9158), .A2(n9331), .A3(n9157), .ZN(n9161) );
  AOI22_X1 U10490 ( .A1(n9159), .A2(n9805), .B1(n9796), .B2(n9356), .ZN(n9160)
         );
  NAND2_X1 U10491 ( .A1(n9161), .A2(n9160), .ZN(n9342) );
  INV_X1 U10492 ( .A(n9342), .ZN(n9171) );
  XNOR2_X1 U10493 ( .A(n9163), .B(n9162), .ZN(n9344) );
  NAND2_X1 U10494 ( .A1(n9344), .A2(n9275), .ZN(n9170) );
  AOI211_X1 U10495 ( .C1(n5882), .C2(n9183), .A(n9291), .B(n9145), .ZN(n9343)
         );
  INV_X1 U10496 ( .A(n9165), .ZN(n9166) );
  AOI22_X1 U10497 ( .A1(n9166), .A2(n9293), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9295), .ZN(n9167) );
  OAI21_X1 U10498 ( .B1(n9436), .B2(n9756), .A(n9167), .ZN(n9168) );
  AOI21_X1 U10499 ( .B1(n9343), .B2(n9764), .A(n9168), .ZN(n9169) );
  OAI211_X1 U10500 ( .C1(n9295), .C2(n9171), .A(n9170), .B(n9169), .ZN(
        P1_U3269) );
  XOR2_X1 U10501 ( .A(n9172), .B(n9173), .Z(n9350) );
  XNOR2_X1 U10502 ( .A(n9174), .B(n9173), .ZN(n9352) );
  NAND2_X1 U10503 ( .A1(n9352), .A2(n9275), .ZN(n9189) );
  INV_X1 U10504 ( .A(n9175), .ZN(n9176) );
  NAND2_X1 U10505 ( .A1(n9293), .A2(n9176), .ZN(n9178) );
  NAND2_X1 U10506 ( .A1(n9295), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U10507 ( .A1(n9178), .A2(n9177), .ZN(n9179) );
  AOI21_X1 U10508 ( .B1(n9211), .B2(n9347), .A(n9179), .ZN(n9180) );
  OAI21_X1 U10509 ( .B1(n9181), .B2(n9216), .A(n9180), .ZN(n9186) );
  INV_X1 U10510 ( .A(n9182), .ZN(n9199) );
  NAND2_X1 U10511 ( .A1(n9199), .A2(n9187), .ZN(n9184) );
  NAND3_X1 U10512 ( .A1(n9184), .A2(n9183), .A3(n9761), .ZN(n9348) );
  NOR2_X1 U10513 ( .A1(n9348), .A2(n9282), .ZN(n9185) );
  AOI211_X1 U10514 ( .C1(n9286), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9188)
         );
  OAI211_X1 U10515 ( .C1(n9350), .C2(n9225), .A(n9189), .B(n9188), .ZN(
        P1_U3270) );
  INV_X1 U10516 ( .A(n9195), .ZN(n9190) );
  XNOR2_X1 U10517 ( .A(n9191), .B(n9190), .ZN(n9359) );
  NAND2_X1 U10518 ( .A1(n9192), .A2(n9193), .ZN(n9194) );
  XOR2_X1 U10519 ( .A(n9195), .B(n9194), .Z(n9361) );
  NAND2_X1 U10520 ( .A1(n9361), .A2(n9275), .ZN(n9205) );
  NAND2_X1 U10521 ( .A1(n9356), .A2(n9211), .ZN(n9198) );
  AOI22_X1 U10522 ( .A1(n9196), .A2(n9293), .B1(n9295), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9197) );
  OAI211_X1 U10523 ( .C1(n9375), .C2(n9216), .A(n9198), .B(n9197), .ZN(n9202)
         );
  INV_X1 U10524 ( .A(n9218), .ZN(n9200) );
  OAI211_X1 U10525 ( .C1(n9444), .C2(n9200), .A(n9199), .B(n9761), .ZN(n9357)
         );
  NOR2_X1 U10526 ( .A1(n9357), .A2(n9282), .ZN(n9201) );
  AOI211_X1 U10527 ( .C1(n9286), .C2(n9203), .A(n9202), .B(n9201), .ZN(n9204)
         );
  OAI211_X1 U10528 ( .C1(n9359), .C2(n9225), .A(n9205), .B(n9204), .ZN(
        P1_U3271) );
  OAI21_X1 U10529 ( .B1(n9207), .B2(n9209), .A(n9206), .ZN(n9208) );
  INV_X1 U10530 ( .A(n9208), .ZN(n9368) );
  XNOR2_X1 U10531 ( .A(n9210), .B(n9209), .ZN(n9370) );
  NAND2_X1 U10532 ( .A1(n9370), .A2(n9275), .ZN(n9224) );
  NAND2_X1 U10533 ( .A1(n9211), .A2(n9365), .ZN(n9215) );
  INV_X1 U10534 ( .A(n9212), .ZN(n9213) );
  AOI22_X1 U10535 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9295), .B1(n9213), .B2(
        n9293), .ZN(n9214) );
  OAI211_X1 U10536 ( .C1(n9217), .C2(n9216), .A(n9215), .B(n9214), .ZN(n9221)
         );
  INV_X1 U10537 ( .A(n9222), .ZN(n9448) );
  INV_X1 U10538 ( .A(n9231), .ZN(n9219) );
  OAI211_X1 U10539 ( .C1(n9448), .C2(n9219), .A(n9761), .B(n9218), .ZN(n9366)
         );
  NOR2_X1 U10540 ( .A1(n9366), .A2(n9282), .ZN(n9220) );
  AOI211_X1 U10541 ( .C1(n9286), .C2(n9222), .A(n9221), .B(n9220), .ZN(n9223)
         );
  OAI211_X1 U10542 ( .C1(n9368), .C2(n9225), .A(n9224), .B(n9223), .ZN(
        P1_U3272) );
  XNOR2_X1 U10543 ( .A(n4383), .B(n9227), .ZN(n9226) );
  AOI22_X1 U10544 ( .A1(n9226), .A2(n9331), .B1(n9796), .B2(n9265), .ZN(n9374)
         );
  XNOR2_X1 U10545 ( .A(n9228), .B(n9227), .ZN(n9377) );
  NAND2_X1 U10546 ( .A1(n9377), .A2(n9275), .ZN(n9236) );
  AOI22_X1 U10547 ( .A1(n9295), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9229), .B2(
        n9293), .ZN(n9230) );
  OAI21_X1 U10548 ( .B1(n9375), .B2(n9279), .A(n9230), .ZN(n9233) );
  OAI211_X1 U10549 ( .C1(n9452), .C2(n4444), .A(n9761), .B(n9231), .ZN(n9373)
         );
  NOR2_X1 U10550 ( .A1(n9373), .A2(n9282), .ZN(n9232) );
  AOI211_X1 U10551 ( .C1(n9286), .C2(n9234), .A(n9233), .B(n9232), .ZN(n9235)
         );
  OAI211_X1 U10552 ( .C1(n9295), .C2(n9374), .A(n9236), .B(n9235), .ZN(
        P1_U3273) );
  XNOR2_X1 U10553 ( .A(n9237), .B(n9240), .ZN(n9382) );
  INV_X1 U10554 ( .A(n9382), .ZN(n9253) );
  OAI21_X1 U10555 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9241) );
  NAND2_X1 U10556 ( .A1(n9241), .A2(n9331), .ZN(n9244) );
  AOI22_X1 U10557 ( .A1(n9364), .A2(n9805), .B1(n9796), .B2(n9242), .ZN(n9243)
         );
  NAND2_X1 U10558 ( .A1(n9244), .A2(n9243), .ZN(n9380) );
  INV_X1 U10559 ( .A(n9245), .ZN(n9456) );
  AOI211_X1 U10560 ( .C1(n9245), .C2(n9256), .A(n9291), .B(n4444), .ZN(n9381)
         );
  NAND2_X1 U10561 ( .A1(n9381), .A2(n9764), .ZN(n9249) );
  INV_X1 U10562 ( .A(n9246), .ZN(n9247) );
  AOI22_X1 U10563 ( .A1(n9295), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9247), .B2(
        n9293), .ZN(n9248) );
  OAI211_X1 U10564 ( .C1(n9456), .C2(n9756), .A(n9249), .B(n9248), .ZN(n9250)
         );
  AOI21_X1 U10565 ( .B1(n9251), .B2(n9380), .A(n9250), .ZN(n9252) );
  OAI21_X1 U10566 ( .B1(n9253), .B2(n9307), .A(n9252), .ZN(P1_U3274) );
  XNOR2_X1 U10567 ( .A(n9254), .B(n9263), .ZN(n9389) );
  INV_X1 U10568 ( .A(n9255), .ZN(n9281) );
  INV_X1 U10569 ( .A(n9256), .ZN(n9257) );
  AOI211_X1 U10570 ( .C1(n9386), .C2(n9281), .A(n9291), .B(n9257), .ZN(n9385)
         );
  INV_X1 U10571 ( .A(n9258), .ZN(n9259) );
  AOI22_X1 U10572 ( .A1(n9295), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9259), .B2(
        n9293), .ZN(n9260) );
  OAI21_X1 U10573 ( .B1(n9261), .B2(n9756), .A(n9260), .ZN(n9268) );
  OAI21_X1 U10574 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9266) );
  AOI222_X1 U10575 ( .A1(n9331), .A2(n9266), .B1(n9265), .B2(n9805), .C1(n9301), .C2(n9796), .ZN(n9388) );
  NOR2_X1 U10576 ( .A1(n9388), .A2(n9295), .ZN(n9267) );
  AOI211_X1 U10577 ( .C1(n9385), .C2(n9764), .A(n9268), .B(n9267), .ZN(n9269)
         );
  OAI21_X1 U10578 ( .B1(n9389), .B2(n9307), .A(n9269), .ZN(P1_U3275) );
  XNOR2_X1 U10579 ( .A(n9270), .B(n9273), .ZN(n9272) );
  AOI22_X1 U10580 ( .A1(n9272), .A2(n9331), .B1(n9796), .B2(n9271), .ZN(n9391)
         );
  XNOR2_X1 U10581 ( .A(n9274), .B(n9273), .ZN(n9394) );
  NAND2_X1 U10582 ( .A1(n9394), .A2(n9275), .ZN(n9288) );
  INV_X1 U10583 ( .A(n9276), .ZN(n9277) );
  AOI22_X1 U10584 ( .A1(n9295), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9277), .B2(
        n9293), .ZN(n9278) );
  OAI21_X1 U10585 ( .B1(n9279), .B2(n9392), .A(n9278), .ZN(n9284) );
  INV_X1 U10586 ( .A(n9285), .ZN(n9461) );
  OAI211_X1 U10587 ( .C1(n9461), .C2(n4652), .A(n9281), .B(n9761), .ZN(n9390)
         );
  NOR2_X1 U10588 ( .A1(n9390), .A2(n9282), .ZN(n9283) );
  AOI211_X1 U10589 ( .C1(n9286), .C2(n9285), .A(n9284), .B(n9283), .ZN(n9287)
         );
  OAI211_X1 U10590 ( .C1(n9295), .C2(n9391), .A(n9288), .B(n9287), .ZN(
        P1_U3276) );
  XNOR2_X1 U10591 ( .A(n9289), .B(n9290), .ZN(n9401) );
  AOI211_X1 U10592 ( .C1(n9398), .C2(n9292), .A(n9291), .B(n4652), .ZN(n9397)
         );
  INV_X1 U10593 ( .A(n9398), .ZN(n9297) );
  AOI22_X1 U10594 ( .A1(n9295), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9294), .B2(
        n9293), .ZN(n9296) );
  OAI21_X1 U10595 ( .B1(n9297), .B2(n9756), .A(n9296), .ZN(n9305) );
  OAI21_X1 U10596 ( .B1(n9300), .B2(n9299), .A(n9298), .ZN(n9303) );
  AOI222_X1 U10597 ( .A1(n9331), .A2(n9303), .B1(n9302), .B2(n9796), .C1(n9301), .C2(n9805), .ZN(n9400) );
  NOR2_X1 U10598 ( .A1(n9400), .A2(n9295), .ZN(n9304) );
  AOI211_X1 U10599 ( .C1(n9397), .C2(n9764), .A(n9305), .B(n9304), .ZN(n9306)
         );
  OAI21_X1 U10600 ( .B1(n9307), .B2(n9401), .A(n9306), .ZN(P1_U3277) );
  AND2_X1 U10601 ( .A1(n9308), .A2(n9311), .ZN(n9414) );
  MUX2_X1 U10602 ( .A(n9309), .B(n9414), .S(n9826), .Z(n9310) );
  OAI21_X1 U10603 ( .B1(n9417), .B2(n9406), .A(n9310), .ZN(P1_U3553) );
  MUX2_X1 U10604 ( .A(n9313), .B(n9418), .S(n9826), .Z(n9314) );
  OAI21_X1 U10605 ( .B1(n9421), .B2(n9406), .A(n9314), .ZN(P1_U3552) );
  OAI22_X1 U10606 ( .A1(n9317), .A2(n9740), .B1(n9316), .B2(n9738), .ZN(n9318)
         );
  INV_X1 U10607 ( .A(n9318), .ZN(n9319) );
  AND2_X1 U10608 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  OAI211_X1 U10609 ( .C1(n9746), .C2(n9323), .A(n9322), .B(n9321), .ZN(n9422)
         );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9422), .S(n9826), .Z(n9324) );
  INV_X1 U10611 ( .A(n9324), .ZN(n9325) );
  OAI21_X1 U10612 ( .B1(n9425), .B2(n9406), .A(n9325), .ZN(P1_U3549) );
  OAI22_X1 U10613 ( .A1(n9327), .A2(n9740), .B1(n9326), .B2(n9738), .ZN(n9329)
         );
  AOI211_X1 U10614 ( .C1(n9331), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9332)
         );
  INV_X1 U10615 ( .A(n9332), .ZN(n9333) );
  AOI21_X1 U10616 ( .B1(n9334), .B2(n9812), .A(n9333), .ZN(n9427) );
  MUX2_X1 U10617 ( .A(n9427), .B(n9335), .S(n9824), .Z(n9336) );
  OAI21_X1 U10618 ( .B1(n9429), .B2(n9406), .A(n9336), .ZN(P1_U3548) );
  AOI211_X1 U10619 ( .C1(n9339), .C2(n9812), .A(n9338), .B(n9337), .ZN(n9430)
         );
  MUX2_X1 U10620 ( .A(n9340), .B(n9430), .S(n9826), .Z(n9341) );
  OAI21_X1 U10621 ( .B1(n5883), .B2(n9406), .A(n9341), .ZN(P1_U3547) );
  AOI211_X1 U10622 ( .C1(n9344), .C2(n9812), .A(n9343), .B(n9342), .ZN(n9433)
         );
  MUX2_X1 U10623 ( .A(n9345), .B(n9433), .S(n9826), .Z(n9346) );
  OAI21_X1 U10624 ( .B1(n9436), .B2(n9406), .A(n9346), .ZN(P1_U3546) );
  AOI22_X1 U10625 ( .A1(n9347), .A2(n9805), .B1(n9796), .B2(n9365), .ZN(n9349)
         );
  OAI211_X1 U10626 ( .C1(n9350), .C2(n9746), .A(n9349), .B(n9348), .ZN(n9351)
         );
  AOI21_X1 U10627 ( .B1(n9352), .B2(n9812), .A(n9351), .ZN(n9437) );
  MUX2_X1 U10628 ( .A(n9353), .B(n9437), .S(n9826), .Z(n9354) );
  OAI21_X1 U10629 ( .B1(n9440), .B2(n9406), .A(n9354), .ZN(P1_U3545) );
  AOI22_X1 U10630 ( .A1(n9356), .A2(n9805), .B1(n9796), .B2(n9355), .ZN(n9358)
         );
  OAI211_X1 U10631 ( .C1(n9359), .C2(n9746), .A(n9358), .B(n9357), .ZN(n9360)
         );
  AOI21_X1 U10632 ( .B1(n9361), .B2(n9812), .A(n9360), .ZN(n9441) );
  MUX2_X1 U10633 ( .A(n9362), .B(n9441), .S(n9826), .Z(n9363) );
  OAI21_X1 U10634 ( .B1(n9444), .B2(n9406), .A(n9363), .ZN(P1_U3544) );
  AOI22_X1 U10635 ( .A1(n9365), .A2(n9805), .B1(n9796), .B2(n9364), .ZN(n9367)
         );
  OAI211_X1 U10636 ( .C1(n9368), .C2(n9746), .A(n9367), .B(n9366), .ZN(n9369)
         );
  AOI21_X1 U10637 ( .B1(n9370), .B2(n9812), .A(n9369), .ZN(n9445) );
  MUX2_X1 U10638 ( .A(n9371), .B(n9445), .S(n9826), .Z(n9372) );
  OAI21_X1 U10639 ( .B1(n9448), .B2(n9406), .A(n9372), .ZN(P1_U3543) );
  OAI211_X1 U10640 ( .C1(n9375), .C2(n9740), .A(n9374), .B(n9373), .ZN(n9376)
         );
  AOI21_X1 U10641 ( .B1(n9377), .B2(n9812), .A(n9376), .ZN(n9449) );
  MUX2_X1 U10642 ( .A(n9378), .B(n9449), .S(n9826), .Z(n9379) );
  OAI21_X1 U10643 ( .B1(n9452), .B2(n9406), .A(n9379), .ZN(P1_U3542) );
  AOI211_X1 U10644 ( .C1(n9382), .C2(n9812), .A(n9381), .B(n9380), .ZN(n9453)
         );
  MUX2_X1 U10645 ( .A(n9383), .B(n9453), .S(n9826), .Z(n9384) );
  OAI21_X1 U10646 ( .B1(n9456), .B2(n9406), .A(n9384), .ZN(P1_U3541) );
  AOI21_X1 U10647 ( .B1(n9806), .B2(n9386), .A(n9385), .ZN(n9387) );
  OAI211_X1 U10648 ( .C1(n9389), .C2(n9773), .A(n9388), .B(n9387), .ZN(n9457)
         );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9457), .S(n9826), .Z(
        P1_U3540) );
  OAI211_X1 U10650 ( .C1(n9392), .C2(n9740), .A(n9391), .B(n9390), .ZN(n9393)
         );
  AOI21_X1 U10651 ( .B1(n9394), .B2(n9812), .A(n9393), .ZN(n9458) );
  MUX2_X1 U10652 ( .A(n9395), .B(n9458), .S(n9826), .Z(n9396) );
  OAI21_X1 U10653 ( .B1(n9461), .B2(n9406), .A(n9396), .ZN(P1_U3539) );
  AOI21_X1 U10654 ( .B1(n9806), .B2(n9398), .A(n9397), .ZN(n9399) );
  OAI211_X1 U10655 ( .C1(n9401), .C2(n9773), .A(n9400), .B(n9399), .ZN(n9462)
         );
  MUX2_X1 U10656 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9462), .S(n9826), .Z(
        P1_U3538) );
  AOI211_X1 U10657 ( .C1(n9404), .C2(n9812), .A(n9403), .B(n9402), .ZN(n9463)
         );
  MUX2_X1 U10658 ( .A(n9682), .B(n9463), .S(n9826), .Z(n9405) );
  OAI21_X1 U10659 ( .B1(n9467), .B2(n9406), .A(n9405), .ZN(P1_U3537) );
  INV_X1 U10660 ( .A(n9806), .ZN(n9790) );
  OAI211_X1 U10661 ( .C1(n9409), .C2(n9790), .A(n9408), .B(n9407), .ZN(n9410)
         );
  AOI21_X1 U10662 ( .B1(n9812), .B2(n9411), .A(n9410), .ZN(n9469) );
  NAND2_X1 U10663 ( .A1(n9824), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9412) );
  OAI21_X1 U10664 ( .B1(n9469), .B2(n9824), .A(n9412), .ZN(P1_U3536) );
  MUX2_X1 U10665 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9413), .S(n9826), .Z(
        P1_U3522) );
  INV_X1 U10666 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9415) );
  MUX2_X1 U10667 ( .A(n9415), .B(n9414), .S(n9816), .Z(n9416) );
  OAI21_X1 U10668 ( .B1(n9417), .B2(n9466), .A(n9416), .ZN(P1_U3521) );
  MUX2_X1 U10669 ( .A(n9419), .B(n9418), .S(n9816), .Z(n9420) );
  OAI21_X1 U10670 ( .B1(n9421), .B2(n9466), .A(n9420), .ZN(P1_U3520) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9422), .S(n9816), .Z(n9423) );
  INV_X1 U10672 ( .A(n9423), .ZN(n9424) );
  OAI21_X1 U10673 ( .B1(n9425), .B2(n9466), .A(n9424), .ZN(P1_U3517) );
  INV_X1 U10674 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9426) );
  MUX2_X1 U10675 ( .A(n9427), .B(n9426), .S(n9814), .Z(n9428) );
  OAI21_X1 U10676 ( .B1(n9429), .B2(n9466), .A(n9428), .ZN(P1_U3516) );
  INV_X1 U10677 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9431) );
  MUX2_X1 U10678 ( .A(n9431), .B(n9430), .S(n9816), .Z(n9432) );
  OAI21_X1 U10679 ( .B1(n5883), .B2(n9466), .A(n9432), .ZN(P1_U3515) );
  INV_X1 U10680 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9434) );
  MUX2_X1 U10681 ( .A(n9434), .B(n9433), .S(n9816), .Z(n9435) );
  OAI21_X1 U10682 ( .B1(n9436), .B2(n9466), .A(n9435), .ZN(P1_U3514) );
  INV_X1 U10683 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9438) );
  MUX2_X1 U10684 ( .A(n9438), .B(n9437), .S(n9816), .Z(n9439) );
  OAI21_X1 U10685 ( .B1(n9440), .B2(n9466), .A(n9439), .ZN(P1_U3513) );
  INV_X1 U10686 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9442) );
  MUX2_X1 U10687 ( .A(n9442), .B(n9441), .S(n9816), .Z(n9443) );
  OAI21_X1 U10688 ( .B1(n9444), .B2(n9466), .A(n9443), .ZN(P1_U3512) );
  INV_X1 U10689 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9446) );
  MUX2_X1 U10690 ( .A(n9446), .B(n9445), .S(n9816), .Z(n9447) );
  OAI21_X1 U10691 ( .B1(n9448), .B2(n9466), .A(n9447), .ZN(P1_U3511) );
  INV_X1 U10692 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9450) );
  MUX2_X1 U10693 ( .A(n9450), .B(n9449), .S(n9816), .Z(n9451) );
  OAI21_X1 U10694 ( .B1(n9452), .B2(n9466), .A(n9451), .ZN(P1_U3510) );
  INV_X1 U10695 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9454) );
  MUX2_X1 U10696 ( .A(n9454), .B(n9453), .S(n9816), .Z(n9455) );
  OAI21_X1 U10697 ( .B1(n9456), .B2(n9466), .A(n9455), .ZN(P1_U3509) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9457), .S(n9816), .Z(
        P1_U3507) );
  MUX2_X1 U10699 ( .A(n9459), .B(n9458), .S(n9816), .Z(n9460) );
  OAI21_X1 U10700 ( .B1(n9461), .B2(n9466), .A(n9460), .ZN(P1_U3504) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9462), .S(n9816), .Z(
        P1_U3501) );
  INV_X1 U10702 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9464) );
  MUX2_X1 U10703 ( .A(n9464), .B(n9463), .S(n9816), .Z(n9465) );
  OAI21_X1 U10704 ( .B1(n9467), .B2(n9466), .A(n9465), .ZN(P1_U3498) );
  NAND2_X1 U10705 ( .A1(n9814), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9468) );
  OAI21_X1 U10706 ( .B1(n9469), .B2(n9814), .A(n9468), .ZN(P1_U3495) );
  MUX2_X1 U10707 ( .A(n9470), .B(P1_D_REG_0__SCAN_IN), .S(n9768), .Z(P1_U3439)
         );
  NOR4_X1 U10708 ( .A1(n9471), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n4945), .ZN(n9472) );
  AOI21_X1 U10709 ( .B1(n9479), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9472), .ZN(
        n9473) );
  OAI21_X1 U10710 ( .B1(n9474), .B2(n6469), .A(n9473), .ZN(P1_U3324) );
  AOI22_X1 U10711 ( .A1(n9476), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9475), .ZN(n9477) );
  OAI21_X1 U10712 ( .B1(n9478), .B2(n6469), .A(n9477), .ZN(P1_U3325) );
  AOI22_X1 U10713 ( .A1(n9480), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9479), .ZN(n9481) );
  OAI21_X1 U10714 ( .B1(n9482), .B2(n6469), .A(n9481), .ZN(P1_U3326) );
  MUX2_X1 U10715 ( .A(n9483), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10716 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U10717 ( .A1(n9485), .A2(n9484), .ZN(n9488) );
  INV_X1 U10718 ( .A(n9486), .ZN(n9487) );
  NAND2_X1 U10719 ( .A1(n9488), .A2(n9487), .ZN(n9496) );
  NAND2_X1 U10720 ( .A1(n9724), .A2(n9489), .ZN(n9495) );
  AOI21_X1 U10721 ( .B1(n9492), .B2(n9491), .A(n9490), .ZN(n9493) );
  NAND2_X1 U10722 ( .A1(n9717), .A2(n9493), .ZN(n9494) );
  OAI211_X1 U10723 ( .C1(n9721), .C2(n9496), .A(n9495), .B(n9494), .ZN(n9497)
         );
  INV_X1 U10724 ( .A(n9497), .ZN(n9499) );
  OAI211_X1 U10725 ( .C1(n9732), .C2(n9500), .A(n9499), .B(n9498), .ZN(
        P1_U3253) );
  INV_X1 U10726 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9515) );
  OAI21_X1 U10727 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9511) );
  INV_X1 U10728 ( .A(n9504), .ZN(n9505) );
  OAI211_X1 U10729 ( .C1(n9507), .C2(n9506), .A(n9717), .B(n9505), .ZN(n9510)
         );
  NAND2_X1 U10730 ( .A1(n9724), .A2(n9508), .ZN(n9509) );
  OAI211_X1 U10731 ( .C1(n9511), .C2(n9721), .A(n9510), .B(n9509), .ZN(n9512)
         );
  INV_X1 U10732 ( .A(n9512), .ZN(n9514) );
  OAI211_X1 U10733 ( .C1(n9732), .C2(n9515), .A(n9514), .B(n9513), .ZN(
        P1_U3250) );
  INV_X1 U10734 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U10735 ( .A1(n9517), .A2(n9516), .ZN(n9520) );
  INV_X1 U10736 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U10737 ( .A1(n9520), .A2(n9519), .ZN(n9528) );
  NAND2_X1 U10738 ( .A1(n9724), .A2(n9521), .ZN(n9527) );
  AOI21_X1 U10739 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9525) );
  NAND2_X1 U10740 ( .A1(n9717), .A2(n9525), .ZN(n9526) );
  OAI211_X1 U10741 ( .C1(n9721), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9529)
         );
  INV_X1 U10742 ( .A(n9529), .ZN(n9531) );
  OAI211_X1 U10743 ( .C1(n9732), .C2(n9532), .A(n9531), .B(n9530), .ZN(
        P1_U3251) );
  INV_X1 U10744 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9548) );
  OAI21_X1 U10745 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9536) );
  INV_X1 U10746 ( .A(n9536), .ZN(n9544) );
  NAND2_X1 U10747 ( .A1(n9724), .A2(n9537), .ZN(n9543) );
  OAI21_X1 U10748 ( .B1(n9540), .B2(n9539), .A(n9538), .ZN(n9541) );
  NAND2_X1 U10749 ( .A1(n9717), .A2(n9541), .ZN(n9542) );
  OAI211_X1 U10750 ( .C1(n9721), .C2(n9544), .A(n9543), .B(n9542), .ZN(n9545)
         );
  INV_X1 U10751 ( .A(n9545), .ZN(n9547) );
  OAI211_X1 U10752 ( .C1(n9732), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3252) );
  XNOR2_X1 U10753 ( .A(n9549), .B(n9555), .ZN(n9567) );
  AND2_X1 U10754 ( .A1(n9550), .A2(n9985), .ZN(n9566) );
  NAND2_X1 U10755 ( .A1(n9566), .A2(n9551), .ZN(n9552) );
  OAI21_X1 U10756 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9560) );
  XNOR2_X1 U10757 ( .A(n9556), .B(n9555), .ZN(n9557) );
  OAI222_X1 U10758 ( .A1(n9920), .A2(n9559), .B1(n9922), .B2(n9558), .C1(n9928), .C2(n9557), .ZN(n9565) );
  AOI211_X1 U10759 ( .C1(n9567), .C2(n9561), .A(n9560), .B(n9565), .ZN(n9563)
         );
  AOI22_X1 U10760 ( .A1(n9936), .A2(n9564), .B1(n9563), .B2(n9562), .ZN(
        P2_U3220) );
  AOI211_X1 U10761 ( .C1(n9567), .C2(n9980), .A(n9566), .B(n9565), .ZN(n9569)
         );
  AOI22_X1 U10762 ( .A1(n10003), .A2(n9569), .B1(n9568), .B2(n10004), .ZN(
        P2_U3472) );
  INV_X1 U10763 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9570) );
  AOI22_X1 U10764 ( .A1(n9988), .A2(n9570), .B1(n9569), .B2(n9986), .ZN(
        P2_U3429) );
  XNOR2_X1 U10765 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10766 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U10767 ( .A1(n4358), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9571) );
  INV_X1 U10768 ( .A(n9571), .ZN(n9574) );
  OR2_X1 U10769 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  MUX2_X1 U10770 ( .A(n9574), .B(n9573), .S(P1_IR_REG_0__SCAN_IN), .Z(n9576)
         );
  NAND2_X1 U10771 ( .A1(n9576), .A2(n9575), .ZN(n9578) );
  AOI22_X1 U10772 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9593), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9577) );
  OAI21_X1 U10773 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(P1_U3243) );
  OAI21_X1 U10774 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9590) );
  INV_X1 U10775 ( .A(n9583), .ZN(n9584) );
  OAI211_X1 U10776 ( .C1(n9586), .C2(n9585), .A(n9717), .B(n9584), .ZN(n9589)
         );
  NAND2_X1 U10777 ( .A1(n9724), .A2(n9587), .ZN(n9588) );
  OAI211_X1 U10778 ( .C1(n9721), .C2(n9590), .A(n9589), .B(n9588), .ZN(n9591)
         );
  INV_X1 U10779 ( .A(n9591), .ZN(n9597) );
  AOI21_X1 U10780 ( .B1(n9593), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9592), .ZN(
        n9594) );
  AND2_X1 U10781 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  NAND2_X1 U10782 ( .A1(n9597), .A2(n9596), .ZN(P1_U3247) );
  INV_X1 U10783 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U10784 ( .A1(n9599), .A2(n9598), .ZN(n9601) );
  NAND2_X1 U10785 ( .A1(n9601), .A2(n9600), .ZN(n9609) );
  NAND2_X1 U10786 ( .A1(n9724), .A2(n9602), .ZN(n9608) );
  AOI21_X1 U10787 ( .B1(n9605), .B2(n9604), .A(n9603), .ZN(n9606) );
  NAND2_X1 U10788 ( .A1(n9717), .A2(n9606), .ZN(n9607) );
  OAI211_X1 U10789 ( .C1(n9721), .C2(n9609), .A(n9608), .B(n9607), .ZN(n9610)
         );
  INV_X1 U10790 ( .A(n9610), .ZN(n9612) );
  OAI211_X1 U10791 ( .C1(n9732), .C2(n9613), .A(n9612), .B(n9611), .ZN(
        P1_U3248) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U10793 ( .A1(n9615), .A2(n9614), .ZN(n9618) );
  INV_X1 U10794 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U10795 ( .A1(n9618), .A2(n9617), .ZN(n9626) );
  NAND2_X1 U10796 ( .A1(n9724), .A2(n9619), .ZN(n9625) );
  AOI21_X1 U10797 ( .B1(n9622), .B2(n9621), .A(n9620), .ZN(n9623) );
  NAND2_X1 U10798 ( .A1(n9717), .A2(n9623), .ZN(n9624) );
  OAI211_X1 U10799 ( .C1(n9721), .C2(n9626), .A(n9625), .B(n9624), .ZN(n9627)
         );
  INV_X1 U10800 ( .A(n9627), .ZN(n9629) );
  OAI211_X1 U10801 ( .C1(n9732), .C2(n9630), .A(n9629), .B(n9628), .ZN(
        P1_U3254) );
  INV_X1 U10802 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9646) );
  OAI21_X1 U10803 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9634) );
  INV_X1 U10804 ( .A(n9634), .ZN(n9642) );
  NAND2_X1 U10805 ( .A1(n9724), .A2(n9635), .ZN(n9641) );
  OAI21_X1 U10806 ( .B1(n9638), .B2(n9637), .A(n9636), .ZN(n9639) );
  NAND2_X1 U10807 ( .A1(n9717), .A2(n9639), .ZN(n9640) );
  OAI211_X1 U10808 ( .C1(n9721), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9643)
         );
  INV_X1 U10809 ( .A(n9643), .ZN(n9645) );
  OAI211_X1 U10810 ( .C1(n9732), .C2(n9646), .A(n9645), .B(n9644), .ZN(
        P1_U3255) );
  INV_X1 U10811 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U10812 ( .A1(n9648), .A2(n9647), .ZN(n9651) );
  INV_X1 U10813 ( .A(n9649), .ZN(n9650) );
  NAND2_X1 U10814 ( .A1(n9651), .A2(n9650), .ZN(n9659) );
  NAND2_X1 U10815 ( .A1(n9724), .A2(n9652), .ZN(n9658) );
  AOI21_X1 U10816 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9656) );
  NAND2_X1 U10817 ( .A1(n9717), .A2(n9656), .ZN(n9657) );
  OAI211_X1 U10818 ( .C1(n9721), .C2(n9659), .A(n9658), .B(n9657), .ZN(n9660)
         );
  INV_X1 U10819 ( .A(n9660), .ZN(n9662) );
  OAI211_X1 U10820 ( .C1(n9732), .C2(n9663), .A(n9662), .B(n9661), .ZN(
        P1_U3256) );
  INV_X1 U10821 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U10822 ( .A1(n9665), .A2(n9664), .ZN(n9668) );
  INV_X1 U10823 ( .A(n9666), .ZN(n9667) );
  NAND2_X1 U10824 ( .A1(n9668), .A2(n9667), .ZN(n9676) );
  NAND2_X1 U10825 ( .A1(n9724), .A2(n9669), .ZN(n9675) );
  AOI21_X1 U10826 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9673) );
  NAND2_X1 U10827 ( .A1(n9717), .A2(n9673), .ZN(n9674) );
  OAI211_X1 U10828 ( .C1(n9721), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9677)
         );
  INV_X1 U10829 ( .A(n9677), .ZN(n9679) );
  OAI211_X1 U10830 ( .C1(n9732), .C2(n9680), .A(n9679), .B(n9678), .ZN(
        P1_U3257) );
  INV_X1 U10831 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9691) );
  AOI211_X1 U10832 ( .C1(n9683), .C2(n9682), .A(n9681), .B(n9721), .ZN(n9687)
         );
  INV_X1 U10833 ( .A(n9717), .ZN(n9692) );
  AOI211_X1 U10834 ( .C1(n9685), .C2(n7444), .A(n9684), .B(n9692), .ZN(n9686)
         );
  AOI211_X1 U10835 ( .C1(n9724), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9690)
         );
  OAI211_X1 U10836 ( .C1(n9732), .C2(n9691), .A(n9690), .B(n9689), .ZN(
        P1_U3258) );
  INV_X1 U10837 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10012) );
  AOI21_X1 U10838 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9702) );
  XOR2_X1 U10839 ( .A(n9696), .B(n9695), .Z(n9699) );
  INV_X1 U10840 ( .A(n9724), .ZN(n9697) );
  OAI22_X1 U10841 ( .A1(n9699), .A2(n9721), .B1(n9698), .B2(n9697), .ZN(n9700)
         );
  AOI21_X1 U10842 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9704) );
  OAI211_X1 U10843 ( .C1(n9732), .C2(n10012), .A(n9704), .B(n9703), .ZN(
        P1_U3259) );
  INV_X1 U10844 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9716) );
  OAI21_X1 U10845 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9713) );
  XNOR2_X1 U10846 ( .A(n9709), .B(n9708), .ZN(n9711) );
  AOI222_X1 U10847 ( .A1(n9713), .A2(n9717), .B1(n9712), .B2(n9711), .C1(n9710), .C2(n9724), .ZN(n9715) );
  OAI211_X1 U10848 ( .C1(n9732), .C2(n9716), .A(n9715), .B(n9714), .ZN(
        P1_U3260) );
  INV_X1 U10849 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10246) );
  OAI211_X1 U10850 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9729)
         );
  AOI21_X1 U10851 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9727) );
  AOI22_X1 U10852 ( .A1(n9727), .A2(n9726), .B1(n9725), .B2(n9724), .ZN(n9728)
         );
  AND2_X1 U10853 ( .A1(n9729), .A2(n9728), .ZN(n9731) );
  OAI211_X1 U10854 ( .C1(n9732), .C2(n10246), .A(n9731), .B(n9730), .ZN(
        P1_U3261) );
  INV_X1 U10855 ( .A(n9733), .ZN(n9734) );
  NOR2_X1 U10856 ( .A1(n9735), .A2(n9734), .ZN(n9748) );
  XNOR2_X1 U10857 ( .A(n9736), .B(n9748), .ZN(n9786) );
  INV_X1 U10858 ( .A(n9737), .ZN(n9751) );
  OAI22_X1 U10859 ( .A1(n9741), .A2(n9740), .B1(n9739), .B2(n9738), .ZN(n9750)
         );
  INV_X1 U10860 ( .A(n9742), .ZN(n9743) );
  NOR2_X1 U10861 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  AOI211_X1 U10862 ( .C1(n9748), .C2(n9747), .A(n9746), .B(n9745), .ZN(n9749)
         );
  AOI211_X1 U10863 ( .C1(n9786), .C2(n9751), .A(n9750), .B(n9749), .ZN(n9783)
         );
  NOR2_X1 U10864 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  AOI21_X1 U10865 ( .B1(n9295), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9754), .ZN(
        n9755) );
  OAI21_X1 U10866 ( .B1(n9756), .B2(n4642), .A(n9755), .ZN(n9757) );
  INV_X1 U10867 ( .A(n9757), .ZN(n9767) );
  INV_X1 U10868 ( .A(n9758), .ZN(n9765) );
  INV_X1 U10869 ( .A(n9759), .ZN(n9762) );
  OAI211_X1 U10870 ( .C1(n9762), .C2(n4642), .A(n9761), .B(n9760), .ZN(n9782)
         );
  INV_X1 U10871 ( .A(n9782), .ZN(n9763) );
  AOI22_X1 U10872 ( .A1(n9786), .A2(n9765), .B1(n9764), .B2(n9763), .ZN(n9766)
         );
  OAI211_X1 U10873 ( .C1(n9295), .C2(n9783), .A(n9767), .B(n9766), .ZN(
        P1_U3285) );
  AND2_X1 U10874 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9768), .ZN(P1_U3294) );
  AND2_X1 U10875 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9768), .ZN(P1_U3295) );
  AND2_X1 U10876 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9768), .ZN(P1_U3296) );
  AND2_X1 U10877 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9768), .ZN(P1_U3297) );
  AND2_X1 U10878 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9768), .ZN(P1_U3298) );
  AND2_X1 U10879 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9768), .ZN(P1_U3299) );
  AND2_X1 U10880 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9768), .ZN(P1_U3300) );
  AND2_X1 U10881 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9768), .ZN(P1_U3301) );
  AND2_X1 U10882 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9768), .ZN(P1_U3302) );
  AND2_X1 U10883 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9768), .ZN(P1_U3303) );
  AND2_X1 U10884 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9768), .ZN(P1_U3304) );
  AND2_X1 U10885 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9768), .ZN(P1_U3305) );
  AND2_X1 U10886 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9768), .ZN(P1_U3306) );
  AND2_X1 U10887 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9768), .ZN(P1_U3307) );
  AND2_X1 U10888 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9768), .ZN(P1_U3308) );
  AND2_X1 U10889 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9768), .ZN(P1_U3309) );
  AND2_X1 U10890 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9768), .ZN(P1_U3310) );
  AND2_X1 U10891 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9768), .ZN(P1_U3311) );
  AND2_X1 U10892 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9768), .ZN(P1_U3312) );
  AND2_X1 U10893 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9768), .ZN(P1_U3313) );
  AND2_X1 U10894 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9768), .ZN(P1_U3314) );
  AND2_X1 U10895 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9768), .ZN(P1_U3315) );
  AND2_X1 U10896 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9768), .ZN(P1_U3316) );
  AND2_X1 U10897 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9768), .ZN(P1_U3317) );
  AND2_X1 U10898 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9768), .ZN(P1_U3318) );
  AND2_X1 U10899 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9768), .ZN(P1_U3319) );
  AND2_X1 U10900 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9768), .ZN(P1_U3320) );
  AND2_X1 U10901 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9768), .ZN(P1_U3321) );
  AND2_X1 U10902 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9768), .ZN(P1_U3322) );
  AND2_X1 U10903 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9768), .ZN(P1_U3323) );
  AOI21_X1 U10904 ( .B1(n9806), .B2(n9770), .A(n9769), .ZN(n9771) );
  OAI211_X1 U10905 ( .C1(n9774), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9775)
         );
  INV_X1 U10906 ( .A(n9775), .ZN(n9818) );
  AOI22_X1 U10907 ( .A1(n9816), .A2(n9818), .B1(n5087), .B2(n9814), .ZN(
        P1_U3465) );
  OAI211_X1 U10908 ( .C1(n9778), .C2(n9790), .A(n9777), .B(n9776), .ZN(n9779)
         );
  AOI21_X1 U10909 ( .B1(n9812), .B2(n9780), .A(n9779), .ZN(n9819) );
  INV_X1 U10910 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10911 ( .A1(n9816), .A2(n9819), .B1(n9781), .B2(n9814), .ZN(
        P1_U3471) );
  OAI21_X1 U10912 ( .B1(n4642), .B2(n9790), .A(n9782), .ZN(n9785) );
  INV_X1 U10913 ( .A(n9783), .ZN(n9784) );
  AOI211_X1 U10914 ( .C1(n9787), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9820)
         );
  AOI22_X1 U10915 ( .A1(n9816), .A2(n9820), .B1(n5219), .B2(n9814), .ZN(
        P1_U3477) );
  OAI21_X1 U10916 ( .B1(n4641), .B2(n9790), .A(n9789), .ZN(n9792) );
  AOI211_X1 U10917 ( .C1(n9812), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9821)
         );
  INV_X1 U10918 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U10919 ( .A1(n9816), .A2(n9821), .B1(n9794), .B2(n9814), .ZN(
        P1_U3480) );
  AOI22_X1 U10920 ( .A1(n9797), .A2(n9806), .B1(n9796), .B2(n9795), .ZN(n9799)
         );
  NAND3_X1 U10921 ( .A1(n9800), .A2(n9799), .A3(n9798), .ZN(n9801) );
  AOI21_X1 U10922 ( .B1(n9802), .B2(n9812), .A(n9801), .ZN(n9823) );
  INV_X1 U10923 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9803) );
  AOI22_X1 U10924 ( .A1(n9816), .A2(n9823), .B1(n9803), .B2(n9814), .ZN(
        P1_U3483) );
  AOI22_X1 U10925 ( .A1(n9807), .A2(n9806), .B1(n9805), .B2(n9804), .ZN(n9809)
         );
  NAND3_X1 U10926 ( .A1(n9810), .A2(n9809), .A3(n9808), .ZN(n9811) );
  AOI21_X1 U10927 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9825) );
  INV_X1 U10928 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10929 ( .A1(n9816), .A2(n9825), .B1(n9815), .B2(n9814), .ZN(
        P1_U3489) );
  AOI22_X1 U10930 ( .A1(n9826), .A2(n9818), .B1(n9817), .B2(n9824), .ZN(
        P1_U3526) );
  AOI22_X1 U10931 ( .A1(n9826), .A2(n9819), .B1(n7849), .B2(n9824), .ZN(
        P1_U3528) );
  AOI22_X1 U10932 ( .A1(n9826), .A2(n9820), .B1(n7853), .B2(n9824), .ZN(
        P1_U3530) );
  AOI22_X1 U10933 ( .A1(n9826), .A2(n9821), .B1(n7839), .B2(n9824), .ZN(
        P1_U3531) );
  INV_X1 U10934 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10935 ( .A1(n9826), .A2(n9823), .B1(n9822), .B2(n9824), .ZN(
        P1_U3532) );
  AOI22_X1 U10936 ( .A1(n9826), .A2(n9825), .B1(n7855), .B2(n9824), .ZN(
        P1_U3534) );
  AOI22_X1 U10937 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9900), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9832) );
  XNOR2_X1 U10938 ( .A(n9828), .B(P2_IR_REG_0__SCAN_IN), .ZN(n9829) );
  OAI21_X1 U10939 ( .B1(n9830), .B2(n6411), .A(n9829), .ZN(n9831) );
  OAI211_X1 U10940 ( .C1(n9871), .C2(n9833), .A(n9832), .B(n9831), .ZN(
        P2_U3182) );
  OAI21_X1 U10941 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9837) );
  NAND2_X1 U10942 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  OAI21_X1 U10943 ( .B1(n9871), .B2(n4350), .A(n9839), .ZN(n9843) );
  INV_X1 U10944 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9840) );
  NOR2_X1 U10945 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  NOR2_X1 U10946 ( .A1(n9843), .A2(n9842), .ZN(n9849) );
  OAI21_X1 U10947 ( .B1(n9845), .B2(n9844), .A(n6411), .ZN(n9846) );
  OR2_X1 U10948 ( .A1(n9847), .A2(n9846), .ZN(n9848) );
  AND2_X1 U10949 ( .A1(n9849), .A2(n9848), .ZN(n9855) );
  OAI21_X1 U10950 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(n9853) );
  NAND2_X1 U10951 ( .A1(n8489), .A2(n9853), .ZN(n9854) );
  OAI211_X1 U10952 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6719), .A(n9855), .B(
        n9854), .ZN(P2_U3184) );
  AOI211_X1 U10953 ( .C1(n9859), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9867)
         );
  AOI21_X1 U10954 ( .B1(n9993), .B2(n9861), .A(n9860), .ZN(n9865) );
  AOI21_X1 U10955 ( .B1(n6016), .B2(n9863), .A(n9862), .ZN(n9864) );
  OAI22_X1 U10956 ( .A1(n9909), .A2(n9865), .B1(n9864), .B2(n9905), .ZN(n9866)
         );
  AOI211_X1 U10957 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9900), .A(n9867), .B(
        n9866), .ZN(n9869) );
  OAI211_X1 U10958 ( .C1(n9871), .C2(n9870), .A(n9869), .B(n9868), .ZN(
        P2_U3187) );
  AOI21_X1 U10959 ( .B1(n9896), .B2(n9873), .A(n9872), .ZN(n9892) );
  OAI21_X1 U10960 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(n9877) );
  AOI22_X1 U10961 ( .A1(n9900), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n9877), .B2(
        n6411), .ZN(n9891) );
  INV_X1 U10962 ( .A(n9878), .ZN(n9879) );
  AOI21_X1 U10963 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n9882) );
  OR2_X1 U10964 ( .A1(n9882), .A2(n9905), .ZN(n9890) );
  INV_X1 U10965 ( .A(n9883), .ZN(n9887) );
  INV_X1 U10966 ( .A(n9884), .ZN(n9886) );
  OAI21_X1 U10967 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9888) );
  NAND2_X1 U10968 ( .A1(n9888), .A2(n8489), .ZN(n9889) );
  NAND4_X1 U10969 ( .A1(n9892), .A2(n9891), .A3(n9890), .A4(n9889), .ZN(
        P2_U3188) );
  INV_X1 U10970 ( .A(n9893), .ZN(n9895) );
  AOI21_X1 U10971 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9914) );
  OAI21_X1 U10972 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9901) );
  AOI22_X1 U10973 ( .A1(n9901), .A2(n6411), .B1(n9900), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n9913) );
  INV_X1 U10974 ( .A(n9902), .ZN(n9903) );
  AOI21_X1 U10975 ( .B1(n9904), .B2(n9903), .A(n4458), .ZN(n9906) );
  OR2_X1 U10976 ( .A1(n9906), .A2(n9905), .ZN(n9912) );
  AOI21_X1 U10977 ( .B1(n9908), .B2(n9907), .A(n4457), .ZN(n9910) );
  OR2_X1 U10978 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  NAND4_X1 U10979 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(
        P2_U3190) );
  XNOR2_X1 U10980 ( .A(n9917), .B(n9915), .ZN(n9927) );
  OAI21_X1 U10981 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9939) );
  NAND2_X1 U10982 ( .A1(n9939), .A2(n9919), .ZN(n9926) );
  OAI22_X1 U10983 ( .A1(n9923), .A2(n9922), .B1(n9921), .B2(n9920), .ZN(n9924)
         );
  INV_X1 U10984 ( .A(n9924), .ZN(n9925) );
  OAI211_X1 U10985 ( .C1(n9928), .C2(n9927), .A(n9926), .B(n9925), .ZN(n9937)
         );
  INV_X1 U10986 ( .A(n9939), .ZN(n9932) );
  OAI22_X1 U10987 ( .A1(n9932), .A2(n9931), .B1(n9930), .B2(n9929), .ZN(n9933)
         );
  AOI211_X1 U10988 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n9934), .A(n9937), .B(
        n9933), .ZN(n9935) );
  AOI22_X1 U10989 ( .A1(n9936), .A2(n6435), .B1(n9935), .B2(n9562), .ZN(
        P2_U3231) );
  INV_X1 U10990 ( .A(n9937), .ZN(n9941) );
  AOI22_X1 U10991 ( .A1(n9939), .A2(n6344), .B1(n9985), .B2(n9938), .ZN(n9940)
         );
  NAND2_X1 U10992 ( .A1(n9941), .A2(n9940), .ZN(n9989) );
  OAI22_X1 U10993 ( .A1(n9986), .A2(P2_REG0_REG_2__SCAN_IN), .B1(n9989), .B2(
        n9988), .ZN(n9942) );
  INV_X1 U10994 ( .A(n9942), .ZN(P2_U3396) );
  INV_X1 U10995 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9947) );
  OAI21_X1 U10996 ( .B1(n9944), .B2(n9967), .A(n9943), .ZN(n9945) );
  AOI21_X1 U10997 ( .B1(n9946), .B2(n9980), .A(n9945), .ZN(n9992) );
  AOI22_X1 U10998 ( .A1(n9988), .A2(n9947), .B1(n9992), .B2(n9986), .ZN(
        P2_U3402) );
  INV_X1 U10999 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U11000 ( .A1(n9948), .A2(n9967), .ZN(n9950) );
  AOI211_X1 U11001 ( .C1(n9980), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9994)
         );
  AOI22_X1 U11002 ( .A1(n9988), .A2(n9952), .B1(n9994), .B2(n9986), .ZN(
        P2_U3405) );
  NOR2_X1 U11003 ( .A1(n9953), .A2(n9967), .ZN(n9955) );
  AOI211_X1 U11004 ( .C1(n9956), .C2(n9980), .A(n9955), .B(n9954), .ZN(n9995)
         );
  AOI22_X1 U11005 ( .A1(n9988), .A2(n6025), .B1(n9995), .B2(n9986), .ZN(
        P2_U3408) );
  INV_X1 U11006 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9961) );
  OAI22_X1 U11007 ( .A1(n9958), .A2(n9969), .B1(n9957), .B2(n9967), .ZN(n9959)
         );
  NOR2_X1 U11008 ( .A1(n9960), .A2(n9959), .ZN(n9997) );
  AOI22_X1 U11009 ( .A1(n9988), .A2(n9961), .B1(n9997), .B2(n9986), .ZN(
        P2_U3411) );
  INV_X1 U11010 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U11011 ( .A1(n9962), .A2(n9967), .ZN(n9964) );
  AOI211_X1 U11012 ( .C1(n9980), .C2(n9965), .A(n9964), .B(n9963), .ZN(n9999)
         );
  AOI22_X1 U11013 ( .A1(n9988), .A2(n9966), .B1(n9999), .B2(n9986), .ZN(
        P2_U3414) );
  INV_X1 U11014 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9973) );
  OAI22_X1 U11015 ( .A1(n9970), .A2(n9969), .B1(n9968), .B2(n9967), .ZN(n9971)
         );
  NOR2_X1 U11016 ( .A1(n9972), .A2(n9971), .ZN(n10000) );
  AOI22_X1 U11017 ( .A1(n9988), .A2(n9973), .B1(n10000), .B2(n9986), .ZN(
        P2_U3420) );
  INV_X1 U11018 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9979) );
  NOR2_X1 U11019 ( .A1(n9975), .A2(n9974), .ZN(n9977) );
  AOI211_X1 U11020 ( .C1(n9985), .C2(n9978), .A(n9977), .B(n9976), .ZN(n10002)
         );
  AOI22_X1 U11021 ( .A1(n9988), .A2(n9979), .B1(n10002), .B2(n9986), .ZN(
        P2_U3423) );
  INV_X1 U11022 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9987) );
  AND2_X1 U11023 ( .A1(n9981), .A2(n9980), .ZN(n9983) );
  AOI211_X1 U11024 ( .C1(n9985), .C2(n9984), .A(n9983), .B(n9982), .ZN(n10005)
         );
  AOI22_X1 U11025 ( .A1(n9988), .A2(n9987), .B1(n10005), .B2(n9986), .ZN(
        P2_U3426) );
  OAI22_X1 U11026 ( .A1(n10004), .A2(n9989), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n10003), .ZN(n9990) );
  INV_X1 U11027 ( .A(n9990), .ZN(P2_U3461) );
  AOI22_X1 U11028 ( .A1(n10003), .A2(n9992), .B1(n9991), .B2(n10004), .ZN(
        P2_U3463) );
  AOI22_X1 U11029 ( .A1(n10003), .A2(n9994), .B1(n9993), .B2(n10004), .ZN(
        P2_U3464) );
  AOI22_X1 U11030 ( .A1(n10003), .A2(n9995), .B1(n6914), .B2(n10004), .ZN(
        P2_U3465) );
  AOI22_X1 U11031 ( .A1(n10003), .A2(n9997), .B1(n9996), .B2(n10004), .ZN(
        P2_U3466) );
  INV_X1 U11032 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U11033 ( .A1(n10003), .A2(n9999), .B1(n9998), .B2(n10004), .ZN(
        P2_U3467) );
  AOI22_X1 U11034 ( .A1(n10003), .A2(n10000), .B1(n7359), .B2(n10004), .ZN(
        P2_U3469) );
  AOI22_X1 U11035 ( .A1(n10003), .A2(n10002), .B1(n10001), .B2(n10004), .ZN(
        P2_U3470) );
  AOI22_X1 U11036 ( .A1(n10003), .A2(n10005), .B1(n7376), .B2(n10004), .ZN(
        P2_U3471) );
  NAND3_X1 U11037 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10008) );
  AND2_X1 U11038 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10006) );
  NOR2_X1 U11039 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10006), .ZN(n10007) );
  INV_X1 U11040 ( .A(n10007), .ZN(n10025) );
  NAND2_X1 U11041 ( .A1(n10009), .A2(n10008), .ZN(n10024) );
  OAI222_X1 U11042 ( .A1(n10009), .A2(n10008), .B1(n10009), .B2(n10025), .C1(
        n10007), .C2(n10024), .ZN(ADD_1068_U5) );
  XOR2_X1 U11043 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11044 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10010) );
  AOI21_X1 U11045 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10010), .ZN(n10032) );
  AOI22_X1 U11046 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10012), .B2(n10011), .ZN(n10035) );
  NOR2_X1 U11047 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10013) );
  AOI21_X1 U11048 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10013), .ZN(n10038) );
  NOR2_X1 U11049 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10014) );
  AOI21_X1 U11050 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10014), .ZN(n10041) );
  NOR2_X1 U11051 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10015) );
  AOI21_X1 U11052 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10015), .ZN(n10044) );
  NOR2_X1 U11053 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10016) );
  AOI21_X1 U11054 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10016), .ZN(n10047) );
  NOR2_X1 U11055 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10017) );
  AOI21_X1 U11056 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10017), .ZN(n10050) );
  NOR2_X1 U11057 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10018) );
  AOI21_X1 U11058 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10018), .ZN(n10053) );
  NOR2_X1 U11059 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10019) );
  AOI21_X1 U11060 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10019), .ZN(n10258) );
  NOR2_X1 U11061 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10020) );
  AOI21_X1 U11062 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10020), .ZN(n10261) );
  NOR2_X1 U11063 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10021) );
  AOI21_X1 U11064 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10021), .ZN(n10264) );
  NOR2_X1 U11065 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10022) );
  AOI21_X1 U11066 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10022), .ZN(n10267) );
  NOR2_X1 U11067 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10023) );
  AOI21_X1 U11068 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10023), .ZN(n10270) );
  NAND2_X1 U11069 ( .A1(n10025), .A2(n10024), .ZN(n10255) );
  NAND2_X1 U11070 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10026) );
  OAI21_X1 U11071 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10026), .ZN(n10254) );
  NOR2_X1 U11072 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  AOI21_X1 U11073 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10253), .ZN(n10273) );
  NAND2_X1 U11074 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10027) );
  OAI21_X1 U11075 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10027), .ZN(n10272) );
  NOR2_X1 U11076 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  AOI21_X1 U11077 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10271), .ZN(n10276) );
  NOR2_X1 U11078 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10028) );
  AOI21_X1 U11079 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10028), .ZN(n10275) );
  NAND2_X1 U11080 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  OAI21_X1 U11081 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10274), .ZN(n10269) );
  NAND2_X1 U11082 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  OAI21_X1 U11083 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10268), .ZN(n10266) );
  NAND2_X1 U11084 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  OAI21_X1 U11085 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10265), .ZN(n10263) );
  NAND2_X1 U11086 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  OAI21_X1 U11087 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10262), .ZN(n10260) );
  NAND2_X1 U11088 ( .A1(n10261), .A2(n10260), .ZN(n10259) );
  OAI21_X1 U11089 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10259), .ZN(n10257) );
  NAND2_X1 U11090 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U11091 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10256), .ZN(n10052) );
  NAND2_X1 U11092 ( .A1(n10053), .A2(n10052), .ZN(n10051) );
  OAI21_X1 U11093 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10051), .ZN(n10049) );
  NAND2_X1 U11094 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  OAI21_X1 U11095 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10048), .ZN(n10046) );
  NAND2_X1 U11096 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  OAI21_X1 U11097 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10045), .ZN(n10043) );
  NAND2_X1 U11098 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  OAI21_X1 U11099 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10042), .ZN(n10040) );
  NAND2_X1 U11100 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  OAI21_X1 U11101 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10039), .ZN(n10037) );
  NAND2_X1 U11102 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  OAI21_X1 U11103 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10036), .ZN(n10034) );
  NAND2_X1 U11104 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  OAI21_X1 U11105 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10033), .ZN(n10031) );
  NAND2_X1 U11106 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  OAI21_X1 U11107 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10030), .ZN(n10245) );
  NAND2_X1 U11108 ( .A1(n10246), .A2(n10245), .ZN(n10247) );
  OAI21_X1 U11109 ( .B1(n10245), .B2(n10246), .A(n10247), .ZN(n10029) );
  XNOR2_X1 U11110 ( .A(n10029), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11111 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(ADD_1068_U56) );
  OAI21_X1 U11112 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(ADD_1068_U57) );
  OAI21_X1 U11113 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(ADD_1068_U58) );
  OAI21_X1 U11114 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(ADD_1068_U59) );
  OAI21_X1 U11115 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(ADD_1068_U60) );
  OAI21_X1 U11116 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(ADD_1068_U61) );
  OAI21_X1 U11117 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(ADD_1068_U62) );
  OAI21_X1 U11118 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(ADD_1068_U63) );
  OAI22_X1 U11119 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        keyinput_f4), .B2(SI_28_), .ZN(n10054) );
  AOI221_X1 U11120 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        SI_28_), .C2(keyinput_f4), .A(n10054), .ZN(n10112) );
  OAI22_X1 U11121 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f49), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n10055) );
  AOI221_X1 U11122 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n10055), .ZN(n10111) );
  AOI22_X1 U11123 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n10056) );
  OAI221_X1 U11124 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_23_), .C2(
        keyinput_f9), .A(n10056), .ZN(n10063) );
  AOI22_X1 U11125 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n10057) );
  OAI221_X1 U11126 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n10057), .ZN(n10062)
         );
  AOI22_X1 U11127 ( .A1(SI_18_), .A2(keyinput_f14), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n10058) );
  OAI221_X1 U11128 ( .B1(SI_18_), .B2(keyinput_f14), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n10058), .ZN(n10061) );
  AOI22_X1 U11129 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10059) );
  OAI221_X1 U11130 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10059), .ZN(n10060)
         );
  NOR4_X1 U11131 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10067) );
  OAI22_X1 U11132 ( .A1(n10065), .A2(keyinput_f5), .B1(keyinput_f22), .B2(
        SI_10_), .ZN(n10064) );
  AOI221_X1 U11133 ( .B1(n10065), .B2(keyinput_f5), .C1(SI_10_), .C2(
        keyinput_f22), .A(n10064), .ZN(n10066) );
  OAI211_X1 U11134 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(
        n10067), .B(n10066), .ZN(n10068) );
  AOI21_X1 U11135 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .A(n10068), .ZN(n10110) );
  OAI22_X1 U11136 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(SI_7_), 
        .B2(keyinput_f25), .ZN(n10069) );
  AOI221_X1 U11137 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f25), .C2(SI_7_), .A(n10069), .ZN(n10076) );
  OAI22_X1 U11138 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        keyinput_f44), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10070) );
  AOI221_X1 U11139 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n10070), .ZN(n10075) );
  OAI22_X1 U11140 ( .A1(SI_13_), .A2(keyinput_f19), .B1(keyinput_f32), .B2(
        SI_0_), .ZN(n10071) );
  AOI221_X1 U11141 ( .B1(SI_13_), .B2(keyinput_f19), .C1(SI_0_), .C2(
        keyinput_f32), .A(n10071), .ZN(n10074) );
  OAI22_X1 U11142 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        keyinput_f27), .B2(SI_5_), .ZN(n10072) );
  AOI221_X1 U11143 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        SI_5_), .C2(keyinput_f27), .A(n10072), .ZN(n10073) );
  NAND4_X1 U11144 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10108) );
  OAI22_X1 U11145 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_f55), .B1(
        keyinput_f16), .B2(SI_16_), .ZN(n10077) );
  AOI221_X1 U11146 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .C1(
        SI_16_), .C2(keyinput_f16), .A(n10077), .ZN(n10084) );
  OAI22_X1 U11147 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        keyinput_f11), .B2(SI_21_), .ZN(n10078) );
  AOI221_X1 U11148 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_21_), .C2(keyinput_f11), .A(n10078), .ZN(n10083) );
  OAI22_X1 U11149 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f12), .B2(SI_20_), .ZN(n10079) );
  AOI221_X1 U11150 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        SI_20_), .C2(keyinput_f12), .A(n10079), .ZN(n10082) );
  OAI22_X1 U11151 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f17), .B2(SI_15_), .ZN(n10080) );
  AOI221_X1 U11152 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        SI_15_), .C2(keyinput_f17), .A(n10080), .ZN(n10081) );
  NAND4_X1 U11153 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n10107) );
  OAI22_X1 U11154 ( .A1(n10222), .A2(keyinput_f46), .B1(n10211), .B2(
        keyinput_f40), .ZN(n10085) );
  AOI221_X1 U11155 ( .B1(n10222), .B2(keyinput_f46), .C1(keyinput_f40), .C2(
        n10211), .A(n10085), .ZN(n10094) );
  OAI22_X1 U11156 ( .A1(n10231), .A2(keyinput_f18), .B1(n7526), .B2(
        keyinput_f1), .ZN(n10086) );
  AOI221_X1 U11157 ( .B1(n10231), .B2(keyinput_f18), .C1(keyinput_f1), .C2(
        n7526), .A(n10086), .ZN(n10093) );
  OAI22_X1 U11158 ( .A1(n10185), .A2(keyinput_f52), .B1(n10088), .B2(
        keyinput_f23), .ZN(n10087) );
  AOI221_X1 U11159 ( .B1(n10185), .B2(keyinput_f52), .C1(keyinput_f23), .C2(
        n10088), .A(n10087), .ZN(n10092) );
  OAI22_X1 U11160 ( .A1(n10090), .A2(keyinput_f6), .B1(n6719), .B2(
        keyinput_f59), .ZN(n10089) );
  AOI221_X1 U11161 ( .B1(n10090), .B2(keyinput_f6), .C1(keyinput_f59), .C2(
        n6719), .A(n10089), .ZN(n10091) );
  NAND4_X1 U11162 ( .A1(n10094), .A2(n10093), .A3(n10092), .A4(n10091), .ZN(
        n10106) );
  OAI22_X1 U11163 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n10095) );
  AOI221_X1 U11164 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        keyinput_f13), .C2(SI_19_), .A(n10095), .ZN(n10104) );
  OAI22_X1 U11165 ( .A1(SI_17_), .A2(keyinput_f15), .B1(keyinput_f28), .B2(
        SI_4_), .ZN(n10096) );
  AOI221_X1 U11166 ( .B1(SI_17_), .B2(keyinput_f15), .C1(SI_4_), .C2(
        keyinput_f28), .A(n10096), .ZN(n10103) );
  OAI22_X1 U11167 ( .A1(n10099), .A2(keyinput_f21), .B1(n10098), .B2(
        keyinput_f54), .ZN(n10097) );
  AOI221_X1 U11168 ( .B1(n10099), .B2(keyinput_f21), .C1(keyinput_f54), .C2(
        n10098), .A(n10097), .ZN(n10102) );
  INV_X1 U11169 ( .A(SI_6_), .ZN(n10232) );
  OAI22_X1 U11170 ( .A1(n10232), .A2(keyinput_f26), .B1(keyinput_f29), .B2(
        SI_3_), .ZN(n10100) );
  AOI221_X1 U11171 ( .B1(n10232), .B2(keyinput_f26), .C1(SI_3_), .C2(
        keyinput_f29), .A(n10100), .ZN(n10101) );
  NAND4_X1 U11172 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10105) );
  NOR4_X1 U11173 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        n10109) );
  NAND4_X1 U11174 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10142) );
  OAI22_X1 U11175 ( .A1(n10153), .A2(keyinput_f45), .B1(n10114), .B2(
        keyinput_f7), .ZN(n10113) );
  AOI221_X1 U11176 ( .B1(n10153), .B2(keyinput_f45), .C1(keyinput_f7), .C2(
        n10114), .A(n10113), .ZN(n10140) );
  INV_X1 U11177 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10117) );
  OAI22_X1 U11178 ( .A1(n10117), .A2(keyinput_f38), .B1(n10116), .B2(
        keyinput_f24), .ZN(n10115) );
  AOI221_X1 U11179 ( .B1(n10117), .B2(keyinput_f38), .C1(keyinput_f24), .C2(
        n10116), .A(n10115), .ZN(n10139) );
  OAI22_X1 U11180 ( .A1(n10119), .A2(keyinput_f48), .B1(n10184), .B2(
        keyinput_f8), .ZN(n10118) );
  AOI221_X1 U11181 ( .B1(n10119), .B2(keyinput_f48), .C1(keyinput_f8), .C2(
        n10184), .A(n10118), .ZN(n10121) );
  XNOR2_X1 U11182 ( .A(keyinput_f0), .B(P2_WR_REG_SCAN_IN), .ZN(n10120) );
  OAI211_X1 U11183 ( .C1(n10123), .C2(keyinput_f10), .A(n10121), .B(n10120), 
        .ZN(n10122) );
  AOI21_X1 U11184 ( .B1(n10123), .B2(keyinput_f10), .A(n10122), .ZN(n10138) );
  AOI22_X1 U11185 ( .A1(n10125), .A2(keyinput_f63), .B1(n6173), .B2(
        keyinput_f50), .ZN(n10124) );
  OAI221_X1 U11186 ( .B1(n10125), .B2(keyinput_f63), .C1(n6173), .C2(
        keyinput_f50), .A(n10124), .ZN(n10136) );
  AOI22_X1 U11187 ( .A1(n10127), .A2(keyinput_f35), .B1(keyinput_f3), .B2(
        n7516), .ZN(n10126) );
  OAI221_X1 U11188 ( .B1(n10127), .B2(keyinput_f35), .C1(n7516), .C2(
        keyinput_f3), .A(n10126), .ZN(n10135) );
  AOI22_X1 U11189 ( .A1(n10130), .A2(keyinput_f61), .B1(n10129), .B2(
        keyinput_f37), .ZN(n10128) );
  OAI221_X1 U11190 ( .B1(n10130), .B2(keyinput_f61), .C1(n10129), .C2(
        keyinput_f37), .A(n10128), .ZN(n10134) );
  XOR2_X1 U11191 ( .A(n6121), .B(keyinput_f56), .Z(n10132) );
  XNOR2_X1 U11192 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10131) );
  NAND2_X1 U11193 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  NOR4_X1 U11194 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  NAND4_X1 U11195 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10141) );
  OAI22_X1 U11196 ( .A1(n10142), .A2(n10141), .B1(keyinput_f30), .B2(SI_2_), 
        .ZN(n10143) );
  AOI21_X1 U11197 ( .B1(keyinput_f30), .B2(SI_2_), .A(n10143), .ZN(n10244) );
  AOI22_X1 U11198 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n10144) );
  OAI221_X1 U11199 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P2_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n10144), .ZN(n10151) );
  AOI22_X1 U11200 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10145) );
  OAI221_X1 U11201 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n10145), .ZN(n10150)
         );
  AOI22_X1 U11202 ( .A1(SI_31_), .A2(keyinput_g1), .B1(SI_11_), .B2(
        keyinput_g21), .ZN(n10146) );
  OAI221_X1 U11203 ( .B1(SI_31_), .B2(keyinput_g1), .C1(SI_11_), .C2(
        keyinput_g21), .A(n10146), .ZN(n10149) );
  AOI22_X1 U11204 ( .A1(SI_22_), .A2(keyinput_g10), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10147) );
  OAI221_X1 U11205 ( .B1(SI_22_), .B2(keyinput_g10), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n10147), .ZN(n10148)
         );
  NOR4_X1 U11206 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10179) );
  XNOR2_X1 U11207 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_g38), .ZN(n10159)
         );
  AOI22_X1 U11208 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        n10153), .B2(keyinput_g45), .ZN(n10152) );
  OAI221_X1 U11209 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        n10153), .C2(keyinput_g45), .A(n10152), .ZN(n10158) );
  AOI22_X1 U11210 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10154) );
  OAI221_X1 U11211 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10154), .ZN(n10157)
         );
  AOI22_X1 U11212 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n10155) );
  OAI221_X1 U11213 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n10155), .ZN(n10156) );
  NOR4_X1 U11214 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10178) );
  AOI22_X1 U11215 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n10160) );
  OAI221_X1 U11216 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_29_), .C2(
        keyinput_g3), .A(n10160), .ZN(n10167) );
  AOI22_X1 U11217 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_9_), 
        .B2(keyinput_g23), .ZN(n10161) );
  OAI221_X1 U11218 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(SI_9_), .C2(keyinput_g23), .A(n10161), .ZN(n10166) );
  AOI22_X1 U11219 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n10162) );
  OAI221_X1 U11220 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_27_), .C2(
        keyinput_g5), .A(n10162), .ZN(n10165) );
  AOI22_X1 U11221 ( .A1(SI_8_), .A2(keyinput_g24), .B1(SI_26_), .B2(
        keyinput_g6), .ZN(n10163) );
  OAI221_X1 U11222 ( .B1(SI_8_), .B2(keyinput_g24), .C1(SI_26_), .C2(
        keyinput_g6), .A(n10163), .ZN(n10164) );
  NOR4_X1 U11223 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10177) );
  AOI22_X1 U11224 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n10168) );
  OAI221_X1 U11225 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n10168), .ZN(n10175)
         );
  AOI22_X1 U11226 ( .A1(SI_7_), .A2(keyinput_g25), .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n10169) );
  OAI221_X1 U11227 ( .B1(SI_7_), .B2(keyinput_g25), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n10169), .ZN(n10174)
         );
  AOI22_X1 U11228 ( .A1(SI_12_), .A2(keyinput_g20), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n10170) );
  OAI221_X1 U11229 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10170), .ZN(n10173)
         );
  AOI22_X1 U11230 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n10171) );
  OAI221_X1 U11231 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n10171), .ZN(n10172)
         );
  NOR4_X1 U11232 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10176) );
  NAND4_X1 U11233 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10242) );
  INV_X1 U11234 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U11235 ( .A1(n10182), .A2(keyinput_g15), .B1(n10181), .B2(
        keyinput_g42), .ZN(n10180) );
  OAI221_X1 U11236 ( .B1(n10182), .B2(keyinput_g15), .C1(n10181), .C2(
        keyinput_g42), .A(n10180), .ZN(n10194) );
  AOI22_X1 U11237 ( .A1(n10185), .A2(keyinput_g52), .B1(keyinput_g8), .B2(
        n10184), .ZN(n10183) );
  OAI221_X1 U11238 ( .B1(n10185), .B2(keyinput_g52), .C1(n10184), .C2(
        keyinput_g8), .A(n10183), .ZN(n10193) );
  INV_X1 U11239 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U11240 ( .A1(n10188), .A2(keyinput_g17), .B1(n10187), .B2(
        keyinput_g36), .ZN(n10186) );
  OAI221_X1 U11241 ( .B1(n10188), .B2(keyinput_g17), .C1(n10187), .C2(
        keyinput_g36), .A(n10186), .ZN(n10192) );
  XNOR2_X1 U11242 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_g43), .ZN(n10190)
         );
  XNOR2_X1 U11243 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10189) );
  NAND2_X1 U11244 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  NOR4_X1 U11245 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10240) );
  AOI22_X1 U11246 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n10195) );
  OAI221_X1 U11247 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n10195), .ZN(n10206) );
  AOI22_X1 U11248 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n10196) );
  OAI221_X1 U11249 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n10196), .ZN(n10205)
         );
  AOI22_X1 U11250 ( .A1(n10199), .A2(keyinput_g11), .B1(keyinput_g27), .B2(
        n10198), .ZN(n10197) );
  OAI221_X1 U11251 ( .B1(n10199), .B2(keyinput_g11), .C1(n10198), .C2(
        keyinput_g27), .A(n10197), .ZN(n10204) );
  INV_X1 U11252 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10202) );
  AOI22_X1 U11253 ( .A1(n10202), .A2(keyinput_g0), .B1(n10201), .B2(
        keyinput_g4), .ZN(n10200) );
  OAI221_X1 U11254 ( .B1(n10202), .B2(keyinput_g0), .C1(n10201), .C2(
        keyinput_g4), .A(n10200), .ZN(n10203) );
  NOR4_X1 U11255 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10239) );
  AOI22_X1 U11256 ( .A1(n10208), .A2(keyinput_g55), .B1(keyinput_g53), .B2(
        n6068), .ZN(n10207) );
  OAI221_X1 U11257 ( .B1(n10208), .B2(keyinput_g55), .C1(n6068), .C2(
        keyinput_g53), .A(n10207), .ZN(n10220) );
  AOI22_X1 U11258 ( .A1(n10211), .A2(keyinput_g40), .B1(keyinput_g19), .B2(
        n10210), .ZN(n10209) );
  OAI221_X1 U11259 ( .B1(n10211), .B2(keyinput_g40), .C1(n10210), .C2(
        keyinput_g19), .A(n10209), .ZN(n10219) );
  AOI22_X1 U11260 ( .A1(n10214), .A2(keyinput_g9), .B1(keyinput_g16), .B2(
        n10213), .ZN(n10212) );
  OAI221_X1 U11261 ( .B1(n10214), .B2(keyinput_g9), .C1(n10213), .C2(
        keyinput_g16), .A(n10212), .ZN(n10218) );
  XNOR2_X1 U11262 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10216) );
  XNOR2_X1 U11263 ( .A(SI_20_), .B(keyinput_g12), .ZN(n10215) );
  NAND2_X1 U11264 ( .A1(n10216), .A2(n10215), .ZN(n10217) );
  NOR4_X1 U11265 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10238) );
  AOI22_X1 U11266 ( .A1(n10223), .A2(keyinput_g13), .B1(n10222), .B2(
        keyinput_g46), .ZN(n10221) );
  OAI221_X1 U11267 ( .B1(n10223), .B2(keyinput_g13), .C1(n10222), .C2(
        keyinput_g46), .A(n10221), .ZN(n10236) );
  INV_X1 U11268 ( .A(SI_18_), .ZN(n10225) );
  AOI22_X1 U11269 ( .A1(n10226), .A2(keyinput_g2), .B1(n10225), .B2(
        keyinput_g14), .ZN(n10224) );
  OAI221_X1 U11270 ( .B1(n10226), .B2(keyinput_g2), .C1(n10225), .C2(
        keyinput_g14), .A(n10224), .ZN(n10235) );
  INV_X1 U11271 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10229) );
  INV_X1 U11272 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10228) );
  AOI22_X1 U11273 ( .A1(n10229), .A2(keyinput_g41), .B1(keyinput_g33), .B2(
        n10228), .ZN(n10227) );
  OAI221_X1 U11274 ( .B1(n10229), .B2(keyinput_g41), .C1(n10228), .C2(
        keyinput_g33), .A(n10227), .ZN(n10234) );
  AOI22_X1 U11275 ( .A1(n10232), .A2(keyinput_g26), .B1(n10231), .B2(
        keyinput_g18), .ZN(n10230) );
  OAI221_X1 U11276 ( .B1(n10232), .B2(keyinput_g26), .C1(n10231), .C2(
        keyinput_g18), .A(n10230), .ZN(n10233) );
  NOR4_X1 U11277 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10237) );
  NAND4_X1 U11278 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  OAI22_X1 U11279 ( .A1(SI_2_), .A2(keyinput_g30), .B1(n10242), .B2(n10241), 
        .ZN(n10243) );
  AOI211_X1 U11280 ( .C1(SI_2_), .C2(keyinput_g30), .A(n10244), .B(n10243), 
        .ZN(n10252) );
  NOR2_X1 U11281 ( .A1(n10246), .A2(n10245), .ZN(n10248) );
  OAI21_X1 U11282 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10248), .A(n10247), 
        .ZN(n10250) );
  XNOR2_X1 U11283 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10249) );
  XNOR2_X1 U11284 ( .A(n10250), .B(n10249), .ZN(n10251) );
  XNOR2_X1 U11285 ( .A(n10252), .B(n10251), .ZN(ADD_1068_U4) );
  AOI21_X1 U11286 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(ADD_1068_U54) );
  OAI21_X1 U11287 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(ADD_1068_U47) );
  OAI21_X1 U11288 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(ADD_1068_U48) );
  OAI21_X1 U11289 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(ADD_1068_U49) );
  OAI21_X1 U11290 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(ADD_1068_U50) );
  OAI21_X1 U11291 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(ADD_1068_U51) );
  AOI21_X1 U11292 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(ADD_1068_U53) );
  OAI21_X1 U11293 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(ADD_1068_U52) );
  AND3_X2 U6231 ( .A1(n5047), .A2(n5046), .A3(n5045), .ZN(n5813) );
  BUF_X1 U4946 ( .A(n5058), .Z(n6495) );
  AND2_X1 U4873 ( .A1(n5857), .A2(n5002), .ZN(n4975) );
  AND2_X1 U4874 ( .A1(n4937), .A2(n4722), .ZN(n4946) );
  CLKBUF_X1 U4880 ( .A(n6712), .Z(n7922) );
  CLKBUF_X1 U4886 ( .A(n5975), .Z(n4357) );
  CLKBUF_X1 U4894 ( .A(n5758), .Z(n4355) );
  CLKBUF_X2 U4919 ( .A(n6420), .Z(n4350) );
endmodule

