

module b17_C_AntiSAT_k_256_9 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9809, n9810, n9811, n9812, n9813, n9815, n9816, n9817, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363;

  NOR2_X1 U11253 ( .A1(n17900), .A2(n18233), .ZN(n17899) );
  NOR2_X1 U11254 ( .A1(n15374), .A2(n15373), .ZN(n15372) );
  NAND2_X1 U11255 ( .A1(n10660), .A2(n10659), .ZN(n13608) );
  NAND2_X1 U11256 ( .A1(n13719), .A2(n13996), .ZN(n13720) );
  OR2_X1 U11257 ( .A1(n17914), .A2(n12275), .ZN(n9871) );
  INV_X1 U11258 ( .A(n10456), .ZN(n12132) );
  CLKBUF_X1 U11259 ( .A(n9835), .Z(n11081) );
  OR2_X1 U11260 ( .A1(n12566), .A2(n12544), .ZN(n12616) );
  NAND3_X2 U11261 ( .A1(n12377), .A2(n12376), .A3(n12375), .ZN(n18367) );
  CLKBUF_X1 U11263 ( .A(n12240), .Z(n9813) );
  INV_X1 U11264 ( .A(n11799), .ZN(n15158) );
  AND2_X1 U11265 ( .A1(n11626), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15101) );
  INV_X1 U11266 ( .A(n14198), .ZN(n17319) );
  INV_X1 U11267 ( .A(n17325), .ZN(n12379) );
  AND2_X1 U11268 ( .A1(n11620), .A2(n10218), .ZN(n15143) );
  CLKBUF_X2 U11269 ( .A(n11636), .Z(n15320) );
  INV_X1 U11270 ( .A(n9874), .ZN(n17318) );
  BUF_X2 U11271 ( .A(n12302), .Z(n17283) );
  CLKBUF_X2 U11272 ( .A(n12183), .Z(n17317) );
  CLKBUF_X2 U11273 ( .A(n12240), .Z(n17310) );
  INV_X2 U11274 ( .A(n12318), .ZN(n17301) );
  CLKBUF_X2 U11275 ( .A(n10610), .Z(n10910) );
  CLKBUF_X2 U11276 ( .A(n10506), .Z(n11074) );
  CLKBUF_X2 U11277 ( .A(n10421), .Z(n9821) );
  BUF_X2 U11278 ( .A(n10359), .Z(n11055) );
  CLKBUF_X1 U11279 ( .A(n12183), .Z(n14174) );
  INV_X1 U11280 ( .A(n9874), .ZN(n14169) );
  NAND2_X1 U11281 ( .A1(n11437), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11510) );
  INV_X1 U11282 ( .A(n12929), .ZN(n12911) );
  INV_X2 U11283 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12414) );
  NAND2_X2 U11284 ( .A1(n10446), .A2(n10448), .ZN(n13009) );
  INV_X1 U11285 ( .A(n10412), .ZN(n10447) );
  BUF_X1 U11288 ( .A(n11440), .Z(n19337) );
  AND2_X1 U11289 ( .A1(n13490), .A2(n10327), .ZN(n9824) );
  AND2_X1 U11290 ( .A1(n10322), .A2(n10334), .ZN(n9835) );
  AND2_X1 U11291 ( .A1(n10322), .A2(n10334), .ZN(n9836) );
  AND2_X1 U11292 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10334) );
  INV_X1 U11293 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10321) );
  OR2_X1 U11294 ( .A1(n18357), .A2(n9811), .ZN(n17445) );
  INV_X1 U11295 ( .A(n17445), .ZN(n9809) );
  INV_X1 U11296 ( .A(n17511), .ZN(n9810) );
  INV_X1 U11297 ( .A(n9810), .ZN(n9811) );
  INV_X1 U11298 ( .A(n9810), .ZN(n9812) );
  INV_X4 U11299 ( .A(n18317), .ZN(n9816) );
  OR2_X1 U11300 ( .A1(n11510), .A2(n21237), .ZN(n11504) );
  AND2_X1 U11301 ( .A1(n11621), .A2(n10218), .ZN(n15064) );
  CLKBUF_X2 U11302 ( .A(n11644), .Z(n15319) );
  NAND2_X1 U11303 ( .A1(n12415), .A2(n18925), .ZN(n12161) );
  OR2_X1 U11304 ( .A1(n10395), .A2(n10394), .ZN(n13193) );
  XNOR2_X1 U11305 ( .A(n12843), .B(n12844), .ZN(n13719) );
  NOR2_X1 U11306 ( .A1(n15475), .A2(n15481), .ZN(n12865) );
  OR2_X1 U11307 ( .A1(n10052), .A2(n10286), .ZN(n10027) );
  OR2_X1 U11308 ( .A1(n12566), .A2(n12536), .ZN(n19442) );
  AND2_X1 U11309 ( .A1(n12566), .A2(n12546), .ZN(n19636) );
  AND2_X1 U11310 ( .A1(n12545), .A2(n12566), .ZN(n12634) );
  INV_X1 U11312 ( .A(n18342), .ZN(n15945) );
  OR2_X1 U11313 ( .A1(n17769), .A2(n10072), .ZN(n12288) );
  NOR2_X1 U11314 ( .A1(n12404), .A2(n12409), .ZN(n15936) );
  INV_X1 U11316 ( .A(n13280), .ZN(n20274) );
  NOR2_X1 U11317 ( .A1(n15363), .A2(n15196), .ZN(n15220) );
  NAND2_X1 U11318 ( .A1(n12526), .A2(n12527), .ZN(n10007) );
  NOR2_X1 U11319 ( .A1(n15767), .A2(n15768), .ZN(n15766) );
  INV_X1 U11320 ( .A(n16460), .ZN(n19124) );
  AND2_X1 U11321 ( .A1(n12578), .A2(n13228), .ZN(n12630) );
  NAND2_X1 U11322 ( .A1(n13445), .A2(n13444), .ZN(n20257) );
  INV_X1 U11324 ( .A(n17780), .ZN(n10072) );
  INV_X1 U11325 ( .A(n13789), .ZN(n15399) );
  INV_X1 U11326 ( .A(n20136), .ZN(n20114) );
  NAND2_X1 U11327 ( .A1(n14420), .A2(n11274), .ZN(n14244) );
  INV_X1 U11328 ( .A(n12307), .ZN(n9815) );
  INV_X1 U11329 ( .A(n9815), .ZN(n9817) );
  NAND2_X1 U11330 ( .A1(n12553), .A2(n12538), .ZN(n19150) );
  NAND2_X2 U11331 ( .A1(n12537), .A2(n12553), .ZN(n12528) );
  NAND3_X1 U11333 ( .A1(n18354), .A2(n17377), .A3(n15945), .ZN(n12402) );
  INV_X2 U11334 ( .A(n14084), .ZN(n10151) );
  OR2_X1 U11335 ( .A1(n14430), .A2(n10161), .ZN(n11103) );
  NAND2_X2 U11336 ( .A1(n11467), .A2(n11466), .ZN(n11492) );
  AOI21_X4 U11337 ( .B1(n16023), .B2(n16022), .A(n18817), .ZN(n17517) );
  NAND2_X1 U11338 ( .A1(n13591), .A2(n10211), .ZN(n13730) );
  NAND2_X2 U11339 ( .A1(n13401), .A2(n13400), .ZN(n13591) );
  NOR2_X2 U11340 ( .A1(n17865), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17854) );
  OAI21_X2 U11341 ( .B1(n12832), .B2(n11953), .A(n11667), .ZN(n13298) );
  AOI211_X2 U11342 ( .C1(n16426), .C2(n16301), .A(n15497), .B(n15496), .ZN(
        n15498) );
  INV_X4 U11343 ( .A(n12379), .ZN(n14185) );
  AOI21_X2 U11344 ( .B1(n10072), .B2(n17648), .A(n16597), .ZN(n17640) );
  NAND2_X2 U11345 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12293), .ZN(
        n17648) );
  OAI211_X2 U11346 ( .C1(n10471), .C2(n10321), .A(n9974), .B(n10455), .ZN(
        n10501) );
  AND2_X4 U11347 ( .A1(n13280), .A2(n13309), .ZN(n13349) );
  AND3_X1 U11348 ( .A1(n12291), .A2(n10061), .A3(n10060), .ZN(n17658) );
  XNOR2_X1 U11349 ( .A(n12134), .B(n12133), .ZN(n14508) );
  NAND2_X1 U11350 ( .A1(n13759), .A2(n10210), .ZN(n13900) );
  NOR2_X1 U11351 ( .A1(n16454), .A2(n12961), .ZN(n15851) );
  AND2_X1 U11352 ( .A1(n15750), .A2(n15753), .ZN(n15864) );
  NAND2_X2 U11353 ( .A1(n20157), .A2(n13353), .ZN(n14564) );
  NAND2_X1 U11354 ( .A1(n17517), .A2(n18367), .ZN(n17511) );
  NAND2_X2 U11355 ( .A1(n18788), .A2(n18197), .ZN(n18288) );
  AND2_X1 U11356 ( .A1(n11519), .A2(n11518), .ZN(n12523) );
  NOR2_X1 U11357 ( .A1(n17581), .A2(n15934), .ZN(n16696) );
  AND2_X1 U11358 ( .A1(n11429), .A2(n11438), .ZN(n15216) );
  INV_X4 U11359 ( .A(n15191), .ZN(n15910) );
  INV_X1 U11360 ( .A(n13306), .ZN(n20966) );
  AND2_X1 U11361 ( .A1(n13181), .A2(n10452), .ZN(n13039) );
  OR2_X1 U11362 ( .A1(n11117), .A2(n12041), .ZN(n10438) );
  NAND2_X1 U11363 ( .A1(n11428), .A2(n11429), .ZN(n11683) );
  AND2_X1 U11364 ( .A1(n20298), .A2(n13019), .ZN(n11160) );
  AND3_X1 U11365 ( .A1(n11453), .A2(n11440), .A3(n11439), .ZN(n11443) );
  AND2_X1 U11366 ( .A1(n11446), .A2(n11439), .ZN(n11450) );
  INV_X2 U11367 ( .A(n13309), .ZN(n20287) );
  NOR2_X1 U11368 ( .A1(n13193), .A2(n13019), .ZN(n12494) );
  OR2_X2 U11370 ( .A1(n10411), .A2(n10410), .ZN(n13280) );
  AND4_X2 U11371 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10412) );
  AND4_X1 U11372 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10437) );
  INV_X1 U11373 ( .A(n14198), .ZN(n17298) );
  CLKBUF_X2 U11374 ( .A(n9825), .Z(n10981) );
  BUF_X1 U11375 ( .A(n12307), .Z(n9822) );
  CLKBUF_X3 U11377 ( .A(n12241), .Z(n17323) );
  CLKBUF_X1 U11378 ( .A(n9829), .Z(n10916) );
  INV_X1 U11379 ( .A(n12229), .ZN(n12246) );
  CLKBUF_X2 U11380 ( .A(n10389), .Z(n11082) );
  BUF_X2 U11381 ( .A(n10708), .Z(n11080) );
  CLKBUF_X2 U11382 ( .A(n10367), .Z(n10915) );
  AND2_X2 U11383 ( .A1(n10327), .A2(n10332), .ZN(n10389) );
  OR2_X2 U11384 ( .A1(n17075), .A2(n12158), .ZN(n17022) );
  AND2_X2 U11385 ( .A1(n10332), .A2(n14894), .ZN(n9839) );
  AND2_X1 U11386 ( .A1(n10333), .A2(n10332), .ZN(n10488) );
  NAND2_X4 U11387 ( .A1(n12414), .A2(n12413), .ZN(n17074) );
  NOR2_X4 U11388 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10332) );
  AND2_X1 U11389 ( .A1(n12983), .A2(n12982), .ZN(n12984) );
  AND2_X1 U11390 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  OR2_X1 U11391 ( .A1(n12932), .A2(n16424), .ZN(n12874) );
  XNOR2_X1 U11393 ( .A(n14623), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14753) );
  NAND2_X1 U11394 ( .A1(n12864), .A2(n12966), .ZN(n15475) );
  NAND2_X1 U11395 ( .A1(n15682), .A2(n10006), .ZN(n16338) );
  AND2_X1 U11396 ( .A1(n9968), .A2(n9967), .ZN(n15802) );
  NAND2_X1 U11397 ( .A1(n16376), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16377) );
  AND2_X1 U11398 ( .A1(n15834), .A2(n15817), .ZN(n16376) );
  OR2_X1 U11399 ( .A1(n15572), .A2(n15788), .ZN(n16345) );
  OR2_X1 U11400 ( .A1(n15344), .A2(n15343), .ZN(n10205) );
  AND2_X1 U11401 ( .A1(n15599), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15834) );
  AND2_X1 U11402 ( .A1(n9880), .A2(n14526), .ZN(n16051) );
  AND2_X1 U11403 ( .A1(n14646), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14658) );
  NAND2_X1 U11404 ( .A1(n10027), .A2(n10025), .ZN(n15595) );
  NAND2_X1 U11405 ( .A1(n10059), .A2(n10057), .ZN(n10052) );
  NAND2_X1 U11406 ( .A1(n13956), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13955) );
  NAND2_X1 U11407 ( .A1(n15348), .A2(n15350), .ZN(n15349) );
  NAND2_X1 U11408 ( .A1(n15961), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16005) );
  AND2_X1 U11409 ( .A1(n10012), .A2(n16403), .ZN(n10014) );
  NAND2_X1 U11410 ( .A1(n15357), .A2(n15221), .ZN(n10197) );
  NAND2_X1 U11411 ( .A1(n10268), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10267) );
  NAND2_X1 U11412 ( .A1(n15359), .A2(n15358), .ZN(n15357) );
  INV_X1 U11413 ( .A(n10269), .ZN(n10266) );
  NAND2_X1 U11414 ( .A1(n9979), .A2(n9977), .ZN(n9976) );
  XNOR2_X1 U11415 ( .A(n15220), .B(n15217), .ZN(n15359) );
  NAND2_X1 U11416 ( .A1(n16185), .A2(n16183), .ZN(n9979) );
  OAI22_X1 U11417 ( .A1(n13717), .A2(n13718), .B1(n13818), .B2(n13996), .ZN(
        n13992) );
  CLKBUF_X1 U11418 ( .A(n12858), .Z(n12860) );
  NAND2_X1 U11419 ( .A1(n10169), .A2(n11223), .ZN(n16185) );
  NAND2_X1 U11420 ( .A1(n12842), .A2(n12841), .ZN(n12844) );
  NAND2_X1 U11421 ( .A1(n12292), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10061) );
  NAND3_X1 U11422 ( .A1(n9971), .A2(n10004), .A3(n12612), .ZN(n12698) );
  NOR2_X1 U11423 ( .A1(n10184), .A2(n9978), .ZN(n9977) );
  INV_X1 U11424 ( .A(n12650), .ZN(n9971) );
  AND4_X1 U11425 ( .A1(n14701), .A2(n14702), .A3(n11254), .A4(n16160), .ZN(
        n11255) );
  AND2_X1 U11426 ( .A1(n12287), .A2(n12288), .ZN(n17693) );
  AND2_X1 U11427 ( .A1(n14705), .A2(n16159), .ZN(n16148) );
  AND2_X1 U11428 ( .A1(n11239), .A2(n9896), .ZN(n10185) );
  AND2_X1 U11429 ( .A1(n12288), .A2(n9994), .ZN(n17765) );
  NOR2_X1 U11430 ( .A1(n11247), .A2(n14308), .ZN(n14713) );
  AND2_X1 U11431 ( .A1(n11220), .A2(n11219), .ZN(n16189) );
  OR2_X1 U11432 ( .A1(n17781), .A2(n17690), .ZN(n12283) );
  OR2_X1 U11433 ( .A1(n17781), .A2(n12289), .ZN(n9994) );
  XNOR2_X1 U11434 ( .A(n11215), .B(n10681), .ZN(n11225) );
  NAND2_X2 U11435 ( .A1(n11215), .A2(n11171), .ZN(n16173) );
  NAND2_X1 U11436 ( .A1(n12279), .A2(n17780), .ZN(n12286) );
  AND2_X1 U11437 ( .A1(n12285), .A2(n10064), .ZN(n9995) );
  NAND2_X1 U11438 ( .A1(n10638), .A2(n9917), .ZN(n11215) );
  NAND2_X1 U11439 ( .A1(n12794), .A2(n12798), .ZN(n16299) );
  NAND2_X1 U11440 ( .A1(n10636), .A2(n10601), .ZN(n11190) );
  NOR2_X1 U11441 ( .A1(n17801), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17818) );
  OAI21_X1 U11442 ( .B1(n13386), .B2(n13385), .A(n13401), .ZN(n19972) );
  NOR2_X1 U11443 ( .A1(n13797), .A2(n13798), .ZN(n15800) );
  OAI22_X1 U11444 ( .A1(n12569), .A2(n15174), .B1(n15181), .B2(n12685), .ZN(
        n12570) );
  AND2_X1 U11445 ( .A1(n10259), .A2(n12551), .ZN(n12631) );
  NAND2_X1 U11446 ( .A1(n17902), .A2(n10072), .ZN(n17901) );
  OAI22_X1 U11447 ( .A1(n12616), .A2(n12592), .B1(n19442), .B2(n12591), .ZN(
        n12593) );
  OAI22_X1 U11448 ( .A1(n19785), .A2(n12598), .B1(n12685), .B2(n15230), .ZN(
        n12599) );
  NAND2_X1 U11449 ( .A1(n12556), .A2(n13119), .ZN(n12615) );
  AND2_X1 U11450 ( .A1(n12578), .A2(n13119), .ZN(n19411) );
  AND2_X1 U11451 ( .A1(n12551), .A2(n12552), .ZN(n12556) );
  NAND2_X1 U11452 ( .A1(n12551), .A2(n12568), .ZN(n12685) );
  NAND2_X1 U11453 ( .A1(n10005), .A2(n12539), .ZN(n12561) );
  OR2_X1 U11454 ( .A1(n12572), .A2(n12573), .ZN(n19785) );
  AOI21_X1 U11455 ( .B1(n13379), .B2(n13378), .A(n9924), .ZN(n13381) );
  CLKBUF_X1 U11456 ( .A(n12516), .Z(n14611) );
  XNOR2_X1 U11457 ( .A(n13328), .B(n10167), .ZN(n13031) );
  NOR2_X1 U11458 ( .A1(n12280), .A2(n10072), .ZN(n17878) );
  INV_X1 U11459 ( .A(n17861), .ZN(n17906) );
  AND2_X1 U11460 ( .A1(n13374), .A2(n13375), .ZN(n13378) );
  NAND2_X1 U11461 ( .A1(n10599), .A2(n10598), .ZN(n20447) );
  NAND2_X1 U11462 ( .A1(n13074), .A2(n13073), .ZN(n13271) );
  NAND2_X2 U11463 ( .A1(n14600), .A2(n13365), .ZN(n14615) );
  OAI21_X1 U11464 ( .B1(n13176), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10495), 
        .ZN(n10498) );
  AND2_X1 U11465 ( .A1(n12928), .A2(n13295), .ZN(n12974) );
  NOR2_X1 U11466 ( .A1(n17915), .A2(n18228), .ZN(n17914) );
  NOR2_X1 U11467 ( .A1(n14560), .A2(n14559), .ZN(n14562) );
  NOR2_X2 U11468 ( .A1(n19325), .A2(n19576), .ZN(n19326) );
  NOR2_X1 U11469 ( .A1(n13814), .A2(n13698), .ZN(n13994) );
  XNOR2_X1 U11470 ( .A(n10581), .B(n20448), .ZN(n20558) );
  NOR2_X2 U11471 ( .A1(n19232), .A2(n19576), .ZN(n15917) );
  NOR2_X1 U11472 ( .A1(n18057), .A2(n18302), .ZN(n18307) );
  NOR2_X1 U11473 ( .A1(n12751), .A2(n12740), .ZN(n12741) );
  INV_X1 U11474 ( .A(n14061), .ZN(n10115) );
  OR2_X1 U11475 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  XNOR2_X1 U11476 ( .A(n10549), .B(n10547), .ZN(n10561) );
  INV_X2 U11477 ( .A(n11321), .ZN(n19117) );
  NAND2_X1 U11478 ( .A1(n10037), .A2(n10036), .ZN(n10549) );
  NAND2_X1 U11479 ( .A1(n12530), .A2(n12529), .ZN(n12553) );
  INV_X1 U11480 ( .A(n12523), .ZN(n12524) );
  OR2_X1 U11481 ( .A1(n16250), .A2(n13981), .ZN(n14061) );
  NAND2_X1 U11482 ( .A1(n9970), .A2(n11505), .ZN(n11509) );
  NAND2_X1 U11483 ( .A1(n15936), .A2(n15935), .ZN(n18760) );
  NAND2_X1 U11484 ( .A1(n12921), .A2(n12919), .ZN(n16523) );
  AOI21_X1 U11485 ( .B1(n10472), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10473), .ZN(n10482) );
  OR2_X1 U11486 ( .A1(n11516), .A2(n11517), .ZN(n11519) );
  NAND2_X1 U11487 ( .A1(n11504), .A2(n11503), .ZN(n11506) );
  NAND2_X1 U11488 ( .A1(n11491), .A2(n11490), .ZN(n12529) );
  NAND2_X1 U11489 ( .A1(n13034), .A2(n10453), .ZN(n10454) );
  AND2_X1 U11490 ( .A1(n10465), .A2(n10464), .ZN(n10467) );
  CLKBUF_X1 U11491 ( .A(n11487), .Z(n15884) );
  AND2_X1 U11492 ( .A1(n13298), .A2(n13297), .ZN(n13300) );
  NAND2_X1 U11493 ( .A1(n11465), .A2(n11612), .ZN(n16495) );
  AND2_X1 U11494 ( .A1(n11613), .A2(n11427), .ZN(n11465) );
  NOR2_X1 U11495 ( .A1(n12660), .A2(n10243), .ZN(n10242) );
  AOI21_X1 U11496 ( .B1(n12020), .B2(n12138), .A(n13039), .ZN(n10453) );
  AND2_X1 U11497 ( .A1(n11426), .A2(n12945), .ZN(n12947) );
  XNOR2_X1 U11498 ( .A(n12436), .B(n12258), .ZN(n12259) );
  AND2_X1 U11499 ( .A1(n10415), .A2(n10457), .ZN(n13018) );
  NOR2_X1 U11500 ( .A1(n12260), .A2(n17507), .ZN(n12264) );
  NOR2_X1 U11501 ( .A1(n15191), .A2(n19237), .ZN(n11438) );
  INV_X1 U11502 ( .A(n10456), .ZN(n12121) );
  OR2_X2 U11503 ( .A1(n11615), .A2(n11616), .ZN(n11978) );
  NAND2_X1 U11504 ( .A1(n10456), .A2(n13349), .ZN(n12040) );
  INV_X1 U11505 ( .A(n17520), .ZN(n12258) );
  NAND2_X2 U11506 ( .A1(n12218), .A2(n10298), .ZN(n17520) );
  AND2_X1 U11507 ( .A1(n11445), .A2(n11446), .ZN(n11455) );
  AND2_X1 U11508 ( .A1(n12494), .A2(n12496), .ZN(n13181) );
  NOR2_X1 U11509 ( .A1(n17772), .A2(n17773), .ZN(n16718) );
  AND4_X1 U11510 ( .A1(n12215), .A2(n12214), .A3(n12213), .A4(n12212), .ZN(
        n12218) );
  INV_X1 U11511 ( .A(n11446), .ZN(n13303) );
  NAND2_X1 U11512 ( .A1(n11352), .A2(n11351), .ZN(n11446) );
  NAND2_X1 U11513 ( .A1(n11340), .A2(n11339), .ZN(n11439) );
  NAND2_X2 U11514 ( .A1(n11375), .A2(n11376), .ZN(n13630) );
  NAND2_X1 U11515 ( .A1(n10009), .A2(n10008), .ZN(n11440) );
  NAND2_X1 U11516 ( .A1(n11362), .A2(n9886), .ZN(n11363) );
  NAND2_X1 U11517 ( .A1(n9890), .A2(n10011), .ZN(n10008) );
  NAND2_X1 U11518 ( .A1(n9891), .A2(n10010), .ZN(n10009) );
  AND4_X1 U11519 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  AND4_X1 U11520 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10435) );
  NAND2_X1 U11521 ( .A1(n11387), .A2(n11386), .ZN(n11388) );
  NAND2_X1 U11522 ( .A1(n10300), .A2(n11381), .ZN(n11389) );
  NAND2_X2 U11523 ( .A1(n10310), .A2(n9870), .ZN(n13353) );
  AND2_X1 U11524 ( .A1(n11385), .A2(n11384), .ZN(n11386) );
  AND3_X1 U11525 ( .A1(n11380), .A2(n11408), .A3(n11379), .ZN(n11381) );
  AND4_X1 U11526 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        n10436) );
  AND4_X1 U11527 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10339) );
  AND4_X1 U11528 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10340) );
  AND4_X1 U11529 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10341) );
  NAND2_X2 U11530 ( .A1(n18980), .A2(n18847), .ZN(n18905) );
  AND4_X1 U11531 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10342) );
  CLKBUF_X1 U11532 ( .A(n10752), .Z(n9843) );
  AND3_X1 U11533 ( .A1(n11396), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11395), .ZN(n10010) );
  CLKBUF_X1 U11534 ( .A(n10752), .Z(n9844) );
  AND3_X1 U11535 ( .A1(n11392), .A2(n11408), .A3(n11390), .ZN(n10011) );
  INV_X2 U11536 ( .A(n12348), .ZN(n17327) );
  BUF_X2 U11537 ( .A(n12246), .Z(n17324) );
  AND2_X2 U11538 ( .A1(n11104), .A2(n20680), .ZN(n16192) );
  INV_X2 U11539 ( .A(n20022), .ZN(n19299) );
  INV_X4 U11540 ( .A(n17022), .ZN(n12247) );
  INV_X2 U11541 ( .A(n17098), .ZN(n17178) );
  INV_X1 U11542 ( .A(n12208), .ZN(n14198) );
  INV_X2 U11543 ( .A(n16684), .ZN(U215) );
  INV_X1 U11544 ( .A(n17098), .ZN(n9819) );
  NOR2_X1 U11545 ( .A1(n12161), .A2(n17074), .ZN(n12245) );
  INV_X1 U11546 ( .A(n17022), .ZN(n9820) );
  NOR2_X1 U11547 ( .A1(n12156), .A2(n17074), .ZN(n12241) );
  CLKBUF_X3 U11548 ( .A(n10488), .Z(n9825) );
  INV_X1 U11549 ( .A(n12163), .ZN(n12158) );
  NAND2_X1 U11550 ( .A1(n12415), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12156) );
  NAND2_X1 U11551 ( .A1(n18925), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12160) );
  AND2_X2 U11552 ( .A1(n10314), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13491) );
  NAND2_X1 U11553 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17075) );
  AND2_X1 U11554 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12163) );
  INV_X1 U11555 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18925) );
  AND2_X2 U11556 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14894) );
  MUX2_X1 U11557 ( .A(n10396), .B(n11162), .S(n13193), .Z(n10399) );
  NAND2_X2 U11558 ( .A1(n10274), .A2(n10002), .ZN(n10273) );
  OAI21_X1 U11559 ( .B1(n14301), .B2(n11256), .A(n11255), .ZN(n14696) );
  NAND2_X1 U11560 ( .A1(n13018), .A2(n10412), .ZN(n13012) );
  NOR2_X2 U11561 ( .A1(n17912), .A2(n17895), .ZN(n17892) );
  NAND2_X2 U11562 ( .A1(n15513), .A2(n15514), .ZN(n15515) );
  NAND2_X2 U11563 ( .A1(n12781), .A2(n15685), .ZN(n15513) );
  OR2_X1 U11564 ( .A1(n10471), .A2(n10470), .ZN(n10481) );
  AOI21_X1 U11565 ( .B1(n10471), .B2(n10467), .A(n10295), .ZN(n10468) );
  XNOR2_X1 U11566 ( .A(n10471), .B(n10468), .ZN(n20413) );
  NAND2_X2 U11567 ( .A1(n10288), .A2(n9885), .ZN(n14338) );
  NAND2_X2 U11568 ( .A1(n15515), .A2(n10289), .ZN(n10288) );
  NAND3_X2 U11569 ( .A1(n13720), .A2(n9973), .A3(n12845), .ZN(n12853) );
  NOR2_X1 U11570 ( .A1(n12848), .A2(n13997), .ZN(n14004) );
  XNOR2_X1 U11571 ( .A(n12698), .B(n12697), .ZN(n12848) );
  AND2_X2 U11572 ( .A1(n13950), .A2(n13973), .ZN(n13974) );
  AND2_X1 U11573 ( .A1(n10501), .A2(n10499), .ZN(n10541) );
  NAND2_X1 U11574 ( .A1(n13031), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13032) );
  NAND2_X2 U11575 ( .A1(n12023), .A2(n10445), .ZN(n12488) );
  NOR2_X4 U11576 ( .A1(n13608), .A2(n13707), .ZN(n13711) );
  AND2_X2 U11577 ( .A1(n11265), .A2(n14755), .ZN(n14622) );
  INV_X1 U11578 ( .A(n9815), .ZN(n9823) );
  NOR2_X1 U11579 ( .A1(n12156), .A2(n12162), .ZN(n12307) );
  AND2_X1 U11580 ( .A1(n13490), .A2(n10327), .ZN(n10367) );
  NAND2_X1 U11581 ( .A1(n12522), .A2(n12523), .ZN(n13374) );
  AND2_X2 U11582 ( .A1(n13491), .A2(n14894), .ZN(n9829) );
  AND2_X2 U11583 ( .A1(n13490), .A2(n10322), .ZN(n10752) );
  AND2_X4 U11584 ( .A1(n10315), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13490) );
  AND2_X2 U11585 ( .A1(n10333), .A2(n10334), .ZN(n10506) );
  NAND2_X4 U11586 ( .A1(n11364), .A2(n11363), .ZN(n11458) );
  OR2_X1 U11588 ( .A1(n12161), .A2(n12159), .ZN(n17098) );
  OR2_X1 U11589 ( .A1(n12162), .A2(n12160), .ZN(n12229) );
  AND2_X1 U11590 ( .A1(n13490), .A2(n10333), .ZN(n9828) );
  AND2_X1 U11591 ( .A1(n13490), .A2(n10333), .ZN(n9832) );
  NAND2_X2 U11592 ( .A1(n15553), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15539) );
  AND2_X2 U11593 ( .A1(n11643), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11942) );
  MUX2_X2 U11594 ( .A(n9898), .B(n14622), .S(n14728), .Z(n14623) );
  AND2_X1 U11596 ( .A1(n13491), .A2(n14894), .ZN(n9830) );
  NAND2_X2 U11597 ( .A1(n9976), .A2(n10182), .ZN(n14301) );
  AND2_X2 U11598 ( .A1(n13490), .A2(n10333), .ZN(n9831) );
  AND2_X1 U11599 ( .A1(n13490), .A2(n10333), .ZN(n11073) );
  AND2_X1 U11600 ( .A1(n13491), .A2(n10327), .ZN(n9833) );
  AND2_X1 U11601 ( .A1(n13491), .A2(n10327), .ZN(n10421) );
  INV_X2 U11602 ( .A(n13516), .ZN(n10546) );
  XNOR2_X2 U11603 ( .A(n11195), .B(n20241), .ZN(n13570) );
  NOR2_X2 U11604 ( .A1(n14548), .A2(n14599), .ZN(n14541) );
  NAND2_X2 U11605 ( .A1(n10600), .A2(n10554), .ZN(n14890) );
  AND2_X1 U11606 ( .A1(n10327), .A2(n10334), .ZN(n9834) );
  AND2_X1 U11607 ( .A1(n10327), .A2(n10334), .ZN(n10359) );
  AND2_X1 U11608 ( .A1(n10334), .A2(n14894), .ZN(n9837) );
  AND2_X2 U11609 ( .A1(n10334), .A2(n14894), .ZN(n9838) );
  AND2_X4 U11610 ( .A1(n10332), .A2(n14894), .ZN(n10366) );
  AND2_X1 U11611 ( .A1(n13491), .A2(n10333), .ZN(n9840) );
  AND2_X2 U11612 ( .A1(n13491), .A2(n10333), .ZN(n9841) );
  AND2_X1 U11613 ( .A1(n13491), .A2(n10322), .ZN(n9845) );
  AND2_X1 U11614 ( .A1(n13491), .A2(n10322), .ZN(n10708) );
  NAND2_X2 U11615 ( .A1(n14443), .A2(n14444), .ZN(n14430) );
  NOR2_X4 U11616 ( .A1(n14457), .A2(n14458), .ZN(n14443) );
  NAND2_X2 U11617 ( .A1(n10374), .A2(n10413), .ZN(n10416) );
  AOI21_X2 U11618 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14627) );
  XNOR2_X1 U11619 ( .A(n10563), .B(n10562), .ZN(n13515) );
  INV_X1 U11620 ( .A(n10677), .ZN(n10040) );
  OR2_X1 U11621 ( .A1(n12860), .A2(n12859), .ZN(n12862) );
  NOR2_X1 U11622 ( .A1(n17075), .A2(n12160), .ZN(n12240) );
  NAND2_X1 U11623 ( .A1(n10412), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10587) );
  INV_X1 U11624 ( .A(n11143), .ZN(n11122) );
  NAND2_X1 U11625 ( .A1(n11477), .A2(n20028), .ZN(n11463) );
  NAND2_X1 U11626 ( .A1(n11273), .A2(n10164), .ZN(n10163) );
  INV_X1 U11627 ( .A(n14431), .ZN(n10164) );
  OR2_X1 U11628 ( .A1(n14059), .A2(n14073), .ZN(n10159) );
  INV_X1 U11629 ( .A(n13951), .ZN(n10149) );
  INV_X1 U11630 ( .A(n12030), .ZN(n11098) );
  OR2_X1 U11631 ( .A1(n12492), .A2(n20964), .ZN(n10812) );
  NOR2_X1 U11632 ( .A1(n11266), .A2(n14745), .ZN(n10043) );
  INV_X1 U11633 ( .A(n11224), .ZN(n11194) );
  NAND2_X1 U11634 ( .A1(n20274), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U11635 ( .A1(n9894), .A2(n10570), .ZN(n10036) );
  INV_X1 U11636 ( .A(n10600), .ZN(n10029) );
  AOI21_X1 U11637 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19980), .A(
        n11600), .ZN(n11610) );
  OR2_X1 U11638 ( .A1(n15220), .A2(n15219), .ZN(n15221) );
  AND2_X1 U11639 ( .A1(n10241), .A2(n13645), .ZN(n10240) );
  INV_X1 U11640 ( .A(n11508), .ZN(n10000) );
  NOR2_X1 U11641 ( .A1(n10056), .A2(n10051), .ZN(n10050) );
  INV_X1 U11642 ( .A(n14281), .ZN(n11593) );
  AND2_X1 U11643 ( .A1(n10291), .A2(n10058), .ZN(n10057) );
  AND2_X1 U11644 ( .A1(n12724), .A2(n10292), .ZN(n10291) );
  AND4_X1 U11645 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11783) );
  INV_X1 U11646 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n21204) );
  NOR2_X1 U11647 ( .A1(n16696), .A2(n12405), .ZN(n15929) );
  AND2_X1 U11648 ( .A1(n12401), .A2(n18773), .ZN(n14103) );
  NAND2_X1 U11649 ( .A1(n20964), .A2(n20965), .ZN(n12030) );
  NAND2_X1 U11650 ( .A1(n13417), .A2(n10580), .ZN(n13545) );
  NAND2_X1 U11651 ( .A1(n12491), .A2(n12490), .ZN(n13200) );
  OR3_X1 U11652 ( .A1(n13276), .A2(n12021), .A3(n20042), .ZN(n13308) );
  INV_X1 U11653 ( .A(n11093), .ZN(n11100) );
  OR2_X1 U11654 ( .A1(n13276), .A2(n13033), .ZN(n15980) );
  NAND2_X1 U11655 ( .A1(n13017), .A2(n13201), .ZN(n13041) );
  NAND2_X1 U11656 ( .A1(n9846), .A2(n11174), .ZN(n20755) );
  NOR2_X1 U11657 ( .A1(n20009), .A2(n12931), .ZN(n12825) );
  AND2_X1 U11658 ( .A1(n9909), .A2(n13640), .ZN(n10211) );
  NAND2_X1 U11659 ( .A1(n10003), .A2(n10264), .ZN(n16400) );
  AOI21_X1 U11660 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(n10264) );
  INV_X1 U11661 ( .A(n16401), .ZN(n10265) );
  NOR2_X1 U11662 ( .A1(n16374), .A2(n10056), .ZN(n10028) );
  CLKBUF_X3 U11663 ( .A(n11988), .Z(n15191) );
  INV_X1 U11664 ( .A(n16553), .ZN(n13295) );
  INV_X1 U11665 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16540) );
  NOR2_X1 U11666 ( .A1(n17581), .A2(n15929), .ZN(n18761) );
  NOR2_X2 U11667 ( .A1(n12313), .A2(n12312), .ZN(n18972) );
  NOR2_X1 U11668 ( .A1(n17658), .A2(n10062), .ZN(n12293) );
  INV_X1 U11669 ( .A(n11997), .ZN(n12018) );
  NAND2_X1 U11670 ( .A1(n17343), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17338) );
  AND2_X2 U11671 ( .A1(n10316), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10322) );
  NAND2_X1 U11672 ( .A1(n10650), .A2(n10649), .ZN(n10662) );
  NAND2_X1 U11673 ( .A1(n10622), .A2(n10621), .ZN(n10637) );
  INV_X1 U11674 ( .A(n12001), .ZN(n10243) );
  AND4_X1 U11675 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11766) );
  NAND2_X1 U11676 ( .A1(n11986), .A2(n15216), .ZN(n11501) );
  NAND2_X1 U11677 ( .A1(n12645), .A2(n12644), .ZN(n12697) );
  NAND2_X1 U11678 ( .A1(n19636), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12547) );
  AOI21_X1 U11679 ( .B1(n19411), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12599), .ZN(n12606) );
  NOR2_X1 U11680 ( .A1(n11617), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11618) );
  NOR2_X1 U11681 ( .A1(n14549), .A2(n10153), .ZN(n10150) );
  NOR2_X1 U11682 ( .A1(n10110), .A2(n14451), .ZN(n10109) );
  INV_X1 U11683 ( .A(n10111), .ZN(n10110) );
  NOR2_X1 U11684 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  INV_X1 U11685 ( .A(n14316), .ZN(n10117) );
  OR2_X1 U11686 ( .A1(n10119), .A2(n14062), .ZN(n10118) );
  INV_X1 U11687 ( .A(n14089), .ZN(n10119) );
  INV_X1 U11688 ( .A(n16182), .ZN(n9978) );
  INV_X1 U11689 ( .A(n10185), .ZN(n10184) );
  INV_X1 U11690 ( .A(n11238), .ZN(n10183) );
  NAND2_X1 U11691 ( .A1(n10638), .A2(n10038), .ZN(n10678) );
  NAND2_X1 U11692 ( .A1(n13349), .A2(n12121), .ZN(n12122) );
  AND2_X1 U11693 ( .A1(n12047), .A2(n12039), .ZN(n10123) );
  INV_X1 U11694 ( .A(n13418), .ZN(n12047) );
  OR2_X1 U11695 ( .A1(n10512), .A2(n10511), .ZN(n11235) );
  OR2_X1 U11696 ( .A1(n10587), .A2(n11191), .ZN(n10495) );
  NOR2_X1 U11697 ( .A1(n13029), .A2(n13030), .ZN(n13189) );
  NAND2_X1 U11698 ( .A1(n12817), .A2(n10306), .ZN(n11452) );
  AND3_X1 U11699 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11610), .A3(
        n13100), .ZN(n12912) );
  NAND2_X1 U11700 ( .A1(n16299), .A2(n12797), .ZN(n12809) );
  AND2_X1 U11701 ( .A1(n10244), .A2(n10242), .ZN(n12659) );
  INV_X1 U11702 ( .A(n12975), .ZN(n10219) );
  AND2_X1 U11703 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  INV_X1 U11704 ( .A(n15392), .ZN(n10209) );
  AND2_X1 U11705 ( .A1(n13466), .A2(n13427), .ZN(n10225) );
  NOR2_X1 U11706 ( .A1(n12666), .A2(n16479), .ZN(n10279) );
  NAND2_X1 U11707 ( .A1(n16374), .A2(n16373), .ZN(n10284) );
  AND2_X1 U11708 ( .A1(n10285), .A2(n10054), .ZN(n10053) );
  NAND2_X1 U11709 ( .A1(n10055), .A2(n12729), .ZN(n10054) );
  NOR2_X1 U11710 ( .A1(n12778), .A2(n10286), .ZN(n10285) );
  INV_X1 U11711 ( .A(n10057), .ZN(n10055) );
  AND2_X1 U11712 ( .A1(n15037), .A2(n10229), .ZN(n15017) );
  AND2_X1 U11713 ( .A1(n10230), .A2(n9955), .ZN(n10229) );
  AND2_X1 U11714 ( .A1(n10228), .A2(n13943), .ZN(n10227) );
  INV_X1 U11715 ( .A(n14019), .ZN(n10228) );
  OR2_X1 U11716 ( .A1(n13805), .A2(n14364), .ZN(n12735) );
  NOR2_X1 U11717 ( .A1(n13830), .A2(n10235), .ZN(n10234) );
  INV_X1 U11718 ( .A(n14038), .ZN(n10235) );
  NAND2_X1 U11719 ( .A1(n9852), .A2(n10016), .ZN(n10013) );
  NAND2_X1 U11720 ( .A1(n9971), .A2(n10004), .ZN(n12829) );
  INV_X1 U11721 ( .A(n11506), .ZN(n9970) );
  AOI21_X1 U11722 ( .B1(n13222), .B2(n11709), .A(n11708), .ZN(n11712) );
  NAND2_X1 U11723 ( .A1(n13268), .A2(n13267), .ZN(n13384) );
  NOR2_X1 U11724 ( .A1(n15261), .A2(n19336), .ZN(n13380) );
  NAND2_X1 U11725 ( .A1(n12560), .A2(n12543), .ZN(n12536) );
  NAND2_X1 U11726 ( .A1(n16502), .A2(n13228), .ZN(n12567) );
  INV_X1 U11727 ( .A(n12566), .ZN(n10005) );
  AND4_X1 U11728 ( .A1(n11356), .A2(n11355), .A3(n11354), .A4(n11353), .ZN(
        n11357) );
  NAND3_X1 U11729 ( .A1(n19971), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19833), 
        .ZN(n13629) );
  INV_X1 U11730 ( .A(n12244), .ZN(n12318) );
  NAND2_X1 U11731 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12414), .ZN(
        n12162) );
  NOR2_X1 U11732 ( .A1(n12162), .A2(n12158), .ZN(n12208) );
  INV_X1 U11733 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U11734 ( .A1(n18367), .A2(n18346), .ZN(n12403) );
  NAND2_X1 U11735 ( .A1(n10102), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10101) );
  INV_X1 U11736 ( .A(n9877), .ZN(n10102) );
  AND2_X1 U11737 ( .A1(n12269), .A2(n12456), .ZN(n12272) );
  AND2_X1 U11738 ( .A1(n12280), .A2(n10077), .ZN(n10076) );
  NOR2_X1 U11739 ( .A1(n17927), .A2(n12271), .ZN(n12274) );
  NAND2_X1 U11740 ( .A1(n10066), .A2(n10065), .ZN(n12262) );
  NAND2_X1 U11741 ( .A1(n9875), .A2(n17969), .ZN(n10066) );
  AND2_X1 U11742 ( .A1(n12412), .A2(n12398), .ZN(n15933) );
  NOR2_X1 U11743 ( .A1(n18354), .A2(n18361), .ZN(n18774) );
  NOR2_X1 U11744 ( .A1(n12367), .A2(n12366), .ZN(n12390) );
  NAND2_X1 U11745 ( .A1(n15933), .A2(n18774), .ZN(n15940) );
  INV_X1 U11746 ( .A(n13349), .ZN(n13059) );
  NAND2_X1 U11747 ( .A1(n12049), .A2(n12121), .ZN(n13333) );
  NOR2_X1 U11748 ( .A1(n13280), .A2(n13309), .ZN(n12496) );
  AND4_X1 U11749 ( .A1(n12495), .A2(n12494), .A3(n20342), .A4(n12493), .ZN(
        n13350) );
  NOR2_X1 U11750 ( .A1(n11105), .A2(n14618), .ZN(n11106) );
  INV_X1 U11751 ( .A(n10810), .ZN(n11099) );
  INV_X1 U11752 ( .A(n10162), .ZN(n10160) );
  OAI21_X1 U11753 ( .B1(n14633), .B2(n12030), .A(n11031), .ZN(n14431) );
  AND2_X1 U11754 ( .A1(n10798), .A2(n10159), .ZN(n10158) );
  NAND2_X1 U11755 ( .A1(n10673), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10682) );
  NOR2_X1 U11756 ( .A1(n10558), .A2(n10303), .ZN(n10559) );
  NOR2_X2 U11757 ( .A1(n14434), .A2(n14233), .ZN(n14418) );
  NAND2_X1 U11758 ( .A1(n10034), .A2(n16173), .ZN(n14670) );
  NAND2_X1 U11759 ( .A1(n11262), .A2(n14728), .ZN(n14669) );
  NAND2_X1 U11760 ( .A1(n14301), .A2(n11255), .ZN(n10032) );
  OR2_X1 U11761 ( .A1(n16173), .A2(n11243), .ZN(n14714) );
  OR2_X1 U11762 ( .A1(n20248), .A2(n14878), .ZN(n16238) );
  NAND2_X1 U11763 ( .A1(n16197), .A2(n16196), .ZN(n16195) );
  OR2_X1 U11764 ( .A1(n14890), .A2(n11194), .ZN(n11187) );
  INV_X1 U11765 ( .A(n20248), .ZN(n16236) );
  NAND2_X1 U11766 ( .A1(n10551), .A2(n10550), .ZN(n10552) );
  INV_X1 U11767 ( .A(n20346), .ZN(n20454) );
  AND2_X1 U11768 ( .A1(n12023), .A2(n12022), .ZN(n13065) );
  NAND2_X1 U11769 ( .A1(n11159), .A2(n11158), .ZN(n13276) );
  INV_X1 U11770 ( .A(n20534), .ZN(n20528) );
  NAND2_X1 U11771 ( .A1(n20556), .A2(n14890), .ZN(n20655) );
  INV_X1 U11772 ( .A(n20800), .ZN(n20757) );
  OR2_X1 U11773 ( .A1(n14890), .A2(n20264), .ZN(n20800) );
  AOI21_X1 U11774 ( .B1(n20952), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20454), 
        .ZN(n20801) );
  AND2_X1 U11775 ( .A1(n20857), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15995) );
  NOR2_X1 U11776 ( .A1(n16521), .A2(n16519), .ZN(n13092) );
  NOR2_X1 U11777 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20018) );
  CLKBUF_X1 U11778 ( .A(n12817), .Z(n12818) );
  NOR2_X1 U11779 ( .A1(n14928), .A2(n19117), .ZN(n10129) );
  OR3_X1 U11780 ( .A1(n10247), .A2(n12740), .A3(P2_EBX_REG_20__SCAN_IN), .ZN(
        n10245) );
  AND2_X1 U11781 ( .A1(n13589), .A2(n13588), .ZN(n13590) );
  NAND2_X1 U11782 ( .A1(n10200), .A2(n15305), .ZN(n10199) );
  INV_X1 U11783 ( .A(n9943), .ZN(n10200) );
  AND2_X1 U11784 ( .A1(n11970), .A2(n11969), .ZN(n14971) );
  AND2_X1 U11785 ( .A1(n13784), .A2(n13760), .ZN(n10210) );
  NOR2_X1 U11786 ( .A1(n15835), .A2(n15836), .ZN(n15822) );
  CLKBUF_X1 U11787 ( .A(n11663), .Z(n13301) );
  NAND2_X1 U11788 ( .A1(n11300), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11323) );
  AND2_X1 U11789 ( .A1(n13617), .A2(n9916), .ZN(n13726) );
  AND2_X1 U11790 ( .A1(n16376), .A2(n16430), .ZN(n16360) );
  AND2_X1 U11791 ( .A1(n13617), .A2(n10240), .ZN(n13648) );
  AND2_X1 U11792 ( .A1(n13551), .A2(n13565), .ZN(n13617) );
  NAND2_X1 U11793 ( .A1(n14026), .A2(n14036), .ZN(n10269) );
  AND2_X1 U11794 ( .A1(n12861), .A2(n12862), .ZN(n16401) );
  INV_X1 U11795 ( .A(n14026), .ZN(n10268) );
  AND2_X1 U11796 ( .A1(n14935), .A2(n9949), .ZN(n14283) );
  INV_X1 U11797 ( .A(n11594), .ZN(n10236) );
  INV_X1 U11798 ( .A(n12646), .ZN(n14364) );
  NAND2_X1 U11799 ( .A1(n14293), .A2(n14292), .ZN(n14294) );
  NAND2_X1 U11800 ( .A1(n15466), .A2(n10046), .ZN(n10048) );
  NOR2_X1 U11801 ( .A1(n14363), .A2(n10047), .ZN(n10046) );
  INV_X1 U11802 ( .A(n15464), .ZN(n10047) );
  NAND2_X1 U11803 ( .A1(n14935), .A2(n9861), .ZN(n14914) );
  AND2_X1 U11804 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15657), .ZN(
        n15644) );
  NOR2_X1 U11805 ( .A1(n15012), .A2(n14996), .ZN(n14998) );
  OR2_X1 U11806 ( .A1(n15539), .A2(n10262), .ZN(n15540) );
  AND2_X1 U11807 ( .A1(n10026), .A2(n15522), .ZN(n10025) );
  NAND3_X1 U11808 ( .A1(n12852), .A2(n12850), .A3(n12851), .ZN(n13956) );
  OR2_X1 U11809 ( .A1(n12854), .A2(n9872), .ZN(n12850) );
  NAND2_X1 U11810 ( .A1(n12843), .A2(n9972), .ZN(n12845) );
  INV_X1 U11811 ( .A(n12844), .ZN(n9972) );
  NAND2_X1 U11812 ( .A1(n12653), .A2(n13701), .ZN(n10280) );
  INV_X1 U11813 ( .A(n11942), .ZN(n13913) );
  AOI21_X1 U11814 ( .B1(n13119), .B2(n13376), .A(n13118), .ZN(n13270) );
  XNOR2_X1 U11815 ( .A(n13300), .B(n11672), .ZN(n13224) );
  OR2_X1 U11816 ( .A1(n19150), .A2(n13072), .ZN(n13074) );
  AND2_X1 U11817 ( .A1(n19972), .A2(n19158), .ZN(n19436) );
  NAND2_X1 U11818 ( .A1(n19972), .A2(n20002), .ZN(n19546) );
  NOR2_X2 U11820 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19971) );
  OR2_X1 U11821 ( .A1(n19972), .A2(n19158), .ZN(n19780) );
  NOR2_X1 U11822 ( .A1(n13789), .A2(n13629), .ZN(n19352) );
  NOR2_X1 U11823 ( .A1(n15399), .A2(n13629), .ZN(n19353) );
  OAI22_X2 U11824 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19965), .B1(n19238), 
        .B2(n20024), .ZN(n19833) );
  INV_X1 U11825 ( .A(n19833), .ZN(n19576) );
  OAI221_X1 U11826 ( .B1(n15938), .B2(n17581), .C1(n15938), .C2(n18338), .A(
        n15937), .ZN(n16023) );
  INV_X1 U11827 ( .A(n18760), .ZN(n15938) );
  INV_X1 U11828 ( .A(n17684), .ZN(n17673) );
  INV_X1 U11829 ( .A(n10101), .ZN(n10099) );
  NOR2_X1 U11830 ( .A1(n17856), .A2(n17859), .ZN(n10103) );
  NOR2_X1 U11831 ( .A1(n17939), .A2(n17940), .ZN(n17920) );
  NAND2_X1 U11832 ( .A1(n16596), .A2(n10072), .ZN(n10071) );
  NAND2_X1 U11833 ( .A1(n16596), .A2(n21268), .ZN(n10073) );
  OAI22_X1 U11834 ( .A1(n17649), .A2(n10070), .B1(n17648), .B2(n10069), .ZN(
        n15961) );
  OR2_X1 U11835 ( .A1(n10073), .A2(n16571), .ZN(n10070) );
  OR2_X1 U11836 ( .A1(n10071), .A2(n16571), .ZN(n10069) );
  NAND2_X1 U11837 ( .A1(n10063), .A2(n9920), .ZN(n10062) );
  INV_X1 U11838 ( .A(n17679), .ZN(n9993) );
  NAND3_X1 U11839 ( .A1(n12172), .A2(n12171), .A3(n12170), .ZN(n15959) );
  OAI21_X1 U11840 ( .B1(n9987), .B2(n12263), .A(n9988), .ZN(n9986) );
  OAI21_X1 U11841 ( .B1(n12407), .B2(n12406), .A(n18761), .ZN(n12408) );
  NOR2_X1 U11842 ( .A1(n18819), .A2(n18822), .ZN(n18967) );
  AND2_X1 U11843 ( .A1(n12137), .A2(n12144), .ZN(n20097) );
  OR2_X1 U11844 ( .A1(n20970), .A2(n12033), .ZN(n20123) );
  INV_X1 U11845 ( .A(n20097), .ZN(n20140) );
  INV_X1 U11846 ( .A(n14600), .ZN(n14609) );
  INV_X1 U11847 ( .A(n14693), .ZN(n20222) );
  AND2_X1 U11848 ( .A1(n14693), .A2(n11166), .ZN(n16169) );
  OR2_X1 U11849 ( .A1(n15980), .A2(n20042), .ZN(n20048) );
  XNOR2_X1 U11850 ( .A(n10035), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14203) );
  NAND2_X1 U11851 ( .A1(n9879), .A2(n10172), .ZN(n10035) );
  INV_X1 U11852 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20687) );
  INV_X1 U11853 ( .A(n10561), .ZN(n10563) );
  CLKBUF_X1 U11854 ( .A(n13516), .Z(n20559) );
  NOR2_X2 U11855 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20680) );
  INV_X1 U11856 ( .A(n20855), .ZN(n20835) );
  OR2_X1 U11857 ( .A1(n16521), .A2(n11987), .ZN(n13079) );
  OR2_X1 U11858 ( .A1(n12927), .A2(n12827), .ZN(n13052) );
  INV_X1 U11859 ( .A(n14284), .ZN(n11327) );
  NAND2_X1 U11860 ( .A1(n10129), .A2(n15471), .ZN(n10128) );
  INV_X1 U11861 ( .A(n14921), .ZN(n10126) );
  NOR2_X1 U11862 ( .A1(n10129), .A2(n15471), .ZN(n14920) );
  CLKBUF_X1 U11863 ( .A(n11324), .Z(n19136) );
  XNOR2_X1 U11864 ( .A(n14289), .B(n14288), .ZN(n19163) );
  AND2_X1 U11865 ( .A1(n14289), .A2(n11985), .ZN(n15405) );
  NAND2_X1 U11866 ( .A1(n19301), .A2(n20022), .ZN(n19256) );
  INV_X1 U11867 ( .A(n19233), .ZN(n19305) );
  NAND2_X1 U11868 ( .A1(n15405), .A2(n19310), .ZN(n14396) );
  NAND2_X1 U11869 ( .A1(n12974), .A2(n20011), .ZN(n19316) );
  NAND2_X1 U11870 ( .A1(n12974), .A2(n12970), .ZN(n19312) );
  AND2_X1 U11871 ( .A1(n12974), .A2(n12973), .ZN(n19310) );
  INV_X1 U11872 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19996) );
  INV_X1 U11873 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19980) );
  INV_X1 U11874 ( .A(n15950), .ZN(n18958) );
  NAND2_X1 U11875 ( .A1(n17371), .A2(n17390), .ZN(n10181) );
  NAND2_X1 U11876 ( .A1(n17119), .A2(n9956), .ZN(n15921) );
  NAND2_X1 U11877 ( .A1(n17121), .A2(n17356), .ZN(n17119) );
  AND2_X1 U11878 ( .A1(n17137), .A2(n9869), .ZN(n17129) );
  NOR2_X1 U11879 ( .A1(n17091), .A2(n17161), .ZN(n17137) );
  NOR2_X1 U11880 ( .A1(n18367), .A2(n10192), .ZN(n10190) );
  AND2_X1 U11881 ( .A1(n17294), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17267) );
  NOR2_X1 U11882 ( .A1(n17297), .A2(n17338), .ZN(n17294) );
  NOR2_X1 U11883 ( .A1(n17352), .A2(n10194), .ZN(n17343) );
  INV_X1 U11884 ( .A(n17371), .ZN(n17356) );
  AOI21_X1 U11885 ( .B1(n11074), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A(n9953), .ZN(n11060) );
  AOI21_X1 U11886 ( .B1(n11074), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n9907), .ZN(n10644) );
  AOI21_X1 U11887 ( .B1(n10910), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(n9908), .ZN(n10612) );
  AND2_X1 U11888 ( .A1(n10414), .A2(n13353), .ZN(n10457) );
  AOI22_X1 U11889 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11628), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11421) );
  OAI21_X1 U11890 ( .B1(n12674), .B2(n12673), .A(n9969), .ZN(n12675) );
  NAND2_X1 U11891 ( .A1(n19636), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n9969) );
  AND3_X1 U11892 ( .A1(n11383), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11382), .ZN(n11387) );
  AND2_X1 U11893 ( .A1(n20952), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11120) );
  AOI21_X1 U11894 ( .B1(n11074), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A(n9938), .ZN(n10962) );
  AOI21_X1 U11895 ( .B1(n11074), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A(n9937), .ZN(n10936) );
  AOI21_X1 U11896 ( .B1(n10916), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n9934), .ZN(n10946) );
  AOI21_X1 U11897 ( .B1(n10366), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A(n9940), .ZN(n10788) );
  NOR2_X1 U11898 ( .A1(n10041), .A2(n10039), .ZN(n10038) );
  INV_X1 U11899 ( .A(n10662), .ZN(n10041) );
  INV_X1 U11900 ( .A(n10637), .ZN(n10039) );
  AOI21_X1 U11901 ( .B1(n11055), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n9881), .ZN(n10510) );
  AOI21_X1 U11902 ( .B1(n9821), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(n9882), .ZN(n10529) );
  OAI211_X1 U11903 ( .C1(n13306), .C2(n10412), .A(n10438), .B(n10439), .ZN(
        n10168) );
  NAND2_X1 U11904 ( .A1(n11122), .A2(n11224), .ZN(n11150) );
  AOI21_X1 U11905 ( .B1(n10752), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A(n9889), .ZN(n10376) );
  AND2_X1 U11906 ( .A1(n11601), .A2(n11602), .ZN(n11600) );
  INV_X1 U11907 ( .A(n15123), .ZN(n10218) );
  NAND2_X1 U11908 ( .A1(n15879), .A2(n11408), .ZN(n15123) );
  NAND2_X1 U11909 ( .A1(n12911), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10206) );
  AND4_X1 U11910 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11785) );
  INV_X1 U11911 ( .A(n11435), .ZN(n12920) );
  NOR2_X1 U11912 ( .A1(n12882), .A2(n11447), .ZN(n12936) );
  INV_X1 U11913 ( .A(n12567), .ZN(n12568) );
  NAND2_X1 U11914 ( .A1(n12413), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12159) );
  NOR2_X1 U11915 ( .A1(n17500), .A2(n12267), .ZN(n12269) );
  NAND2_X1 U11916 ( .A1(n12257), .A2(n17520), .ZN(n12260) );
  NAND2_X1 U11917 ( .A1(n12402), .A2(n15944), .ZN(n12398) );
  AOI22_X1 U11918 ( .A1(n10708), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U11919 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9832), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10409) );
  NOR2_X1 U11920 ( .A1(n10163), .A2(n14421), .ZN(n10162) );
  NOR2_X1 U11921 ( .A1(n14583), .A2(n10156), .ZN(n10155) );
  INV_X1 U11922 ( .A(n10157), .ZN(n10156) );
  NOR2_X1 U11923 ( .A1(n14525), .A2(n10909), .ZN(n10157) );
  AOI21_X1 U11924 ( .B1(n10916), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n9952), .ZN(n10883) );
  OR2_X1 U11925 ( .A1(n10844), .A2(n14477), .ZN(n10859) );
  AOI21_X1 U11926 ( .B1(n11074), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n9939), .ZN(n10836) );
  INV_X1 U11927 ( .A(n14083), .ZN(n10154) );
  AOI21_X1 U11928 ( .B1(n10916), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n9935), .ZN(n10729) );
  NAND2_X1 U11929 ( .A1(n10703), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10719) );
  AOI21_X1 U11930 ( .B1(n11075), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A(n9936), .ZN(n10711) );
  NAND2_X1 U11931 ( .A1(n10638), .A2(n10637), .ZN(n10661) );
  AND2_X1 U11932 ( .A1(n10627), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10652) );
  OR2_X1 U11933 ( .A1(n10597), .A2(n10596), .ZN(n11206) );
  OR2_X1 U11934 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10176) );
  NOR2_X1 U11935 ( .A1(n10113), .A2(n10112), .ZN(n10111) );
  INV_X1 U11936 ( .A(n14518), .ZN(n10112) );
  INV_X1 U11937 ( .A(n14459), .ZN(n10113) );
  NAND2_X1 U11938 ( .A1(n11250), .A2(n11249), .ZN(n11256) );
  NAND2_X1 U11939 ( .A1(n10107), .A2(n9887), .ZN(n10106) );
  INV_X1 U11940 ( .A(n16273), .ZN(n10107) );
  NAND2_X1 U11941 ( .A1(n11182), .A2(n11181), .ZN(n10167) );
  INV_X1 U11942 ( .A(n10587), .ZN(n10545) );
  NOR2_X1 U11943 ( .A1(n10494), .A2(n10493), .ZN(n11191) );
  AND3_X1 U11944 ( .A1(n10540), .A2(n10539), .A3(n10538), .ZN(n10547) );
  NAND2_X1 U11945 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U11946 ( .A1(n9975), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9974) );
  INV_X1 U11947 ( .A(n11150), .ZN(n11154) );
  NAND2_X1 U11948 ( .A1(n10587), .A2(n10586), .ZN(n11157) );
  NAND2_X1 U11949 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10331) );
  INV_X1 U11950 ( .A(n20447), .ZN(n20264) );
  AOI21_X1 U11951 ( .B1(n20967), .B2(n16289), .A(n15999), .ZN(n20273) );
  OR2_X1 U11952 ( .A1(n12935), .A2(n12934), .ZN(n15877) );
  INV_X1 U11953 ( .A(n12003), .ZN(n12907) );
  OR2_X1 U11954 ( .A1(n16294), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12798) );
  INV_X1 U11955 ( .A(n15507), .ZN(n10138) );
  INV_X1 U11956 ( .A(n12738), .ZN(n10247) );
  NOR2_X1 U11957 ( .A1(n10253), .A2(n10256), .ZN(n10252) );
  INV_X1 U11958 ( .A(n12009), .ZN(n10256) );
  INV_X1 U11959 ( .A(n10254), .ZN(n10253) );
  NOR2_X1 U11960 ( .A1(n12761), .A2(n10255), .ZN(n10254) );
  INV_X1 U11961 ( .A(n12732), .ZN(n10255) );
  NAND2_X1 U11962 ( .A1(n12723), .A2(n12732), .ZN(n12763) );
  NOR2_X1 U11963 ( .A1(n12717), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U11964 ( .A1(n12730), .A2(n12794), .ZN(n12723) );
  NAND2_X1 U11965 ( .A1(n12701), .A2(n12705), .ZN(n10250) );
  NOR3_X1 U11966 ( .A1(n12667), .A2(n12647), .A3(n10251), .ZN(n12707) );
  NOR2_X1 U11967 ( .A1(n12667), .A2(n12647), .ZN(n12702) );
  AND3_X1 U11968 ( .A1(n10242), .A2(n12652), .A3(n10244), .ZN(n12668) );
  NAND2_X1 U11969 ( .A1(n12669), .A2(n12668), .ZN(n12667) );
  NAND2_X1 U11970 ( .A1(n10218), .A2(n11637), .ZN(n11799) );
  AND2_X1 U11972 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11622), .ZN(
        n15145) );
  INV_X1 U11973 ( .A(n14940), .ZN(n10220) );
  NAND2_X1 U11974 ( .A1(n15349), .A2(n10195), .ZN(n15265) );
  INV_X1 U11975 ( .A(n15388), .ZN(n10208) );
  AND2_X1 U11976 ( .A1(n15038), .A2(n13787), .ZN(n10232) );
  INV_X1 U11977 ( .A(n15216), .ZN(n15261) );
  NOR2_X1 U11978 ( .A1(n11285), .A2(n10141), .ZN(n10140) );
  INV_X1 U11979 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U11980 ( .A1(n16389), .A2(n10132), .ZN(n10131) );
  INV_X1 U11981 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U11982 ( .A1(n19127), .A2(n10144), .ZN(n10147) );
  INV_X1 U11983 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U11984 ( .A1(n14345), .A2(n12011), .ZN(n14293) );
  INV_X1 U11985 ( .A(n14911), .ZN(n10237) );
  OR2_X1 U11986 ( .A1(n16299), .A2(n14364), .ZN(n12801) );
  NOR2_X1 U11987 ( .A1(n15501), .A2(n10290), .ZN(n10289) );
  INV_X1 U11988 ( .A(n15376), .ZN(n10223) );
  OR2_X1 U11989 ( .A1(n10261), .A2(n15669), .ZN(n10260) );
  NAND2_X1 U11990 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10261) );
  AND2_X1 U11991 ( .A1(n15000), .A2(n14986), .ZN(n10239) );
  AND2_X1 U11992 ( .A1(n10232), .A2(n10231), .ZN(n10230) );
  INV_X1 U11993 ( .A(n15026), .ZN(n10231) );
  AOI21_X1 U11994 ( .B1(n10023), .B2(n15768), .A(n10022), .ZN(n10021) );
  INV_X1 U11995 ( .A(n15583), .ZN(n10022) );
  OR2_X1 U11996 ( .A1(n10028), .A2(n10286), .ZN(n10026) );
  AND2_X1 U11997 ( .A1(n13616), .A2(n13584), .ZN(n10241) );
  AND2_X1 U11998 ( .A1(n15831), .A2(n15605), .ZN(n10292) );
  INV_X1 U11999 ( .A(n16404), .ZN(n10058) );
  NOR2_X1 U12000 ( .A1(n12846), .A2(n14004), .ZN(n12849) );
  INV_X1 U12001 ( .A(n14004), .ZN(n12854) );
  AND3_X1 U12002 ( .A1(n11750), .A2(n11749), .A3(n11748), .ZN(n12643) );
  AND4_X1 U12003 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11749) );
  AND4_X1 U12004 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11750) );
  AND3_X1 U12005 ( .A1(n11705), .A2(n11704), .A3(n11703), .ZN(n12837) );
  AND4_X1 U12006 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11704) );
  AND4_X1 U12007 ( .A1(n11702), .A2(n11701), .A3(n11700), .A4(n11699), .ZN(
        n11703) );
  AND4_X1 U12008 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11705) );
  AND2_X1 U12009 ( .A1(n19237), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13376) );
  NOR2_X1 U12010 ( .A1(n13252), .A2(n11712), .ZN(n13699) );
  NOR2_X1 U12011 ( .A1(n15261), .A2(n15903), .ZN(n13267) );
  AND2_X1 U12012 ( .A1(n13264), .A2(n15895), .ZN(n19468) );
  INV_X1 U12013 ( .A(n12685), .ZN(n19721) );
  INV_X1 U12014 ( .A(n12245), .ZN(n12337) );
  NAND2_X1 U12015 ( .A1(n9997), .A2(n9996), .ZN(n12280) );
  NOR2_X1 U12016 ( .A1(n12275), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9996) );
  INV_X1 U12017 ( .A(n17914), .ZN(n9997) );
  INV_X1 U12018 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14477) );
  INV_X1 U12019 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20065) );
  AND2_X1 U12020 ( .A1(n16082), .A2(n14538), .ZN(n14540) );
  AND3_X1 U12021 ( .A1(n12096), .A2(n12101), .A3(n12095), .ZN(n14545) );
  NAND2_X1 U12022 ( .A1(n12483), .A2(n10162), .ZN(n10161) );
  NAND2_X1 U12023 ( .A1(n11049), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11051) );
  INV_X1 U12024 ( .A(n11032), .ZN(n11049) );
  AND2_X1 U12025 ( .A1(n10928), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10929) );
  NAND2_X1 U12026 ( .A1(n10891), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10892) );
  INV_X1 U12027 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10904) );
  NOR2_X1 U12028 ( .A1(n10859), .A2(n14692), .ZN(n10860) );
  AND2_X1 U12029 ( .A1(n10860), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10891) );
  CLKBUF_X1 U12030 ( .A(n14548), .Z(n14598) );
  NAND2_X1 U12031 ( .A1(n10831), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10844) );
  NOR2_X1 U12032 ( .A1(n14084), .A2(n14083), .ZN(n14473) );
  NOR2_X1 U12033 ( .A1(n10817), .A2(n16114), .ZN(n10831) );
  NAND2_X1 U12034 ( .A1(n10799), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10817) );
  NOR2_X1 U12035 ( .A1(n10768), .A2(n14323), .ZN(n10799) );
  AND2_X1 U12036 ( .A1(n13974), .A2(n10159), .ZN(n14048) );
  AND2_X1 U12037 ( .A1(n14058), .A2(n14060), .ZN(n14074) );
  NOR2_X1 U12038 ( .A1(n21212), .A2(n10720), .ZN(n10738) );
  AND3_X1 U12039 ( .A1(n10701), .A2(n10700), .A3(n10699), .ZN(n13737) );
  NOR2_X1 U12040 ( .A1(n10682), .A2(n20076), .ZN(n10703) );
  AOI21_X1 U12041 ( .B1(n11214), .B2(n10761), .A(n10676), .ZN(n13707) );
  AND2_X1 U12042 ( .A1(n10652), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10673) );
  INV_X1 U12043 ( .A(n13576), .ZN(n10634) );
  AND2_X1 U12044 ( .A1(n13347), .A2(n10580), .ZN(n10148) );
  NOR2_X1 U12045 ( .A1(n10176), .A2(n10174), .ZN(n10173) );
  INV_X1 U12046 ( .A(n11267), .ZN(n10174) );
  INV_X1 U12047 ( .A(n10176), .ZN(n10175) );
  AND2_X1 U12048 ( .A1(n10043), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10042) );
  AND2_X1 U12049 ( .A1(n12129), .A2(n12128), .ZN(n14233) );
  NAND2_X1 U12050 ( .A1(n14807), .A2(n9945), .ZN(n14434) );
  INV_X1 U12051 ( .A(n14432), .ZN(n10108) );
  NAND2_X1 U12052 ( .A1(n14807), .A2(n10109), .ZN(n14453) );
  OAI21_X1 U12053 ( .B1(n11275), .B2(n11276), .A(n14728), .ZN(n14638) );
  NAND2_X1 U12054 ( .A1(n14807), .A2(n10111), .ZN(n14461) );
  AND2_X1 U12055 ( .A1(n14807), .A2(n14518), .ZN(n14520) );
  NOR2_X1 U12056 ( .A1(n14806), .A2(n14805), .ZN(n14807) );
  OR2_X1 U12057 ( .A1(n14533), .A2(n14527), .ZN(n14806) );
  NAND2_X1 U12058 ( .A1(n10121), .A2(n10120), .ZN(n16083) );
  INV_X1 U12059 ( .A(n14545), .ZN(n10120) );
  NOR2_X1 U12060 ( .A1(n16083), .A2(n16084), .ZN(n16082) );
  NAND2_X1 U12061 ( .A1(n11256), .A2(n11255), .ZN(n10033) );
  INV_X1 U12062 ( .A(n14053), .ZN(n10114) );
  NOR2_X1 U12063 ( .A1(n14876), .A2(n14218), .ZN(n14868) );
  NAND2_X1 U12064 ( .A1(n11244), .A2(n14714), .ZN(n14308) );
  AND2_X1 U12065 ( .A1(n12083), .A2(n12082), .ZN(n14316) );
  NAND2_X1 U12066 ( .A1(n10115), .A2(n10116), .ZN(n14319) );
  NOR2_X1 U12067 ( .A1(n14061), .A2(n10118), .ZN(n14317) );
  NOR2_X1 U12068 ( .A1(n14061), .A2(n14062), .ZN(n14090) );
  AND2_X1 U12069 ( .A1(n12074), .A2(n12073), .ZN(n13981) );
  AOI21_X1 U12070 ( .B1(n10185), .B2(n10183), .A(n9883), .ZN(n10182) );
  NAND2_X1 U12071 ( .A1(n13930), .A2(n11238), .ZN(n10186) );
  NOR2_X1 U12072 ( .A1(n16274), .A2(n10104), .ZN(n16248) );
  NAND2_X1 U12073 ( .A1(n10105), .A2(n13862), .ZN(n10104) );
  INV_X1 U12074 ( .A(n10106), .ZN(n10105) );
  NAND2_X1 U12075 ( .A1(n16195), .A2(n11213), .ZN(n16191) );
  OR2_X1 U12076 ( .A1(n16274), .A2(n16273), .ZN(n16276) );
  INV_X1 U12077 ( .A(n11196), .ZN(n9981) );
  INV_X1 U12078 ( .A(n13569), .ZN(n10178) );
  AND3_X1 U12079 ( .A1(n13042), .A2(n10123), .A3(n10122), .ZN(n13579) );
  INV_X1 U12080 ( .A(n13547), .ZN(n10122) );
  INV_X1 U12081 ( .A(n10552), .ZN(n10031) );
  INV_X1 U12082 ( .A(n10553), .ZN(n10030) );
  OR3_X1 U12083 ( .A1(n13200), .A2(n13199), .A3(n13198), .ZN(n13507) );
  NAND2_X1 U12084 ( .A1(n11190), .A2(n14890), .ZN(n20426) );
  NAND2_X1 U12085 ( .A1(n9846), .A2(n20265), .ZN(n20649) );
  NOR2_X1 U12086 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20273), .ZN(n20346) );
  OR2_X1 U12087 ( .A1(n9846), .A2(n20265), .ZN(n20679) );
  OR2_X1 U12088 ( .A1(n9846), .A2(n11174), .ZN(n20728) );
  INV_X1 U12089 ( .A(n20649), .ZN(n20527) );
  INV_X1 U12090 ( .A(n10448), .ZN(n20323) );
  NAND2_X1 U12091 ( .A1(n16192), .A2(n20270), .ZN(n20338) );
  NAND2_X1 U12092 ( .A1(n16192), .A2(n20271), .ZN(n20340) );
  INV_X1 U12093 ( .A(n15877), .ZN(n16517) );
  OR2_X1 U12094 ( .A1(n12818), .A2(n12824), .ZN(n12931) );
  NAND2_X1 U12095 ( .A1(n12791), .A2(n15360), .ZN(n16294) );
  OR2_X1 U12096 ( .A1(n12779), .A2(n12782), .ZN(n12786) );
  NOR2_X1 U12097 ( .A1(n12786), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12791) );
  INV_X1 U12098 ( .A(n16310), .ZN(n10137) );
  OAI21_X1 U12099 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(n14965) );
  NAND2_X1 U12100 ( .A1(n10138), .A2(n10137), .ZN(n10135) );
  NAND2_X1 U12101 ( .A1(n19117), .A2(n10138), .ZN(n10134) );
  INV_X1 U12102 ( .A(n14982), .ZN(n10136) );
  NAND2_X1 U12103 ( .A1(n14987), .A2(n12794), .ZN(n12737) );
  NOR3_X1 U12104 ( .A1(n12751), .A2(n10247), .A3(n12740), .ZN(n12744) );
  AND2_X1 U12105 ( .A1(n15037), .A2(n15038), .ZN(n15040) );
  OR2_X1 U12106 ( .A1(n12749), .A2(n12748), .ZN(n12751) );
  NOR2_X1 U12107 ( .A1(n11315), .A2(n15588), .ZN(n11318) );
  NAND2_X1 U12108 ( .A1(n12710), .A2(n11998), .ZN(n12794) );
  NOR3_X2 U12109 ( .A1(n12667), .A2(n10248), .A3(n12647), .ZN(n12714) );
  NAND2_X1 U12110 ( .A1(n10249), .A2(n12709), .ZN(n10248) );
  INV_X1 U12111 ( .A(n10250), .ZN(n10249) );
  NOR3_X1 U12112 ( .A1(n12667), .A2(n12647), .A3(n10250), .ZN(n12710) );
  NOR2_X1 U12113 ( .A1(n11303), .A2(n13659), .ZN(n11305) );
  NAND2_X1 U12114 ( .A1(n10244), .A2(n12001), .ZN(n12661) );
  OR2_X1 U12115 ( .A1(n12918), .A2(n11611), .ZN(n16521) );
  AND2_X1 U12116 ( .A1(n13562), .A2(n13561), .ZN(n13588) );
  INV_X1 U12117 ( .A(n11978), .ZN(n14286) );
  CLKBUF_X2 U12118 ( .A(n11670), .Z(n14285) );
  NAND2_X1 U12119 ( .A1(n15428), .A2(n9864), .ZN(n11983) );
  AND2_X1 U12120 ( .A1(n15267), .A2(n15305), .ZN(n10202) );
  INV_X1 U12121 ( .A(n15337), .ZN(n10203) );
  NAND2_X1 U12122 ( .A1(n15428), .A2(n9933), .ZN(n14942) );
  NAND2_X1 U12123 ( .A1(n15428), .A2(n15427), .ZN(n14939) );
  AND2_X1 U12124 ( .A1(n14999), .A2(n9950), .ZN(n14973) );
  INV_X1 U12125 ( .A(n14971), .ZN(n10238) );
  NAND2_X1 U12126 ( .A1(n14999), .A2(n9860), .ZN(n15449) );
  AND2_X1 U12127 ( .A1(n15170), .A2(n15195), .ZN(n15171) );
  XNOR2_X1 U12128 ( .A(n15170), .B(n15195), .ZN(n15374) );
  OR2_X1 U12129 ( .A1(n13924), .A2(n9911), .ZN(n15387) );
  AND2_X1 U12130 ( .A1(n13899), .A2(n13898), .ZN(n13925) );
  NAND2_X1 U12131 ( .A1(n11769), .A2(n11768), .ZN(n13959) );
  AND2_X1 U12132 ( .A1(n13399), .A2(n13398), .ZN(n13400) );
  NAND2_X1 U12133 ( .A1(n11450), .A2(n19198), .ZN(n13790) );
  NAND2_X1 U12134 ( .A1(n11435), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19239) );
  INV_X1 U12135 ( .A(n12999), .ZN(n13789) );
  XNOR2_X1 U12136 ( .A(n11289), .B(n11288), .ZN(n14378) );
  NAND2_X1 U12137 ( .A1(n11286), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11291) );
  AND2_X1 U12138 ( .A1(n11300), .A2(n10139), .ZN(n11296) );
  AND2_X1 U12139 ( .A1(n9859), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10139) );
  NAND2_X1 U12140 ( .A1(n11300), .A2(n9859), .ZN(n11297) );
  NOR2_X1 U12141 ( .A1(n11299), .A2(n15538), .ZN(n11300) );
  INV_X1 U12142 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19017) );
  NOR2_X1 U12143 ( .A1(n11301), .A2(n19017), .ZN(n11320) );
  INV_X1 U12144 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15588) );
  NOR2_X1 U12145 ( .A1(n11313), .A2(n16359), .ZN(n11316) );
  AND2_X1 U12146 ( .A1(n11311), .A2(n10130), .ZN(n11314) );
  AND2_X1 U12147 ( .A1(n9858), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10130) );
  NAND2_X1 U12148 ( .A1(n11314), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U12149 ( .A1(n11311), .A2(n9858), .ZN(n11312) );
  NOR2_X1 U12150 ( .A1(n11308), .A2(n15610), .ZN(n11311) );
  NAND2_X1 U12151 ( .A1(n11311), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11310) );
  INV_X1 U12152 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15610) );
  AND2_X1 U12153 ( .A1(n9915), .A2(n13552), .ZN(n10224) );
  NAND2_X1 U12154 ( .A1(n10145), .A2(n10146), .ZN(n11308) );
  AND2_X1 U12155 ( .A1(n9853), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10145) );
  AND2_X1 U12156 ( .A1(n10146), .A2(n9853), .ZN(n11309) );
  NAND2_X1 U12157 ( .A1(n10146), .A2(n10147), .ZN(n11306) );
  AND2_X1 U12158 ( .A1(n13426), .A2(n13427), .ZN(n13467) );
  NOR2_X1 U12159 ( .A1(n11304), .A2(n19127), .ZN(n11307) );
  AND2_X1 U12160 ( .A1(n11526), .A2(n11525), .ZN(n13403) );
  NOR2_X1 U12161 ( .A1(n13402), .A2(n13403), .ZN(n13426) );
  NAND2_X1 U12162 ( .A1(n12666), .A2(n16479), .ZN(n10278) );
  NOR2_X1 U12163 ( .A1(n10279), .A2(n10277), .ZN(n10276) );
  INV_X1 U12164 ( .A(n12522), .ZN(n12525) );
  NAND2_X1 U12165 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U12166 ( .A1(n12532), .A2(n12531), .ZN(n12538) );
  NOR2_X1 U12168 ( .A1(n15615), .A2(n12967), .ZN(n10272) );
  OR2_X1 U12169 ( .A1(n14944), .A2(n14364), .ZN(n12806) );
  XNOR2_X1 U12170 ( .A(n12801), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15491) );
  AND2_X1 U12171 ( .A1(n14969), .A2(n14257), .ZN(n15352) );
  OR3_X1 U12172 ( .A1(n14964), .A2(n14364), .A3(n14262), .ZN(n15490) );
  AND2_X1 U12173 ( .A1(n14998), .A2(n10221), .ZN(n14969) );
  AND2_X1 U12174 ( .A1(n9941), .A2(n10222), .ZN(n10221) );
  INV_X1 U12175 ( .A(n14968), .ZN(n10222) );
  NAND2_X1 U12176 ( .A1(n14998), .A2(n9941), .ZN(n15379) );
  NAND2_X1 U12177 ( .A1(n14999), .A2(n10239), .ZN(n15447) );
  NAND2_X1 U12178 ( .A1(n14998), .A2(n14984), .ZN(n15377) );
  INV_X1 U12179 ( .A(n10283), .ZN(n10282) );
  OAI21_X1 U12180 ( .B1(n12778), .B2(n10284), .A(n12777), .ZN(n10283) );
  AND2_X1 U12181 ( .A1(n14999), .A2(n15000), .ZN(n15001) );
  NAND2_X1 U12182 ( .A1(n13944), .A2(n9946), .ZN(n15012) );
  INV_X1 U12183 ( .A(n15015), .ZN(n10226) );
  NAND2_X1 U12184 ( .A1(n13944), .A2(n10227), .ZN(n15014) );
  OR2_X1 U12185 ( .A1(n12767), .A2(n15718), .ZN(n15548) );
  OAI21_X1 U12186 ( .B1(n15767), .B2(n10020), .A(n10018), .ZN(n15546) );
  INV_X1 U12187 ( .A(n10021), .ZN(n10020) );
  AOI21_X1 U12188 ( .B1(n10021), .B2(n15527), .A(n10019), .ZN(n10018) );
  INV_X1 U12189 ( .A(n15528), .ZN(n10019) );
  NAND2_X1 U12190 ( .A1(n15037), .A2(n10230), .ZN(n15024) );
  CLKBUF_X1 U12191 ( .A(n15553), .Z(n15554) );
  NAND2_X1 U12192 ( .A1(n13944), .A2(n13943), .ZN(n14020) );
  NAND2_X1 U12193 ( .A1(n10017), .A2(n10021), .ZN(n15571) );
  NAND2_X1 U12194 ( .A1(n15767), .A2(n10023), .ZN(n10017) );
  NOR2_X1 U12195 ( .A1(n13876), .A2(n13875), .ZN(n13944) );
  AND2_X1 U12196 ( .A1(n13726), .A2(n13727), .ZN(n13742) );
  NAND2_X1 U12197 ( .A1(n13742), .A2(n13741), .ZN(n13876) );
  OAI21_X1 U12198 ( .B1(n15778), .B2(n15525), .A(n15780), .ZN(n15767) );
  AOI21_X1 U12199 ( .B1(n19062), .B2(n16471), .A(n9954), .ZN(n9965) );
  NAND2_X1 U12200 ( .A1(n16377), .A2(n15803), .ZN(n9967) );
  INV_X1 U12201 ( .A(n16360), .ZN(n9968) );
  AND2_X1 U12202 ( .A1(n13617), .A2(n10241), .ZN(n13646) );
  NAND2_X1 U12203 ( .A1(n9849), .A2(n10292), .ZN(n15812) );
  AND2_X1 U12204 ( .A1(n10234), .A2(n15852), .ZN(n10233) );
  NAND2_X1 U12205 ( .A1(n14039), .A2(n14038), .ZN(n13828) );
  INV_X1 U12206 ( .A(n14002), .ZN(n9973) );
  OAI21_X1 U12207 ( .B1(n12523), .B2(n10216), .A(n10215), .ZN(n13411) );
  NAND2_X1 U12208 ( .A1(n10007), .A2(n9919), .ZN(n10215) );
  AND2_X1 U12209 ( .A1(n11612), .A2(n11613), .ZN(n16519) );
  OAI211_X1 U12210 ( .C1(n11978), .C2(n19007), .A(n11669), .B(n11668), .ZN(
        n13297) );
  XNOR2_X1 U12211 ( .A(n13271), .B(n13272), .ZN(n13269) );
  OR2_X1 U12212 ( .A1(n11712), .A2(n11710), .ZN(n13251) );
  CLKBUF_X1 U12213 ( .A(n11619), .Z(n11620) );
  AND2_X1 U12214 ( .A1(n10198), .A2(n13399), .ZN(n13386) );
  OR2_X1 U12215 ( .A1(n13381), .A2(n13380), .ZN(n10198) );
  NAND2_X1 U12216 ( .A1(n13385), .A2(n13386), .ZN(n13401) );
  NAND3_X1 U12217 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12815) );
  AND2_X1 U12218 ( .A1(n19981), .A2(n19990), .ZN(n19635) );
  AND2_X1 U12219 ( .A1(n19981), .A2(n15906), .ZN(n19968) );
  AND2_X1 U12220 ( .A1(n13372), .A2(n19971), .ZN(n19722) );
  INV_X1 U12221 ( .A(n19697), .ZN(n19759) );
  NAND2_X1 U12222 ( .A1(n11403), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11411) );
  AND2_X1 U12223 ( .A1(n11359), .A2(n11358), .ZN(n11362) );
  OR2_X1 U12224 ( .A1(n19972), .A2(n20002), .ZN(n19697) );
  INV_X1 U12225 ( .A(n19352), .ZN(n19358) );
  INV_X1 U12226 ( .A(n19353), .ZN(n19359) );
  INV_X1 U12227 ( .A(n19342), .ZN(n19354) );
  INV_X1 U12228 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20017) );
  NOR2_X1 U12229 ( .A1(n16747), .A2(n16746), .ZN(n16745) );
  NOR2_X1 U12230 ( .A1(n16779), .A2(n16778), .ZN(n16777) );
  AND2_X1 U12231 ( .A1(n10081), .A2(n9928), .ZN(n16789) );
  NAND2_X1 U12232 ( .A1(n16974), .A2(n10085), .ZN(n10082) );
  OR2_X1 U12233 ( .A1(n16809), .A2(n10083), .ZN(n10081) );
  NAND2_X1 U12234 ( .A1(n10085), .A2(n10084), .ZN(n10083) );
  INV_X1 U12235 ( .A(n17701), .ZN(n10084) );
  NOR2_X1 U12236 ( .A1(n17749), .A2(n16719), .ZN(n16847) );
  NOR2_X1 U12237 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16850), .ZN(n16840) );
  AND3_X1 U12238 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16730), .A3(n17087), 
        .ZN(n16902) );
  NOR2_X1 U12239 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17014), .ZN(n17001) );
  AOI21_X1 U12240 ( .B1(n18761), .B2(n18760), .A(n16710), .ZN(n17021) );
  NOR2_X1 U12241 ( .A1(n16812), .A2(n10188), .ZN(n10187) );
  NOR2_X1 U12242 ( .A1(n12210), .A2(n9982), .ZN(n12214) );
  NAND2_X1 U12243 ( .A1(n12209), .A2(n9888), .ZN(n9982) );
  OAI21_X1 U12244 ( .B1(n15940), .B2(n18958), .A(n14104), .ZN(n16021) );
  AOI21_X1 U12245 ( .B1(n15930), .B2(n18811), .A(n18970), .ZN(n17526) );
  NOR2_X1 U12246 ( .A1(n18817), .A2(n18763), .ZN(n17580) );
  NOR2_X1 U12247 ( .A1(n12476), .A2(n17989), .ZN(n16575) );
  NOR2_X1 U12248 ( .A1(n10094), .A2(n10095), .ZN(n10093) );
  INV_X1 U12249 ( .A(n17749), .ZN(n12473) );
  NAND2_X1 U12250 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17749) );
  AND2_X1 U12251 ( .A1(n10097), .A2(n10103), .ZN(n17783) );
  NOR2_X1 U12252 ( .A1(n17894), .A2(n10101), .ZN(n10097) );
  AND2_X1 U12253 ( .A1(n17891), .A2(n10103), .ZN(n17844) );
  AND2_X1 U12254 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17030) );
  AND2_X1 U12255 ( .A1(n16571), .A2(n12295), .ZN(n16004) );
  NOR2_X1 U12256 ( .A1(n17648), .A2(n17780), .ZN(n16599) );
  NAND2_X1 U12257 ( .A1(n12283), .A2(n12282), .ZN(n12287) );
  NOR2_X1 U12258 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17725), .ZN(
        n17712) );
  INV_X1 U12259 ( .A(n9994), .ZN(n17724) );
  OAI211_X1 U12260 ( .C1(n18125), .C2(n10076), .A(n10074), .B(n9914), .ZN(
        n12284) );
  NAND2_X1 U12261 ( .A1(n17854), .A2(n9998), .ZN(n17801) );
  AND2_X1 U12262 ( .A1(n21056), .A2(n18150), .ZN(n9998) );
  NAND2_X1 U12263 ( .A1(n17493), .A2(n18808), .ZN(n18167) );
  NOR2_X1 U12264 ( .A1(n18346), .A2(n18342), .ZN(n18773) );
  OAI21_X1 U12265 ( .B1(n12412), .B2(n12411), .A(n12410), .ZN(n18772) );
  NOR2_X1 U12266 ( .A1(n12468), .A2(n17899), .ZN(n18191) );
  INV_X1 U12267 ( .A(n18241), .ZN(n17902) );
  INV_X1 U12268 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18228) );
  INV_X1 U12269 ( .A(n18361), .ZN(n17377) );
  AOI21_X1 U12270 ( .B1(n12435), .B2(n12428), .A(n15928), .ZN(n15950) );
  AND2_X1 U12271 ( .A1(n15928), .A2(n15927), .ZN(n18763) );
  INV_X1 U12272 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18793) );
  NOR2_X1 U12273 ( .A1(n18969), .A2(n15940), .ZN(n18784) );
  NOR2_X2 U12274 ( .A1(n12324), .A2(n12323), .ZN(n18335) );
  INV_X1 U12275 ( .A(n18972), .ZN(n18338) );
  INV_X1 U12276 ( .A(n12390), .ZN(n18357) );
  NAND2_X1 U12277 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20972) );
  NOR2_X2 U12278 ( .A1(n12146), .A2(n12139), .ZN(n20127) );
  INV_X1 U12279 ( .A(n12144), .ZN(n12139) );
  INV_X1 U12280 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21212) );
  INV_X1 U12281 ( .A(n20098), .ZN(n20110) );
  INV_X1 U12282 ( .A(n20126), .ZN(n20100) );
  INV_X1 U12283 ( .A(n20127), .ZN(n20107) );
  AND2_X1 U12284 ( .A1(n13666), .A2(n13665), .ZN(n20136) );
  AND2_X1 U12285 ( .A1(n20123), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20126) );
  NAND2_X1 U12286 ( .A1(n13042), .A2(n12039), .ZN(n13419) );
  AND2_X1 U12287 ( .A1(n20157), .A2(n20342), .ZN(n20152) );
  NAND2_X2 U12288 ( .A1(n13352), .A2(n13351), .ZN(n20157) );
  OR2_X1 U12289 ( .A1(n13348), .A2(n20042), .ZN(n13352) );
  INV_X1 U12290 ( .A(n20152), .ZN(n20146) );
  INV_X1 U12291 ( .A(n14602), .ZN(n14610) );
  INV_X1 U12292 ( .A(n14082), .ZN(n14314) );
  NAND2_X1 U12293 ( .A1(n12498), .A2(n12497), .ZN(n14600) );
  NAND2_X1 U12294 ( .A1(n13200), .A2(n13201), .ZN(n12498) );
  OR2_X1 U12295 ( .A1(n14609), .A2(n13365), .ZN(n14082) );
  INV_X1 U12296 ( .A(n20172), .ZN(n20973) );
  NOR2_X1 U12297 ( .A1(n13279), .A2(n16016), .ZN(n20170) );
  NOR2_X1 U12298 ( .A1(n20195), .A2(n13309), .ZN(n20192) );
  INV_X1 U12299 ( .A(n13520), .ZN(n20218) );
  INV_X1 U12300 ( .A(n20192), .ZN(n13520) );
  AND2_X1 U12301 ( .A1(n13306), .A2(n16015), .ZN(n13307) );
  INV_X1 U12302 ( .A(n12483), .ZN(n12484) );
  OR2_X1 U12303 ( .A1(n11272), .A2(n11273), .ZN(n11274) );
  INV_X1 U12304 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14656) );
  NAND2_X1 U12305 ( .A1(n20048), .A2(n11163), .ZN(n14693) );
  XNOR2_X1 U12306 ( .A(n9980), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14744) );
  NAND2_X1 U12307 ( .A1(n10170), .A2(n10171), .ZN(n9980) );
  INV_X1 U12308 ( .A(n13601), .ZN(n20236) );
  INV_X1 U12309 ( .A(n20250), .ZN(n20237) );
  NOR2_X1 U12310 ( .A1(n16236), .A2(n13600), .ZN(n20243) );
  OR2_X1 U12311 ( .A1(n13332), .A2(n13038), .ZN(n20248) );
  NOR2_X1 U12312 ( .A1(n13041), .A2(n15965), .ZN(n13332) );
  INV_X1 U12313 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20945) );
  NOR2_X1 U12314 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13205) );
  OR2_X1 U12315 ( .A1(n13276), .A2(n20694), .ZN(n14906) );
  INV_X1 U12316 ( .A(n20425), .ZN(n20443) );
  OAI21_X1 U12317 ( .B1(n20471), .B2(n20455), .A(n20765), .ZN(n20473) );
  OAI211_X1 U12318 ( .C1(n20583), .C2(n20694), .A(n20624), .B(n20568), .ZN(
        n20586) );
  INV_X1 U12319 ( .A(n20628), .ZN(n20645) );
  OAI21_X1 U12320 ( .B1(n20658), .B2(n20657), .A(n20801), .ZN(n20676) );
  OAI211_X1 U12321 ( .C1(n20785), .C2(n20766), .A(n20765), .B(n20764), .ZN(
        n20789) );
  INV_X1 U12322 ( .A(n20702), .ZN(n20808) );
  NAND2_X1 U12323 ( .A1(n20757), .A2(n20527), .ZN(n20838) );
  INV_X1 U12324 ( .A(n20838), .ZN(n20851) );
  NAND2_X1 U12325 ( .A1(n20757), .A2(n20756), .ZN(n20855) );
  AND3_X1 U12326 ( .A1(n15989), .A2(n15988), .A3(n15987), .ZN(n16003) );
  INV_X1 U12327 ( .A(n14906), .ZN(n15999) );
  INV_X1 U12328 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20857) );
  INV_X2 U12329 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20964) );
  NAND2_X1 U12330 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16289) );
  INV_X1 U12331 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20694) );
  INV_X1 U12332 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20968) );
  NOR2_X1 U12334 ( .A1(n16309), .A2(n16310), .ZN(n16308) );
  NOR2_X1 U12335 ( .A1(n14982), .A2(n19117), .ZN(n16309) );
  INV_X1 U12336 ( .A(n12553), .ZN(n12554) );
  INV_X1 U12337 ( .A(n19149), .ZN(n19135) );
  AND2_X1 U12338 ( .A1(n11952), .A2(n11951), .ZN(n13731) );
  INV_X1 U12339 ( .A(n13726), .ZN(n13635) );
  CLKBUF_X1 U12340 ( .A(n15368), .Z(n15370) );
  NAND2_X1 U12341 ( .A1(n15395), .A2(n19355), .ZN(n15397) );
  AND2_X2 U12342 ( .A1(n13077), .A2(n13295), .ZN(n15395) );
  NAND2_X1 U12343 ( .A1(n19198), .A2(n9999), .ZN(n16319) );
  NOR2_X1 U12344 ( .A1(n13790), .A2(n15399), .ZN(n19169) );
  NOR2_X1 U12345 ( .A1(n19210), .A2(n19223), .ZN(n19207) );
  NAND2_X1 U12346 ( .A1(n16319), .A2(n13790), .ZN(n19200) );
  INV_X1 U12347 ( .A(n19198), .ZN(n19222) );
  INV_X1 U12348 ( .A(n19227), .ZN(n19210) );
  NOR2_X1 U12349 ( .A1(n13271), .A2(n13076), .ZN(n19158) );
  OAI21_X1 U12350 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(n19236) );
  OR2_X1 U12351 ( .A1(n19305), .A2(n13080), .ZN(n13101) );
  INV_X1 U12352 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U12353 ( .A1(n14025), .A2(n10269), .ZN(n10263) );
  INV_X1 U12354 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19127) );
  INV_X1 U12355 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13659) );
  AND2_X1 U12356 ( .A1(n16429), .A2(n12870), .ZN(n16426) );
  NAND2_X1 U12357 ( .A1(n12828), .A2(n15910), .ZN(n16421) );
  NAND2_X1 U12358 ( .A1(n13052), .A2(n12866), .ZN(n16429) );
  INV_X1 U12359 ( .A(n16420), .ZN(n16419) );
  INV_X1 U12360 ( .A(n16426), .ZN(n16393) );
  INV_X1 U12361 ( .A(n16415), .ZN(n16424) );
  INV_X1 U12362 ( .A(n16429), .ZN(n16411) );
  INV_X1 U12363 ( .A(n16421), .ZN(n16414) );
  OR2_X1 U12364 ( .A1(n14371), .A2(n14380), .ZN(n14372) );
  OR2_X1 U12365 ( .A1(n15475), .A2(n10270), .ZN(n14369) );
  NAND2_X1 U12366 ( .A1(n10272), .A2(n10271), .ZN(n10270) );
  NOR2_X1 U12367 ( .A1(n15481), .A2(n14355), .ZN(n10271) );
  NAND2_X1 U12368 ( .A1(n10048), .A2(n10304), .ZN(n14368) );
  NOR2_X1 U12369 ( .A1(n14365), .A2(n14364), .ZN(n14366) );
  NAND2_X1 U12370 ( .A1(n15540), .A2(n15689), .ZN(n10006) );
  AND2_X1 U12371 ( .A1(n15756), .A2(n15755), .ZN(n15775) );
  NAND2_X1 U12372 ( .A1(n9966), .A2(n9963), .ZN(n15805) );
  INV_X1 U12373 ( .A(n9964), .ZN(n9963) );
  NAND2_X1 U12374 ( .A1(n15802), .A2(n15847), .ZN(n9966) );
  OAI21_X1 U12375 ( .B1(n19182), .B2(n16469), .A(n9965), .ZN(n9964) );
  NAND2_X1 U12376 ( .A1(n10052), .A2(n10028), .ZN(n10024) );
  INV_X1 U12377 ( .A(n15834), .ZN(n15848) );
  NOR2_X1 U12378 ( .A1(n13966), .A2(n13957), .ZN(n16462) );
  INV_X1 U12379 ( .A(n19310), .ZN(n16469) );
  AOI211_X1 U12380 ( .C1(n15750), .C2(n13238), .A(n13241), .B(n15864), .ZN(
        n16467) );
  NAND2_X1 U12381 ( .A1(n10280), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13654) );
  OR2_X1 U12382 ( .A1(n10280), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13655) );
  INV_X1 U12383 ( .A(n19316), .ZN(n16475) );
  INV_X1 U12384 ( .A(n19158), .ZN(n20002) );
  XNOR2_X1 U12385 ( .A(n13120), .B(n13270), .ZN(n19990) );
  INV_X1 U12386 ( .A(n13269), .ZN(n13120) );
  INV_X1 U12387 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16512) );
  INV_X1 U12388 ( .A(n19990), .ZN(n15906) );
  XNOR2_X1 U12389 ( .A(n13382), .B(n13383), .ZN(n19981) );
  AND2_X1 U12390 ( .A1(n13097), .A2(n13096), .ZN(n19966) );
  INV_X1 U12391 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15903) );
  INV_X1 U12392 ( .A(n19461), .ZN(n19463) );
  INV_X1 U12393 ( .A(n19534), .ZN(n19539) );
  OAI21_X1 U12394 ( .B1(n13628), .B2(n19471), .A(n13627), .ZN(n19540) );
  INV_X1 U12395 ( .A(n19550), .ZN(n19570) );
  NOR2_X1 U12396 ( .A1(n19973), .A2(n19546), .ZN(n19594) );
  NOR2_X2 U12397 ( .A1(n19780), .A2(n19602), .ZN(n19658) );
  NOR2_X2 U12398 ( .A1(n19697), .A2(n19602), .ZN(n19682) );
  INV_X1 U12399 ( .A(n19840), .ZN(n19703) );
  NAND2_X1 U12400 ( .A1(n19759), .A2(n19758), .ZN(n19811) );
  NOR2_X1 U12401 ( .A1(n19780), .A2(n19973), .ZN(n19808) );
  OAI21_X1 U12402 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(n19819) );
  INV_X1 U12403 ( .A(n19811), .ZN(n19817) );
  INV_X1 U12404 ( .A(n19327), .ZN(n19835) );
  AND2_X1 U12405 ( .A1(n11432), .A2(n19354), .ZN(n19827) );
  OAI22_X1 U12406 ( .A1(n13792), .A2(n19359), .B1(n13791), .B2(n19358), .ZN(
        n19840) );
  INV_X1 U12407 ( .A(n19484), .ZN(n19839) );
  AND2_X1 U12408 ( .A1(n13630), .A2(n19354), .ZN(n19850) );
  NOR2_X2 U12409 ( .A1(n19697), .A2(n19973), .ZN(n19879) );
  OAI22_X1 U12410 ( .A1(n20336), .A2(n19359), .B1(n15450), .B2(n19358), .ZN(
        n19878) );
  INV_X1 U12411 ( .A(n19808), .ZN(n19883) );
  INV_X1 U12412 ( .A(n20012), .ZN(n16539) );
  AND2_X1 U12413 ( .A1(n16547), .A2(n16546), .ZN(n16550) );
  OAI21_X1 U12414 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n19237), .ZN(n20024) );
  INV_X1 U12415 ( .A(n16550), .ZN(n19885) );
  INV_X1 U12416 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19897) );
  INV_X2 U12417 ( .A(n20036), .ZN(n20039) );
  NAND2_X1 U12418 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19897), .ZN(n20036) );
  INV_X1 U12419 ( .A(n18057), .ZN(n18959) );
  OR2_X1 U12420 ( .A1(n16754), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12421 ( .A1(n16751), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n10088) );
  XNOR2_X1 U12422 ( .A(n16738), .B(n10091), .ZN(n10090) );
  INV_X1 U12423 ( .A(n16739), .ZN(n10091) );
  NOR2_X1 U12424 ( .A1(n18898), .A2(n16785), .ZN(n16756) );
  NOR2_X1 U12425 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16810), .ZN(n16800) );
  NOR2_X1 U12426 ( .A1(n16809), .A2(n17701), .ZN(n16808) );
  NOR2_X1 U12427 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16831), .ZN(n16818) );
  NOR2_X1 U12428 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16874), .ZN(n16859) );
  CLKBUF_X1 U12429 ( .A(n16729), .Z(n16974) );
  NOR2_X1 U12430 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16947), .ZN(n16946) );
  INV_X1 U12431 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17050) );
  NAND2_X1 U12432 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17087), .ZN(n17059) );
  INV_X1 U12433 ( .A(n18825), .ZN(n17066) );
  INV_X1 U12434 ( .A(n17059), .ZN(n17071) );
  INV_X1 U12435 ( .A(n17028), .ZN(n17084) );
  INV_X1 U12436 ( .A(n17047), .ZN(n17083) );
  NAND4_X1 U12437 ( .A1(n18317), .A2(n18985), .A3(n18825), .A4(n18815), .ZN(
        n17087) );
  AND2_X1 U12438 ( .A1(n10190), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U12439 ( .A1(n14108), .A2(n10191), .ZN(n17185) );
  AND2_X1 U12440 ( .A1(n14108), .A2(n9959), .ZN(n17197) );
  INV_X1 U12441 ( .A(n17211), .ZN(n14108) );
  NAND2_X1 U12442 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17225), .ZN(n17211) );
  NOR3_X1 U12443 ( .A1(n16906), .A2(n17252), .A3(n17228), .ZN(n17225) );
  INV_X1 U12444 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17252) );
  AND2_X1 U12445 ( .A1(n17267), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17280) );
  NOR2_X1 U12446 ( .A1(n17357), .A2(n17360), .ZN(n17353) );
  NAND2_X1 U12447 ( .A1(n17353), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U12448 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12376) );
  NAND2_X1 U12449 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17361), .ZN(n17357) );
  NOR2_X1 U12450 ( .A1(n17370), .A2(n17073), .ZN(n17361) );
  INV_X1 U12451 ( .A(n17370), .ZN(n17367) );
  NAND4_X1 U12452 ( .A1(n18967), .A2(n18338), .A3(n16711), .A4(n16021), .ZN(
        n17370) );
  INV_X1 U12453 ( .A(n17391), .ZN(n17387) );
  INV_X1 U12454 ( .A(n17409), .ZN(n17405) );
  AND2_X1 U12455 ( .A1(n17462), .A2(n17516), .ZN(n17495) );
  NOR2_X1 U12456 ( .A1(n12193), .A2(n12192), .ZN(n17507) );
  NAND2_X1 U12457 ( .A1(n17483), .A2(n16024), .ZN(n17515) );
  NAND2_X1 U12458 ( .A1(n18787), .A2(n17517), .ZN(n17512) );
  INV_X1 U12459 ( .A(n18367), .ZN(n17519) );
  INV_X1 U12460 ( .A(n17515), .ZN(n17522) );
  NOR2_X1 U12461 ( .A1(n17576), .A2(n17568), .ZN(n17561) );
  INV_X1 U12462 ( .A(n17578), .ZN(n17568) );
  BUF_X1 U12463 ( .A(n17561), .Z(n20977) );
  OAI211_X1 U12464 ( .C1(n18972), .C2(n18973), .A(n17581), .B(n17580), .ZN(
        n17619) );
  INV_X1 U12465 ( .A(n17629), .ZN(n17623) );
  INV_X1 U12466 ( .A(n17619), .ZN(n17629) );
  AND2_X1 U12467 ( .A1(n17673), .A2(n9929), .ZN(n16578) );
  INV_X1 U12468 ( .A(n18364), .ZN(n18705) );
  NAND2_X1 U12469 ( .A1(n17673), .A2(n9847), .ZN(n17635) );
  NAND2_X1 U12470 ( .A1(n17673), .A2(n9857), .ZN(n17661) );
  AND2_X1 U12471 ( .A1(n16718), .A2(n9912), .ZN(n17703) );
  NAND2_X1 U12472 ( .A1(n16718), .A2(n12473), .ZN(n17734) );
  INV_X1 U12473 ( .A(n17846), .ZN(n17831) );
  NOR2_X1 U12474 ( .A1(n17894), .A2(n10098), .ZN(n10096) );
  NAND2_X1 U12475 ( .A1(n10099), .A2(n9922), .ZN(n10098) );
  INV_X1 U12476 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17773) );
  NOR2_X1 U12477 ( .A1(n18928), .A2(n17882), .ZN(n17846) );
  NAND2_X1 U12478 ( .A1(n10103), .A2(n10100), .ZN(n17813) );
  NOR2_X1 U12479 ( .A1(n17894), .A2(n9877), .ZN(n10100) );
  NAND2_X1 U12480 ( .A1(n17993), .A2(n17829), .ZN(n17882) );
  NAND2_X1 U12481 ( .A1(n17986), .A2(n15959), .ZN(n17877) );
  INV_X1 U12482 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17912) );
  INV_X1 U12483 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17940) );
  INV_X1 U12484 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17980) );
  INV_X1 U12485 ( .A(n17985), .ZN(n17977) );
  NOR2_X2 U12486 ( .A1(n18057), .A2(n17975), .ZN(n17983) );
  INV_X1 U12487 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18928) );
  INV_X1 U12488 ( .A(n17983), .ZN(n17998) );
  OAI22_X1 U12489 ( .A1(n17649), .A2(n10073), .B1(n17648), .B2(n10071), .ZN(
        n10068) );
  NAND2_X1 U12490 ( .A1(n10062), .A2(n9992), .ZN(n9990) );
  AND2_X1 U12491 ( .A1(n10060), .A2(n9992), .ZN(n9991) );
  NAND2_X1 U12492 ( .A1(n10061), .A2(n12291), .ZN(n17659) );
  NAND2_X1 U12493 ( .A1(n12280), .A2(n18189), .ZN(n18241) );
  INV_X1 U12494 ( .A(n18221), .ZN(n18236) );
  INV_X1 U12495 ( .A(n9986), .ZN(n17953) );
  INV_X1 U12496 ( .A(n12263), .ZN(n10078) );
  INV_X1 U12497 ( .A(n18963), .ZN(n18808) );
  AND2_X1 U12498 ( .A1(n10067), .A2(n9850), .ZN(n17970) );
  INV_X1 U12499 ( .A(n18788), .ZN(n18768) );
  INV_X1 U12500 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18802) );
  AOI211_X1 U12501 ( .C1(n18967), .C2(n18785), .A(n18334), .B(n15941), .ZN(
        n18947) );
  INV_X1 U12502 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18767) );
  INV_X1 U12503 ( .A(n18947), .ZN(n18945) );
  OAI21_X1 U12505 ( .B1(n14508), .B2(n20140), .A(n12152), .ZN(n12153) );
  OAI21_X1 U12506 ( .B1(n14203), .B2(n20048), .A(n9893), .ZN(P1_U2968) );
  NOR4_X1 U12507 ( .A1(n14229), .A2(n14228), .A3(n14227), .A4(n14226), .ZN(
        n14230) );
  AOI211_X1 U12508 ( .C1(n19163), .C2(n16306), .A(n14295), .B(n10213), .ZN(
        n14296) );
  NAND2_X1 U12509 ( .A1(n14291), .A2(n10214), .ZN(n10213) );
  AOI21_X1 U12510 ( .B1(n11325), .B2(n14357), .A(n19888), .ZN(n11326) );
  INV_X1 U12511 ( .A(n10125), .ZN(n14922) );
  OAI21_X1 U12512 ( .B1(n14920), .B2(n10127), .A(n10126), .ZN(n10125) );
  NAND2_X1 U12513 ( .A1(n10128), .A2(n19136), .ZN(n10127) );
  AOI211_X1 U12514 ( .C1(n9962), .C2(P2_REIP_REG_18__SCAN_IN), .A(n15030), .B(
        n15029), .ZN(n15031) );
  AOI21_X1 U12515 ( .B1(n14399), .B2(n15847), .A(n14398), .ZN(n14400) );
  INV_X1 U12516 ( .A(n10179), .ZN(P3_U2675) );
  AOI21_X1 U12517 ( .B1(n15921), .B2(P3_EBX_REG_28__SCAN_IN), .A(n10180), .ZN(
        n10179) );
  OAI21_X1 U12518 ( .B1(n17121), .B2(n15922), .A(n10181), .ZN(n10180) );
  INV_X1 U12519 ( .A(n17267), .ZN(n17293) );
  INV_X1 U12520 ( .A(n17294), .ZN(n17315) );
  AND2_X1 U12521 ( .A1(n9848), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9847) );
  BUF_X1 U12522 ( .A(n11439), .Z(n19347) );
  INV_X1 U12523 ( .A(n12242), .ZN(n12348) );
  NOR2_X2 U12524 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15942), .ZN(
        n12242) );
  AND2_X1 U12525 ( .A1(n9857), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9848) );
  INV_X1 U12526 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17347) );
  AND2_X1 U12527 ( .A1(n10059), .A2(n10058), .ZN(n9849) );
  INV_X1 U12528 ( .A(n12211), .ZN(n17322) );
  NOR2_X2 U12529 ( .A1(n17074), .A2(n12158), .ZN(n12211) );
  INV_X1 U12530 ( .A(n11617), .ZN(n11988) );
  INV_X1 U12531 ( .A(n12729), .ZN(n10056) );
  NAND2_X1 U12532 ( .A1(n10151), .A2(n10152), .ZN(n14471) );
  NOR2_X1 U12533 ( .A1(n15539), .A2(n10261), .ZN(n15511) );
  NAND2_X1 U12534 ( .A1(n11453), .A2(n11446), .ZN(n11615) );
  OR2_X1 U12535 ( .A1(n17520), .A2(n18927), .ZN(n9850) );
  NAND2_X1 U12536 ( .A1(n10204), .A2(n9943), .ZN(n9851) );
  AND2_X1 U12537 ( .A1(n12704), .A2(n9947), .ZN(n9852) );
  NAND2_X1 U12538 ( .A1(n12566), .A2(n19150), .ZN(n12572) );
  INV_X1 U12539 ( .A(n10068), .ZN(n15960) );
  AND2_X1 U12540 ( .A1(n10147), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9853) );
  INV_X1 U12541 ( .A(n13119), .ZN(n13228) );
  AND2_X1 U12542 ( .A1(n14695), .A2(n9960), .ZN(n9854) );
  AND2_X1 U12543 ( .A1(n12473), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9855) );
  NAND2_X1 U12544 ( .A1(n13019), .A2(n13309), .ZN(n12041) );
  AND2_X1 U12545 ( .A1(n14039), .A2(n10234), .ZN(n13829) );
  NOR2_X1 U12546 ( .A1(n13924), .A2(n13925), .ZN(n9856) );
  AND2_X1 U12547 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U12548 ( .A1(n13759), .A2(n13760), .ZN(n13783) );
  AND2_X1 U12549 ( .A1(n10131), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9858) );
  AOI21_X1 U12550 ( .B1(n14982), .B2(n10137), .A(n19117), .ZN(n10133) );
  INV_X1 U12551 ( .A(n10153), .ZN(n10152) );
  NAND2_X1 U12552 ( .A1(n14472), .A2(n10154), .ZN(n10153) );
  INV_X2 U12553 ( .A(n15127), .ZN(n11643) );
  AND2_X1 U12554 ( .A1(n10140), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9859) );
  AND2_X1 U12555 ( .A1(n10239), .A2(n11968), .ZN(n9860) );
  AND2_X1 U12556 ( .A1(n9942), .A2(n10237), .ZN(n9861) );
  AND2_X1 U12557 ( .A1(n9933), .A2(n10219), .ZN(n9862) );
  AND2_X1 U12558 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9863) );
  INV_X1 U12559 ( .A(n10212), .ZN(n13637) );
  AND2_X1 U12560 ( .A1(n9862), .A2(n14915), .ZN(n9864) );
  AND2_X1 U12561 ( .A1(n9863), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9865) );
  AND2_X1 U12562 ( .A1(n15715), .A2(n12863), .ZN(n9866) );
  AND2_X1 U12563 ( .A1(n9866), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9867) );
  AND2_X1 U12564 ( .A1(n10187), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n9868) );
  AND2_X1 U12565 ( .A1(n9868), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12566 ( .A1(n13968), .A2(n13969), .ZN(n10016) );
  INV_X2 U12567 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11408) );
  AND4_X1 U12568 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n9870) );
  NAND2_X1 U12569 ( .A1(n13274), .A2(n13273), .ZN(n13383) );
  NAND2_X1 U12570 ( .A1(n15599), .A2(n15715), .ZN(n15572) );
  AND2_X1 U12571 ( .A1(n12696), .A2(n12695), .ZN(n9872) );
  AND4_X1 U12572 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n9873) );
  INV_X1 U12573 ( .A(n11304), .ZN(n10146) );
  OR2_X1 U12574 ( .A1(n12159), .A2(n12156), .ZN(n9874) );
  OR2_X1 U12575 ( .A1(n18292), .A2(n12259), .ZN(n9875) );
  NAND2_X1 U12576 ( .A1(n10288), .A2(n15500), .ZN(n14253) );
  INV_X1 U12577 ( .A(n17300), .ZN(n17272) );
  NAND2_X1 U12578 ( .A1(n10186), .A2(n10185), .ZN(n14724) );
  NAND2_X1 U12579 ( .A1(n14534), .A2(n14536), .ZN(n14524) );
  XOR2_X1 U12580 ( .A(n15467), .B(n15466), .Z(n9876) );
  NAND2_X1 U12581 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9877) );
  NOR2_X1 U12582 ( .A1(n12156), .A2(n17075), .ZN(n12244) );
  AND2_X1 U12583 ( .A1(n14534), .A2(n10155), .ZN(n14515) );
  AND2_X1 U12584 ( .A1(n15428), .A2(n9862), .ZN(n9878) );
  NAND2_X1 U12585 ( .A1(n14629), .A2(n10042), .ZN(n9879) );
  NAND2_X1 U12586 ( .A1(n14534), .A2(n10157), .ZN(n9880) );
  AND2_X1 U12587 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n9881) );
  AND2_X1 U12588 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12589 ( .A1(n10013), .A2(n14029), .ZN(n16402) );
  NAND2_X1 U12590 ( .A1(n10052), .A2(n12729), .ZN(n16372) );
  NAND2_X1 U12591 ( .A1(n10186), .A2(n11239), .ZN(n13986) );
  INV_X1 U12592 ( .A(n11439), .ZN(n11429) );
  NAND2_X1 U12593 ( .A1(n12723), .A2(n10252), .ZN(n12745) );
  NAND2_X1 U12594 ( .A1(n12865), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14354) );
  AND2_X1 U12595 ( .A1(n16173), .A2(n16256), .ZN(n9883) );
  AND2_X1 U12596 ( .A1(n9849), .A2(n15605), .ZN(n9884) );
  XNOR2_X1 U12597 ( .A(n10197), .B(n15243), .ZN(n15348) );
  AND2_X2 U12598 ( .A1(n15874), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11621) );
  AND3_X1 U12599 ( .A1(n15491), .A2(n15500), .A3(n15488), .ZN(n9885) );
  NAND2_X1 U12600 ( .A1(n10263), .A2(n10267), .ZN(n16399) );
  NAND2_X1 U12601 ( .A1(n9990), .A2(n9989), .ZN(n16597) );
  OAI21_X1 U12602 ( .B1(n12848), .B2(n12646), .A(n19128), .ZN(n12670) );
  AND3_X1 U12603 ( .A1(n11361), .A2(n11408), .A3(n11360), .ZN(n9886) );
  OAI21_X1 U12604 ( .B1(n13382), .B2(n13383), .A(n13384), .ZN(n13385) );
  NAND2_X1 U12605 ( .A1(n10204), .A2(n15337), .ZN(n15332) );
  AND2_X1 U12606 ( .A1(n16259), .A2(n16258), .ZN(n9887) );
  NAND2_X1 U12607 ( .A1(n12566), .A2(n12534), .ZN(n12619) );
  OR2_X1 U12608 ( .A1(n9874), .A2(n9983), .ZN(n9888) );
  INV_X1 U12609 ( .A(n10002), .ZN(n12526) );
  NAND2_X1 U12610 ( .A1(n11508), .A2(n11509), .ZN(n10002) );
  AND2_X1 U12611 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n9889) );
  AND2_X1 U12612 ( .A1(n11393), .A2(n11391), .ZN(n9890) );
  AND2_X1 U12613 ( .A1(n11397), .A2(n11394), .ZN(n9891) );
  AND2_X1 U12614 ( .A1(n12723), .A2(n10254), .ZN(n9892) );
  INV_X1 U12615 ( .A(n20028), .ZN(n11435) );
  NAND2_X1 U12616 ( .A1(n15599), .A2(n9866), .ZN(n15563) );
  AND2_X1 U12617 ( .A1(n11271), .A2(n11270), .ZN(n9893) );
  AND2_X1 U12618 ( .A1(n15352), .A2(n15351), .ZN(n14935) );
  NAND2_X1 U12619 ( .A1(n13974), .A2(n14059), .ZN(n14058) );
  XNOR2_X1 U12620 ( .A(n12829), .B(n12830), .ZN(n12843) );
  NAND2_X1 U12621 ( .A1(n11443), .A2(n13303), .ZN(n12942) );
  NAND2_X1 U12622 ( .A1(n10568), .A2(n11170), .ZN(n9894) );
  INV_X1 U12623 ( .A(n12701), .ZN(n10251) );
  OR2_X1 U12624 ( .A1(n12751), .A2(n10245), .ZN(n9895) );
  OR2_X1 U12625 ( .A1(n16173), .A2(n16256), .ZN(n9896) );
  AND2_X1 U12626 ( .A1(n10570), .A2(n20968), .ZN(n9897) );
  AND2_X1 U12627 ( .A1(n14629), .A2(n14754), .ZN(n9898) );
  AND2_X1 U12628 ( .A1(n10007), .A2(n13265), .ZN(n9899) );
  NOR2_X1 U12629 ( .A1(n16742), .A2(n10086), .ZN(n9900) );
  NAND2_X1 U12630 ( .A1(n17901), .A2(n10076), .ZN(n9901) );
  NOR2_X1 U12631 ( .A1(n17780), .A2(n18125), .ZN(n10075) );
  AND2_X2 U12632 ( .A1(n11617), .A2(n19825), .ZN(n11664) );
  INV_X1 U12633 ( .A(n11497), .ZN(n11585) );
  INV_X2 U12634 ( .A(n11585), .ZN(n14276) );
  NOR2_X2 U12635 ( .A1(n15883), .A2(n19237), .ZN(n11497) );
  INV_X1 U12636 ( .A(n12288), .ZN(n17697) );
  AND2_X1 U12637 ( .A1(n17137), .A2(n9868), .ZN(n9902) );
  NAND2_X1 U12638 ( .A1(n11320), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U12639 ( .A1(n15037), .A2(n10232), .ZN(n13786) );
  NOR2_X1 U12640 ( .A1(n15799), .A2(n13853), .ZN(n13852) );
  AND2_X1 U12641 ( .A1(n17137), .A2(n10187), .ZN(n9903) );
  AND2_X1 U12642 ( .A1(n17137), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12643 ( .A1(n17901), .A2(n12280), .ZN(n17800) );
  AND2_X1 U12644 ( .A1(n10072), .A2(n18025), .ZN(n9905) );
  AND2_X1 U12645 ( .A1(n11311), .A2(n10131), .ZN(n9906) );
  NAND2_X1 U12647 ( .A1(n13711), .A2(n13710), .ZN(n13709) );
  AND2_X1 U12648 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n9907) );
  AND2_X1 U12649 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n9908) );
  XNOR2_X1 U12650 ( .A(n12670), .B(n13997), .ZN(n13993) );
  AND2_X1 U12651 ( .A1(n13590), .A2(n13644), .ZN(n9909) );
  OR2_X1 U12652 ( .A1(n10209), .A2(n13925), .ZN(n9910) );
  OR2_X1 U12653 ( .A1(n9910), .A2(n10208), .ZN(n9911) );
  NAND2_X1 U12654 ( .A1(n9979), .A2(n16182), .ZN(n13930) );
  NAND2_X1 U12655 ( .A1(n12857), .A2(n13955), .ZN(n14025) );
  NAND2_X1 U12656 ( .A1(n10016), .A2(n12704), .ZN(n14028) );
  AND2_X1 U12657 ( .A1(n9855), .A2(n10093), .ZN(n9912) );
  OR2_X1 U12658 ( .A1(n9911), .A2(n15382), .ZN(n9913) );
  OR2_X1 U12659 ( .A1(n17780), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9914) );
  AND2_X1 U12660 ( .A1(n13852), .A2(n15784), .ZN(n15037) );
  INV_X1 U12661 ( .A(n15500), .ZN(n10287) );
  AND2_X1 U12662 ( .A1(n10225), .A2(n13433), .ZN(n9915) );
  AND2_X1 U12663 ( .A1(n17854), .A2(n21056), .ZN(n17837) );
  AND2_X1 U12664 ( .A1(n10412), .A2(n10448), .ZN(n11162) );
  NAND2_X1 U12665 ( .A1(n13720), .A2(n12845), .ZN(n14001) );
  AND2_X1 U12666 ( .A1(n10240), .A2(n13636), .ZN(n9916) );
  AND2_X1 U12667 ( .A1(n12286), .A2(n9995), .ZN(n17769) );
  AND2_X1 U12668 ( .A1(n10038), .A2(n10040), .ZN(n9917) );
  INV_X1 U12669 ( .A(n15527), .ZN(n10023) );
  AND2_X1 U12670 ( .A1(n10024), .A2(n16373), .ZN(n9918) );
  AND2_X1 U12671 ( .A1(n11519), .A2(n11509), .ZN(n9919) );
  NAND2_X1 U12672 ( .A1(n12470), .A2(n10072), .ZN(n9920) );
  NAND2_X1 U12673 ( .A1(n12883), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n9921) );
  INV_X1 U12674 ( .A(n10207), .ZN(n15391) );
  OR2_X1 U12675 ( .A1(n13924), .A2(n9910), .ZN(n10207) );
  NAND4_X1 U12676 ( .A1(n9873), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n12612) );
  INV_X1 U12677 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21100) );
  AND2_X1 U12678 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9922) );
  AND2_X1 U12679 ( .A1(n14108), .A2(n10190), .ZN(n9923) );
  NAND2_X1 U12680 ( .A1(n11300), .A2(n10140), .ZN(n10143) );
  NOR2_X1 U12681 ( .A1(n13377), .A2(n13376), .ZN(n9924) );
  AND2_X1 U12682 ( .A1(n15017), .A2(n15016), .ZN(n14999) );
  AND2_X1 U12683 ( .A1(n10155), .A2(n14517), .ZN(n9925) );
  AND2_X1 U12684 ( .A1(n10252), .A2(n9921), .ZN(n9926) );
  AND2_X1 U12685 ( .A1(n10116), .A2(n10114), .ZN(n9927) );
  INV_X1 U12686 ( .A(n14029), .ZN(n10015) );
  AND2_X1 U12687 ( .A1(n10082), .A2(n10080), .ZN(n9928) );
  AND2_X1 U12688 ( .A1(n9847), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9929) );
  AND2_X1 U12689 ( .A1(n10149), .A2(n10702), .ZN(n9930) );
  AND2_X1 U12690 ( .A1(n9912), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9931) );
  INV_X1 U12691 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15598) );
  NAND4_X2 U12692 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n12646) );
  INV_X1 U12693 ( .A(n11628), .ZN(n15127) );
  NAND2_X1 U12694 ( .A1(n11787), .A2(n11786), .ZN(n14039) );
  AND2_X1 U12695 ( .A1(n11286), .A2(n9863), .ZN(n9932) );
  AND2_X1 U12696 ( .A1(n13426), .A2(n9915), .ZN(n13431) );
  AND2_X1 U12697 ( .A1(n13617), .A2(n13616), .ZN(n13583) );
  INV_X1 U12698 ( .A(n16306), .ZN(n19143) );
  AND2_X1 U12699 ( .A1(n19305), .A2(n16542), .ZN(n16306) );
  AND2_X1 U12700 ( .A1(n13426), .A2(n10225), .ZN(n13432) );
  AND2_X1 U12701 ( .A1(n13426), .A2(n10224), .ZN(n13551) );
  NAND2_X1 U12702 ( .A1(n13411), .A2(n13410), .ZN(n13402) );
  NAND2_X1 U12703 ( .A1(n13591), .A2(n9909), .ZN(n13638) );
  INV_X1 U12704 ( .A(n17685), .ZN(n10085) );
  AND2_X1 U12705 ( .A1(n15427), .A2(n10220), .ZN(n9933) );
  AND2_X1 U12706 ( .A1(n13190), .A2(n13280), .ZN(n12020) );
  AND2_X1 U12707 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n9934) );
  AND2_X1 U12708 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n9935) );
  AND2_X1 U12709 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9936) );
  AND2_X1 U12710 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n9937) );
  AND2_X1 U12711 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n9938) );
  AND2_X1 U12712 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9939) );
  AND2_X1 U12713 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n9940) );
  AND2_X1 U12714 ( .A1(n10223), .A2(n14984), .ZN(n9941) );
  AND2_X1 U12715 ( .A1(n14938), .A2(n12869), .ZN(n9942) );
  NOR2_X1 U12716 ( .A1(n15333), .A2(n10203), .ZN(n9943) );
  INV_X1 U12717 ( .A(n16373), .ZN(n10286) );
  INV_X1 U12718 ( .A(n16403), .ZN(n10051) );
  NOR2_X1 U12719 ( .A1(n16808), .A2(n16729), .ZN(n9944) );
  AND2_X1 U12720 ( .A1(n10109), .A2(n10108), .ZN(n9945) );
  AND2_X1 U12721 ( .A1(n15308), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11916) );
  NOR3_X1 U12722 ( .A1(n12751), .A2(n10245), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n10246) );
  INV_X1 U12723 ( .A(n10121), .ZN(n14546) );
  NOR2_X1 U12724 ( .A1(n14556), .A2(n14475), .ZN(n10121) );
  AND2_X1 U12725 ( .A1(n10227), .A2(n10226), .ZN(n9946) );
  NOR2_X1 U12726 ( .A1(n11294), .A2(n15482), .ZN(n11286) );
  INV_X1 U12727 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U12728 ( .A1(n19103), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9947) );
  NAND2_X1 U12729 ( .A1(n13591), .A2(n13590), .ZN(n10212) );
  NOR2_X1 U12730 ( .A1(n16274), .A2(n10106), .ZN(n9948) );
  AND2_X1 U12731 ( .A1(n9861), .A2(n10236), .ZN(n9949) );
  AND2_X1 U12732 ( .A1(n9860), .A2(n10238), .ZN(n9950) );
  BUF_X1 U12733 ( .A(n11629), .Z(n15128) );
  XOR2_X1 U12734 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n12474), .Z(
        n16729) );
  INV_X1 U12735 ( .A(n16974), .ZN(n10080) );
  INV_X1 U12736 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10315) );
  INV_X1 U12737 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10142) );
  OR2_X1 U12738 ( .A1(n17991), .A2(n17981), .ZN(n10067) );
  INV_X1 U12739 ( .A(n13701), .ZN(n10277) );
  INV_X1 U12740 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14323) );
  AND2_X1 U12741 ( .A1(n17673), .A2(n9848), .ZN(n9951) );
  AND2_X1 U12742 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n9952) );
  AND2_X1 U12743 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n9953) );
  AND2_X1 U12744 ( .A1(n16460), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U12745 ( .A1(n11962), .A2(n11961), .ZN(n9955) );
  NOR2_X1 U12746 ( .A1(n17970), .A2(n17969), .ZN(n17968) );
  OR2_X1 U12747 ( .A1(n17373), .A2(n14193), .ZN(n9956) );
  AND2_X1 U12748 ( .A1(n9985), .A2(n9984), .ZN(n17932) );
  AND2_X1 U12749 ( .A1(n10079), .A2(n10078), .ZN(n9957) );
  OR2_X1 U12750 ( .A1(n17962), .A2(n18280), .ZN(n10079) );
  NOR2_X1 U12751 ( .A1(n17962), .A2(n18280), .ZN(n9987) );
  INV_X1 U12752 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17337) );
  INV_X1 U12753 ( .A(n18957), .ZN(n18981) );
  INV_X1 U12754 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10092) );
  INV_X1 U12755 ( .A(n16560), .ZN(n10077) );
  AND2_X1 U12756 ( .A1(n16718), .A2(n9855), .ZN(n9958) );
  INV_X1 U12757 ( .A(n11615), .ZN(n9999) );
  INV_X1 U12758 ( .A(n19136), .ZN(n19888) );
  AND3_X1 U12759 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(P3_EBX_REG_17__SCAN_IN), .ZN(n9959) );
  AND2_X1 U12760 ( .A1(n11257), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9960) );
  NAND2_X1 U12761 ( .A1(n17920), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17894) );
  INV_X1 U12762 ( .A(n10192), .ZN(n10191) );
  NAND2_X1 U12763 ( .A1(n9959), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n10192) );
  INV_X1 U12764 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10044) );
  INV_X1 U12765 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9992) );
  INV_X1 U12766 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10193) );
  INV_X1 U12767 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10060) );
  INV_X1 U12768 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10188) );
  INV_X1 U12769 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10064) );
  INV_X1 U12770 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U12771 ( .A1(n10272), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9961) );
  INV_X1 U12772 ( .A(n19042), .ZN(n19155) );
  NOR3_X2 U12773 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18820), .A3(
        n18554), .ZN(n18526) );
  CLKBUF_X1 U12774 ( .A(n19152), .Z(n9962) );
  NAND2_X1 U12775 ( .A1(n9962), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12776 ( .A1(n9962), .A2(n19825), .ZN(n19042) );
  NOR4_X1 U12777 ( .A1(n16460), .A2(n19136), .A3(n20019), .A4(n16537), .ZN(
        n19152) );
  NOR3_X4 U12778 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18791), .A3(
        n18554), .ZN(n18598) );
  NOR2_X2 U12779 ( .A1(n20343), .A2(n20287), .ZN(n20809) );
  OR3_X1 U12780 ( .A1(n20694), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20273), 
        .ZN(n20343) );
  NAND2_X2 U12781 ( .A1(n16400), .A2(n12862), .ZN(n15599) );
  NAND2_X4 U12782 ( .A1(n10273), .A2(n10007), .ZN(n16502) );
  NOR2_X1 U12783 ( .A1(n16502), .A2(n12559), .ZN(n12546) );
  NAND2_X1 U12784 ( .A1(n10471), .A2(n10465), .ZN(n10472) );
  INV_X1 U12785 ( .A(n10465), .ZN(n9975) );
  XNOR2_X2 U12786 ( .A(n10501), .B(n10500), .ZN(n10573) );
  NAND2_X2 U12787 ( .A1(n13032), .A2(n10165), .ZN(n11188) );
  NAND2_X2 U12788 ( .A1(n13329), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13328) );
  NAND2_X2 U12789 ( .A1(n14630), .A2(n14638), .ZN(n14629) );
  NAND2_X1 U12791 ( .A1(n13597), .A2(n11203), .ZN(n16197) );
  OAI211_X2 U12792 ( .C1(n13570), .C2(n9981), .A(n13598), .B(n10177), .ZN(
        n13597) );
  INV_X2 U12793 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12415) );
  INV_X2 U12794 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12413) );
  NAND2_X1 U12795 ( .A1(n9987), .A2(n9988), .ZN(n9985) );
  AOI21_X1 U12796 ( .B1(n9988), .B2(n12263), .A(n12266), .ZN(n9984) );
  INV_X1 U12797 ( .A(n17954), .ZN(n9988) );
  NAND3_X1 U12798 ( .A1(n12291), .A2(n9991), .A3(n10061), .ZN(n9989) );
  NOR2_X2 U12799 ( .A1(n9993), .A2(n9905), .ZN(n12291) );
  AND2_X2 U12800 ( .A1(n12286), .A2(n9901), .ZN(n17781) );
  XNOR2_X1 U12801 ( .A(n12274), .B(n12273), .ZN(n17915) );
  NAND2_X1 U12802 ( .A1(n17818), .A2(n12278), .ZN(n12279) );
  NOR2_X2 U12803 ( .A1(n12877), .A2(n20028), .ZN(n11986) );
  NAND3_X1 U12804 ( .A1(n9999), .A2(n11429), .A3(n11451), .ZN(n12877) );
  AND3_X2 U12805 ( .A1(n13630), .A2(n11440), .A3(n11458), .ZN(n11451) );
  INV_X1 U12806 ( .A(n12853), .ZN(n12847) );
  NAND2_X1 U12807 ( .A1(n12528), .A2(n11495), .ZN(n12527) );
  AOI22_X2 U12808 ( .A1(n12528), .A2(n10001), .B1(n11509), .B2(n10000), .ZN(
        n12522) );
  AND2_X1 U12809 ( .A1(n11509), .A2(n11495), .ZN(n10001) );
  NAND3_X1 U12810 ( .A1(n12857), .A2(n13955), .A3(n10267), .ZN(n10003) );
  XNOR2_X2 U12811 ( .A(n10004), .B(n12650), .ZN(n13652) );
  NAND2_X2 U12812 ( .A1(n12611), .A2(n12610), .ZN(n10004) );
  NOR2_X2 U12813 ( .A1(n12561), .A2(n12552), .ZN(n12633) );
  NAND2_X4 U12814 ( .A1(n13369), .A2(n13374), .ZN(n12566) );
  INV_X1 U12815 ( .A(n11440), .ZN(n11445) );
  NAND3_X1 U12816 ( .A1(n13968), .A2(n14029), .A3(n13969), .ZN(n10012) );
  OAI21_X2 U12817 ( .B1(n9852), .B2(n10015), .A(n10014), .ZN(n10059) );
  XNOR2_X1 U12818 ( .A(n10498), .B(n10497), .ZN(n10553) );
  NAND2_X2 U12819 ( .A1(n10029), .A2(n20447), .ZN(n10636) );
  NAND2_X2 U12820 ( .A1(n10030), .A2(n10031), .ZN(n10600) );
  NAND3_X1 U12821 ( .A1(n10033), .A2(n14695), .A3(n10032), .ZN(n14676) );
  NAND3_X1 U12822 ( .A1(n10033), .A2(n9854), .A3(n10032), .ZN(n10034) );
  NAND2_X1 U12823 ( .A1(n10573), .A2(n20968), .ZN(n10569) );
  NAND2_X1 U12824 ( .A1(n10573), .A2(n9897), .ZN(n10037) );
  AND2_X1 U12825 ( .A1(n14629), .A2(n10043), .ZN(n11268) );
  INV_X2 U12826 ( .A(n16173), .ZN(n14728) );
  NAND2_X1 U12827 ( .A1(n13993), .A2(n13992), .ZN(n12672) );
  INV_X2 U12828 ( .A(n11453), .ZN(n11998) );
  NAND2_X2 U12829 ( .A1(n11389), .A2(n11388), .ZN(n11453) );
  NAND3_X1 U12830 ( .A1(n11451), .A2(n11450), .A3(n11998), .ZN(n12817) );
  NAND2_X1 U12831 ( .A1(n10045), .A2(n15465), .ZN(n14353) );
  NAND2_X1 U12832 ( .A1(n15466), .A2(n15464), .ZN(n10045) );
  NAND2_X1 U12833 ( .A1(n10049), .A2(n10053), .ZN(n10281) );
  NAND2_X1 U12834 ( .A1(n16402), .A2(n10050), .ZN(n10049) );
  INV_X1 U12835 ( .A(n12292), .ZN(n17680) );
  NAND2_X1 U12836 ( .A1(n12292), .A2(n10072), .ZN(n10063) );
  NAND2_X1 U12837 ( .A1(n12285), .A2(n12286), .ZN(n17770) );
  NOR2_X2 U12838 ( .A1(n12161), .A2(n17075), .ZN(n17325) );
  NAND3_X1 U12839 ( .A1(n10067), .A2(n9850), .A3(n9875), .ZN(n10065) );
  INV_X1 U12840 ( .A(n10067), .ZN(n17984) );
  XNOR2_X1 U12841 ( .A(n12259), .B(n18292), .ZN(n17969) );
  NOR2_X1 U12842 ( .A1(n17649), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12295) );
  NAND2_X1 U12843 ( .A1(n17902), .A2(n10075), .ZN(n10074) );
  NAND2_X1 U12844 ( .A1(n10081), .A2(n10082), .ZN(n16801) );
  NAND2_X1 U12845 ( .A1(n10089), .A2(n9900), .ZN(P3_U2641) );
  NAND3_X1 U12846 ( .A1(n16744), .A2(n10088), .A3(n10087), .ZN(n10086) );
  NAND2_X1 U12847 ( .A1(n10090), .A2(n17066), .ZN(n10089) );
  NOR2_X1 U12848 ( .A1(n16745), .A2(n16974), .ZN(n16738) );
  NAND2_X1 U12849 ( .A1(n16718), .A2(n9931), .ZN(n17684) );
  INV_X1 U12850 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10094) );
  INV_X1 U12851 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U12852 ( .A1(n10103), .A2(n10096), .ZN(n17772) );
  NAND2_X1 U12853 ( .A1(n10115), .A2(n9927), .ZN(n14560) );
  NAND2_X1 U12854 ( .A1(n13042), .A2(n10123), .ZN(n13548) );
  NAND2_X1 U12855 ( .A1(n12036), .A2(n10124), .ZN(n12039) );
  NAND3_X1 U12856 ( .A1(n10456), .A2(n13349), .A3(n13669), .ZN(n10124) );
  NAND2_X1 U12857 ( .A1(n11286), .A2(n9865), .ZN(n11289) );
  INV_X1 U12858 ( .A(n11286), .ZN(n11290) );
  INV_X1 U12859 ( .A(n10143), .ZN(n11322) );
  NAND3_X1 U12860 ( .A1(n10148), .A2(n10560), .A3(n13346), .ZN(n13417) );
  NAND2_X1 U12861 ( .A1(n13346), .A2(n13347), .ZN(n13414) );
  NAND2_X1 U12862 ( .A1(n10560), .A2(n10580), .ZN(n13415) );
  NAND3_X1 U12863 ( .A1(n13711), .A2(n13710), .A3(n10702), .ZN(n13735) );
  AND3_X2 U12864 ( .A1(n13711), .A2(n13710), .A3(n9930), .ZN(n13950) );
  NAND2_X1 U12865 ( .A1(n10151), .A2(n10150), .ZN(n14548) );
  NAND2_X1 U12866 ( .A1(n14534), .A2(n9925), .ZN(n14457) );
  NAND2_X1 U12867 ( .A1(n13974), .A2(n10158), .ZN(n14049) );
  INV_X1 U12868 ( .A(n14049), .ZN(n10816) );
  NOR2_X1 U12869 ( .A1(n14430), .A2(n10160), .ZN(n14419) );
  NOR2_X1 U12870 ( .A1(n14430), .A2(n14431), .ZN(n11272) );
  OR2_X2 U12871 ( .A1(n14430), .A2(n10163), .ZN(n14420) );
  NAND2_X1 U12872 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
  INV_X1 U12873 ( .A(n13328), .ZN(n10166) );
  NOR2_X1 U12874 ( .A1(n10441), .A2(n10168), .ZN(n10442) );
  NOR2_X1 U12875 ( .A1(n10460), .A2(n10168), .ZN(n10462) );
  NAND2_X1 U12876 ( .A1(n16191), .A2(n11221), .ZN(n10169) );
  NAND2_X1 U12877 ( .A1(n14622), .A2(n11267), .ZN(n10170) );
  INV_X1 U12878 ( .A(n11268), .ZN(n10171) );
  AOI22_X1 U12879 ( .A1(n11268), .A2(n10175), .B1(n14622), .B2(n10173), .ZN(
        n10172) );
  NAND2_X1 U12880 ( .A1(n11196), .A2(n10178), .ZN(n10177) );
  NAND2_X1 U12881 ( .A1(n13568), .A2(n11196), .ZN(n13599) );
  NAND2_X1 U12882 ( .A1(n13570), .A2(n13569), .ZN(n13568) );
  NAND2_X1 U12883 ( .A1(n14108), .A2(n10189), .ZN(n17161) );
  NAND3_X1 U12884 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U12885 ( .A1(n10197), .A2(n10196), .ZN(n10195) );
  INV_X1 U12886 ( .A(n15243), .ZN(n10196) );
  NAND2_X1 U12887 ( .A1(n10205), .A2(n15267), .ZN(n10204) );
  INV_X1 U12888 ( .A(n10205), .ZN(n15342) );
  NAND2_X1 U12889 ( .A1(n10201), .A2(n10199), .ZN(n15328) );
  NAND2_X1 U12890 ( .A1(n10205), .A2(n10202), .ZN(n10201) );
  OAI22_X2 U12891 ( .A1(n11475), .A2(n19237), .B1(n11476), .B2(n10206), .ZN(
        n11514) );
  AOI21_X1 U12892 ( .B1(n11514), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11496), .ZN(n11505) );
  NOR2_X2 U12893 ( .A1(n13924), .A2(n9913), .ZN(n15170) );
  INV_X1 U12894 ( .A(n13900), .ZN(n13923) );
  INV_X1 U12895 ( .A(n11519), .ZN(n10216) );
  NOR2_X4 U12896 ( .A1(n15123), .A2(n10217), .ZN(n15157) );
  INV_X1 U12897 ( .A(n10257), .ZN(n10217) );
  NAND2_X1 U12898 ( .A1(n14039), .A2(n10233), .ZN(n15835) );
  NAND2_X1 U12899 ( .A1(n14935), .A2(n9942), .ZN(n14912) );
  AND2_X1 U12900 ( .A1(n14935), .A2(n14938), .ZN(n14936) );
  NAND2_X1 U12901 ( .A1(n12821), .A2(n11998), .ZN(n10244) );
  INV_X1 U12902 ( .A(n10246), .ZN(n14987) );
  NAND2_X1 U12903 ( .A1(n12723), .A2(n9926), .ZN(n12749) );
  AND2_X4 U12904 ( .A1(n10257), .A2(n15879), .ZN(n15308) );
  AND2_X4 U12905 ( .A1(n10257), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11638) );
  NOR2_X4 U12906 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10257) );
  NOR2_X1 U12907 ( .A1(n16502), .A2(n13119), .ZN(n10259) );
  AND2_X2 U12908 ( .A1(n15599), .A2(n9867), .ZN(n15553) );
  NOR2_X2 U12909 ( .A1(n15539), .A2(n10260), .ZN(n15503) );
  INV_X1 U12910 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10262) );
  NOR2_X1 U12911 ( .A1(n15475), .A2(n9961), .ZN(n15468) );
  AOI21_X1 U12912 ( .B1(n9899), .B2(n10273), .A(n10302), .ZN(n13268) );
  INV_X1 U12913 ( .A(n12527), .ZN(n10274) );
  NAND2_X1 U12914 ( .A1(n12653), .A2(n10276), .ZN(n10275) );
  NAND2_X1 U12915 ( .A1(n10275), .A2(n10278), .ZN(n13717) );
  NAND2_X1 U12916 ( .A1(n10281), .A2(n10282), .ZN(n15683) );
  NAND2_X1 U12917 ( .A1(n15515), .A2(n12785), .ZN(n15499) );
  INV_X1 U12918 ( .A(n12785), .ZN(n10290) );
  NOR2_X2 U12919 ( .A1(n14338), .A2(n12806), .ZN(n14341) );
  OAI21_X1 U12920 ( .B1(n13268), .B2(n13267), .A(n13384), .ZN(n13382) );
  INV_X1 U12921 ( .A(n10636), .ZN(n10638) );
  NAND2_X1 U12922 ( .A1(n15800), .A2(n15801), .ZN(n15799) );
  AOI21_X1 U12923 ( .B1(n19163), .B2(n19310), .A(n14372), .ZN(n14375) );
  NAND2_X1 U12924 ( .A1(n10816), .A2(n10815), .ZN(n14084) );
  CLKBUF_X1 U12925 ( .A(n13176), .Z(n20684) );
  AOI21_X1 U12926 ( .B1(n13278), .B2(n20287), .A(n13277), .ZN(n13279) );
  NAND2_X1 U12927 ( .A1(n10397), .A2(n13003), .ZN(n10398) );
  NAND2_X1 U12928 ( .A1(n12699), .A2(n9872), .ZN(n12858) );
  XNOR2_X1 U12929 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12896) );
  AND2_X1 U12930 ( .A1(n19347), .A2(n19354), .ZN(n19868) );
  NAND2_X1 U12931 ( .A1(n12853), .A2(n12849), .ZN(n12851) );
  BUF_X8 U12932 ( .A(n10401), .Z(n11075) );
  AND2_X4 U12933 ( .A1(n10322), .A2(n10332), .ZN(n10401) );
  NAND2_X1 U12934 ( .A1(n10541), .A2(n20413), .ZN(n10544) );
  NAND2_X1 U12935 ( .A1(n11449), .A2(n11448), .ZN(n11476) );
  NAND2_X1 U12936 ( .A1(n12936), .A2(n13630), .ZN(n11449) );
  AND2_X1 U12937 ( .A1(n11683), .A2(n11988), .ZN(n12941) );
  NAND2_X2 U12938 ( .A1(n20287), .A2(n13280), .ZN(n13306) );
  NAND2_X1 U12939 ( .A1(n11374), .A2(n11408), .ZN(n11375) );
  OAI21_X1 U12940 ( .B1(n12615), .B2(n12587), .A(n12586), .ZN(n12597) );
  NAND2_X1 U12941 ( .A1(n12595), .A2(n12594), .ZN(n12596) );
  NAND2_X1 U12942 ( .A1(n16502), .A2(n12543), .ZN(n12544) );
  AND4_X1 U12943 ( .A1(n12603), .A2(n12602), .A3(n12601), .A4(n12600), .ZN(
        n12604) );
  AOI22_X1 U12944 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11361) );
  CLKBUF_X1 U12945 ( .A(n13719), .Z(n13721) );
  AND2_X1 U12946 ( .A1(n14396), .A2(n14395), .ZN(n10293) );
  NOR2_X1 U12947 ( .A1(n20620), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10294) );
  NOR2_X1 U12948 ( .A1(n10466), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10295) );
  INV_X1 U12949 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14355) );
  AND2_X1 U12950 ( .A1(n10545), .A2(n11177), .ZN(n10296) );
  AND4_X1 U12951 ( .A1(n12679), .A2(n12678), .A3(n12677), .A4(n12676), .ZN(
        n10297) );
  AND2_X1 U12952 ( .A1(n12217), .A2(n12216), .ZN(n10298) );
  AND2_X1 U12953 ( .A1(n12018), .A2(n12017), .ZN(n10299) );
  AND2_X1 U12954 ( .A1(n11378), .A2(n11377), .ZN(n10300) );
  INV_X1 U12955 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20865) );
  CLKBUF_X1 U12956 ( .A(n16687), .Z(n16688) );
  OR2_X1 U12957 ( .A1(n18963), .A2(n17493), .ZN(n10301) );
  NOR2_X1 U12958 ( .A1(n13266), .A2(n13376), .ZN(n10302) );
  INV_X1 U12959 ( .A(n14841), .ZN(n11257) );
  INV_X1 U12960 ( .A(n20270), .ZN(n20271) );
  AND2_X2 U12961 ( .A1(n12510), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20270)
         );
  AND2_X1 U12962 ( .A1(n10574), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10303) );
  INV_X1 U12963 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18233) );
  AND2_X1 U12964 ( .A1(n14362), .A2(n15465), .ZN(n10304) );
  NOR2_X1 U12965 ( .A1(n14392), .A2(n14391), .ZN(n10305) );
  NAND2_X1 U12966 ( .A1(n12941), .A2(n12942), .ZN(n11477) );
  NOR2_X1 U12967 ( .A1(n13353), .A2(n20964), .ZN(n10651) );
  INV_X2 U12968 ( .A(n19256), .ZN(n19288) );
  INV_X1 U12969 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11285) );
  AND2_X1 U12970 ( .A1(n11617), .A2(n11458), .ZN(n10306) );
  INV_X1 U12971 ( .A(n11664), .ZN(n11809) );
  INV_X1 U12972 ( .A(n11626), .ZN(n15121) );
  AND4_X1 U12973 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n10307) );
  NAND2_X1 U12974 ( .A1(n17827), .A2(n17993), .ZN(n17700) );
  INV_X1 U12975 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13100) );
  AND4_X1 U12976 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n10308) );
  AND3_X1 U12977 ( .A1(n11927), .A2(n11926), .A3(n11925), .ZN(n13639) );
  INV_X1 U12978 ( .A(n13639), .ZN(n13640) );
  AND2_X1 U12979 ( .A1(n12804), .A2(n14342), .ZN(n10309) );
  NAND2_X1 U12980 ( .A1(n17367), .A2(n18367), .ZN(n17365) );
  AND4_X1 U12981 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10310) );
  AND4_X1 U12982 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10311) );
  AND2_X1 U12983 ( .A1(n13501), .A2(n13500), .ZN(n10312) );
  AND4_X1 U12984 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10313) );
  AND3_X1 U12985 ( .A1(n11125), .A2(n11124), .A3(n11123), .ZN(n11130) );
  OAI22_X1 U12986 ( .A1(n19442), .A2(n12541), .B1(n12620), .B2(n12540), .ZN(
        n12542) );
  AOI22_X1 U12987 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19636), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U12988 ( .A1(n19573), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12548) );
  OR2_X1 U12989 ( .A1(n10648), .A2(n10647), .ZN(n11227) );
  INV_X1 U12990 ( .A(n12654), .ZN(n11595) );
  NAND2_X1 U12991 ( .A1(n12948), .A2(n11425), .ZN(n11448) );
  AND4_X1 U12992 ( .A1(n12638), .A2(n12637), .A3(n12636), .A4(n12635), .ZN(
        n12639) );
  NAND2_X1 U12993 ( .A1(n10447), .A2(n13353), .ZN(n10397) );
  INV_X1 U12994 ( .A(n11638), .ZN(n15120) );
  NAND2_X1 U12995 ( .A1(n12883), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12001) );
  OAI21_X1 U12996 ( .B1(n12846), .B2(n12646), .A(n19112), .ZN(n12703) );
  AOI22_X1 U12997 ( .A1(n11636), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U12998 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U12999 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11626), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U13000 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11330) );
  OAI21_X1 U13001 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n12415), .A(
        n12417), .ZN(n12418) );
  AND2_X1 U13002 ( .A1(n11140), .A2(n11139), .ZN(n11142) );
  AND2_X1 U13003 ( .A1(n10797), .A2(n14047), .ZN(n10798) );
  INV_X1 U13004 ( .A(n13737), .ZN(n10702) );
  OR2_X1 U13005 ( .A1(n10536), .A2(n10535), .ZN(n11177) );
  OR2_X1 U13006 ( .A1(n10672), .A2(n10671), .ZN(n11226) );
  OR2_X1 U13007 ( .A1(n10620), .A2(n10619), .ZN(n11205) );
  INV_X1 U13008 ( .A(n11162), .ZN(n11117) );
  XNOR2_X1 U13009 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11602) );
  INV_X1 U13010 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U13011 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  OAI21_X1 U13012 ( .B1(n9872), .B2(n12699), .A(n12858), .ZN(n12846) );
  AOI22_X1 U13013 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11368) );
  INV_X1 U13014 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16505) );
  NAND2_X1 U13015 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12197) );
  INV_X1 U13016 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21237) );
  AOI21_X1 U13017 ( .B1(n20945), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11142), .ZN(n11153) );
  OR2_X1 U13018 ( .A1(n11012), .A2(n14640), .ZN(n11014) );
  INV_X1 U13019 ( .A(n11095), .ZN(n11068) );
  INV_X1 U13020 ( .A(n13609), .ZN(n10659) );
  AND2_X1 U13021 ( .A1(n10557), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10574) );
  OR2_X1 U13022 ( .A1(n10522), .A2(n10521), .ZN(n11176) );
  NAND3_X1 U13023 ( .A1(n10447), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13280), 
        .ZN(n11143) );
  INV_X1 U13024 ( .A(n11175), .ZN(n10562) );
  NAND2_X1 U13025 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20006), .ZN(
        n12654) );
  OR2_X1 U13026 ( .A1(n15214), .A2(n15218), .ZN(n15240) );
  AND4_X1 U13027 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11748) );
  AND2_X1 U13028 ( .A1(n10305), .A2(n14394), .ZN(n14395) );
  AND2_X1 U13029 ( .A1(n15490), .A2(n12803), .ZN(n14342) );
  AND2_X1 U13030 ( .A1(n12883), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U13031 ( .A1(n13396), .A2(n19825), .ZN(n13373) );
  OR2_X1 U13032 ( .A1(n12918), .A2(n12915), .ZN(n12916) );
  INV_X1 U13033 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n21243) );
  AND2_X1 U13034 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12270), .ZN(
        n12271) );
  AND2_X1 U13035 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12265), .ZN(
        n12266) );
  INV_X1 U13036 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17282) );
  INV_X1 U13037 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n21140) );
  AOI221_X1 U13038 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11153), 
        .C1(n13208), .C2(n11153), .A(n11152), .ZN(n12027) );
  INV_X1 U13039 ( .A(n10973), .ZN(n10974) );
  OR2_X1 U13040 ( .A1(n12032), .A2(n20221), .ZN(n12033) );
  AND2_X1 U13041 ( .A1(n12087), .A2(n12086), .ZN(n14053) );
  OR2_X1 U13042 ( .A1(n16044), .A2(n12030), .ZN(n10956) );
  OR2_X1 U13043 ( .A1(n11051), .A2(n11050), .ZN(n11105) );
  OR2_X1 U13044 ( .A1(n11014), .A2(n11013), .ZN(n11032) );
  NOR2_X1 U13045 ( .A1(n10416), .A2(n20968), .ZN(n11095) );
  INV_X1 U13046 ( .A(n10812), .ZN(n10761) );
  NOR2_X1 U13047 ( .A1(n11170), .A2(n11194), .ZN(n11171) );
  AND2_X1 U13048 ( .A1(n12513), .A2(n13309), .ZN(n11224) );
  NAND2_X1 U13049 ( .A1(n12027), .A2(n11157), .ZN(n11158) );
  INV_X1 U13050 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15974) );
  NAND2_X1 U13051 ( .A1(n10585), .A2(n10584), .ZN(n20448) );
  NOR2_X1 U13052 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16512), .ZN(
        n11599) );
  AND3_X1 U13053 ( .A1(n11575), .A2(n11574), .A3(n11573), .ZN(n15376) );
  AND2_X1 U13054 ( .A1(n15260), .A2(n15266), .ZN(n15284) );
  AND2_X1 U13055 ( .A1(n15142), .A2(n15141), .ZN(n15192) );
  NOR2_X1 U13056 ( .A1(n14927), .A2(n14364), .ZN(n14340) );
  AND2_X1 U13057 ( .A1(n15668), .A2(n15676), .ZN(n15657) );
  AND2_X1 U13058 ( .A1(n16431), .A2(n15796), .ZN(n15715) );
  NOR2_X1 U13059 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12413), .ZN(
        n12429) );
  NOR2_X1 U13060 ( .A1(n12200), .A2(n12199), .ZN(n12205) );
  NAND2_X1 U13061 ( .A1(n16578), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12476) );
  INV_X1 U13062 ( .A(n17818), .ZN(n17819) );
  INV_X1 U13063 ( .A(n18167), .ZN(n18190) );
  NOR2_X1 U13064 ( .A1(n10974), .A2(n14656), .ZN(n10975) );
  AND2_X1 U13065 ( .A1(n12109), .A2(n12108), .ZN(n14527) );
  INV_X1 U13066 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16114) );
  INV_X1 U13067 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16121) );
  INV_X1 U13068 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20076) );
  AND2_X1 U13069 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10602), .ZN(
        n10627) );
  OR2_X1 U13070 ( .A1(n13002), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12146) );
  AND2_X1 U13071 ( .A1(n12105), .A2(n12104), .ZN(n14531) );
  OR2_X1 U13072 ( .A1(n10792), .A2(n16121), .ZN(n10768) );
  OR2_X1 U13073 ( .A1(n10719), .A2(n20065), .ZN(n10720) );
  INV_X1 U13074 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11269) );
  OR2_X1 U13075 ( .A1(n13041), .A2(n13061), .ZN(n20244) );
  OR2_X1 U13076 ( .A1(n20417), .A2(n20948), .ZN(n20799) );
  OR2_X1 U13077 ( .A1(n14890), .A2(n20447), .ZN(n20534) );
  INV_X1 U13078 ( .A(n11174), .ZN(n20265) );
  NOR2_X1 U13079 ( .A1(n20622), .A2(n20454), .ZN(n20765) );
  INV_X1 U13080 ( .A(n20680), .ZN(n20948) );
  INV_X1 U13081 ( .A(n19147), .ZN(n19126) );
  AOI221_X1 U13082 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11610), 
        .C1(n13100), .C2(n11610), .A(n11599), .ZN(n12918) );
  AND2_X1 U13083 ( .A1(n13782), .A2(n13781), .ZN(n13785) );
  OAI21_X1 U13084 ( .B1(n12998), .B2(n12997), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12999) );
  INV_X1 U13085 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14270) );
  INV_X1 U13086 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13217) );
  OR3_X1 U13087 ( .A1(n19371), .A2(n19369), .A3(n19574), .ZN(n19398) );
  INV_X1 U13088 ( .A(n19436), .ZN(n19581) );
  INV_X1 U13089 ( .A(n19635), .ZN(n19602) );
  OR2_X1 U13090 ( .A1(n19981), .A2(n19990), .ZN(n19973) );
  NOR2_X1 U13091 ( .A1(n20017), .A2(n16540), .ZN(n19238) );
  NOR2_X1 U13092 ( .A1(n17654), .A2(n16769), .ZN(n16768) );
  NOR2_X1 U13093 ( .A1(n17718), .A2(n16822), .ZN(n16821) );
  NOR2_X1 U13094 ( .A1(n16839), .A2(n16838), .ZN(n16837) );
  NOR2_X1 U13095 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16916), .ZN(n16905) );
  NOR2_X1 U13096 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16941), .ZN(n16924) );
  NOR2_X1 U13097 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16987), .ZN(n16964) );
  INV_X1 U13098 ( .A(n17054), .ZN(n17076) );
  NOR4_X1 U13099 ( .A1(n17489), .A2(n17463), .A3(n17626), .A4(n17552), .ZN(
        n17375) );
  NOR2_X1 U13100 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18819), .ZN(n17827) );
  NOR2_X1 U13101 ( .A1(n17715), .A2(n16561), .ZN(n18002) );
  NOR2_X1 U13102 ( .A1(n10094), .A2(n16728), .ZN(n16727) );
  NOR2_X1 U13103 ( .A1(n17989), .A2(n17748), .ZN(n17747) );
  OAI21_X1 U13104 ( .B1(n16006), .B2(n10072), .A(n16005), .ZN(n16007) );
  NAND2_X1 U13105 ( .A1(n15959), .A2(n12272), .ZN(n17780) );
  NOR2_X1 U13106 ( .A1(n12277), .A2(n17809), .ZN(n18132) );
  INV_X1 U13107 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18280) );
  INV_X1 U13108 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18292) );
  NOR2_X2 U13109 ( .A1(n15936), .A2(n12408), .ZN(n18788) );
  INV_X1 U13110 ( .A(n18674), .ZN(n18626) );
  NOR2_X1 U13111 ( .A1(n12335), .A2(n12334), .ZN(n18354) );
  AOI22_X1 U13112 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12377) );
  INV_X1 U13113 ( .A(n16000), .ZN(n20967) );
  NAND2_X1 U13114 ( .A1(n10975), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11012) );
  AND2_X1 U13115 ( .A1(n10929), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10973) );
  NOR2_X1 U13116 ( .A1(n10892), .A2(n10904), .ZN(n10928) );
  XNOR2_X1 U13117 ( .A(n11106), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13666) );
  INV_X1 U13118 ( .A(n16104), .ZN(n20089) );
  INV_X1 U13119 ( .A(n14564), .ZN(n20153) );
  INV_X1 U13120 ( .A(n13345), .ZN(n20203) );
  NAND2_X1 U13122 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n10738), .ZN(
        n10792) );
  INV_X1 U13123 ( .A(n20048), .ZN(n20225) );
  OR2_X1 U13124 ( .A1(n14811), .A2(n14221), .ZN(n14800) );
  AND2_X1 U13125 ( .A1(n16224), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14849) );
  NAND2_X1 U13126 ( .A1(n13205), .A2(n20968), .ZN(n11167) );
  INV_X1 U13127 ( .A(n20244), .ZN(n14878) );
  INV_X2 U13128 ( .A(n20252), .ZN(n20221) );
  INV_X1 U13129 ( .A(n20254), .ZN(n20234) );
  INV_X1 U13130 ( .A(n16238), .ZN(n14856) );
  OAI22_X1 U13131 ( .A1(n20279), .A2(n20278), .B1(n20562), .B2(n20450), .ZN(
        n20347) );
  INV_X1 U13132 ( .A(n20351), .ZN(n20374) );
  OAI21_X1 U13133 ( .B1(n20384), .B2(n20383), .A(n20382), .ZN(n20409) );
  NOR2_X2 U13134 ( .A1(n20426), .A2(n20755), .ZN(n20442) );
  NOR2_X2 U13135 ( .A1(n20426), .A2(n20649), .ZN(n20472) );
  NOR2_X2 U13136 ( .A1(n20534), .A2(n20728), .ZN(n20522) );
  NOR2_X2 U13137 ( .A1(n20534), .A2(n20755), .ZN(n20552) );
  INV_X1 U13138 ( .A(n20564), .ZN(n20585) );
  INV_X1 U13139 ( .A(n20679), .ZN(n20557) );
  NOR2_X2 U13140 ( .A1(n20655), .A2(n20728), .ZN(n20644) );
  NOR2_X2 U13141 ( .A1(n20655), .A2(n20755), .ZN(n20675) );
  INV_X1 U13142 ( .A(n20695), .ZN(n20722) );
  NOR2_X2 U13143 ( .A1(n20800), .A2(n20679), .ZN(n20751) );
  INV_X1 U13144 ( .A(n20761), .ZN(n20788) );
  INV_X1 U13145 ( .A(n20713), .ZN(n20826) );
  INV_X1 U13146 ( .A(n20720), .ZN(n20840) );
  AND2_X1 U13147 ( .A1(n15995), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13201) );
  INV_X1 U13148 ( .A(n20972), .ZN(n16015) );
  INV_X1 U13149 ( .A(n20917), .ZN(n20902) );
  INV_X1 U13150 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20874) );
  AOI21_X1 U13151 ( .B1(n16539), .B2(n12826), .A(n12825), .ZN(n12927) );
  AND2_X1 U13152 ( .A1(n20019), .A2(n12016), .ZN(n19102) );
  INV_X1 U13153 ( .A(n19155), .ZN(n19115) );
  INV_X1 U13154 ( .A(n15395), .ZN(n15368) );
  INV_X1 U13155 ( .A(n15397), .ZN(n15383) );
  NOR2_X1 U13156 ( .A1(n13790), .A2(n13789), .ZN(n19168) );
  AND2_X1 U13157 ( .A1(n19198), .A2(n13303), .ZN(n19223) );
  INV_X2 U13158 ( .A(n13101), .ZN(n19306) );
  INV_X1 U13159 ( .A(n15692), .ZN(n16340) );
  AND2_X1 U13160 ( .A1(n16429), .A2(n13235), .ZN(n16420) );
  NOR2_X1 U13161 ( .A1(n16461), .A2(n12964), .ZN(n15855) );
  AND2_X1 U13162 ( .A1(n13816), .A2(n13815), .ZN(n19309) );
  INV_X1 U13163 ( .A(n19318), .ZN(n15847) );
  INV_X1 U13164 ( .A(n19312), .ZN(n16471) );
  NAND2_X1 U13165 ( .A1(n16523), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19965) );
  NOR2_X2 U13166 ( .A1(n19602), .A2(n19546), .ZN(n19400) );
  OR2_X1 U13167 ( .A1(n19414), .A2(n19576), .ZN(n19432) );
  INV_X1 U13168 ( .A(n19968), .ZN(n19694) );
  AND2_X1 U13169 ( .A1(n19436), .A2(n19968), .ZN(n19512) );
  OR2_X1 U13170 ( .A1(n19981), .A2(n15906), .ZN(n19755) );
  AND2_X1 U13171 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13370), .ZN(
        n19609) );
  NOR2_X1 U13172 ( .A1(n19581), .A2(n19973), .ZN(n19624) );
  OAI21_X1 U13173 ( .B1(n15916), .B2(n15915), .A(n15914), .ZN(n19683) );
  NOR2_X2 U13174 ( .A1(n19780), .A2(n19694), .ZN(n19717) );
  AND2_X1 U13175 ( .A1(n19695), .A2(n19691), .ZN(n19716) );
  AND2_X1 U13176 ( .A1(n19756), .A2(n19752), .ZN(n19775) );
  INV_X1 U13177 ( .A(n19755), .ZN(n19758) );
  AND2_X1 U13178 ( .A1(n19355), .A2(n19354), .ZN(n19875) );
  AND3_X1 U13179 ( .A1(n19897), .A2(n19948), .A3(n19902), .ZN(n20027) );
  INV_X1 U13180 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19908) );
  INV_X1 U13181 ( .A(n17021), .ZN(n18985) );
  NOR2_X1 U13182 ( .A1(n18784), .A2(n18288), .ZN(n18035) );
  NOR2_X1 U13183 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16795), .ZN(n16776) );
  NOR2_X1 U13184 ( .A1(n18889), .A2(n16836), .ZN(n16825) );
  NOR2_X1 U13185 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16892), .ZN(n16878) );
  NOR2_X1 U13186 ( .A1(n18875), .A2(n16904), .ZN(n16897) );
  INV_X1 U13187 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17812) );
  INV_X1 U13188 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17297) );
  INV_X1 U13189 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n12475) );
  NOR2_X1 U13190 ( .A1(n18810), .A2(n16716), .ZN(n17054) );
  INV_X1 U13191 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16988) );
  NAND2_X1 U13192 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17405), .ZN(n17404) );
  NOR2_X1 U13193 ( .A1(n17545), .A2(n17441), .ZN(n17436) );
  NAND2_X1 U13194 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17458), .ZN(n17454) );
  INV_X1 U13195 ( .A(n12257), .ZN(n12436) );
  INV_X1 U13196 ( .A(n17512), .ZN(n17521) );
  INV_X1 U13197 ( .A(n17631), .ZN(n17620) );
  NOR2_X1 U13198 ( .A1(n18972), .A2(n17623), .ZN(n17624) );
  OAI21_X1 U13199 ( .B1(n17989), .B2(n17700), .A(n18364), .ZN(n17843) );
  INV_X1 U13200 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17660) );
  INV_X1 U13201 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18066) );
  NOR2_X1 U13202 ( .A1(n18191), .A2(n18133), .ZN(n17817) );
  AOI21_X1 U13203 ( .B1(n18958), .B2(n15951), .A(n18817), .ZN(n17825) );
  INV_X1 U13204 ( .A(n17877), .ZN(n17903) );
  INV_X1 U13205 ( .A(n17993), .ZN(n17946) );
  NOR2_X1 U13206 ( .A1(n18972), .A2(n16697), .ZN(n17986) );
  NOR2_X1 U13207 ( .A1(n9816), .A2(n21268), .ZN(n16604) );
  NOR2_X1 U13208 ( .A1(n16561), .A2(n18095), .ZN(n18008) );
  INV_X1 U13209 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17764) );
  INV_X1 U13210 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21056) );
  AOI21_X1 U13211 ( .B1(n18178), .B2(n18177), .A(n18302), .ZN(n18213) );
  NAND2_X1 U13212 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17992), .ZN(
        n17991) );
  NAND2_X1 U13213 ( .A1(n12475), .A2(n18333), .ZN(n18674) );
  INV_X1 U13214 ( .A(n18451), .ZN(n18457) );
  INV_X1 U13215 ( .A(n18474), .ZN(n18480) );
  INV_X1 U13216 ( .A(n18521), .ZN(n18527) );
  INV_X1 U13217 ( .A(n18660), .ZN(n18667) );
  INV_X1 U13218 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18819) );
  INV_X1 U13219 ( .A(n18973), .ZN(n18836) );
  INV_X1 U13220 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18838) );
  INV_X1 U13221 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20965) );
  INV_X1 U13222 ( .A(n12153), .ZN(n12154) );
  OR2_X1 U13223 ( .A1(n13666), .A2(n13664), .ZN(n16104) );
  NOR2_X1 U13224 ( .A1(n12519), .A2(n12518), .ZN(n12520) );
  INV_X1 U13225 ( .A(n16051), .ZN(n14590) );
  INV_X1 U13226 ( .A(n20186), .ZN(n20172) );
  INV_X1 U13227 ( .A(n20170), .ZN(n20188) );
  NOR2_X1 U13228 ( .A1(n13308), .A2(n13307), .ZN(n13521) );
  OAI21_X1 U13229 ( .B1(n14766), .B2(n20048), .A(n11282), .ZN(n11283) );
  INV_X1 U13230 ( .A(n16092), .ZN(n14700) );
  INV_X1 U13231 ( .A(n16169), .ZN(n20230) );
  OR2_X1 U13232 ( .A1(n11167), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20252) );
  OR2_X1 U13233 ( .A1(n13041), .A2(n13040), .ZN(n20254) );
  OR2_X1 U13234 ( .A1(n13041), .A2(n13037), .ZN(n20250) );
  INV_X1 U13235 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20952) );
  INV_X1 U13236 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13208) );
  OR2_X1 U13237 ( .A1(n20426), .A2(n20679), .ZN(n20351) );
  OR2_X1 U13238 ( .A1(n20426), .A2(n20728), .ZN(n20403) );
  AOI22_X1 U13239 ( .A1(n20381), .A2(n20383), .B1(n10294), .B2(n20622), .ZN(
        n20412) );
  AOI22_X1 U13240 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20421), .B1(n20420), 
        .B2(n20424), .ZN(n20446) );
  NAND2_X1 U13241 ( .A1(n20528), .A2(n20557), .ZN(n20499) );
  AOI22_X1 U13242 ( .A1(n20505), .A2(n20502), .B1(n10294), .B2(n20686), .ZN(
        n20526) );
  NAND2_X1 U13243 ( .A1(n20528), .A2(n20527), .ZN(n20564) );
  NAND2_X1 U13244 ( .A1(n20939), .A2(n20557), .ZN(n20617) );
  AOI22_X1 U13245 ( .A1(n20627), .A2(n20623), .B1(n20622), .B2(n20621), .ZN(
        n20648) );
  OR2_X1 U13246 ( .A1(n20655), .A2(n20649), .ZN(n20695) );
  AOI22_X1 U13247 ( .A1(n20692), .A2(n20689), .B1(n20686), .B2(n20685), .ZN(
        n20727) );
  NAND2_X1 U13248 ( .A1(n20757), .A2(n20729), .ZN(n20761) );
  INV_X1 U13249 ( .A(n20842), .ZN(n20784) );
  INV_X1 U13250 ( .A(n20707), .ZN(n20825) );
  INV_X1 U13251 ( .A(n13201), .ZN(n20042) );
  NOR2_X1 U13252 ( .A1(n20867), .A2(n20976), .ZN(n20933) );
  INV_X1 U13253 ( .A(n20961), .ZN(n20919) );
  NAND2_X1 U13254 ( .A1(n20865), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20961) );
  AND2_X1 U13255 ( .A1(n13092), .A2(n13295), .ZN(n20019) );
  INV_X1 U13256 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19007) );
  NAND2_X1 U13257 ( .A1(n20019), .A2(n11614), .ZN(n19149) );
  INV_X1 U13258 ( .A(n19102), .ZN(n19145) );
  INV_X1 U13259 ( .A(n9962), .ZN(n19110) );
  AND2_X1 U13260 ( .A1(n13296), .A2(n13295), .ZN(n19198) );
  NAND2_X1 U13261 ( .A1(n13301), .A2(n19198), .ZN(n19227) );
  INV_X1 U13262 ( .A(n19200), .ZN(n19231) );
  OR2_X1 U13263 ( .A1(n19301), .A2(n19239), .ZN(n19268) );
  NAND2_X1 U13264 ( .A1(n19236), .A2(n20027), .ZN(n19301) );
  OR2_X1 U13265 ( .A1(n13079), .A2(n15910), .ZN(n19233) );
  INV_X1 U13266 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16359) );
  INV_X1 U13267 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16389) );
  NAND2_X1 U13268 ( .A1(n12974), .A2(n20010), .ZN(n19318) );
  OR2_X1 U13269 ( .A1(n18992), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19324) );
  INV_X1 U13270 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20006) );
  INV_X1 U13271 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19336) );
  AOI211_X2 U13272 ( .C1(n15900), .C2(n15899), .A(n15898), .B(n19576), .ZN(
        n19364) );
  NAND2_X1 U13273 ( .A1(n19635), .A2(n19436), .ZN(n19435) );
  OR2_X1 U13274 ( .A1(n19546), .A2(n19694), .ZN(n19461) );
  INV_X1 U13275 ( .A(n19512), .ZN(n19523) );
  OR2_X1 U13276 ( .A1(n19546), .A2(n19755), .ZN(n19534) );
  INV_X1 U13277 ( .A(n19569), .ZN(n19559) );
  INV_X1 U13278 ( .A(n19594), .ZN(n19601) );
  INV_X1 U13279 ( .A(n19624), .ZN(n19632) );
  INV_X1 U13280 ( .A(n19658), .ZN(n19654) );
  AOI211_X2 U13281 ( .C1(n15909), .C2(n15915), .A(n15908), .B(n19576), .ZN(
        n19687) );
  INV_X1 U13282 ( .A(n19717), .ZN(n19714) );
  NAND2_X1 U13283 ( .A1(n19759), .A2(n19968), .ZN(n19750) );
  INV_X1 U13284 ( .A(n19772), .ZN(n19779) );
  INV_X1 U13285 ( .A(n19846), .ZN(n19799) );
  INV_X1 U13286 ( .A(n19878), .ZN(n19823) );
  INV_X1 U13287 ( .A(n19804), .ZN(n19861) );
  OR2_X1 U13288 ( .A1(n19891), .A2(n20017), .ZN(n16553) );
  INV_X1 U13289 ( .A(n19959), .ZN(n19892) );
  CLKBUF_X1 U13290 ( .A(n19950), .Z(n19947) );
  NAND2_X1 U13291 ( .A1(n18928), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18822) );
  NAND2_X1 U13292 ( .A1(n18035), .A2(n17825), .ZN(n16697) );
  INV_X1 U13293 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17859) );
  NOR2_X1 U13294 ( .A1(n17096), .A2(n17095), .ZN(n17115) );
  INV_X1 U13295 ( .A(n17365), .ZN(n17371) );
  AND2_X1 U13296 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17399), .ZN(n17398) );
  INV_X1 U13297 ( .A(n9811), .ZN(n17483) );
  NOR2_X1 U13298 ( .A1(n12182), .A2(n12181), .ZN(n17500) );
  INV_X1 U13299 ( .A(n20978), .ZN(n17548) );
  OR2_X1 U13300 ( .A1(n18928), .A2(n17994), .ZN(n17570) );
  NAND2_X1 U13301 ( .A1(n17580), .A2(n17526), .ZN(n17578) );
  INV_X1 U13302 ( .A(n17624), .ZN(n17627) );
  AND2_X1 U13303 ( .A1(n12481), .A2(n12480), .ZN(n12482) );
  NAND2_X1 U13304 ( .A1(n10077), .A2(n17874), .ZN(n17792) );
  INV_X1 U13305 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18169) );
  INV_X1 U13306 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18212) );
  OAI21_X1 U13307 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18966), .A(n16697), 
        .ZN(n17993) );
  INV_X1 U13308 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17989) );
  NAND3_X1 U13309 ( .A1(n18315), .A2(n18808), .A3(n15959), .ZN(n18221) );
  INV_X1 U13310 ( .A(n18315), .ZN(n18302) );
  AND2_X1 U13311 ( .A1(n18983), .A2(n16692), .ZN(n18966) );
  INV_X1 U13312 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18798) );
  INV_X1 U13313 ( .A(n18644), .ZN(n18637) );
  INV_X1 U13314 ( .A(n18657), .ZN(n18736) );
  INV_X1 U13315 ( .A(n18967), .ZN(n18817) );
  INV_X1 U13316 ( .A(n18917), .ZN(n18915) );
  INV_X1 U13317 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18845) );
  NOR2_X1 U13318 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13000), .ZN(n16670)
         );
  INV_X1 U13319 ( .A(n16647), .ZN(n16652) );
  INV_X1 U13320 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19911) );
  OR2_X1 U13321 ( .A1(n11284), .A2(n11283), .ZN(P1_U2971) );
  OAI21_X1 U13322 ( .B1(n16595), .B2(n17877), .A(n12482), .ZN(P3_U2799) );
  NOR2_X4 U13323 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10333) );
  AND2_X2 U13324 ( .A1(n13491), .A2(n10333), .ZN(n10365) );
  NAND2_X1 U13325 ( .A1(n10365), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10320) );
  NAND2_X1 U13326 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10319) );
  NAND2_X1 U13327 ( .A1(n10708), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10318) );
  NAND2_X1 U13328 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10317) );
  AND2_X2 U13329 ( .A1(n10321), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10327) );
  NAND2_X1 U13330 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10326) );
  NAND2_X1 U13331 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10325) );
  NAND2_X1 U13332 ( .A1(n10359), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10324) );
  NAND2_X1 U13333 ( .A1(n10366), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10323) );
  NAND2_X1 U13334 ( .A1(n10421), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10330) );
  NAND2_X1 U13335 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10329) );
  NAND2_X1 U13336 ( .A1(n10506), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10328) );
  AND2_X2 U13337 ( .A1(n13490), .A2(n14894), .ZN(n10610) );
  NAND2_X1 U13338 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10338) );
  NAND2_X1 U13339 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U13340 ( .A1(n10488), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10336) );
  AND2_X2 U13341 ( .A1(n10334), .A2(n14894), .ZN(n10360) );
  NAND2_X1 U13342 ( .A1(n10360), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10335) );
  AOI22_X1 U13343 ( .A1(n9845), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13344 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13345 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13346 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13347 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9832), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13348 ( .A1(n9833), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13349 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10506), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13350 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10347) );
  INV_X1 U13351 ( .A(n10397), .ZN(n10374) );
  AOI22_X1 U13352 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10389), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13353 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9837), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13354 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9840), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13355 ( .A1(n9830), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10506), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13356 ( .A1(n9845), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13357 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13358 ( .A1(n10421), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10401), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13359 ( .A1(n10359), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10355) );
  AND2_X2 U13360 ( .A1(n10313), .A2(n10311), .ZN(n10446) );
  AOI22_X1 U13361 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9836), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13362 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10421), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13363 ( .A1(n9834), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10389), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13364 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9838), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10361) );
  NAND4_X1 U13365 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10373) );
  AOI22_X1 U13366 ( .A1(n10708), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13367 ( .A1(n9832), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9829), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13368 ( .A1(n10367), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13369 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10506), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U13370 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10372) );
  OR2_X2 U13371 ( .A1(n10373), .A2(n10372), .ZN(n10448) );
  INV_X1 U13372 ( .A(n13009), .ZN(n10413) );
  AOI22_X1 U13373 ( .A1(n9845), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13374 ( .A1(n9832), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9833), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13375 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13376 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10384) );
  AOI22_X1 U13377 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9836), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13378 ( .A1(n9834), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13379 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10506), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13380 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10379) );
  NAND4_X1 U13381 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10383) );
  OR2_X2 U13382 ( .A1(n10384), .A2(n10383), .ZN(n13019) );
  NAND2_X1 U13383 ( .A1(n10416), .A2(n13019), .ZN(n10400) );
  INV_X2 U13384 ( .A(n10446), .ZN(n12492) );
  NAND2_X1 U13385 ( .A1(n10448), .A2(n12492), .ZN(n10396) );
  AOI22_X1 U13386 ( .A1(n9845), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13387 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9836), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13388 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9834), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13389 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9839), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U13390 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10395) );
  AOI22_X1 U13391 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9832), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13392 ( .A1(n9833), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13393 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10506), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13394 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10390) );
  NAND4_X1 U13395 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10394) );
  NAND2_X1 U13396 ( .A1(n13353), .A2(n12492), .ZN(n13003) );
  NAND3_X1 U13397 ( .A1(n10400), .A2(n10399), .A3(n10398), .ZN(n10444) );
  AOI22_X1 U13398 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13399 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10359), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13400 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10402) );
  NAND4_X1 U13401 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10411) );
  AOI22_X1 U13402 ( .A1(n9833), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13403 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10506), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13404 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10406) );
  NAND4_X1 U13405 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10410) );
  NAND2_X1 U13406 ( .A1(n10444), .A2(n20274), .ZN(n13024) );
  NAND2_X1 U13407 ( .A1(n10413), .A2(n10412), .ZN(n10415) );
  NAND2_X1 U13408 ( .A1(n20323), .A2(n12492), .ZN(n10414) );
  NAND2_X1 U13409 ( .A1(n13012), .A2(n10416), .ZN(n10443) );
  NAND2_X1 U13410 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10420) );
  NAND2_X1 U13411 ( .A1(n10708), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13412 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13413 ( .A1(n10359), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10417) );
  NAND2_X1 U13414 ( .A1(n10610), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13415 ( .A1(n9832), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10424) );
  NAND2_X1 U13416 ( .A1(n9833), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U13417 ( .A1(n10506), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U13418 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10429) );
  NAND2_X1 U13419 ( .A1(n10365), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10428) );
  NAND2_X1 U13420 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10427) );
  NAND2_X1 U13421 ( .A1(n9839), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10426) );
  NAND2_X1 U13422 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10433) );
  NAND2_X1 U13423 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10431) );
  NAND2_X1 U13424 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10430) );
  NAND4_X4 U13425 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n13309) );
  NAND2_X1 U13426 ( .A1(n13280), .A2(n13193), .ZN(n10439) );
  INV_X1 U13427 ( .A(n12494), .ZN(n10440) );
  NAND2_X1 U13428 ( .A1(n20274), .A2(n13309), .ZN(n13668) );
  NAND2_X1 U13429 ( .A1(n10440), .A2(n13668), .ZN(n10441) );
  NAND3_X1 U13430 ( .A1(n13024), .A2(n10443), .A3(n10442), .ZN(n13029) );
  NAND2_X1 U13431 ( .A1(n13029), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10465) );
  INV_X1 U13432 ( .A(n10444), .ZN(n12023) );
  NOR2_X1 U13433 ( .A1(n11117), .A2(n13280), .ZN(n12022) );
  AND2_X1 U13434 ( .A1(n20287), .A2(n12022), .ZN(n10445) );
  INV_X2 U13435 ( .A(n13193), .ZN(n20298) );
  AND2_X1 U13436 ( .A1(n10446), .A2(n13353), .ZN(n10450) );
  NOR2_X1 U13437 ( .A1(n10447), .A2(n12513), .ZN(n10449) );
  AND3_X2 U13438 ( .A1(n11160), .A2(n10450), .A3(n10449), .ZN(n13190) );
  NAND2_X1 U13439 ( .A1(n13190), .A2(n13349), .ZN(n12485) );
  AND2_X2 U13440 ( .A1(n12488), .A2(n12485), .ZN(n13034) );
  INV_X1 U13441 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n10451) );
  XNOR2_X1 U13442 ( .A(n10451), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12138) );
  NOR2_X1 U13443 ( .A1(n13003), .A2(n12513), .ZN(n10452) );
  NAND2_X2 U13444 ( .A1(n10454), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10471) );
  MUX2_X1 U13445 ( .A(n11167), .B(n15995), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10455) );
  INV_X1 U13446 ( .A(n12496), .ZN(n13663) );
  INV_X1 U13447 ( .A(n12041), .ZN(n10456) );
  AND2_X1 U13448 ( .A1(n13663), .A2(n12121), .ZN(n13055) );
  NAND2_X1 U13449 ( .A1(n13009), .A2(n13019), .ZN(n10459) );
  INV_X1 U13450 ( .A(n10457), .ZN(n10458) );
  AOI22_X1 U13451 ( .A1(n13055), .A2(n10459), .B1(n10458), .B2(n20966), .ZN(
        n10463) );
  NAND2_X1 U13452 ( .A1(n12494), .A2(n10446), .ZN(n13026) );
  NAND4_X1 U13453 ( .A1(n13026), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13205), 
        .A4(n13668), .ZN(n10460) );
  NAND3_X1 U13454 ( .A1(n13012), .A2(n10416), .A3(n13309), .ZN(n10461) );
  NAND4_X1 U13455 ( .A1(n13024), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10499) );
  NAND2_X1 U13456 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10475) );
  OAI21_X1 U13457 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10475), .ZN(n20620) );
  OR2_X1 U13458 ( .A1(n15995), .A2(n20687), .ZN(n10469) );
  OAI21_X1 U13459 ( .B1(n11167), .B2(n20620), .A(n10469), .ZN(n10466) );
  INV_X1 U13460 ( .A(n10466), .ZN(n10464) );
  AND2_X1 U13461 ( .A1(n10469), .A2(n10316), .ZN(n10470) );
  NAND2_X1 U13462 ( .A1(n10544), .A2(n10481), .ZN(n10479) );
  NOR2_X1 U13463 ( .A1(n15995), .A2(n15974), .ZN(n10473) );
  INV_X1 U13464 ( .A(n11167), .ZN(n10477) );
  INV_X1 U13465 ( .A(n10475), .ZN(n10474) );
  NAND2_X1 U13466 ( .A1(n10474), .A2(n15974), .ZN(n20651) );
  NAND2_X1 U13467 ( .A1(n10475), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10476) );
  NAND2_X1 U13468 ( .A1(n20651), .A2(n10476), .ZN(n20277) );
  NAND2_X1 U13469 ( .A1(n10477), .A2(n20277), .ZN(n10480) );
  NAND2_X1 U13470 ( .A1(n10482), .A2(n10480), .ZN(n10478) );
  NAND2_X1 U13471 ( .A1(n10479), .A2(n10478), .ZN(n10581) );
  NAND4_X1 U13472 ( .A1(n10544), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10483) );
  NAND2_X1 U13473 ( .A1(n10581), .A2(n10483), .ZN(n13176) );
  AOI22_X1 U13474 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13475 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9836), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10486) );
  INV_X1 U13476 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21213) );
  AOI22_X1 U13477 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13478 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13479 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10494) );
  AOI22_X1 U13480 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13481 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13482 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13483 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10489) );
  NAND4_X1 U13484 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10493) );
  INV_X1 U13485 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10496) );
  OAI22_X1 U13486 ( .A1(n11191), .A2(n10586), .B1(n11143), .B2(n10496), .ZN(
        n10497) );
  INV_X1 U13487 ( .A(n10499), .ZN(n10500) );
  AOI22_X1 U13488 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13489 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13490 ( .A1(n9832), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11075), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13491 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10502) );
  NAND4_X1 U13492 ( .A1(n10505), .A2(n10504), .A3(n10503), .A4(n10502), .ZN(
        n10512) );
  AOI22_X1 U13493 ( .A1(n10708), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13494 ( .A1(n9830), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13495 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10507) );
  NAND4_X1 U13496 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10511) );
  INV_X1 U13497 ( .A(n11235), .ZN(n10523) );
  AOI22_X1 U13498 ( .A1(n9824), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13499 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9832), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13500 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13501 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10513) );
  NAND4_X1 U13502 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10522) );
  AOI22_X1 U13503 ( .A1(n9845), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13504 ( .A1(n10752), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9835), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13505 ( .A1(n10389), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13506 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10517) );
  NAND4_X1 U13507 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10521) );
  XNOR2_X1 U13508 ( .A(n10523), .B(n11176), .ZN(n10524) );
  NAND2_X1 U13509 ( .A1(n10524), .A2(n10545), .ZN(n10568) );
  NAND2_X1 U13510 ( .A1(n10545), .A2(n11235), .ZN(n11170) );
  INV_X1 U13511 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n21187) );
  AOI21_X1 U13512 ( .B1(n10412), .B2(n11235), .A(n20968), .ZN(n10526) );
  NAND2_X1 U13513 ( .A1(n20274), .A2(n11176), .ZN(n10525) );
  OAI211_X1 U13514 ( .C1(n11143), .C2(n21187), .A(n10526), .B(n10525), .ZN(
        n10570) );
  NAND2_X1 U13515 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10540) );
  OR2_X1 U13516 ( .A1(n10587), .A2(n11235), .ZN(n10539) );
  INV_X1 U13517 ( .A(n10586), .ZN(n10537) );
  AOI22_X1 U13518 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9841), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13519 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13520 ( .A1(n9835), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10527) );
  NAND4_X1 U13521 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10536) );
  AOI22_X1 U13522 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13523 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13524 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13525 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10531) );
  NAND4_X1 U13526 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10535) );
  NAND2_X1 U13527 ( .A1(n10537), .A2(n11177), .ZN(n10538) );
  INV_X1 U13528 ( .A(n20413), .ZN(n10543) );
  INV_X1 U13529 ( .A(n10541), .ZN(n10542) );
  NAND2_X1 U13530 ( .A1(n10543), .A2(n10542), .ZN(n20352) );
  NAND2_X1 U13531 ( .A1(n20352), .A2(n10544), .ZN(n13516) );
  AOI21_X2 U13532 ( .B1(n10546), .B2(n20968), .A(n10296), .ZN(n11175) );
  NAND2_X1 U13533 ( .A1(n10561), .A2(n11175), .ZN(n10551) );
  INV_X1 U13534 ( .A(n10547), .ZN(n10548) );
  NAND2_X1 U13535 ( .A1(n10553), .A2(n10552), .ZN(n10554) );
  INV_X1 U13536 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13447) );
  XNOR2_X1 U13537 ( .A(n13447), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20137) );
  NAND2_X1 U13538 ( .A1(n20964), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10810) );
  OAI21_X1 U13539 ( .B1(n20137), .B2(n12030), .A(n10810), .ZN(n10555) );
  AOI21_X1 U13540 ( .B1(n11100), .B2(P1_EAX_REG_2__SCAN_IN), .A(n10555), .ZN(
        n10556) );
  INV_X1 U13541 ( .A(n10556), .ZN(n10558) );
  INV_X1 U13542 ( .A(n13003), .ZN(n10557) );
  OAI21_X2 U13543 ( .B1(n14890), .B2(n10812), .A(n10559), .ZN(n10560) );
  NAND2_X1 U13544 ( .A1(n11099), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13545 ( .A1(n13515), .A2(n10761), .ZN(n10567) );
  AOI22_X1 U13546 ( .A1(n11100), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20964), .ZN(n10565) );
  NAND2_X1 U13547 ( .A1(n10574), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10564) );
  AND2_X1 U13548 ( .A1(n10565), .A2(n10564), .ZN(n10566) );
  NAND2_X1 U13549 ( .A1(n10567), .A2(n10566), .ZN(n13347) );
  NAND2_X1 U13550 ( .A1(n10569), .A2(n10568), .ZN(n10571) );
  XNOR2_X2 U13551 ( .A(n10571), .B(n10570), .ZN(n11174) );
  NAND2_X1 U13552 ( .A1(n11174), .A2(n10446), .ZN(n10572) );
  NAND2_X1 U13553 ( .A1(n10572), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13355) );
  INV_X1 U13554 ( .A(n10574), .ZN(n10625) );
  NAND2_X1 U13555 ( .A1(n10651), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13556 ( .A1(n20964), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10575) );
  OAI211_X1 U13557 ( .C1(n10625), .C2(n10321), .A(n10576), .B(n10575), .ZN(
        n10577) );
  AOI21_X1 U13558 ( .B1(n10573), .B2(n10761), .A(n10577), .ZN(n10578) );
  OR2_X1 U13559 ( .A1(n13355), .A2(n10578), .ZN(n13356) );
  INV_X1 U13560 ( .A(n10578), .ZN(n13357) );
  OR2_X1 U13561 ( .A1(n13357), .A2(n12030), .ZN(n10579) );
  NAND2_X1 U13562 ( .A1(n13356), .A2(n10579), .ZN(n13346) );
  NAND2_X1 U13563 ( .A1(n10472), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10585) );
  NOR3_X1 U13564 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15974), .A3(
        n20687), .ZN(n20535) );
  NAND2_X1 U13565 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20535), .ZN(
        n20533) );
  NAND2_X1 U13566 ( .A1(n20945), .A2(n20533), .ZN(n10582) );
  NAND3_X1 U13567 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20795) );
  INV_X1 U13568 ( .A(n20795), .ZN(n20802) );
  NAND2_X1 U13569 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20802), .ZN(
        n20796) );
  NAND2_X1 U13570 ( .A1(n10582), .A2(n20796), .ZN(n20560) );
  OAI22_X1 U13571 ( .A1(n11167), .A2(n20560), .B1(n15995), .B2(n20945), .ZN(
        n10583) );
  INV_X1 U13572 ( .A(n10583), .ZN(n10584) );
  NAND2_X1 U13573 ( .A1(n20558), .A2(n20968), .ZN(n10599) );
  AOI22_X1 U13574 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13575 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9836), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10590) );
  INV_X1 U13576 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n21175) );
  AOI22_X1 U13577 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13578 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10588) );
  NAND4_X1 U13579 ( .A1(n10591), .A2(n10590), .A3(n10589), .A4(n10588), .ZN(
        n10597) );
  AOI22_X1 U13580 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13581 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13582 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13583 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13584 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10596) );
  AOI22_X1 U13585 ( .A1(n11157), .A2(n11206), .B1(n11122), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10598) );
  NAND2_X1 U13586 ( .A1(n10600), .A2(n20264), .ZN(n10601) );
  NAND2_X1 U13587 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10603) );
  INV_X1 U13588 ( .A(n10603), .ZN(n10602) );
  INV_X1 U13589 ( .A(n10627), .ZN(n10629) );
  INV_X1 U13590 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10604) );
  NAND2_X1 U13591 ( .A1(n10604), .A2(n10603), .ZN(n10605) );
  NAND2_X1 U13592 ( .A1(n10629), .A2(n10605), .ZN(n13693) );
  AOI22_X1 U13593 ( .A1(n13693), .A2(n11098), .B1(n11099), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13594 ( .A1(n11100), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10606) );
  OAI211_X1 U13595 ( .C1(n10625), .C2(n10315), .A(n10607), .B(n10606), .ZN(
        n10608) );
  INV_X1 U13596 ( .A(n10608), .ZN(n10609) );
  OAI21_X1 U13597 ( .B1(n11190), .B2(n10812), .A(n10609), .ZN(n13544) );
  NAND2_X1 U13598 ( .A1(n13545), .A2(n13544), .ZN(n13543) );
  INV_X1 U13599 ( .A(n13543), .ZN(n10635) );
  AOI22_X1 U13600 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13601 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13602 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10611) );
  NAND4_X1 U13603 ( .A1(n10614), .A2(n10613), .A3(n10612), .A4(n10611), .ZN(
        n10620) );
  AOI22_X1 U13604 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9831), .B1(n9821), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13605 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9835), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13606 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13607 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9830), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10615) );
  NAND4_X1 U13608 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10619) );
  NAND2_X1 U13609 ( .A1(n11157), .A2(n11205), .ZN(n10622) );
  NAND2_X1 U13610 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10621) );
  XNOR2_X1 U13611 ( .A(n10636), .B(n10637), .ZN(n11197) );
  NAND2_X1 U13612 ( .A1(n20964), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10624) );
  NAND2_X1 U13613 ( .A1(n11100), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10623) );
  OAI211_X1 U13614 ( .C1(n10625), .C2(n13208), .A(n10624), .B(n10623), .ZN(
        n10626) );
  NAND2_X1 U13615 ( .A1(n10626), .A2(n12030), .ZN(n10632) );
  INV_X1 U13616 ( .A(n10652), .ZN(n10653) );
  INV_X1 U13617 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13618 ( .A1(n10629), .A2(n10628), .ZN(n10630) );
  NAND2_X1 U13619 ( .A1(n10653), .A2(n10630), .ZN(n20229) );
  NAND2_X1 U13620 ( .A1(n20229), .A2(n11098), .ZN(n10631) );
  NAND2_X1 U13621 ( .A1(n10632), .A2(n10631), .ZN(n10633) );
  AOI21_X1 U13622 ( .B1(n11197), .B2(n10761), .A(n10633), .ZN(n13576) );
  NAND2_X1 U13623 ( .A1(n10635), .A2(n10634), .ZN(n13610) );
  INV_X1 U13624 ( .A(n13610), .ZN(n10660) );
  AOI22_X1 U13625 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13626 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13627 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10640) );
  INV_X1 U13628 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n21162) );
  AOI22_X1 U13629 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10639) );
  NAND4_X1 U13630 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10648) );
  AOI22_X1 U13631 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13632 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13633 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9837), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U13634 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10647) );
  NAND2_X1 U13635 ( .A1(n11157), .A2(n11227), .ZN(n10650) );
  NAND2_X1 U13636 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10649) );
  XNOR2_X1 U13637 ( .A(n10661), .B(n10662), .ZN(n11204) );
  INV_X1 U13638 ( .A(n10651), .ZN(n11093) );
  INV_X1 U13639 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10657) );
  INV_X1 U13640 ( .A(n10673), .ZN(n10655) );
  INV_X1 U13641 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20101) );
  NAND2_X1 U13642 ( .A1(n10653), .A2(n20101), .ZN(n10654) );
  NAND2_X1 U13643 ( .A1(n10655), .A2(n10654), .ZN(n20105) );
  AOI22_X1 U13644 ( .A1(n20105), .A2(n11098), .B1(n11099), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10656) );
  OAI21_X1 U13645 ( .B1(n11093), .B2(n10657), .A(n10656), .ZN(n10658) );
  AOI21_X1 U13646 ( .B1(n11204), .B2(n10761), .A(n10658), .ZN(n13609) );
  AOI22_X1 U13647 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9840), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13648 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13649 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13650 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10663) );
  NAND4_X1 U13651 ( .A1(n10666), .A2(n10665), .A3(n10664), .A4(n10663), .ZN(
        n10672) );
  AOI22_X1 U13652 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13653 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9836), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13654 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13655 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10667) );
  NAND4_X1 U13656 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(
        n10671) );
  AOI22_X1 U13657 ( .A1(n11157), .A2(n11226), .B1(n11122), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13658 ( .A1(n10678), .A2(n10677), .ZN(n11214) );
  INV_X1 U13659 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10675) );
  OAI21_X1 U13660 ( .B1(n10673), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10682), .ZN(n20093) );
  AOI22_X1 U13661 ( .A1(n20093), .A2(n11098), .B1(n11099), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10674) );
  OAI21_X1 U13662 ( .B1(n11093), .B2(n10675), .A(n10674), .ZN(n10676) );
  NAND2_X1 U13663 ( .A1(n11157), .A2(n11235), .ZN(n10680) );
  NAND2_X1 U13664 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10679) );
  NAND2_X1 U13665 ( .A1(n10680), .A2(n10679), .ZN(n10681) );
  NAND2_X1 U13666 ( .A1(n11225), .A2(n10761), .ZN(n10688) );
  INV_X1 U13667 ( .A(n10682), .ZN(n10684) );
  INV_X1 U13668 ( .A(n10703), .ZN(n10683) );
  OAI21_X1 U13669 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10684), .A(
        n10683), .ZN(n20083) );
  NAND2_X1 U13670 ( .A1(n11098), .A2(n20083), .ZN(n10685) );
  OAI21_X1 U13671 ( .B1(n20076), .B2(n10810), .A(n10685), .ZN(n10686) );
  AOI21_X1 U13672 ( .B1(n11100), .B2(P1_EAX_REG_7__SCAN_IN), .A(n10686), .ZN(
        n10687) );
  NAND2_X1 U13673 ( .A1(n10688), .A2(n10687), .ZN(n13710) );
  NAND2_X1 U13674 ( .A1(n11100), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13675 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13676 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13677 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13678 ( .A1(n9830), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10689) );
  NAND4_X1 U13679 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10698) );
  AOI22_X1 U13680 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9841), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13681 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13682 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13683 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10693) );
  NAND4_X1 U13684 ( .A1(n10696), .A2(n10695), .A3(n10694), .A4(n10693), .ZN(
        n10697) );
  OAI21_X1 U13685 ( .B1(n10698), .B2(n10697), .A(n10761), .ZN(n10700) );
  XNOR2_X1 U13686 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10703), .ZN(
        n14497) );
  AOI22_X1 U13687 ( .A1(n11098), .A2(n14497), .B1(n11099), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10699) );
  XNOR2_X1 U13688 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10719), .ZN(
        n20068) );
  INV_X1 U13689 ( .A(n20068), .ZN(n13989) );
  NAND2_X1 U13690 ( .A1(n11100), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13691 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13692 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13693 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13694 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10704) );
  NAND4_X1 U13695 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10714) );
  AOI22_X1 U13696 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13697 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13698 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U13699 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  OAI21_X1 U13700 ( .B1(n10714), .B2(n10713), .A(n10761), .ZN(n10716) );
  NAND2_X1 U13701 ( .A1(n11099), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10715) );
  NAND3_X1 U13702 ( .A1(n10717), .A2(n10716), .A3(n10715), .ZN(n10718) );
  AOI21_X1 U13703 ( .B1(n13989), .B2(n11098), .A(n10718), .ZN(n13951) );
  NAND2_X1 U13704 ( .A1(n10720), .A2(n21212), .ZN(n10722) );
  INV_X1 U13705 ( .A(n10738), .ZN(n10721) );
  NAND2_X1 U13706 ( .A1(n10722), .A2(n10721), .ZN(n14732) );
  NAND2_X1 U13707 ( .A1(n14732), .A2(n11098), .ZN(n10737) );
  AOI22_X1 U13708 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13709 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13710 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13711 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10723) );
  NAND4_X1 U13712 ( .A1(n10726), .A2(n10725), .A3(n10724), .A4(n10723), .ZN(
        n10732) );
  AOI22_X1 U13713 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9840), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13714 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13715 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10727) );
  NAND4_X1 U13716 ( .A1(n10730), .A2(n10729), .A3(n10728), .A4(n10727), .ZN(
        n10731) );
  OAI21_X1 U13717 ( .B1(n10732), .B2(n10731), .A(n10761), .ZN(n10734) );
  NAND2_X1 U13718 ( .A1(n11100), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10733) );
  OAI211_X1 U13719 ( .C1(n10810), .C2(n21212), .A(n10734), .B(n10733), .ZN(
        n10735) );
  INV_X1 U13720 ( .A(n10735), .ZN(n10736) );
  NAND2_X1 U13721 ( .A1(n10737), .A2(n10736), .ZN(n13973) );
  INV_X1 U13722 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14066) );
  OR2_X1 U13723 ( .A1(n11093), .A2(n14066), .ZN(n10740) );
  OAI21_X1 U13724 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10738), .A(
        n10792), .ZN(n16181) );
  AOI22_X1 U13725 ( .A1(n11098), .A2(n16181), .B1(n11099), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13726 ( .A1(n10740), .A2(n10739), .ZN(n14059) );
  AOI22_X1 U13727 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13728 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10915), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13729 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13730 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10741) );
  NAND4_X1 U13731 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n10750) );
  AOI22_X1 U13732 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13733 ( .A1(n11081), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13734 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13735 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10745) );
  NAND4_X1 U13736 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10749) );
  NOR2_X1 U13737 ( .A1(n10750), .A2(n10749), .ZN(n10751) );
  NOR2_X1 U13738 ( .A1(n10812), .A2(n10751), .ZN(n14073) );
  XNOR2_X1 U13739 ( .A(n10799), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14720) );
  NAND2_X1 U13740 ( .A1(n11100), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13741 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9840), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13742 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13743 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13744 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9837), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10753) );
  NAND4_X1 U13745 ( .A1(n10756), .A2(n10755), .A3(n10754), .A4(n10753), .ZN(
        n10763) );
  AOI22_X1 U13746 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13747 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13748 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13749 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10757) );
  NAND4_X1 U13750 ( .A1(n10760), .A2(n10759), .A3(n10758), .A4(n10757), .ZN(
        n10762) );
  OAI21_X1 U13751 ( .B1(n10763), .B2(n10762), .A(n10761), .ZN(n10765) );
  NAND2_X1 U13752 ( .A1(n11099), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10764) );
  NAND3_X1 U13753 ( .A1(n10766), .A2(n10765), .A3(n10764), .ZN(n10767) );
  AOI21_X1 U13754 ( .B1(n14720), .B2(n11098), .A(n10767), .ZN(n14050) );
  INV_X1 U13755 ( .A(n14050), .ZN(n10797) );
  XNOR2_X1 U13756 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10768), .ZN(
        n14333) );
  AOI22_X1 U13757 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13758 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13759 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13760 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10769) );
  NAND4_X1 U13761 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10778) );
  AOI22_X1 U13762 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13763 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13764 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13765 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10773) );
  NAND4_X1 U13766 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10777) );
  NOR2_X1 U13767 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  OAI22_X1 U13768 ( .A1(n10812), .A2(n10779), .B1(n10810), .B2(n14323), .ZN(
        n10780) );
  AOI21_X1 U13769 ( .B1(n11100), .B2(P1_EAX_REG_13__SCAN_IN), .A(n10780), .ZN(
        n10781) );
  OAI21_X1 U13770 ( .B1(n14333), .B2(n12030), .A(n10781), .ZN(n14299) );
  AOI22_X1 U13771 ( .A1(n10365), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13772 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10915), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13773 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9831), .B1(
        n11075), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13774 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10910), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10782) );
  NAND4_X1 U13775 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10791) );
  AOI22_X1 U13776 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13777 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10916), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13778 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10786) );
  NAND4_X1 U13779 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10790) );
  NOR2_X1 U13780 ( .A1(n10791), .A2(n10790), .ZN(n10796) );
  INV_X1 U13781 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14080) );
  OR2_X1 U13782 ( .A1(n11093), .A2(n14080), .ZN(n10795) );
  XNOR2_X1 U13783 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10792), .ZN(
        n16168) );
  OAI22_X1 U13784 ( .A1(n16168), .A2(n12030), .B1(n10810), .B2(n16121), .ZN(
        n10793) );
  INV_X1 U13785 ( .A(n10793), .ZN(n10794) );
  OAI211_X1 U13786 ( .C1(n10796), .C2(n10812), .A(n10795), .B(n10794), .ZN(
        n14075) );
  AND2_X1 U13787 ( .A1(n14299), .A2(n14075), .ZN(n14047) );
  XNOR2_X1 U13788 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n10817), .ZN(
        n16163) );
  AOI22_X1 U13789 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13790 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13791 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13792 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10800) );
  NAND4_X1 U13793 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10809) );
  AOI22_X1 U13794 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11080), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13795 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13796 ( .A1(n11081), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13797 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10804) );
  NAND4_X1 U13798 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10808) );
  NOR2_X1 U13799 ( .A1(n10809), .A2(n10808), .ZN(n10811) );
  OAI22_X1 U13800 ( .A1(n10812), .A2(n10811), .B1(n10810), .B2(n16114), .ZN(
        n10813) );
  AOI21_X1 U13801 ( .B1(n11100), .B2(P1_EAX_REG_15__SCAN_IN), .A(n10813), .ZN(
        n10814) );
  OAI21_X1 U13802 ( .B1(n16163), .B2(n12030), .A(n10814), .ZN(n10815) );
  INV_X1 U13803 ( .A(n10815), .ZN(n14069) );
  XNOR2_X1 U13804 ( .A(n10831), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16103) );
  AOI22_X1 U13805 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13806 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13807 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13808 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10818) );
  NAND4_X1 U13809 ( .A1(n10821), .A2(n10820), .A3(n10819), .A4(n10818), .ZN(
        n10827) );
  AOI22_X1 U13810 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9840), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13811 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13812 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13813 ( .A1(n10916), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13814 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10826) );
  OAI21_X1 U13815 ( .B1(n10827), .B2(n10826), .A(n11095), .ZN(n10829) );
  AOI22_X1 U13816 ( .A1(n11100), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20964), .ZN(n10828) );
  AOI21_X1 U13817 ( .B1(n10829), .B2(n10828), .A(n11098), .ZN(n10830) );
  AOI21_X1 U13818 ( .B1(n16103), .B2(n11098), .A(n10830), .ZN(n14083) );
  XNOR2_X1 U13819 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10844), .ZN(
        n16155) );
  AOI22_X1 U13820 ( .A1(n11100), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n11099), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13821 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13822 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13823 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13824 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9837), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10832) );
  NAND4_X1 U13825 ( .A1(n10835), .A2(n10834), .A3(n10833), .A4(n10832), .ZN(
        n10841) );
  AOI22_X1 U13826 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9841), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13827 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13828 ( .A1(n10916), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10837) );
  NAND4_X1 U13829 ( .A1(n10839), .A2(n10838), .A3(n10837), .A4(n10836), .ZN(
        n10840) );
  OAI21_X1 U13830 ( .B1(n10841), .B2(n10840), .A(n11095), .ZN(n10842) );
  OAI211_X1 U13831 ( .C1(n16155), .C2(n12030), .A(n10843), .B(n10842), .ZN(
        n14472) );
  INV_X1 U13832 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14692) );
  XNOR2_X1 U13833 ( .A(n10859), .B(n14692), .ZN(n14691) );
  AOI22_X1 U13834 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13835 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13836 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13837 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10845) );
  NAND4_X1 U13838 ( .A1(n10848), .A2(n10847), .A3(n10846), .A4(n10845), .ZN(
        n10854) );
  AOI22_X1 U13839 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13840 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U13841 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13842 ( .A1(n10916), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10849) );
  NAND4_X1 U13843 ( .A1(n10852), .A2(n10851), .A3(n10850), .A4(n10849), .ZN(
        n10853) );
  NOR2_X1 U13844 ( .A1(n10854), .A2(n10853), .ZN(n10857) );
  AOI21_X1 U13845 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14692), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10855) );
  AOI21_X1 U13846 ( .B1(n10651), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10855), .ZN(
        n10856) );
  OAI21_X1 U13847 ( .B1(n11068), .B2(n10857), .A(n10856), .ZN(n10858) );
  OAI21_X1 U13848 ( .B1(n14691), .B2(n12030), .A(n10858), .ZN(n14549) );
  INV_X1 U13849 ( .A(n10891), .ZN(n10862) );
  OR2_X1 U13850 ( .A1(n10860), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10861) );
  NAND2_X1 U13851 ( .A1(n10862), .A2(n10861), .ZN(n16147) );
  AOI22_X1 U13852 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13853 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13854 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13855 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10863) );
  NAND4_X1 U13856 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n10872) );
  AOI22_X1 U13857 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9840), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13858 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13859 ( .A1(n10916), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13860 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10867) );
  NAND4_X1 U13861 ( .A1(n10870), .A2(n10869), .A3(n10868), .A4(n10867), .ZN(
        n10871) );
  NOR2_X1 U13862 ( .A1(n10872), .A2(n10871), .ZN(n10875) );
  OAI21_X1 U13863 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20965), .A(
        n20964), .ZN(n10874) );
  NAND2_X1 U13864 ( .A1(n11100), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n10873) );
  OAI211_X1 U13865 ( .C1(n11068), .C2(n10875), .A(n10874), .B(n10873), .ZN(
        n10876) );
  OAI21_X1 U13866 ( .B1(n16147), .B2(n12030), .A(n10876), .ZN(n14599) );
  INV_X1 U13867 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14684) );
  XNOR2_X1 U13868 ( .A(n10891), .B(n14684), .ZN(n16071) );
  AOI22_X1 U13869 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13870 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9844), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13871 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10915), .B1(
        n10401), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13872 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9831), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10877) );
  NAND4_X1 U13873 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n10886) );
  AOI22_X1 U13874 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10910), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13875 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11055), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13876 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10881) );
  NAND4_X1 U13877 ( .A1(n10884), .A2(n10883), .A3(n10882), .A4(n10881), .ZN(
        n10885) );
  OR2_X1 U13878 ( .A1(n10886), .A2(n10885), .ZN(n10889) );
  INV_X1 U13879 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14593) );
  NAND2_X1 U13880 ( .A1(n20964), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10887) );
  OAI211_X1 U13881 ( .C1(n11093), .C2(n14593), .A(n12030), .B(n10887), .ZN(
        n10888) );
  AOI21_X1 U13882 ( .B1(n11095), .B2(n10889), .A(n10888), .ZN(n10890) );
  AOI21_X1 U13883 ( .B1(n16071), .B2(n11098), .A(n10890), .ZN(n14543) );
  AND2_X2 U13884 ( .A1(n14541), .A2(n14543), .ZN(n14534) );
  AND2_X1 U13885 ( .A1(n10892), .A2(n10904), .ZN(n10893) );
  OR2_X1 U13886 ( .A1(n10893), .A2(n10928), .ZN(n16066) );
  AOI22_X1 U13887 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9840), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13888 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13889 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13890 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9837), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10894) );
  NAND4_X1 U13891 ( .A1(n10897), .A2(n10896), .A3(n10895), .A4(n10894), .ZN(
        n10903) );
  AOI22_X1 U13892 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13893 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13894 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13895 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10898) );
  NAND4_X1 U13896 ( .A1(n10901), .A2(n10900), .A3(n10899), .A4(n10898), .ZN(
        n10902) );
  NOR2_X1 U13897 ( .A1(n10903), .A2(n10902), .ZN(n10907) );
  OAI21_X1 U13898 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n10904), .A(n12030), 
        .ZN(n10905) );
  AOI21_X1 U13899 ( .B1(n10651), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10905), .ZN(
        n10906) );
  OAI21_X1 U13900 ( .B1(n11068), .B2(n10907), .A(n10906), .ZN(n10908) );
  OAI21_X1 U13901 ( .B1(n16066), .B2(n12030), .A(n10908), .ZN(n10909) );
  INV_X1 U13902 ( .A(n10909), .ZN(n14536) );
  INV_X1 U13903 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14672) );
  XNOR2_X1 U13904 ( .A(n10928), .B(n14672), .ZN(n16050) );
  NAND2_X1 U13905 ( .A1(n16050), .A2(n11098), .ZN(n10927) );
  AOI22_X1 U13906 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13907 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13908 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13909 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9837), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10911) );
  NAND4_X1 U13910 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(
        n10922) );
  AOI22_X1 U13911 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13912 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13913 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13914 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10917) );
  NAND4_X1 U13915 ( .A1(n10920), .A2(n10919), .A3(n10918), .A4(n10917), .ZN(
        n10921) );
  NOR2_X1 U13916 ( .A1(n10922), .A2(n10921), .ZN(n10925) );
  AOI21_X1 U13917 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14672), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10923) );
  AOI21_X1 U13918 ( .B1(n10651), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10923), .ZN(
        n10924) );
  OAI21_X1 U13919 ( .B1(n11068), .B2(n10925), .A(n10924), .ZN(n10926) );
  NAND2_X1 U13920 ( .A1(n10927), .A2(n10926), .ZN(n14525) );
  NOR2_X1 U13921 ( .A1(n10929), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10930) );
  OR2_X1 U13922 ( .A1(n10973), .A2(n10930), .ZN(n16044) );
  AOI22_X1 U13923 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9840), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13924 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13925 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13926 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U13927 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10940) );
  AOI22_X1 U13928 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13929 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9830), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13930 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9837), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U13931 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10939) );
  NOR2_X1 U13932 ( .A1(n10940), .A2(n10939), .ZN(n10967) );
  AOI22_X1 U13933 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9841), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13934 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13935 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13936 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10941) );
  NAND4_X1 U13937 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10950) );
  AOI22_X1 U13938 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11075), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13939 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13940 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10945) );
  NAND4_X1 U13941 ( .A1(n10948), .A2(n10947), .A3(n10946), .A4(n10945), .ZN(
        n10949) );
  NOR2_X1 U13942 ( .A1(n10950), .A2(n10949), .ZN(n10968) );
  XNOR2_X1 U13943 ( .A(n10967), .B(n10968), .ZN(n10954) );
  NAND2_X1 U13944 ( .A1(n20964), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10951) );
  NAND2_X1 U13945 ( .A1(n12030), .A2(n10951), .ZN(n10952) );
  AOI21_X1 U13946 ( .B1(n10651), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10952), .ZN(
        n10953) );
  OAI21_X1 U13947 ( .B1(n11068), .B2(n10954), .A(n10953), .ZN(n10955) );
  NAND2_X1 U13948 ( .A1(n10956), .A2(n10955), .ZN(n14583) );
  XOR2_X1 U13949 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n10973), .Z(
        n16033) );
  AOI22_X1 U13950 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13951 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13952 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13953 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10957) );
  NAND4_X1 U13954 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n10966) );
  AOI22_X1 U13955 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13956 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13957 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9837), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10961) );
  NAND4_X1 U13958 ( .A1(n10964), .A2(n10963), .A3(n10962), .A4(n10961), .ZN(
        n10965) );
  OR2_X1 U13959 ( .A1(n10966), .A2(n10965), .ZN(n10979) );
  NOR2_X1 U13960 ( .A1(n10968), .A2(n10967), .ZN(n10980) );
  XOR2_X1 U13961 ( .A(n10979), .B(n10980), .Z(n10971) );
  NAND2_X1 U13962 ( .A1(n11100), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n10969) );
  OAI211_X1 U13963 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14656), .A(n10969), 
        .B(n12030), .ZN(n10970) );
  AOI21_X1 U13964 ( .B1(n10971), .B2(n11095), .A(n10970), .ZN(n10972) );
  AOI21_X1 U13965 ( .B1(n16033), .B2(n11098), .A(n10972), .ZN(n14517) );
  INV_X1 U13966 ( .A(n10975), .ZN(n10977) );
  INV_X1 U13967 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13968 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13969 ( .A1(n11012), .A2(n10978), .ZN(n14652) );
  NAND2_X1 U13970 ( .A1(n10980), .A2(n10979), .ZN(n11006) );
  AOI22_X1 U13971 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U13972 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U13973 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13974 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10982) );
  NAND4_X1 U13975 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n10991) );
  AOI22_X1 U13976 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U13977 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U13978 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U13979 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10986) );
  NAND4_X1 U13980 ( .A1(n10989), .A2(n10988), .A3(n10987), .A4(n10986), .ZN(
        n10990) );
  NOR2_X1 U13981 ( .A1(n10991), .A2(n10990), .ZN(n11007) );
  XNOR2_X1 U13982 ( .A(n11006), .B(n11007), .ZN(n10994) );
  OAI21_X1 U13983 ( .B1(n20965), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20964), .ZN(n10993) );
  NAND2_X1 U13984 ( .A1(n11100), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n10992) );
  OAI211_X1 U13985 ( .C1(n10994), .C2(n11068), .A(n10993), .B(n10992), .ZN(
        n10995) );
  OAI21_X1 U13986 ( .B1(n14652), .B2(n12030), .A(n10995), .ZN(n14458) );
  XNOR2_X1 U13987 ( .A(n11012), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14644) );
  AOI22_X1 U13988 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U13989 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13990 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13991 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10996) );
  NAND4_X1 U13992 ( .A1(n10999), .A2(n10998), .A3(n10997), .A4(n10996), .ZN(
        n11005) );
  AOI22_X1 U13993 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U13994 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13995 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13996 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10360), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11000) );
  NAND4_X1 U13997 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11004) );
  OR2_X1 U13998 ( .A1(n11005), .A2(n11004), .ZN(n11026) );
  NOR2_X1 U13999 ( .A1(n11007), .A2(n11006), .ZN(n11027) );
  XOR2_X1 U14000 ( .A(n11026), .B(n11027), .Z(n11010) );
  INV_X1 U14001 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U14002 ( .A1(n11100), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n11008) );
  OAI211_X1 U14003 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14640), .A(n11008), 
        .B(n12030), .ZN(n11009) );
  AOI21_X1 U14004 ( .B1(n11010), .B2(n11095), .A(n11009), .ZN(n11011) );
  AOI21_X1 U14005 ( .B1(n14644), .B2(n11098), .A(n11011), .ZN(n14444) );
  INV_X1 U14006 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11013) );
  NAND2_X1 U14007 ( .A1(n11014), .A2(n11013), .ZN(n11015) );
  NAND2_X1 U14008 ( .A1(n11032), .A2(n11015), .ZN(n14633) );
  AOI22_X1 U14009 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14010 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10910), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14011 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11075), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14012 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9838), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11016) );
  NAND4_X1 U14013 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11025) );
  AOI22_X1 U14014 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9844), .B1(n9841), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14015 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9831), .B1(n9821), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14016 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14017 ( .A1(n10916), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11020) );
  NAND4_X1 U14018 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11024) );
  NOR2_X1 U14019 ( .A1(n11025), .A2(n11024), .ZN(n11044) );
  NAND2_X1 U14020 ( .A1(n11027), .A2(n11026), .ZN(n11043) );
  XNOR2_X1 U14021 ( .A(n11044), .B(n11043), .ZN(n11030) );
  AOI21_X1 U14022 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20964), .A(
        n11098), .ZN(n11029) );
  NAND2_X1 U14023 ( .A1(n11100), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11028) );
  OAI211_X1 U14024 ( .C1(n11030), .C2(n11068), .A(n11029), .B(n11028), .ZN(
        n11031) );
  XOR2_X1 U14025 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n11049), .Z(
        n14235) );
  AOI22_X1 U14026 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10365), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14027 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14028 ( .A1(n10401), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14029 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11033) );
  NAND4_X1 U14030 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n11042) );
  AOI22_X1 U14031 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14032 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14033 ( .A1(n11082), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U14034 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9837), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11037) );
  NAND4_X1 U14035 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n11041) );
  OR2_X1 U14036 ( .A1(n11042), .A2(n11041), .ZN(n11053) );
  NOR2_X1 U14037 ( .A1(n11044), .A2(n11043), .ZN(n11054) );
  XOR2_X1 U14038 ( .A(n11053), .B(n11054), .Z(n11047) );
  INV_X1 U14039 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14241) );
  NAND2_X1 U14040 ( .A1(n11100), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11045) );
  OAI211_X1 U14041 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14241), .A(n11045), 
        .B(n12030), .ZN(n11046) );
  AOI21_X1 U14042 ( .B1(n11047), .B2(n11095), .A(n11046), .ZN(n11048) );
  AOI21_X1 U14043 ( .B1(n14235), .B2(n11098), .A(n11048), .ZN(n11273) );
  INV_X1 U14044 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U14045 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  NAND2_X1 U14046 ( .A1(n11105), .A2(n11052), .ZN(n14625) );
  NAND2_X1 U14047 ( .A1(n11054), .A2(n11053), .ZN(n11071) );
  AOI22_X1 U14048 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14049 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9821), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14050 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11055), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14051 ( .A1(n9825), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9837), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U14052 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11065) );
  AOI22_X1 U14053 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14054 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U14055 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9839), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11061) );
  NAND4_X1 U14056 ( .A1(n11063), .A2(n11062), .A3(n11061), .A4(n11060), .ZN(
        n11064) );
  NOR2_X1 U14057 ( .A1(n11065), .A2(n11064), .ZN(n11072) );
  XNOR2_X1 U14058 ( .A(n11071), .B(n11072), .ZN(n11069) );
  AOI21_X1 U14059 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20964), .A(
        n11098), .ZN(n11067) );
  NAND2_X1 U14060 ( .A1(n11100), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11066) );
  OAI211_X1 U14061 ( .C1(n11069), .C2(n11068), .A(n11067), .B(n11066), .ZN(
        n11070) );
  OAI21_X1 U14062 ( .B1(n14625), .B2(n12030), .A(n11070), .ZN(n14421) );
  XNOR2_X1 U14063 ( .A(n11105), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14616) );
  NOR2_X1 U14064 ( .A1(n11072), .A2(n11071), .ZN(n11090) );
  AOI22_X1 U14065 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10916), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14066 ( .A1(n10915), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10366), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14067 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14068 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11074), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11076) );
  NAND4_X1 U14069 ( .A1(n11079), .A2(n11078), .A3(n11077), .A4(n11076), .ZN(
        n11088) );
  AOI22_X1 U14070 ( .A1(n11080), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9841), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14071 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11081), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14072 ( .A1(n11055), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11082), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14073 ( .A1(n10910), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9837), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11083) );
  NAND4_X1 U14074 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11087) );
  NOR2_X1 U14075 ( .A1(n11088), .A2(n11087), .ZN(n11089) );
  XNOR2_X1 U14076 ( .A(n11090), .B(n11089), .ZN(n11096) );
  INV_X1 U14077 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n11092) );
  OAI21_X1 U14078 ( .B1(n20965), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n20964), .ZN(n11091) );
  OAI21_X1 U14079 ( .B1(n11093), .B2(n11092), .A(n11091), .ZN(n11094) );
  AOI21_X1 U14080 ( .B1(n11096), .B2(n11095), .A(n11094), .ZN(n11097) );
  AOI21_X1 U14081 ( .B1(n14616), .B2(n11098), .A(n11097), .ZN(n12483) );
  AOI22_X1 U14082 ( .A1(n11100), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11099), .ZN(n11101) );
  INV_X1 U14083 ( .A(n11101), .ZN(n11102) );
  XNOR2_X2 U14084 ( .A(n11103), .B(n11102), .ZN(n14387) );
  NAND3_X1 U14085 ( .A1(n20968), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16285) );
  INV_X1 U14086 ( .A(n16285), .ZN(n11104) );
  NAND2_X1 U14087 ( .A1(n14387), .A2(n16192), .ZN(n11271) );
  INV_X1 U14088 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14618) );
  XNOR2_X1 U14089 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14090 ( .A1(n11120), .A2(n11121), .ZN(n11108) );
  NAND2_X1 U14091 ( .A1(n20687), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11107) );
  NAND2_X1 U14092 ( .A1(n11108), .A2(n11107), .ZN(n11113) );
  MUX2_X1 U14093 ( .A(n15974), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11112) );
  NAND2_X1 U14094 ( .A1(n11113), .A2(n11112), .ZN(n11110) );
  NAND2_X1 U14095 ( .A1(n15974), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14096 ( .A1(n11110), .A2(n11109), .ZN(n11140) );
  XNOR2_X1 U14097 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11139) );
  NAND3_X1 U14098 ( .A1(n13208), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11153), .ZN(n11151) );
  NAND2_X1 U14099 ( .A1(n20323), .A2(n13280), .ZN(n11111) );
  NAND2_X1 U14100 ( .A1(n11111), .A2(n20287), .ZN(n11138) );
  XNOR2_X1 U14101 ( .A(n11113), .B(n11112), .ZN(n12026) );
  INV_X1 U14102 ( .A(n12026), .ZN(n11131) );
  NAND2_X1 U14103 ( .A1(n11157), .A2(n11131), .ZN(n11137) );
  AND2_X1 U14104 ( .A1(n10321), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11114) );
  NOR2_X1 U14105 ( .A1(n11120), .A2(n11114), .ZN(n11116) );
  NAND2_X1 U14106 ( .A1(n11157), .A2(n11116), .ZN(n11115) );
  NAND2_X1 U14107 ( .A1(n11115), .A2(n11150), .ZN(n11119) );
  OAI211_X1 U14108 ( .C1(n11117), .C2(n20274), .A(n11138), .B(n11116), .ZN(
        n11118) );
  NAND2_X1 U14109 ( .A1(n11119), .A2(n11118), .ZN(n11129) );
  INV_X1 U14110 ( .A(n11129), .ZN(n11135) );
  NAND2_X1 U14111 ( .A1(n11157), .A2(n13309), .ZN(n11125) );
  XNOR2_X1 U14112 ( .A(n11121), .B(n11120), .ZN(n12024) );
  NAND2_X1 U14113 ( .A1(n11122), .A2(n12024), .ZN(n11124) );
  NAND2_X1 U14114 ( .A1(n20323), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11123) );
  INV_X1 U14115 ( .A(n11130), .ZN(n11134) );
  INV_X1 U14116 ( .A(n11157), .ZN(n11127) );
  INV_X1 U14117 ( .A(n12024), .ZN(n11126) );
  AOI21_X1 U14118 ( .B1(n11127), .B2(n11224), .A(n11126), .ZN(n11128) );
  OAI21_X1 U14119 ( .B1(n11130), .B2(n11129), .A(n11128), .ZN(n11133) );
  OAI211_X1 U14120 ( .C1(n11131), .C2(n11143), .A(n11137), .B(n11138), .ZN(
        n11132) );
  OAI211_X1 U14121 ( .C1(n11135), .C2(n11134), .A(n11133), .B(n11132), .ZN(
        n11136) );
  OAI21_X1 U14122 ( .B1(n11138), .B2(n11137), .A(n11136), .ZN(n11145) );
  NOR2_X1 U14123 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  NOR2_X1 U14124 ( .A1(n11142), .A2(n11141), .ZN(n11146) );
  NAND2_X1 U14125 ( .A1(n11151), .A2(n11146), .ZN(n12025) );
  NAND2_X1 U14126 ( .A1(n12025), .A2(n11143), .ZN(n11144) );
  NAND2_X1 U14127 ( .A1(n11145), .A2(n11144), .ZN(n11149) );
  INV_X1 U14128 ( .A(n11146), .ZN(n11147) );
  AOI22_X1 U14129 ( .A1(n11154), .A2(n11147), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20968), .ZN(n11148) );
  OAI211_X1 U14130 ( .C1(n11151), .C2(n11150), .A(n11149), .B(n11148), .ZN(
        n11156) );
  INV_X1 U14131 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20263) );
  NOR2_X1 U14132 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20263), .ZN(
        n11152) );
  NAND2_X1 U14133 ( .A1(n12027), .A2(n11154), .ZN(n11155) );
  NAND2_X1 U14134 ( .A1(n11156), .A2(n11155), .ZN(n11159) );
  INV_X1 U14135 ( .A(n11160), .ZN(n11161) );
  AOI21_X1 U14136 ( .B1(n10416), .B2(n20274), .A(n11161), .ZN(n13010) );
  NAND3_X1 U14137 ( .A1(n13010), .A2(n11162), .A3(n13018), .ZN(n13033) );
  NAND2_X1 U14138 ( .A1(n20948), .A2(n11167), .ZN(n20971) );
  NAND2_X1 U14139 ( .A1(n20971), .A2(n20968), .ZN(n11163) );
  NAND2_X1 U14140 ( .A1(n20968), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14141 ( .A1(n20965), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11164) );
  AND2_X1 U14142 ( .A1(n11165), .A2(n11164), .ZN(n13359) );
  INV_X1 U14143 ( .A(n13359), .ZN(n11166) );
  INV_X1 U14144 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20918) );
  NOR2_X1 U14145 ( .A1(n20252), .A2(n20918), .ZN(n14227) );
  AOI21_X1 U14146 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14227), .ZN(n11168) );
  OAI21_X1 U14147 ( .B1(n13666), .B2(n20230), .A(n11168), .ZN(n11169) );
  INV_X1 U14148 ( .A(n11169), .ZN(n11270) );
  NOR2_X1 U14149 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11267) );
  NAND2_X1 U14150 ( .A1(n20274), .A2(n13019), .ZN(n11183) );
  OAI21_X1 U14151 ( .B1(n13306), .B2(n11176), .A(n11183), .ZN(n11172) );
  INV_X1 U14152 ( .A(n11172), .ZN(n11173) );
  OAI21_X2 U14153 ( .B1(n11174), .B2(n11194), .A(n11173), .ZN(n13329) );
  NAND2_X1 U14154 ( .A1(n11175), .A2(n13309), .ZN(n11182) );
  NAND2_X1 U14155 ( .A1(n11176), .A2(n11177), .ZN(n11192) );
  OAI21_X1 U14156 ( .B1(n11177), .B2(n11176), .A(n11192), .ZN(n11178) );
  INV_X1 U14157 ( .A(n11178), .ZN(n11180) );
  NAND3_X1 U14158 ( .A1(n20298), .A2(n12513), .A3(n13019), .ZN(n11179) );
  AOI21_X1 U14159 ( .B1(n20966), .B2(n11180), .A(n11179), .ZN(n11181) );
  INV_X1 U14160 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20261) );
  XNOR2_X2 U14161 ( .A(n11188), .B(n20261), .ZN(n13445) );
  XNOR2_X1 U14162 ( .A(n11192), .B(n11191), .ZN(n11185) );
  INV_X1 U14163 ( .A(n11183), .ZN(n11184) );
  AOI21_X1 U14164 ( .B1(n11185), .B2(n20966), .A(n11184), .ZN(n11186) );
  NAND2_X1 U14165 ( .A1(n11187), .A2(n11186), .ZN(n13444) );
  NAND2_X1 U14166 ( .A1(n11188), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11189) );
  NAND2_X2 U14167 ( .A1(n20257), .A2(n11189), .ZN(n11195) );
  INV_X1 U14168 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20241) );
  NAND2_X1 U14169 ( .A1(n11192), .A2(n11191), .ZN(n11208) );
  XNOR2_X1 U14170 ( .A(n11208), .B(n11206), .ZN(n11193) );
  OAI22_X1 U14171 ( .A1(n11190), .A2(n11194), .B1(n13306), .B2(n11193), .ZN(
        n13569) );
  NAND2_X1 U14172 ( .A1(n11195), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11196) );
  NAND2_X1 U14173 ( .A1(n11197), .A2(n11224), .ZN(n11201) );
  NAND2_X1 U14174 ( .A1(n11208), .A2(n11206), .ZN(n11198) );
  XNOR2_X1 U14175 ( .A(n11198), .B(n11205), .ZN(n11199) );
  NAND2_X1 U14176 ( .A1(n11199), .A2(n20966), .ZN(n11200) );
  NAND2_X1 U14177 ( .A1(n11201), .A2(n11200), .ZN(n11202) );
  INV_X1 U14178 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13603) );
  XNOR2_X1 U14179 ( .A(n11202), .B(n13603), .ZN(n13598) );
  NAND2_X1 U14180 ( .A1(n11202), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U14181 ( .A1(n11204), .A2(n11224), .ZN(n11211) );
  AND2_X1 U14182 ( .A1(n11206), .A2(n11205), .ZN(n11207) );
  NAND2_X1 U14183 ( .A1(n11208), .A2(n11207), .ZN(n11229) );
  XNOR2_X1 U14184 ( .A(n11229), .B(n11227), .ZN(n11209) );
  NAND2_X1 U14185 ( .A1(n11209), .A2(n20966), .ZN(n11210) );
  NAND2_X1 U14186 ( .A1(n11211), .A2(n11210), .ZN(n11212) );
  INV_X1 U14187 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16279) );
  XNOR2_X1 U14188 ( .A(n11212), .B(n16279), .ZN(n16196) );
  NAND2_X1 U14189 ( .A1(n11212), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11213) );
  NAND3_X1 U14190 ( .A1(n11215), .A2(n11224), .A3(n11214), .ZN(n11220) );
  INV_X1 U14191 ( .A(n11229), .ZN(n11216) );
  NAND2_X1 U14192 ( .A1(n11216), .A2(n11227), .ZN(n11217) );
  XNOR2_X1 U14193 ( .A(n11217), .B(n11226), .ZN(n11218) );
  NAND2_X1 U14194 ( .A1(n11218), .A2(n20966), .ZN(n11219) );
  INV_X1 U14195 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16188) );
  NAND2_X1 U14196 ( .A1(n16189), .A2(n16188), .ZN(n11221) );
  INV_X1 U14197 ( .A(n16189), .ZN(n11222) );
  NAND2_X1 U14198 ( .A1(n11222), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14199 ( .A1(n11225), .A2(n11224), .ZN(n11232) );
  NAND2_X1 U14200 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  OR2_X1 U14201 ( .A1(n11229), .A2(n11228), .ZN(n11234) );
  XNOR2_X1 U14202 ( .A(n11234), .B(n11235), .ZN(n11230) );
  NAND2_X1 U14203 ( .A1(n11230), .A2(n20966), .ZN(n11231) );
  NAND2_X1 U14204 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  OR2_X1 U14205 ( .A1(n11233), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16183) );
  NAND2_X1 U14206 ( .A1(n11233), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16182) );
  INV_X1 U14207 ( .A(n11234), .ZN(n11236) );
  NAND3_X1 U14208 ( .A1(n11236), .A2(n20966), .A3(n11235), .ZN(n11237) );
  NAND2_X1 U14209 ( .A1(n16173), .A2(n11237), .ZN(n13931) );
  OR2_X1 U14210 ( .A1(n13931), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11238) );
  NAND2_X1 U14211 ( .A1(n13931), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11239) );
  INV_X1 U14212 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16256) );
  INV_X1 U14213 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U14214 ( .A1(n14728), .A2(n12089), .ZN(n16150) );
  NAND2_X1 U14215 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11240) );
  NAND2_X1 U14216 ( .A1(n16150), .A2(n11240), .ZN(n14705) );
  INV_X1 U14217 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11241) );
  NAND2_X1 U14218 ( .A1(n16173), .A2(n11241), .ZN(n16159) );
  OAI21_X1 U14219 ( .B1(n14728), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16148), .ZN(n11242) );
  INV_X1 U14220 ( .A(n11242), .ZN(n11250) );
  INV_X1 U14221 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U14222 ( .A1(n16173), .A2(n11243), .ZN(n11244) );
  INV_X1 U14223 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11245) );
  NAND2_X1 U14224 ( .A1(n16173), .A2(n11245), .ZN(n14306) );
  NAND2_X1 U14225 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11246) );
  NAND2_X1 U14226 ( .A1(n16173), .A2(n11246), .ZN(n14304) );
  NAND2_X1 U14227 ( .A1(n14306), .A2(n14304), .ZN(n11247) );
  INV_X1 U14228 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14209) );
  NAND2_X1 U14229 ( .A1(n16173), .A2(n14209), .ZN(n11248) );
  NAND2_X1 U14230 ( .A1(n14713), .A2(n11248), .ZN(n14703) );
  INV_X1 U14231 ( .A(n14703), .ZN(n11249) );
  NAND2_X1 U14232 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14305) );
  INV_X1 U14233 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14727) );
  INV_X1 U14234 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11251) );
  NAND2_X1 U14235 ( .A1(n14727), .A2(n11251), .ZN(n11252) );
  NAND2_X1 U14236 ( .A1(n14728), .A2(n11252), .ZN(n14302) );
  AND2_X1 U14237 ( .A1(n14305), .A2(n14302), .ZN(n14701) );
  NAND2_X1 U14238 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11253) );
  AND2_X1 U14239 ( .A1(n14714), .A2(n11253), .ZN(n14702) );
  OAI21_X1 U14240 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n14728), .ZN(n11254) );
  NAND2_X1 U14241 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16160) );
  XNOR2_X1 U14242 ( .A(n16173), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14695) );
  NAND2_X1 U14243 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14841) );
  INV_X1 U14244 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14833) );
  INV_X1 U14245 ( .A(n14696), .ZN(n11261) );
  INV_X1 U14246 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11260) );
  INV_X1 U14247 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11258) );
  INV_X1 U14248 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14687) );
  NAND2_X1 U14249 ( .A1(n11258), .A2(n14687), .ZN(n14842) );
  INV_X1 U14250 ( .A(n14842), .ZN(n11259) );
  NAND4_X1 U14251 ( .A1(n11261), .A2(n11260), .A3(n14833), .A4(n11259), .ZN(
        n11262) );
  NAND3_X1 U14252 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U14253 ( .A1(n11275), .A2(n14779), .ZN(n11264) );
  NAND2_X1 U14254 ( .A1(n11263), .A2(n16173), .ZN(n14646) );
  NAND3_X1 U14255 ( .A1(n11264), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14646), .ZN(n14630) );
  INV_X1 U14256 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14797) );
  INV_X1 U14257 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14786) );
  INV_X1 U14258 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14812) );
  NAND3_X1 U14259 ( .A1(n14797), .A2(n14786), .A3(n14812), .ZN(n11276) );
  INV_X1 U14260 ( .A(n14629), .ZN(n11265) );
  NOR2_X1 U14261 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14755) );
  AND2_X1 U14262 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U14263 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11266) );
  INV_X1 U14264 ( .A(n16192), .ZN(n14699) );
  NOR2_X1 U14265 ( .A1(n14244), .A2(n14699), .ZN(n11284) );
  NAND2_X1 U14266 ( .A1(n16173), .A2(n14779), .ZN(n14637) );
  NAND2_X1 U14267 ( .A1(n11275), .A2(n14637), .ZN(n11279) );
  OAI21_X1 U14268 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n11276), .A(
        n11279), .ZN(n11278) );
  INV_X1 U14269 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14771) );
  MUX2_X1 U14270 ( .A(n14771), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n16173), .Z(n11277) );
  OAI211_X1 U14271 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n11279), .A(
        n11278), .B(n11277), .ZN(n11280) );
  INV_X1 U14272 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12124) );
  XNOR2_X1 U14273 ( .A(n11280), .B(n12124), .ZN(n14766) );
  NAND2_X1 U14274 ( .A1(n20221), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14760) );
  OAI21_X1 U14275 ( .B1(n14693), .B2(n14241), .A(n14760), .ZN(n11281) );
  AOI21_X1 U14276 ( .B1(n14235), .B2(n16169), .A(n11281), .ZN(n11282) );
  INV_X1 U14277 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U14278 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11305), .ZN(
        n11304) );
  NAND2_X1 U14279 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n11316), .ZN(
        n11315) );
  NAND2_X1 U14280 ( .A1(n11318), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11301) );
  NAND2_X1 U14281 ( .A1(n11296), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11294) );
  INV_X1 U14282 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15482) );
  INV_X1 U14283 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12868) );
  INV_X1 U14284 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15469) );
  AND2_X1 U14285 ( .A1(n11291), .A2(n15469), .ZN(n11287) );
  NOR2_X1 U14286 ( .A1(n9932), .A2(n11287), .ZN(n15471) );
  INV_X1 U14287 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14280) );
  OAI22_X2 U14288 ( .A1(n14378), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19237), 
        .B2(n14280), .ZN(n11321) );
  INV_X1 U14289 ( .A(n11291), .ZN(n11292) );
  AOI21_X1 U14290 ( .B1(n12868), .B2(n11290), .A(n11292), .ZN(n14930) );
  AOI21_X1 U14291 ( .B1(n15482), .B2(n11294), .A(n11286), .ZN(n15485) );
  OR2_X1 U14292 ( .A1(n11296), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14293 ( .A1(n11294), .A2(n11293), .ZN(n15494) );
  INV_X1 U14294 ( .A(n15494), .ZN(n16293) );
  AND2_X1 U14295 ( .A1(n11297), .A2(n14270), .ZN(n11295) );
  NOR2_X1 U14296 ( .A1(n11296), .A2(n11295), .ZN(n14954) );
  NAND2_X1 U14297 ( .A1(n10143), .A2(n10142), .ZN(n11298) );
  AND2_X1 U14298 ( .A1(n11298), .A2(n11297), .ZN(n15507) );
  OAI21_X1 U14299 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11300), .A(
        n11323), .ZN(n16344) );
  AOI21_X1 U14300 ( .B1(n15538), .B2(n11299), .A(n11300), .ZN(n15536) );
  AOI21_X1 U14301 ( .B1(n19017), .B2(n11301), .A(n11320), .ZN(n19016) );
  AND2_X1 U14302 ( .A1(n11315), .A2(n15588), .ZN(n11302) );
  OR2_X1 U14303 ( .A1(n11302), .A2(n11318), .ZN(n19036) );
  INV_X1 U14304 ( .A(n19036), .ZN(n11317) );
  AOI21_X1 U14305 ( .B1(n16359), .B2(n11313), .A(n11316), .ZN(n19051) );
  AOI21_X1 U14306 ( .B1(n15598), .B2(n11312), .A(n11314), .ZN(n19058) );
  AOI21_X1 U14307 ( .B1(n16389), .B2(n11310), .A(n9906), .ZN(n19069) );
  AOI21_X1 U14308 ( .B1(n15610), .B2(n11308), .A(n11311), .ZN(n19090) );
  AOI21_X1 U14309 ( .B1(n14031), .B2(n11306), .A(n11309), .ZN(n19100) );
  AOI21_X1 U14310 ( .B1(n19127), .B2(n11304), .A(n11307), .ZN(n19133) );
  AOI21_X1 U14311 ( .B1(n13659), .B2(n11303), .A(n11305), .ZN(n13696) );
  INV_X1 U14312 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19153) );
  AOI22_X1 U14313 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13217), .B1(n19153), 
        .B2(n19237), .ZN(n19140) );
  INV_X1 U14314 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13218) );
  AOI22_X1 U14315 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13218), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19237), .ZN(n15050) );
  NOR2_X1 U14316 ( .A1(n19140), .A2(n15050), .ZN(n15049) );
  OAI21_X1 U14317 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11303), .ZN(n14245) );
  NAND2_X1 U14318 ( .A1(n15049), .A2(n14245), .ZN(n13694) );
  NOR2_X1 U14319 ( .A1(n13696), .A2(n13694), .ZN(n13810) );
  OAI21_X1 U14320 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11305), .A(
        n11304), .ZN(n13809) );
  NAND2_X1 U14321 ( .A1(n13810), .A2(n13809), .ZN(n19131) );
  NOR2_X1 U14322 ( .A1(n19133), .A2(n19131), .ZN(n19116) );
  OAI21_X1 U14323 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11307), .A(
        n11306), .ZN(n19118) );
  NAND2_X1 U14324 ( .A1(n19116), .A2(n19118), .ZN(n19099) );
  NOR2_X1 U14325 ( .A1(n19100), .A2(n19099), .ZN(n13825) );
  OAI21_X1 U14326 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11309), .A(
        n11308), .ZN(n16410) );
  NAND2_X1 U14327 ( .A1(n13825), .A2(n16410), .ZN(n19089) );
  NOR2_X1 U14328 ( .A1(n19090), .A2(n19089), .ZN(n19082) );
  OAI21_X1 U14329 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11311), .A(
        n11310), .ZN(n19083) );
  NAND2_X1 U14330 ( .A1(n19082), .A2(n19083), .ZN(n19068) );
  NOR2_X1 U14331 ( .A1(n19069), .A2(n19068), .ZN(n13799) );
  OAI21_X1 U14332 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9906), .A(
        n11312), .ZN(n16382) );
  NAND2_X1 U14333 ( .A1(n13799), .A2(n16382), .ZN(n19057) );
  NOR2_X1 U14334 ( .A1(n19058), .A2(n19057), .ZN(n13849) );
  OAI21_X1 U14335 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11314), .A(
        n11313), .ZN(n16371) );
  NAND2_X1 U14336 ( .A1(n13849), .A2(n16371), .ZN(n19050) );
  NOR2_X1 U14337 ( .A1(n19051), .A2(n19050), .ZN(n15036) );
  OAI21_X1 U14338 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11316), .A(
        n11315), .ZN(n16352) );
  NAND2_X1 U14339 ( .A1(n15036), .A2(n16352), .ZN(n19034) );
  NOR2_X1 U14340 ( .A1(n11317), .A2(n19034), .ZN(n15022) );
  OR2_X1 U14341 ( .A1(n11318), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11319) );
  NAND2_X1 U14342 ( .A1(n11301), .A2(n11319), .ZN(n15577) );
  NAND2_X1 U14343 ( .A1(n15022), .A2(n15577), .ZN(n19014) );
  NOR2_X1 U14344 ( .A1(n19016), .A2(n19014), .ZN(n15008) );
  OAI21_X1 U14345 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11320), .A(
        n11299), .ZN(n15552) );
  NAND2_X1 U14346 ( .A1(n15008), .A2(n15552), .ZN(n14992) );
  OAI21_X1 U14347 ( .B1(n15536), .B2(n14992), .A(n11321), .ZN(n14979) );
  AND2_X1 U14348 ( .A1(n16344), .A2(n14979), .ZN(n14982) );
  AOI21_X1 U14349 ( .B1(n11285), .B2(n11323), .A(n11322), .ZN(n16310) );
  NOR2_X1 U14350 ( .A1(n19117), .A2(n14965), .ZN(n14955) );
  NOR2_X1 U14351 ( .A1(n14954), .A2(n14955), .ZN(n14953) );
  NOR2_X1 U14352 ( .A1(n19117), .A2(n14953), .ZN(n16292) );
  NOR2_X1 U14353 ( .A1(n16293), .A2(n16292), .ZN(n16291) );
  NOR2_X1 U14354 ( .A1(n19117), .A2(n16291), .ZN(n14949) );
  NOR2_X1 U14355 ( .A1(n15485), .A2(n14949), .ZN(n14948) );
  NOR2_X1 U14356 ( .A1(n19117), .A2(n14948), .ZN(n14929) );
  NOR2_X1 U14357 ( .A1(n14930), .A2(n14929), .ZN(n14928) );
  NOR2_X1 U14358 ( .A1(n14920), .A2(n19117), .ZN(n11325) );
  XOR2_X1 U14359 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9932), .Z(n14357) );
  NOR2_X1 U14360 ( .A1(n11325), .A2(n14357), .ZN(n14284) );
  NOR4_X1 U14361 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n16540), .ZN(n11324) );
  NAND2_X1 U14362 ( .A1(n11327), .A2(n11326), .ZN(n12019) );
  AND2_X4 U14363 ( .A1(n11621), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11628) );
  INV_X1 U14364 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11328) );
  AND2_X2 U14365 ( .A1(n11328), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11619) );
  INV_X2 U14366 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15879) );
  AND2_X4 U14367 ( .A1(n11619), .A2(n15879), .ZN(n11636) );
  AOI22_X1 U14368 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14369 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11331) );
  AND2_X4 U14370 ( .A1(n11619), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11634) );
  AND2_X2 U14371 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11637) );
  AND2_X4 U14372 ( .A1(n11637), .A2(n15879), .ZN(n11644) );
  AND2_X4 U14373 ( .A1(n11621), .A2(n15879), .ZN(n11626) );
  AND2_X4 U14374 ( .A1(n11637), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11629) );
  AOI22_X1 U14375 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11329) );
  NAND4_X1 U14376 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11333) );
  NAND2_X1 U14377 ( .A1(n11333), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11340) );
  AOI22_X1 U14378 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14379 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14380 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14381 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U14382 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  NAND2_X1 U14383 ( .A1(n11338), .A2(n11408), .ZN(n11339) );
  AOI22_X1 U14384 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14385 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14386 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14387 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11341) );
  NAND4_X1 U14388 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11345) );
  NAND2_X1 U14389 ( .A1(n11345), .A2(n11408), .ZN(n11352) );
  AOI22_X1 U14390 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14391 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14392 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14393 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11346) );
  NAND4_X1 U14394 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(
        n11350) );
  NAND2_X1 U14395 ( .A1(n11350), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11351) );
  AOI22_X1 U14396 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14397 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14398 ( .A1(n11636), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11353) );
  NAND2_X1 U14399 ( .A1(n11357), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11364) );
  AOI22_X1 U14400 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14401 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14402 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14403 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14404 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14405 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11365) );
  NAND4_X1 U14406 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n11369) );
  NAND2_X1 U14407 ( .A1(n11369), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11376) );
  AOI22_X1 U14408 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14409 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14410 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11626), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14411 ( .A1(n11636), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11370) );
  NAND4_X1 U14412 ( .A1(n11373), .A2(n11372), .A3(n11371), .A4(n11370), .ZN(
        n11374) );
  NOR2_X1 U14413 ( .A1(n11458), .A2(n13630), .ZN(n11398) );
  AOI22_X1 U14414 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14415 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14416 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14417 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14418 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14419 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14420 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14421 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14422 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14423 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14424 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14425 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14426 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14427 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14428 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14429 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14430 ( .A1(n11450), .A2(n11398), .A3(n11998), .A4(n19337), .ZN(
        n11461) );
  INV_X1 U14431 ( .A(n11461), .ZN(n11412) );
  AOI22_X1 U14432 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14433 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14434 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14435 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U14436 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11403) );
  AOI22_X1 U14437 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14438 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14439 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11644), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14440 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11404) );
  NAND4_X1 U14441 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11409) );
  NAND2_X1 U14442 ( .A1(n11409), .A2(n11408), .ZN(n11410) );
  NAND2_X2 U14443 ( .A1(n11411), .A2(n11410), .ZN(n11432) );
  INV_X4 U14444 ( .A(n11432), .ZN(n20028) );
  NAND2_X1 U14445 ( .A1(n11412), .A2(n20028), .ZN(n11613) );
  AOI22_X1 U14446 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11636), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14447 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14448 ( .A1(n11628), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11413) );
  NAND4_X1 U14449 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11417) );
  NAND2_X1 U14450 ( .A1(n11417), .A2(n11408), .ZN(n11424) );
  AOI22_X1 U14451 ( .A1(n15308), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14452 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11629), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11419) );
  NAND4_X1 U14453 ( .A1(n11421), .A2(n11420), .A3(n11419), .A4(n11418), .ZN(
        n11422) );
  NAND2_X1 U14454 ( .A1(n11422), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11423) );
  NAND2_X2 U14455 ( .A1(n11424), .A2(n11423), .ZN(n11617) );
  INV_X1 U14457 ( .A(n12904), .ZN(n11426) );
  INV_X1 U14458 ( .A(n13630), .ZN(n11425) );
  NAND3_X1 U14460 ( .A1(n12947), .A2(n12883), .A3(n11450), .ZN(n11427) );
  INV_X1 U14461 ( .A(n11453), .ZN(n11428) );
  NAND2_X1 U14462 ( .A1(n11683), .A2(n13630), .ZN(n11459) );
  NAND3_X1 U14463 ( .A1(n11453), .A2(n11429), .A3(n20028), .ZN(n11430) );
  NAND2_X1 U14464 ( .A1(n11430), .A2(n11425), .ZN(n11431) );
  NAND2_X1 U14465 ( .A1(n11459), .A2(n11431), .ZN(n11434) );
  NAND2_X2 U14466 ( .A1(n11617), .A2(n11432), .ZN(n12929) );
  NAND2_X2 U14467 ( .A1(n12904), .A2(n12929), .ZN(n12939) );
  NAND2_X1 U14468 ( .A1(n12939), .A2(n11455), .ZN(n11433) );
  NOR2_X2 U14469 ( .A1(n11434), .A2(n11433), .ZN(n12971) );
  NAND2_X1 U14470 ( .A1(n12971), .A2(n12945), .ZN(n11487) );
  NAND2_X1 U14471 ( .A1(n11986), .A2(n15191), .ZN(n11436) );
  NAND3_X1 U14472 ( .A1(n11465), .A2(n11487), .A3(n11436), .ZN(n11437) );
  CLKBUF_X3 U14473 ( .A(n11501), .Z(n11591) );
  INV_X1 U14474 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14356) );
  NAND3_X2 U14475 ( .A1(n12948), .A2(n12911), .A3(n12945), .ZN(n15883) );
  AOI22_X1 U14476 ( .A1(n14276), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11441) );
  OAI21_X1 U14477 ( .B1(n11591), .B2(n14356), .A(n11441), .ZN(n11442) );
  AOI21_X1 U14478 ( .B1(n11593), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11442), .ZN(n11594) );
  INV_X1 U14479 ( .A(n11683), .ZN(n11663) );
  NAND2_X1 U14480 ( .A1(n11663), .A2(n19337), .ZN(n11444) );
  INV_X1 U14481 ( .A(n11443), .ZN(n11456) );
  NAND2_X1 U14482 ( .A1(n11444), .A2(n11456), .ZN(n12882) );
  NAND2_X1 U14483 ( .A1(n11683), .A2(n11445), .ZN(n12879) );
  NAND2_X1 U14484 ( .A1(n12879), .A2(n19355), .ZN(n11447) );
  INV_X1 U14485 ( .A(n12942), .ZN(n12948) );
  NAND2_X1 U14486 ( .A1(n11452), .A2(n12877), .ZN(n12972) );
  NAND2_X1 U14487 ( .A1(n11428), .A2(n19347), .ZN(n11454) );
  NAND2_X1 U14488 ( .A1(n11455), .A2(n11454), .ZN(n11457) );
  NAND2_X1 U14489 ( .A1(n11457), .A2(n11456), .ZN(n11460) );
  NAND3_X1 U14490 ( .A1(n11460), .A2(n11459), .A3(n11458), .ZN(n11462) );
  NAND3_X1 U14491 ( .A1(n11462), .A2(n11461), .A3(n20028), .ZN(n12951) );
  OAI211_X1 U14492 ( .C1(n12972), .C2(n12920), .A(n11463), .B(n12951), .ZN(
        n11464) );
  INV_X1 U14493 ( .A(n11464), .ZN(n11475) );
  NAND2_X1 U14494 ( .A1(n11514), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11467) );
  INV_X1 U14495 ( .A(n11986), .ZN(n11612) );
  AOI22_X1 U14496 ( .A1(n16495), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20018), .ZN(n11466) );
  INV_X1 U14497 ( .A(n11510), .ZN(n11468) );
  NAND2_X1 U14498 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11474) );
  INV_X1 U14499 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14500 ( .A1(n11497), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14501 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11469) );
  OAI211_X1 U14502 ( .C1(n11501), .C2(n11471), .A(n11470), .B(n11469), .ZN(
        n11472) );
  INV_X1 U14503 ( .A(n11472), .ZN(n11473) );
  AND2_X2 U14504 ( .A1(n11474), .A2(n11473), .ZN(n11493) );
  XNOR2_X2 U14505 ( .A(n11492), .B(n11493), .ZN(n12537) );
  INV_X1 U14506 ( .A(n11476), .ZN(n11478) );
  NAND2_X1 U14507 ( .A1(n11475), .A2(n11479), .ZN(n11480) );
  NAND2_X1 U14508 ( .A1(n11480), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11486) );
  NAND2_X1 U14509 ( .A1(n11497), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11483) );
  AND2_X1 U14510 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11481) );
  NOR2_X1 U14511 ( .A1(n20018), .A2(n11481), .ZN(n11482) );
  OAI211_X1 U14512 ( .C1(n11501), .C2(n19007), .A(n11483), .B(n11482), .ZN(
        n11484) );
  INV_X1 U14513 ( .A(n11484), .ZN(n11485) );
  OAI211_X1 U14514 ( .C1(n11510), .C2(n13217), .A(n11486), .B(n11485), .ZN(
        n12530) );
  NAND2_X1 U14515 ( .A1(n11514), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11491) );
  NAND2_X1 U14516 ( .A1(n20018), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11488) );
  OAI211_X1 U14517 ( .C1(n15884), .C2(n19237), .A(n11585), .B(n11488), .ZN(
        n11489) );
  INV_X1 U14518 ( .A(n11489), .ZN(n11490) );
  INV_X1 U14519 ( .A(n11492), .ZN(n11494) );
  NAND2_X1 U14520 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  OAI21_X1 U14521 ( .B1(n16505), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16540), 
        .ZN(n11496) );
  INV_X1 U14522 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14523 ( .A1(n11497), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11499) );
  NAND2_X1 U14524 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11498) );
  OAI211_X1 U14525 ( .C1(n11501), .C2(n11500), .A(n11499), .B(n11498), .ZN(
        n11502) );
  INV_X1 U14526 ( .A(n11502), .ZN(n11503) );
  INV_X1 U14527 ( .A(n11505), .ZN(n11507) );
  NAND2_X1 U14528 ( .A1(n11507), .A2(n11506), .ZN(n11508) );
  INV_X1 U14529 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11513) );
  OR2_X1 U14530 ( .A1(n11510), .A2(n16479), .ZN(n11512) );
  AOI22_X1 U14531 ( .A1(n11497), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11511) );
  OAI211_X1 U14532 ( .C1(n11591), .C2(n11513), .A(n11512), .B(n11511), .ZN(
        n11516) );
  INV_X1 U14533 ( .A(n11514), .ZN(n11515) );
  INV_X1 U14534 ( .A(n20018), .ZN(n16543) );
  OAI22_X1 U14535 ( .A1(n11515), .A2(n11408), .B1(n16543), .B2(n19980), .ZN(
        n11517) );
  NAND2_X1 U14536 ( .A1(n11517), .A2(n11516), .ZN(n11518) );
  INV_X1 U14537 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U14538 ( .A1(n14276), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11521) );
  INV_X1 U14539 ( .A(n11591), .ZN(n14277) );
  NAND2_X1 U14540 ( .A1(n14277), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11520) );
  OAI211_X1 U14541 ( .C1(n14281), .C2(n13996), .A(n11521), .B(n11520), .ZN(
        n13410) );
  INV_X1 U14542 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13997) );
  OR2_X1 U14543 ( .A1(n14281), .A2(n13997), .ZN(n11526) );
  INV_X1 U14544 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U14545 ( .A1(n14276), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U14546 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11522) );
  OAI211_X1 U14547 ( .C1(n11591), .C2(n11753), .A(n11523), .B(n11522), .ZN(
        n11524) );
  INV_X1 U14548 ( .A(n11524), .ZN(n11525) );
  INV_X1 U14549 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13966) );
  OR2_X1 U14550 ( .A1(n14281), .A2(n13966), .ZN(n11532) );
  INV_X1 U14551 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U14552 ( .A1(n14276), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14553 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11527) );
  OAI211_X1 U14554 ( .C1(n11591), .C2(n11529), .A(n11528), .B(n11527), .ZN(
        n11530) );
  INV_X1 U14555 ( .A(n11530), .ZN(n11531) );
  NAND2_X1 U14556 ( .A1(n11532), .A2(n11531), .ZN(n13427) );
  INV_X1 U14557 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n11535) );
  INV_X1 U14558 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14036) );
  OR2_X1 U14559 ( .A1(n14281), .A2(n14036), .ZN(n11534) );
  AOI22_X1 U14560 ( .A1(n14276), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11533) );
  OAI211_X1 U14561 ( .C1(n11591), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        n13466) );
  INV_X1 U14562 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13838) );
  INV_X1 U14563 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21138) );
  OR2_X1 U14564 ( .A1(n14281), .A2(n21138), .ZN(n11537) );
  AOI22_X1 U14565 ( .A1(n14276), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11536) );
  OAI211_X1 U14566 ( .C1(n11591), .C2(n13838), .A(n11537), .B(n11536), .ZN(
        n13433) );
  INV_X1 U14567 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15608) );
  INV_X1 U14568 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21159) );
  OR2_X1 U14569 ( .A1(n14281), .A2(n21159), .ZN(n11539) );
  AOI22_X1 U14570 ( .A1(n14276), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11538) );
  OAI211_X1 U14571 ( .C1(n11591), .C2(n15608), .A(n11539), .B(n11538), .ZN(
        n13552) );
  INV_X1 U14572 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11845) );
  INV_X1 U14573 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12718) );
  OR2_X1 U14574 ( .A1(n14281), .A2(n12718), .ZN(n11541) );
  AOI22_X1 U14575 ( .A1(n14276), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11540) );
  OAI211_X1 U14576 ( .C1(n11591), .C2(n11845), .A(n11541), .B(n11540), .ZN(
        n13565) );
  INV_X1 U14577 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11862) );
  INV_X1 U14578 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15818) );
  OR2_X1 U14579 ( .A1(n14281), .A2(n15818), .ZN(n11543) );
  AOI22_X1 U14580 ( .A1(n14276), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11542) );
  OAI211_X1 U14581 ( .C1(n11591), .C2(n11862), .A(n11543), .B(n11542), .ZN(
        n13616) );
  INV_X1 U14582 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11883) );
  INV_X1 U14583 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12734) );
  OR2_X1 U14584 ( .A1(n14281), .A2(n12734), .ZN(n11545) );
  AOI22_X1 U14585 ( .A1(n14276), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11544) );
  OAI211_X1 U14586 ( .C1(n11591), .C2(n11883), .A(n11545), .B(n11544), .ZN(
        n13584) );
  INV_X1 U14587 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11903) );
  INV_X1 U14588 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15803) );
  OR2_X1 U14589 ( .A1(n14281), .A2(n15803), .ZN(n11547) );
  AOI22_X1 U14590 ( .A1(n14276), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11546) );
  OAI211_X1 U14591 ( .C1(n11591), .C2(n11903), .A(n11547), .B(n11546), .ZN(
        n13645) );
  INV_X1 U14592 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11930) );
  INV_X1 U14593 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12774) );
  OR2_X1 U14594 ( .A1(n14281), .A2(n12774), .ZN(n11549) );
  AOI22_X1 U14595 ( .A1(n14276), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11548) );
  OAI211_X1 U14596 ( .C1(n11591), .C2(n11930), .A(n11549), .B(n11548), .ZN(
        n13636) );
  INV_X1 U14597 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15788) );
  OR2_X1 U14598 ( .A1(n14281), .A2(n15788), .ZN(n11554) );
  INV_X1 U14599 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U14600 ( .A1(n14276), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14601 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11550) );
  OAI211_X1 U14602 ( .C1(n11591), .C2(n11956), .A(n11551), .B(n11550), .ZN(
        n11552) );
  INV_X1 U14603 ( .A(n11552), .ZN(n11553) );
  NAND2_X1 U14604 ( .A1(n11554), .A2(n11553), .ZN(n13727) );
  INV_X1 U14605 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15769) );
  INV_X1 U14606 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15573) );
  OR2_X1 U14607 ( .A1(n14281), .A2(n15573), .ZN(n11556) );
  AOI22_X1 U14608 ( .A1(n14276), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11555) );
  OAI211_X1 U14609 ( .C1(n11591), .C2(n15769), .A(n11556), .B(n11555), .ZN(
        n13741) );
  INV_X1 U14610 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19925) );
  NAND2_X1 U14611 ( .A1(n14276), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14612 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11557) );
  OAI211_X1 U14613 ( .C1(n11591), .C2(n19925), .A(n11558), .B(n11557), .ZN(
        n11559) );
  AOI21_X1 U14614 ( .B1(n11593), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11559), .ZN(n13875) );
  INV_X1 U14615 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15576) );
  INV_X1 U14616 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15740) );
  OR2_X1 U14617 ( .A1(n14281), .A2(n15740), .ZN(n11561) );
  AOI22_X1 U14618 ( .A1(n14276), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11560) );
  OAI211_X1 U14619 ( .C1(n11591), .C2(n15576), .A(n11561), .B(n11560), .ZN(
        n13943) );
  INV_X1 U14620 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19928) );
  NAND2_X1 U14621 ( .A1(n14276), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14622 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14623 ( .C1(n11591), .C2(n19928), .A(n11563), .B(n11562), .ZN(
        n11564) );
  AOI21_X1 U14624 ( .B1(n11593), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11564), .ZN(n14019) );
  INV_X1 U14625 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19930) );
  NAND2_X1 U14626 ( .A1(n14276), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14627 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11565) );
  OAI211_X1 U14628 ( .C1(n11591), .C2(n19930), .A(n11566), .B(n11565), .ZN(
        n11567) );
  AOI21_X1 U14629 ( .B1(n11593), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11567), .ZN(n15015) );
  INV_X1 U14630 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19932) );
  NAND2_X1 U14631 ( .A1(n14276), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14632 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11568) );
  OAI211_X1 U14633 ( .C1(n11591), .C2(n19932), .A(n11569), .B(n11568), .ZN(
        n11570) );
  AOI21_X1 U14634 ( .B1(n11593), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11570), .ZN(n14996) );
  INV_X1 U14635 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n11966) );
  INV_X1 U14636 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15689) );
  OR2_X1 U14637 ( .A1(n14281), .A2(n15689), .ZN(n11572) );
  AOI22_X1 U14638 ( .A1(n14276), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11571) );
  OAI211_X1 U14639 ( .C1(n11591), .C2(n11966), .A(n11572), .B(n11571), .ZN(
        n14984) );
  INV_X1 U14640 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15669) );
  OR2_X1 U14641 ( .A1(n14281), .A2(n15669), .ZN(n11575) );
  AOI22_X1 U14642 ( .A1(n14276), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11574) );
  NAND2_X1 U14643 ( .A1(n14277), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11573) );
  INV_X1 U14644 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19937) );
  NAND2_X1 U14645 ( .A1(n14276), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U14646 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11576) );
  OAI211_X1 U14647 ( .C1(n11591), .C2(n19937), .A(n11577), .B(n11576), .ZN(
        n11578) );
  AOI21_X1 U14648 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n11593), .A(
        n11578), .ZN(n14968) );
  INV_X1 U14649 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19939) );
  INV_X1 U14650 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14262) );
  OR2_X1 U14651 ( .A1(n14281), .A2(n14262), .ZN(n11580) );
  AOI22_X1 U14652 ( .A1(n14276), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11579) );
  OAI211_X1 U14653 ( .C1(n11591), .C2(n19939), .A(n11580), .B(n11579), .ZN(
        n14257) );
  INV_X1 U14654 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19941) );
  INV_X1 U14655 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15646) );
  OR2_X1 U14656 ( .A1(n14281), .A2(n15646), .ZN(n11582) );
  AOI22_X1 U14657 ( .A1(n14276), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11581) );
  OAI211_X1 U14658 ( .C1(n11591), .C2(n19941), .A(n11582), .B(n11581), .ZN(
        n15351) );
  INV_X1 U14659 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n14943) );
  INV_X1 U14660 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15481) );
  OR2_X1 U14661 ( .A1(n14281), .A2(n15481), .ZN(n11584) );
  AOI22_X1 U14662 ( .A1(n14277), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11583) );
  OAI211_X1 U14663 ( .C1(n14943), .C2(n11585), .A(n11584), .B(n11583), .ZN(
        n14938) );
  INV_X1 U14664 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n11588) );
  INV_X1 U14665 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12967) );
  OR2_X1 U14666 ( .A1(n14281), .A2(n12967), .ZN(n11587) );
  AOI22_X1 U14667 ( .A1(n14276), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11586) );
  OAI211_X1 U14668 ( .C1(n11591), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        n12869) );
  INV_X1 U14669 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19945) );
  NAND2_X1 U14670 ( .A1(n14276), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11590) );
  NAND2_X1 U14671 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11589) );
  OAI211_X1 U14672 ( .C1(n11591), .C2(n19945), .A(n11590), .B(n11589), .ZN(
        n11592) );
  AOI21_X1 U14673 ( .B1(n11593), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11592), .ZN(n14911) );
  AOI21_X1 U14674 ( .B1(n11594), .B2(n14914), .A(n14283), .ZN(n15329) );
  INV_X1 U14675 ( .A(n15329), .ZN(n14397) );
  NAND2_X1 U14676 ( .A1(n12896), .A2(n11595), .ZN(n11597) );
  NAND2_X1 U14677 ( .A1(n19996), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11596) );
  NAND2_X1 U14678 ( .A1(n11597), .A2(n11596), .ZN(n11609) );
  MUX2_X1 U14679 ( .A(n16505), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11608) );
  NAND2_X1 U14680 ( .A1(n11609), .A2(n11608), .ZN(n11607) );
  NAND2_X1 U14681 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n16505), .ZN(
        n11598) );
  NAND2_X1 U14682 ( .A1(n11607), .A2(n11598), .ZN(n11601) );
  XNOR2_X1 U14683 ( .A(n12896), .B(n12654), .ZN(n12899) );
  INV_X1 U14684 ( .A(n11600), .ZN(n11606) );
  INV_X1 U14685 ( .A(n11601), .ZN(n11604) );
  INV_X1 U14686 ( .A(n11602), .ZN(n11603) );
  NAND2_X1 U14687 ( .A1(n11604), .A2(n11603), .ZN(n11605) );
  NAND2_X1 U14688 ( .A1(n11606), .A2(n11605), .ZN(n12003) );
  OAI21_X1 U14689 ( .B1(n11609), .B2(n11608), .A(n11607), .ZN(n12903) );
  NOR3_X1 U14690 ( .A1(n12003), .A2(n12903), .A3(n12912), .ZN(n12813) );
  AND2_X1 U14691 ( .A1(n12899), .A2(n12813), .ZN(n11611) );
  NAND2_X1 U14692 ( .A1(n16540), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19891) );
  NAND2_X1 U14693 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20026) );
  INV_X1 U14694 ( .A(n20026), .ZN(n20023) );
  OR2_X1 U14695 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20023), .ZN(n12014) );
  NOR2_X1 U14696 ( .A1(n12929), .A2(n12014), .ZN(n11614) );
  INV_X1 U14697 ( .A(n11618), .ZN(n11616) );
  INV_X1 U14698 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11650) );
  NOR2_X1 U14699 ( .A1(n19355), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11670) );
  INV_X2 U14700 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U14701 ( .A1(n14285), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11649) );
  NAND2_X1 U14702 ( .A1(n11998), .A2(n11618), .ZN(n11953) );
  NAND2_X1 U14703 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11625) );
  NAND2_X1 U14704 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11624) );
  INV_X1 U14705 ( .A(n12815), .ZN(n11622) );
  NOR2_X1 U14706 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12815), .ZN(
        n11687) );
  AOI22_X1 U14707 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n15144), .ZN(n11623) );
  AND3_X1 U14708 ( .A1(n11625), .A2(n11624), .A3(n11623), .ZN(n11633) );
  INV_X1 U14709 ( .A(n15121), .ZN(n11627) );
  NAND2_X1 U14710 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11632) );
  AND2_X2 U14711 ( .A1(n11643), .A2(n11408), .ZN(n15150) );
  NAND2_X1 U14712 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11631) );
  AND2_X4 U14713 ( .A1(n15128), .A2(n11408), .ZN(n15151) );
  NAND2_X1 U14714 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11630) );
  INV_X1 U14715 ( .A(n11634), .ZN(n15119) );
  INV_X1 U14716 ( .A(n15119), .ZN(n11635) );
  AND2_X4 U14717 ( .A1(n11635), .A2(n11408), .ZN(n15156) );
  AND2_X2 U14718 ( .A1(n15320), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15109) );
  AOI22_X1 U14719 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n15156), .B1(
        n15109), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14720 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11642) );
  AND2_X4 U14721 ( .A1(n15318), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15159) );
  NAND2_X1 U14722 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U14723 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11640) );
  AND2_X4 U14724 ( .A1(n15318), .A2(n11408), .ZN(n15160) );
  NAND2_X1 U14725 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11639) );
  AND4_X1 U14726 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11646) );
  AND2_X2 U14727 ( .A1(n15319), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15110) );
  AOI22_X1 U14728 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11645) );
  INV_X1 U14729 ( .A(n12612), .ZN(n12830) );
  OR2_X1 U14730 ( .A1(n11953), .A2(n12830), .ZN(n11648) );
  OAI211_X1 U14731 ( .C1(n11978), .C2(n11650), .A(n11649), .B(n11648), .ZN(
        n11651) );
  INV_X1 U14732 ( .A(n11651), .ZN(n13814) );
  AOI22_X1 U14733 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14734 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11916), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14735 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15145), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14736 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15150), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11652) );
  NAND4_X1 U14737 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(
        n11661) );
  AOI22_X1 U14738 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15064), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14739 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14740 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15159), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14741 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11687), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14742 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11660) );
  NOR2_X1 U14743 ( .A1(n11661), .A2(n11660), .ZN(n12832) );
  INV_X1 U14744 ( .A(n11953), .ZN(n11662) );
  NAND2_X1 U14745 ( .A1(n13301), .A2(n11664), .ZN(n11707) );
  OAI22_X1 U14746 ( .A1(n19355), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n20006), 
        .B2(n19825), .ZN(n11665) );
  INV_X1 U14747 ( .A(n11665), .ZN(n11666) );
  AND2_X1 U14748 ( .A1(n11707), .A2(n11666), .ZN(n11667) );
  AOI21_X1 U14749 ( .B1(n15910), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11669) );
  NAND2_X1 U14750 ( .A1(n13303), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14751 ( .A1(n11670), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11671) );
  OAI21_X1 U14752 ( .B1(n11978), .B2(n11471), .A(n11671), .ZN(n11686) );
  INV_X1 U14753 ( .A(n11686), .ZN(n11672) );
  AOI22_X1 U14754 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15150), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14755 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15145), .ZN(n11675) );
  AOI22_X1 U14756 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11687), .ZN(n11674) );
  AOI22_X1 U14757 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14758 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11682) );
  AOI22_X1 U14759 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n15143), .B1(
        n15064), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14760 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14761 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n15160), .B1(
        n11916), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14762 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15159), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14763 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  NOR2_X1 U14764 ( .A1(n11682), .A2(n11681), .ZN(n12831) );
  OR2_X1 U14765 ( .A1(n12831), .A2(n11953), .ZN(n11685) );
  NAND2_X1 U14766 ( .A1(n11683), .A2(n19355), .ZN(n12886) );
  MUX2_X1 U14767 ( .A(n19996), .B(n12886), .S(n19825), .Z(n11684) );
  AND2_X1 U14768 ( .A1(n11685), .A2(n11684), .ZN(n13223) );
  NAND2_X1 U14769 ( .A1(n13224), .A2(n13223), .ZN(n13222) );
  OR2_X1 U14770 ( .A1(n13300), .A2(n11686), .ZN(n11709) );
  NAND2_X1 U14771 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11690) );
  NAND2_X1 U14772 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11689) );
  AOI22_X1 U14773 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n11687), .ZN(n11688) );
  AND3_X1 U14774 ( .A1(n11690), .A2(n11689), .A3(n11688), .ZN(n11694) );
  NAND2_X1 U14775 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11693) );
  NAND2_X1 U14776 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11692) );
  NAND2_X1 U14777 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11691) );
  AOI22_X1 U14778 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11698) );
  NAND2_X1 U14779 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11697) );
  NAND2_X1 U14780 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11696) );
  NAND2_X1 U14781 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11695) );
  NAND2_X1 U14782 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11702) );
  NAND2_X1 U14783 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14784 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11700) );
  NAND2_X1 U14785 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11699) );
  OR2_X1 U14786 ( .A1(n11953), .A2(n12837), .ZN(n11706) );
  OAI211_X1 U14787 ( .C1(n19825), .C2(n16505), .A(n11707), .B(n11706), .ZN(
        n11708) );
  AND3_X1 U14788 ( .A1(n13222), .A2(n11709), .A3(n11708), .ZN(n11710) );
  AOI22_X1 U14789 ( .A1(n14285), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11711) );
  OAI21_X1 U14790 ( .B1(n11978), .B2(n11500), .A(n11711), .ZN(n13250) );
  NOR2_X1 U14791 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  NAND2_X1 U14792 ( .A1(n14286), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14793 ( .A1(n11664), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11731) );
  NAND2_X1 U14794 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11716) );
  NAND2_X1 U14795 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U14796 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U14797 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11713) );
  AND4_X1 U14798 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11727) );
  AOI22_X1 U14799 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n15143), .B1(
        n15064), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U14800 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U14801 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U14802 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11717) );
  AND4_X1 U14803 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11726) );
  AOI22_X1 U14804 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15151), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11725) );
  INV_X1 U14805 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15223) );
  NAND2_X1 U14806 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11722) );
  AOI22_X1 U14807 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n15144), .ZN(n11721) );
  OAI211_X1 U14808 ( .C1(n11799), .C2(n15223), .A(n11722), .B(n11721), .ZN(
        n11723) );
  AOI21_X1 U14809 ( .B1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n15150), .A(
        n11723), .ZN(n11724) );
  NAND4_X1 U14810 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n12609) );
  INV_X1 U14811 ( .A(n12609), .ZN(n11728) );
  OR2_X1 U14812 ( .A1(n11953), .A2(n11728), .ZN(n11730) );
  NAND2_X1 U14813 ( .A1(n14285), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14814 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n13700) );
  NAND2_X1 U14815 ( .A1(n13699), .A2(n13700), .ZN(n13698) );
  AOI22_X1 U14816 ( .A1(n14285), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14817 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14818 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11738) );
  NAND2_X1 U14819 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11737) );
  INV_X1 U14820 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U14821 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11734) );
  AOI22_X1 U14822 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .B2(n15144), .ZN(n11733) );
  OAI211_X1 U14823 ( .C1(n11799), .C2(n15269), .A(n11734), .B(n11733), .ZN(
        n11735) );
  INV_X1 U14824 ( .A(n11735), .ZN(n11736) );
  NAND2_X1 U14825 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14826 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14827 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14828 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11740) );
  AOI22_X1 U14829 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n15143), .B1(
        n15064), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14830 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14831 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14832 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11744) );
  OR2_X1 U14833 ( .A1(n11953), .A2(n12643), .ZN(n11751) );
  OAI211_X1 U14834 ( .C1(n11978), .C2(n11753), .A(n11752), .B(n11751), .ZN(
        n13995) );
  NAND2_X1 U14835 ( .A1(n13994), .A2(n13995), .ZN(n11769) );
  NAND2_X1 U14836 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11756) );
  NAND2_X1 U14837 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11755) );
  AOI22_X1 U14838 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n15144), .ZN(n11754) );
  AND3_X1 U14839 ( .A1(n11756), .A2(n11755), .A3(n11754), .ZN(n11760) );
  NAND2_X1 U14840 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U14841 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U14842 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11757) );
  AOI22_X1 U14843 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n15101), .B1(
        n15156), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14844 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U14845 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14846 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11762) );
  NAND2_X1 U14847 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11761) );
  AOI22_X1 U14848 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11765) );
  NAND4_X1 U14849 ( .A1(n10308), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n12006) );
  INV_X1 U14850 ( .A(n12006), .ZN(n12694) );
  OR2_X1 U14851 ( .A1(n11953), .A2(n12694), .ZN(n11768) );
  AOI22_X1 U14852 ( .A1(n14285), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11770) );
  OAI21_X1 U14853 ( .B1(n11978), .B2(n11529), .A(n11770), .ZN(n13958) );
  NAND2_X1 U14854 ( .A1(n13959), .A2(n13958), .ZN(n11787) );
  NAND2_X1 U14855 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U14856 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11772) );
  INV_X1 U14857 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19363) );
  AOI22_X1 U14858 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n15144), .ZN(n11771) );
  AND3_X1 U14859 ( .A1(n11773), .A2(n11772), .A3(n11771), .ZN(n11777) );
  NAND2_X1 U14860 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U14861 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11775) );
  NAND2_X1 U14862 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11774) );
  AOI22_X1 U14863 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n15156), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14864 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U14865 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U14866 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14867 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11778) );
  AOI22_X1 U14868 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11782) );
  OR2_X1 U14869 ( .A1(n11953), .A2(n14364), .ZN(n11786) );
  AOI22_X1 U14870 ( .A1(n14285), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11788) );
  OAI21_X1 U14871 ( .B1(n11978), .B2(n11535), .A(n11788), .ZN(n14038) );
  AOI22_X1 U14872 ( .A1(n14285), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11664), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11807) );
  NAND2_X1 U14873 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U14874 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U14875 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U14876 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11789) );
  AND4_X1 U14877 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11804) );
  AOI22_X1 U14878 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15064), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U14879 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U14880 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U14881 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11793) );
  AND4_X1 U14882 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11803) );
  AOI22_X1 U14883 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15151), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11802) );
  INV_X1 U14884 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19526) );
  NAND2_X1 U14885 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11798) );
  AOI22_X1 U14886 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15144), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11797) );
  OAI211_X1 U14887 ( .C1(n19526), .C2(n11799), .A(n11798), .B(n11797), .ZN(
        n11800) );
  AOI21_X1 U14888 ( .B1(n15150), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11800), .ZN(n11801) );
  NAND4_X1 U14889 ( .A1(n11804), .A2(n11803), .A3(n11802), .A4(n11801), .ZN(
        n13440) );
  INV_X1 U14890 ( .A(n13440), .ZN(n11805) );
  OR2_X1 U14891 ( .A1(n11953), .A2(n11805), .ZN(n11806) );
  OAI211_X1 U14892 ( .C1(n11978), .C2(n13838), .A(n11807), .B(n11806), .ZN(
        n11808) );
  INV_X1 U14893 ( .A(n11808), .ZN(n13830) );
  OAI22_X1 U14894 ( .A1(n11978), .A2(n15608), .B1(n11809), .B2(n21159), .ZN(
        n11810) );
  INV_X1 U14895 ( .A(n11810), .ZN(n11827) );
  INV_X1 U14896 ( .A(n15143), .ZN(n13745) );
  INV_X1 U14897 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U14898 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11812) );
  AOI22_X1 U14899 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15144), .ZN(n11811) );
  OAI211_X1 U14900 ( .C1(n13745), .C2(n15174), .A(n11812), .B(n11811), .ZN(
        n11813) );
  INV_X1 U14901 ( .A(n11813), .ZN(n11817) );
  NAND2_X1 U14902 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14903 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U14904 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11814) );
  AND4_X1 U14905 ( .A1(n11817), .A2(n11816), .A3(n11815), .A4(n11814), .ZN(
        n11825) );
  AOI22_X1 U14906 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n15156), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14907 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U14908 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U14909 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U14910 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11818) );
  AND4_X1 U14911 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11823) );
  AOI22_X1 U14912 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11822) );
  NAND4_X1 U14913 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n13559) );
  AOI22_X1 U14914 ( .A1(n11662), .A2(n13559), .B1(n14285), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n11826) );
  NAND2_X1 U14915 ( .A1(n11827), .A2(n11826), .ZN(n15852) );
  AOI22_X1 U14916 ( .A1(n14285), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11844) );
  INV_X1 U14917 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15204) );
  NAND2_X1 U14918 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11829) );
  AOI22_X1 U14919 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n15144), .ZN(n11828) );
  OAI211_X1 U14920 ( .C1(n13745), .C2(n15204), .A(n11829), .B(n11828), .ZN(
        n11830) );
  INV_X1 U14921 ( .A(n11830), .ZN(n11834) );
  NAND2_X1 U14922 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11833) );
  NAND2_X1 U14923 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11832) );
  NAND2_X1 U14924 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11831) );
  AND4_X1 U14925 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11842) );
  AOI22_X1 U14926 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U14927 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11837) );
  NAND2_X1 U14928 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U14929 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11835) );
  AND4_X1 U14930 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11841) );
  AOI22_X1 U14931 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n15109), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14932 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n15110), .B1(
        n15151), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11839) );
  NAND4_X1 U14933 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n13560) );
  INV_X1 U14934 ( .A(n13560), .ZN(n13556) );
  OR2_X1 U14935 ( .A1(n11953), .A2(n13556), .ZN(n11843) );
  OAI211_X1 U14936 ( .C1(n11978), .C2(n11845), .A(n11844), .B(n11843), .ZN(
        n11846) );
  INV_X1 U14937 ( .A(n11846), .ZN(n15836) );
  NAND2_X1 U14938 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11848) );
  AOI22_X1 U14939 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n15144), .ZN(n11847) );
  OAI211_X1 U14940 ( .C1(n13745), .C2(n15223), .A(n11848), .B(n11847), .ZN(
        n11849) );
  INV_X1 U14941 ( .A(n11849), .ZN(n11853) );
  NAND2_X1 U14942 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11852) );
  NAND2_X1 U14943 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11851) );
  NAND2_X1 U14944 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11850) );
  AND4_X1 U14945 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n11861) );
  AOI22_X1 U14946 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n15156), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14947 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n15157), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U14948 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U14949 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U14950 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11854) );
  AND4_X1 U14951 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11859) );
  AOI22_X1 U14952 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11858) );
  NAND4_X1 U14953 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n13586) );
  INV_X1 U14954 ( .A(n13586), .ZN(n13614) );
  OAI22_X1 U14955 ( .A1(n11978), .A2(n11862), .B1(n11953), .B2(n13614), .ZN(
        n11863) );
  INV_X1 U14956 ( .A(n11863), .ZN(n11865) );
  AOI22_X1 U14957 ( .A1(n14285), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U14958 ( .A1(n11865), .A2(n11864), .ZN(n15821) );
  NAND2_X1 U14959 ( .A1(n15822), .A2(n15821), .ZN(n13797) );
  AOI22_X1 U14960 ( .A1(n14285), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11882) );
  INV_X1 U14961 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U14962 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11867) );
  AOI22_X1 U14963 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n15144), .ZN(n11866) );
  OAI211_X1 U14964 ( .C1(n13745), .C2(n15245), .A(n11867), .B(n11866), .ZN(
        n11868) );
  INV_X1 U14965 ( .A(n11868), .ZN(n11872) );
  NAND2_X1 U14966 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11871) );
  NAND2_X1 U14967 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U14968 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11869) );
  AND4_X1 U14969 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11880) );
  AOI22_X1 U14970 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U14971 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11875) );
  NAND2_X1 U14972 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11874) );
  NAND2_X1 U14973 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11873) );
  AND4_X1 U14974 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11879) );
  AOI22_X1 U14975 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n15156), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14976 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n15151), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U14977 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n13587) );
  INV_X1 U14978 ( .A(n13587), .ZN(n13592) );
  OR2_X1 U14979 ( .A1(n11953), .A2(n13592), .ZN(n11881) );
  OAI211_X1 U14980 ( .C1(n11978), .C2(n11883), .A(n11882), .B(n11881), .ZN(
        n11884) );
  INV_X1 U14981 ( .A(n11884), .ZN(n13798) );
  AOI22_X1 U14982 ( .A1(n14285), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U14983 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11886) );
  AOI22_X1 U14984 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n15144), .ZN(n11885) );
  OAI211_X1 U14985 ( .C1(n13745), .C2(n15269), .A(n11886), .B(n11885), .ZN(
        n11887) );
  INV_X1 U14986 ( .A(n11887), .ZN(n11891) );
  NAND2_X1 U14987 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U14988 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U14989 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11888) );
  AND4_X1 U14990 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11899) );
  AOI22_X1 U14991 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n15156), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U14992 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n15157), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U14993 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U14994 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U14995 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11892) );
  AND4_X1 U14996 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11897) );
  AOI22_X1 U14997 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U14998 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n13644) );
  INV_X1 U14999 ( .A(n13644), .ZN(n11900) );
  OR2_X1 U15000 ( .A1(n11953), .A2(n11900), .ZN(n11901) );
  OAI211_X1 U15001 ( .C1(n11978), .C2(n11903), .A(n11902), .B(n11901), .ZN(
        n15801) );
  AOI22_X1 U15002 ( .A1(n14285), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11929) );
  NAND2_X1 U15003 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U15004 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11906) );
  NAND2_X1 U15005 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15006 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11904) );
  AND4_X1 U15007 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11927) );
  NAND2_X1 U15008 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11915) );
  NAND2_X1 U15009 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11914) );
  INV_X1 U15010 ( .A(n15157), .ZN(n11910) );
  INV_X1 U15011 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12689) );
  NAND2_X1 U15012 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11909) );
  AOI22_X1 U15013 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n15144), .ZN(n11908) );
  OAI211_X1 U15014 ( .C1(n11910), .C2(n12689), .A(n11909), .B(n11908), .ZN(
        n11911) );
  INV_X1 U15015 ( .A(n11911), .ZN(n11913) );
  NAND2_X1 U15016 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11912) );
  AND4_X1 U15017 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11926) );
  INV_X1 U15018 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15111) );
  INV_X1 U15019 ( .A(n15159), .ZN(n11918) );
  INV_X1 U15020 ( .A(n11916), .ZN(n11917) );
  INV_X1 U15021 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15100) );
  OAI22_X1 U15022 ( .A1(n15111), .A2(n11918), .B1(n11917), .B2(n15100), .ZN(
        n11924) );
  INV_X1 U15023 ( .A(n15160), .ZN(n11922) );
  INV_X1 U15024 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11921) );
  NAND2_X1 U15025 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15026 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11919) );
  OAI211_X1 U15027 ( .C1(n11922), .C2(n11921), .A(n11920), .B(n11919), .ZN(
        n11923) );
  NOR2_X1 U15028 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  OR2_X1 U15029 ( .A1(n11953), .A2(n13639), .ZN(n11928) );
  OAI211_X1 U15030 ( .C1(n11978), .C2(n11930), .A(n11929), .B(n11928), .ZN(
        n11931) );
  INV_X1 U15031 ( .A(n11931), .ZN(n13853) );
  AOI22_X1 U15032 ( .A1(n14285), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U15033 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15034 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U15035 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U15036 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11932) );
  NAND4_X1 U15037 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11941) );
  AOI22_X1 U15038 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n15157), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U15039 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15040 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15041 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11936) );
  NAND4_X1 U15042 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11940) );
  NOR2_X1 U15043 ( .A1(n11941), .A2(n11940), .ZN(n11952) );
  INV_X1 U15044 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11944) );
  INV_X1 U15045 ( .A(n15150), .ZN(n13912) );
  INV_X1 U15046 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11943) );
  OAI22_X1 U15047 ( .A1(n13913), .A2(n11944), .B1(n13912), .B2(n11943), .ZN(
        n11950) );
  NAND2_X1 U15048 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11948) );
  AOI22_X1 U15049 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n15144), .ZN(n11947) );
  NAND2_X1 U15050 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11946) );
  NAND2_X1 U15051 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11945) );
  NAND4_X1 U15052 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11949) );
  NOR2_X1 U15053 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  OR2_X1 U15054 ( .A1(n11953), .A2(n13731), .ZN(n11954) );
  OAI211_X1 U15055 ( .C1(n11978), .C2(n11956), .A(n11955), .B(n11954), .ZN(
        n15784) );
  AOI22_X1 U15056 ( .A1(n14285), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11957) );
  OAI21_X1 U15057 ( .B1(n11978), .B2(n15769), .A(n11957), .ZN(n15038) );
  AOI22_X1 U15058 ( .A1(n14285), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11958) );
  OAI21_X1 U15059 ( .B1(n11978), .B2(n19925), .A(n11958), .ZN(n13787) );
  NAND2_X1 U15060 ( .A1(n14286), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U15061 ( .A1(n14285), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11959) );
  AND2_X1 U15062 ( .A1(n11960), .A2(n11959), .ZN(n15026) );
  NAND2_X1 U15063 ( .A1(n14286), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15064 ( .A1(n14285), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15065 ( .A1(n14285), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11963) );
  OAI21_X1 U15066 ( .B1(n11978), .B2(n19930), .A(n11963), .ZN(n15016) );
  AOI22_X1 U15067 ( .A1(n14285), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11964) );
  OAI21_X1 U15068 ( .B1(n11978), .B2(n19932), .A(n11964), .ZN(n15000) );
  AOI22_X1 U15069 ( .A1(n14285), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11965) );
  OAI21_X1 U15070 ( .B1(n11978), .B2(n11966), .A(n11965), .ZN(n14986) );
  INV_X1 U15071 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19935) );
  AOI22_X1 U15072 ( .A1(n14285), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11967) );
  OAI21_X1 U15073 ( .B1(n11978), .B2(n19935), .A(n11967), .ZN(n11968) );
  INV_X1 U15074 ( .A(n11968), .ZN(n15446) );
  NAND2_X1 U15075 ( .A1(n14286), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15076 ( .A1(n14285), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U15077 ( .A1(n14285), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11971) );
  OAI21_X1 U15078 ( .B1(n11978), .B2(n19939), .A(n11971), .ZN(n14259) );
  AND2_X2 U15079 ( .A1(n14973), .A2(n14259), .ZN(n15428) );
  AOI22_X1 U15080 ( .A1(n14285), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11972) );
  OAI21_X1 U15081 ( .B1(n11978), .B2(n19941), .A(n11972), .ZN(n15427) );
  NAND2_X1 U15082 ( .A1(n14286), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15083 ( .A1(n14285), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11973) );
  AND2_X1 U15084 ( .A1(n11974), .A2(n11973), .ZN(n14940) );
  NAND2_X1 U15085 ( .A1(n14286), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15086 ( .A1(n14285), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11975) );
  AND2_X1 U15087 ( .A1(n11976), .A2(n11975), .ZN(n12975) );
  AOI22_X1 U15088 ( .A1(n14285), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11977) );
  OAI21_X1 U15089 ( .B1(n11978), .B2(n19945), .A(n11977), .ZN(n14915) );
  INV_X1 U15090 ( .A(n11983), .ZN(n11982) );
  NAND2_X1 U15091 ( .A1(n14286), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15092 ( .A1(n14285), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11664), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11979) );
  AND2_X1 U15093 ( .A1(n11980), .A2(n11979), .ZN(n11984) );
  INV_X1 U15094 ( .A(n11984), .ZN(n11981) );
  NAND2_X1 U15095 ( .A1(n11982), .A2(n11981), .ZN(n14289) );
  NAND2_X1 U15096 ( .A1(n11983), .A2(n11984), .ZN(n11985) );
  NAND2_X1 U15097 ( .A1(n11986), .A2(n13295), .ZN(n11987) );
  NAND2_X2 U15098 ( .A1(n20039), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19948) );
  INV_X1 U15099 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18990) );
  NAND2_X1 U15100 ( .A1(n18990), .A2(n19908), .ZN(n19902) );
  NAND2_X1 U15101 ( .A1(n20027), .A2(n20026), .ZN(n13087) );
  NOR2_X1 U15102 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13087), .ZN(n16542) );
  INV_X1 U15103 ( .A(n16542), .ZN(n11989) );
  AND2_X1 U15104 ( .A1(n19305), .A2(n11989), .ZN(n14290) );
  INV_X1 U15105 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n11990) );
  NAND2_X1 U15106 ( .A1(n11990), .A2(n12014), .ZN(n11991) );
  NOR2_X1 U15107 ( .A1(n13079), .A2(n11991), .ZN(n11992) );
  OR2_X2 U15108 ( .A1(n14290), .A2(n11992), .ZN(n19147) );
  NAND2_X1 U15109 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19147), .ZN(n11994) );
  NAND2_X1 U15110 ( .A1(n19971), .A2(n16540), .ZN(n18992) );
  INV_X2 U15111 ( .A(n19324), .ZN(n16460) );
  NAND2_X1 U15112 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20017), .ZN(n19368) );
  NOR2_X1 U15113 ( .A1(n19891), .A2(n19368), .ZN(n16537) );
  AOI22_X1 U15114 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19115), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n9962), .ZN(n11993) );
  NAND2_X1 U15115 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  AOI21_X1 U15116 ( .B1(n15405), .B2(n16306), .A(n11995), .ZN(n11996) );
  OAI21_X1 U15117 ( .B1(n14397), .B2(n19149), .A(n11996), .ZN(n11997) );
  INV_X1 U15118 ( .A(n12912), .ZN(n12819) );
  MUX2_X1 U15119 ( .A(n12819), .B(n12612), .S(n12911), .Z(n12000) );
  INV_X1 U15120 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11999) );
  INV_X4 U15121 ( .A(n11998), .ZN(n12883) );
  MUX2_X1 U15122 ( .A(n12000), .B(n11999), .S(n12883), .Z(n12669) );
  MUX2_X1 U15123 ( .A(n12837), .B(n12903), .S(n12929), .Z(n12821) );
  INV_X1 U15124 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12655) );
  INV_X1 U15125 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U15126 ( .A1(n12655), .A2(n13121), .ZN(n12002) );
  MUX2_X1 U15127 ( .A(n12831), .B(n12002), .S(n12883), .Z(n12660) );
  MUX2_X1 U15128 ( .A(n12609), .B(n12907), .S(n12929), .Z(n12005) );
  INV_X1 U15129 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12004) );
  MUX2_X1 U15130 ( .A(n12005), .B(n12004), .S(n12883), .Z(n12652) );
  MUX2_X1 U15131 ( .A(n12643), .B(P2_EBX_REG_5__SCAN_IN), .S(n12883), .Z(
        n12647) );
  INV_X1 U15132 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19111) );
  MUX2_X1 U15133 ( .A(n12006), .B(n19111), .S(n12883), .Z(n12701) );
  INV_X1 U15134 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12007) );
  MUX2_X1 U15135 ( .A(n12646), .B(n12007), .S(n12883), .Z(n12705) );
  NAND2_X1 U15136 ( .A1(n12883), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12709) );
  INV_X1 U15137 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U15138 ( .A1(n12714), .A2(n12008), .ZN(n12717) );
  INV_X1 U15139 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13619) );
  NAND2_X1 U15140 ( .A1(n12720), .A2(n13619), .ZN(n12730) );
  NAND2_X1 U15141 ( .A1(n12883), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12732) );
  OAI21_X1 U15142 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n12883), .ZN(n12009) );
  AND2_X1 U15143 ( .A1(n12883), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12748) );
  AND2_X1 U15144 ( .A1(n12883), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U15145 ( .A1(n12883), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12738) );
  INV_X1 U15146 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15393) );
  NAND2_X1 U15147 ( .A1(n12883), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12010) );
  NAND2_X1 U15148 ( .A1(n12737), .A2(n12010), .ZN(n12779) );
  AND2_X1 U15149 ( .A1(n12883), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12782) );
  INV_X1 U15150 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15360) );
  NAND2_X1 U15151 ( .A1(n12883), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12797) );
  AND2_X1 U15152 ( .A1(n12883), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12808) );
  OR2_X2 U15153 ( .A1(n12809), .A2(n12808), .ZN(n14345) );
  NAND2_X1 U15154 ( .A1(n12883), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14346) );
  INV_X1 U15155 ( .A(n14346), .ZN(n12011) );
  INV_X1 U15156 ( .A(n14293), .ZN(n12013) );
  NAND2_X1 U15157 ( .A1(n12883), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12012) );
  XNOR2_X1 U15158 ( .A(n12013), .B(n12012), .ZN(n14350) );
  NAND2_X1 U15159 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12014), .ZN(n12015) );
  NOR2_X1 U15160 ( .A1(n12929), .A2(n12015), .ZN(n12016) );
  NAND2_X1 U15161 ( .A1(n14350), .A2(n19102), .ZN(n12017) );
  NAND2_X1 U15162 ( .A1(n12019), .A2(n10299), .ZN(P2_U2825) );
  INV_X1 U15163 ( .A(n12020), .ZN(n12021) );
  AND2_X1 U15164 ( .A1(n13065), .A2(n13201), .ZN(n12029) );
  NOR3_X1 U15165 ( .A1(n12026), .A2(n12025), .A3(n12024), .ZN(n12028) );
  NOR2_X1 U15166 ( .A1(n12028), .A2(n12027), .ZN(n13064) );
  NAND2_X1 U15167 ( .A1(n12029), .A2(n13064), .ZN(n13056) );
  NAND2_X1 U15168 ( .A1(n13308), .A2(n13056), .ZN(n20970) );
  NOR2_X1 U15169 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16000) );
  NAND2_X1 U15170 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16000), .ZN(n15997) );
  NAND2_X1 U15171 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20968), .ZN(n12031) );
  OAI22_X1 U15172 ( .A1(n20968), .A2(n15997), .B1(n12031), .B2(n12030), .ZN(
        n12032) );
  NAND2_X1 U15173 ( .A1(n20123), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13664) );
  NAND2_X1 U15174 ( .A1(n14387), .A2(n20089), .ZN(n12155) );
  INV_X1 U15175 ( .A(n13019), .ZN(n20307) );
  NAND2_X1 U15176 ( .A1(n20307), .A2(n13280), .ZN(n12049) );
  AOI22_X1 U15177 ( .A1(n13333), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13059), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14406) );
  INV_X1 U15178 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20249) );
  NAND2_X1 U15179 ( .A1(n12049), .A2(n20249), .ZN(n12035) );
  INV_X1 U15180 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13669) );
  NAND2_X1 U15181 ( .A1(n13349), .A2(n13669), .ZN(n12034) );
  NAND3_X1 U15182 ( .A1(n12035), .A2(n12132), .A3(n12034), .ZN(n12036) );
  NAND2_X1 U15183 ( .A1(n12049), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12038) );
  INV_X1 U15184 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U15185 ( .A1(n12132), .A2(n13389), .ZN(n12037) );
  NAND2_X1 U15186 ( .A1(n12038), .A2(n12037), .ZN(n13334) );
  XNOR2_X1 U15187 ( .A(n12039), .B(n13334), .ZN(n13043) );
  NAND2_X1 U15188 ( .A1(n13043), .A2(n13349), .ZN(n13042) );
  OR2_X1 U15189 ( .A1(n12040), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U15190 ( .A1(n12049), .A2(n20261), .ZN(n12044) );
  INV_X1 U15191 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12042) );
  NAND2_X1 U15192 ( .A1(n13349), .A2(n12042), .ZN(n12043) );
  NAND3_X1 U15193 ( .A1(n12044), .A2(n12132), .A3(n12043), .ZN(n12045) );
  AND2_X1 U15194 ( .A1(n12046), .A2(n12045), .ZN(n13418) );
  MUX2_X1 U15195 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12048) );
  OAI21_X1 U15196 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13333), .A(
        n12048), .ZN(n13547) );
  INV_X1 U15197 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U15198 ( .A1(n12050), .A2(n13059), .ZN(n12101) );
  NAND2_X1 U15199 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13059), .ZN(
        n12051) );
  AND2_X1 U15200 ( .A1(n12101), .A2(n12051), .ZN(n12053) );
  MUX2_X1 U15201 ( .A(n12040), .B(n12049), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12052) );
  NAND2_X1 U15202 ( .A1(n12053), .A2(n12052), .ZN(n13578) );
  NAND2_X1 U15203 ( .A1(n13579), .A2(n13578), .ZN(n16274) );
  INV_X1 U15204 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20156) );
  NAND2_X1 U15205 ( .A1(n13349), .A2(n20156), .ZN(n12055) );
  NAND2_X1 U15206 ( .A1(n12132), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12054) );
  NAND3_X1 U15207 ( .A1(n12055), .A2(n12049), .A3(n12054), .ZN(n12056) );
  OAI21_X1 U15208 ( .B1(n12122), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12056), .ZN(
        n16273) );
  NAND2_X1 U15209 ( .A1(n13059), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12057) );
  AND2_X1 U15210 ( .A1(n12101), .A2(n12057), .ZN(n12059) );
  MUX2_X1 U15211 ( .A(n12040), .B(n12049), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12058) );
  NAND2_X1 U15212 ( .A1(n12059), .A2(n12058), .ZN(n16259) );
  INV_X1 U15213 ( .A(n12122), .ZN(n12079) );
  INV_X1 U15214 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20150) );
  NAND2_X1 U15215 ( .A1(n12079), .A2(n20150), .ZN(n12063) );
  NAND2_X1 U15216 ( .A1(n13349), .A2(n20150), .ZN(n12061) );
  NAND2_X1 U15217 ( .A1(n12121), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12060) );
  NAND3_X1 U15218 ( .A1(n12061), .A2(n12049), .A3(n12060), .ZN(n12062) );
  AND2_X1 U15219 ( .A1(n12063), .A2(n12062), .ZN(n16258) );
  NAND2_X1 U15220 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13059), .ZN(
        n12064) );
  AND2_X1 U15221 ( .A1(n12101), .A2(n12064), .ZN(n12066) );
  MUX2_X1 U15222 ( .A(n12040), .B(n12049), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12065) );
  NAND2_X1 U15223 ( .A1(n12066), .A2(n12065), .ZN(n13862) );
  INV_X1 U15224 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20144) );
  NAND2_X1 U15225 ( .A1(n12079), .A2(n20144), .ZN(n12070) );
  NAND2_X1 U15226 ( .A1(n13349), .A2(n20144), .ZN(n12068) );
  NAND2_X1 U15227 ( .A1(n12121), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12067) );
  NAND3_X1 U15228 ( .A1(n12068), .A2(n12049), .A3(n12067), .ZN(n12069) );
  AND2_X1 U15229 ( .A1(n12070), .A2(n12069), .ZN(n16247) );
  NAND2_X1 U15230 ( .A1(n16248), .A2(n16247), .ZN(n16250) );
  OR2_X1 U15231 ( .A1(n12040), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U15232 ( .A1(n12049), .A2(n14727), .ZN(n12072) );
  INV_X1 U15233 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13983) );
  NAND2_X1 U15234 ( .A1(n13349), .A2(n13983), .ZN(n12071) );
  NAND3_X1 U15235 ( .A1(n12072), .A2(n12132), .A3(n12071), .ZN(n12073) );
  MUX2_X1 U15236 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12075) );
  OAI21_X1 U15237 ( .B1(n13333), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12075), .ZN(n14062) );
  NAND2_X1 U15238 ( .A1(n13059), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12076) );
  AND2_X1 U15239 ( .A1(n12101), .A2(n12076), .ZN(n12078) );
  MUX2_X1 U15240 ( .A(n12040), .B(n12049), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12077) );
  NAND2_X1 U15241 ( .A1(n12078), .A2(n12077), .ZN(n14089) );
  INV_X1 U15242 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U15243 ( .A1(n12079), .A2(n14320), .ZN(n12083) );
  NAND2_X1 U15244 ( .A1(n13349), .A2(n14320), .ZN(n12081) );
  NAND2_X1 U15245 ( .A1(n12132), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12080) );
  NAND3_X1 U15246 ( .A1(n12081), .A2(n12049), .A3(n12080), .ZN(n12082) );
  OR2_X1 U15247 ( .A1(n12040), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12087) );
  NAND2_X1 U15248 ( .A1(n12049), .A2(n14209), .ZN(n12085) );
  INV_X1 U15249 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14055) );
  NAND2_X1 U15250 ( .A1(n13349), .A2(n14055), .ZN(n12084) );
  NAND3_X1 U15251 ( .A1(n12085), .A2(n12132), .A3(n12084), .ZN(n12086) );
  MUX2_X1 U15252 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12088) );
  OAI21_X1 U15253 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13333), .A(
        n12088), .ZN(n14559) );
  OR2_X1 U15254 ( .A1(n12040), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U15255 ( .A1(n12049), .A2(n12089), .ZN(n12091) );
  INV_X1 U15256 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16101) );
  NAND2_X1 U15257 ( .A1(n13349), .A2(n16101), .ZN(n12090) );
  NAND3_X1 U15258 ( .A1(n12091), .A2(n12121), .A3(n12090), .ZN(n12092) );
  NAND2_X1 U15259 ( .A1(n12093), .A2(n12092), .ZN(n14554) );
  NAND2_X1 U15260 ( .A1(n14562), .A2(n14554), .ZN(n14556) );
  MUX2_X1 U15261 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12094) );
  OAI21_X1 U15262 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13333), .A(
        n12094), .ZN(n14475) );
  MUX2_X1 U15263 ( .A(n12040), .B(n12049), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12096) );
  NAND2_X1 U15264 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n13059), .ZN(
        n12095) );
  INV_X1 U15265 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21209) );
  NAND2_X1 U15266 ( .A1(n13349), .A2(n21209), .ZN(n12098) );
  NAND2_X1 U15267 ( .A1(n12132), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12097) );
  NAND3_X1 U15268 ( .A1(n12098), .A2(n12049), .A3(n12097), .ZN(n12099) );
  OAI21_X1 U15269 ( .B1(n12122), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12099), .ZN(
        n16084) );
  NAND2_X1 U15270 ( .A1(n13059), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12100) );
  AND2_X1 U15271 ( .A1(n12101), .A2(n12100), .ZN(n12103) );
  MUX2_X1 U15272 ( .A(n12040), .B(n12049), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12102) );
  NAND2_X1 U15273 ( .A1(n12103), .A2(n12102), .ZN(n14538) );
  MUX2_X1 U15274 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12105) );
  OR2_X1 U15275 ( .A1(n13333), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U15276 ( .A1(n14540), .A2(n14531), .ZN(n14533) );
  OR2_X1 U15277 ( .A1(n12040), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12109) );
  INV_X1 U15278 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U15279 ( .A1(n12049), .A2(n14823), .ZN(n12107) );
  INV_X1 U15280 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16046) );
  NAND2_X1 U15281 ( .A1(n13349), .A2(n16046), .ZN(n12106) );
  NAND3_X1 U15282 ( .A1(n12107), .A2(n12132), .A3(n12106), .ZN(n12108) );
  MUX2_X1 U15283 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12110) );
  OAI21_X1 U15284 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13333), .A(
        n12110), .ZN(n14805) );
  OR2_X1 U15285 ( .A1(n12040), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12114) );
  NAND2_X1 U15286 ( .A1(n12049), .A2(n14797), .ZN(n12112) );
  INV_X1 U15287 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U15288 ( .A1(n13349), .A2(n14521), .ZN(n12111) );
  NAND3_X1 U15289 ( .A1(n12112), .A2(n12132), .A3(n12111), .ZN(n12113) );
  NAND2_X1 U15290 ( .A1(n12114), .A2(n12113), .ZN(n14518) );
  MUX2_X1 U15291 ( .A(n12122), .B(n12132), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12116) );
  OR2_X1 U15292 ( .A1(n13333), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12115) );
  AND2_X1 U15293 ( .A1(n12116), .A2(n12115), .ZN(n14459) );
  OR2_X1 U15294 ( .A1(n12040), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12120) );
  INV_X1 U15295 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U15296 ( .A1(n12049), .A2(n14778), .ZN(n12118) );
  INV_X1 U15297 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14513) );
  NAND2_X1 U15298 ( .A1(n13349), .A2(n14513), .ZN(n12117) );
  NAND3_X1 U15299 ( .A1(n12118), .A2(n12132), .A3(n12117), .ZN(n12119) );
  AND2_X1 U15300 ( .A1(n12120), .A2(n12119), .ZN(n14451) );
  MUX2_X1 U15301 ( .A(n12122), .B(n12121), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12123) );
  OAI21_X1 U15302 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13333), .A(
        n12123), .ZN(n14432) );
  OR2_X1 U15303 ( .A1(n12040), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U15304 ( .A1(n12049), .A2(n12124), .ZN(n12127) );
  INV_X1 U15305 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U15306 ( .A1(n13349), .A2(n12125), .ZN(n12126) );
  NAND3_X1 U15307 ( .A1(n12127), .A2(n12132), .A3(n12126), .ZN(n12128) );
  OR2_X1 U15308 ( .A1(n13333), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12131) );
  INV_X1 U15309 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U15310 ( .A1(n13349), .A2(n14511), .ZN(n12130) );
  NAND2_X1 U15311 ( .A1(n12131), .A2(n12130), .ZN(n14402) );
  OAI22_X1 U15312 ( .A1(n14402), .A2(n10456), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12040), .ZN(n14417) );
  NAND2_X1 U15313 ( .A1(n14418), .A2(n14417), .ZN(n14416) );
  MUX2_X1 U15314 ( .A(n14406), .B(n12132), .S(n14416), .Z(n12134) );
  AOI22_X1 U15315 ( .A1(n13333), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13059), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12133) );
  NAND2_X1 U15316 ( .A1(n13309), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12143) );
  AND2_X1 U15317 ( .A1(n20972), .A2(n20965), .ZN(n12135) );
  NOR2_X1 U15318 ( .A1(n12143), .A2(n12135), .ZN(n12137) );
  NAND2_X1 U15319 ( .A1(n20123), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13667) );
  INV_X1 U15320 ( .A(n13667), .ZN(n12136) );
  AND2_X1 U15321 ( .A1(n13280), .A2(n12136), .ZN(n12144) );
  NAND2_X1 U15322 ( .A1(n12138), .A2(n20865), .ZN(n16016) );
  INV_X1 U15323 ( .A(n16016), .ZN(n15991) );
  OAI21_X1 U15324 ( .B1(n13309), .B2(n15991), .A(n20972), .ZN(n13002) );
  INV_X1 U15325 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20914) );
  INV_X1 U15326 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20911) );
  INV_X1 U15327 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20898) );
  INV_X1 U15328 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20900) );
  INV_X1 U15329 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20887) );
  NAND4_X1 U15330 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14499)
         );
  INV_X1 U15331 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21118) );
  NAND3_X1 U15332 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14495) );
  NOR2_X1 U15333 ( .A1(n21118), .A2(n14495), .ZN(n20069) );
  NAND2_X1 U15334 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20069), .ZN(n14010) );
  NOR3_X1 U15335 ( .A1(n20887), .A2(n14499), .A3(n14010), .ZN(n14326) );
  INV_X1 U15336 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20893) );
  NAND2_X1 U15337 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14327) );
  NOR2_X1 U15338 ( .A1(n20893), .A2(n14327), .ZN(n14486) );
  NAND3_X1 U15339 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14326), .A3(n14486), 
        .ZN(n16097) );
  NAND3_X1 U15340 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n16076) );
  NOR4_X1 U15341 ( .A1(n20898), .A2(n20900), .A3(n16097), .A4(n16076), .ZN(
        n16067) );
  AND2_X1 U15342 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n16036) );
  NAND4_X1 U15343 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n16067), .A4(n16036), .ZN(n16026) );
  INV_X1 U15344 ( .A(n16026), .ZN(n12140) );
  NAND3_X1 U15345 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(n12140), .ZN(n14449) );
  NOR2_X1 U15346 ( .A1(n20911), .A2(n14449), .ZN(n14435) );
  NAND2_X1 U15347 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14435), .ZN(n14236) );
  NOR2_X1 U15348 ( .A1(n20914), .A2(n14236), .ZN(n14422) );
  INV_X1 U15349 ( .A(n14422), .ZN(n12141) );
  INV_X1 U15350 ( .A(n20123), .ZN(n16045) );
  AOI21_X1 U15351 ( .B1(n20127), .B2(n12141), .A(n16045), .ZN(n14425) );
  INV_X1 U15352 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20916) );
  INV_X1 U15353 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n12147) );
  OAI21_X1 U15354 ( .B1(n20916), .B2(n12147), .A(n20127), .ZN(n12142) );
  NAND2_X1 U15355 ( .A1(n14425), .A2(n12142), .ZN(n14409) );
  INV_X1 U15356 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12150) );
  AND2_X1 U15357 ( .A1(n12144), .A2(n12143), .ZN(n12145) );
  AND2_X2 U15358 ( .A1(n12146), .A2(n12145), .ZN(n20125) );
  NAND3_X1 U15359 ( .A1(n20127), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14422), 
        .ZN(n14408) );
  NOR3_X1 U15360 ( .A1(n14408), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12147), 
        .ZN(n12148) );
  AOI21_X1 U15361 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(n20125), .A(n12148), .ZN(
        n12149) );
  OAI21_X1 U15362 ( .B1(n20100), .B2(n12150), .A(n12149), .ZN(n12151) );
  AOI21_X1 U15363 ( .B1(n14409), .B2(P1_REIP_REG_31__SCAN_IN), .A(n12151), 
        .ZN(n12152) );
  NAND2_X1 U15364 ( .A1(n12155), .A2(n12154), .ZN(P1_U2809) );
  AOI22_X1 U15365 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15366 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12211), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15367 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12157) );
  OAI21_X1 U15368 ( .B1(n9874), .B2(n21204), .A(n12157), .ZN(n12169) );
  AOI22_X1 U15369 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12167) );
  NOR2_X2 U15370 ( .A1(n12160), .A2(n17074), .ZN(n17326) );
  AOI22_X1 U15371 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12166) );
  NOR2_X1 U15372 ( .A1(n12160), .A2(n12159), .ZN(n12183) );
  AOI22_X1 U15373 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12165) );
  NOR2_X2 U15374 ( .A1(n12162), .A2(n12161), .ZN(n12302) );
  NAND2_X1 U15375 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12163), .ZN(
        n15942) );
  AOI22_X1 U15376 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12164) );
  NAND4_X1 U15377 ( .A1(n12167), .A2(n12166), .A3(n12165), .A4(n12164), .ZN(
        n12168) );
  AOI211_X1 U15378 ( .C1(n17178), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12169), .B(n12168), .ZN(n12170) );
  INV_X2 U15379 ( .A(n12337), .ZN(n17303) );
  AOI22_X1 U15380 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15381 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15382 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15383 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12173) );
  NAND4_X1 U15384 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12182) );
  AOI22_X1 U15385 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15386 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15387 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15388 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12177) );
  NAND4_X1 U15389 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(
        n12181) );
  AOI22_X1 U15390 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15391 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12186) );
  INV_X2 U15392 ( .A(n17322), .ZN(n17302) );
  AOI22_X1 U15393 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15394 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12184) );
  NAND4_X1 U15395 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12193) );
  AOI22_X1 U15396 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15397 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15398 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15399 ( .A1(n12302), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15400 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12192) );
  AOI22_X1 U15401 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12194) );
  OAI21_X1 U15402 ( .B1(n14198), .B2(n17282), .A(n12194), .ZN(n12195) );
  INV_X1 U15403 ( .A(n12195), .ZN(n12206) );
  AOI22_X1 U15404 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12196) );
  INV_X1 U15405 ( .A(n12196), .ZN(n12200) );
  AOI22_X1 U15406 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12302), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U15407 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  AOI22_X1 U15408 ( .A1(n12244), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12241), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15409 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12211), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15410 ( .A1(n12246), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15411 ( .A1(n12242), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12240), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12201) );
  NAND3_X1 U15412 ( .A1(n12206), .A2(n12205), .A3(n10307), .ZN(n12257) );
  AOI22_X1 U15413 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17326), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12302), .ZN(n12215) );
  AOI22_X1 U15414 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9820), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n12244), .ZN(n12207) );
  OAI21_X1 U15415 ( .B1(n12229), .B2(n21243), .A(n12207), .ZN(n12210) );
  AOI22_X1 U15416 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12241), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n12208), .ZN(n12209) );
  AOI22_X1 U15417 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12242), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15418 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12211), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15419 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n9819), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15420 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12240), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15421 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15422 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12227) );
  INV_X4 U15423 ( .A(n12337), .ZN(n17320) );
  INV_X1 U15424 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n21190) );
  AOI22_X1 U15425 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12219) );
  OAI21_X1 U15426 ( .B1(n17300), .B2(n21190), .A(n12219), .ZN(n12225) );
  AOI22_X1 U15427 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15428 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15429 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12246), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15430 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U15431 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12224) );
  AOI211_X1 U15432 ( .C1(n17320), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n12225), .B(n12224), .ZN(n12226) );
  NAND3_X1 U15433 ( .A1(n12228), .A2(n12227), .A3(n12226), .ZN(n12449) );
  NAND2_X1 U15434 ( .A1(n12264), .A2(n12449), .ZN(n12267) );
  AOI22_X1 U15435 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15436 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12238) );
  INV_X1 U15437 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U15438 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12230) );
  OAI21_X1 U15439 ( .B1(n17022), .B2(n17344), .A(n12230), .ZN(n12236) );
  AOI22_X1 U15440 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15441 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15442 ( .A1(n17317), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15443 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12231) );
  NAND4_X1 U15444 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12235) );
  AOI211_X1 U15445 ( .C1(n17324), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n12236), .B(n12235), .ZN(n12237) );
  NAND3_X1 U15446 ( .A1(n12239), .A2(n12238), .A3(n12237), .ZN(n12456) );
  XNOR2_X1 U15447 ( .A(n12258), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17981) );
  AOI22_X1 U15448 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12211), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15449 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12255) );
  INV_X1 U15450 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21178) );
  AOI22_X1 U15451 ( .A1(n12242), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12241), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12243) );
  OAI21_X1 U15452 ( .B1(n14198), .B2(n21178), .A(n12243), .ZN(n12253) );
  AOI22_X1 U15453 ( .A1(n12245), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12244), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15454 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12302), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15455 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12246), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15456 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9820), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12248) );
  NAND4_X1 U15457 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12252) );
  AOI211_X1 U15458 ( .C1(n17317), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n12253), .B(n12252), .ZN(n12254) );
  NAND3_X1 U15459 ( .A1(n12256), .A2(n12255), .A3(n12254), .ZN(n17992) );
  INV_X1 U15460 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18927) );
  INV_X1 U15461 ( .A(n17507), .ZN(n12437) );
  XOR2_X1 U15462 ( .A(n12437), .B(n12260), .Z(n12261) );
  XNOR2_X1 U15463 ( .A(n12262), .B(n12261), .ZN(n17962) );
  NOR2_X1 U15464 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  INV_X1 U15465 ( .A(n12449), .ZN(n17503) );
  XNOR2_X1 U15466 ( .A(n17503), .B(n12264), .ZN(n12265) );
  XNOR2_X1 U15467 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12265), .ZN(
        n17954) );
  INV_X1 U15468 ( .A(n17500), .ZN(n12438) );
  XOR2_X1 U15469 ( .A(n12438), .B(n12267), .Z(n17934) );
  NOR2_X1 U15470 ( .A1(n17932), .A2(n17934), .ZN(n12268) );
  NAND2_X1 U15471 ( .A1(n17932), .A2(n17934), .ZN(n17933) );
  OAI21_X1 U15472 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12268), .A(
        n17933), .ZN(n17926) );
  INV_X1 U15473 ( .A(n12456), .ZN(n17496) );
  XNOR2_X1 U15474 ( .A(n17496), .B(n12269), .ZN(n12270) );
  XNOR2_X1 U15475 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12270), .ZN(
        n17928) );
  NOR2_X1 U15476 ( .A1(n17926), .A2(n17928), .ZN(n17927) );
  OAI21_X1 U15477 ( .B1(n12272), .B2(n15959), .A(n17780), .ZN(n12273) );
  NOR2_X1 U15478 ( .A1(n12274), .A2(n12273), .ZN(n12275) );
  NAND2_X1 U15479 ( .A1(n17878), .A2(n18212), .ZN(n17865) );
  INV_X1 U15480 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18150) );
  INV_X1 U15481 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12277) );
  INV_X1 U15482 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12276) );
  AND2_X1 U15483 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  NAND2_X1 U15484 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18196) );
  NOR2_X1 U15485 ( .A1(n21056), .A2(n18196), .ZN(n18175) );
  NAND3_X1 U15486 ( .A1(n18175), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17802) );
  NOR2_X1 U15487 ( .A1(n18169), .A2(n17802), .ZN(n18123) );
  NAND2_X1 U15488 ( .A1(n18123), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16560) );
  NAND2_X1 U15489 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12289) );
  INV_X1 U15490 ( .A(n12289), .ZN(n18105) );
  INV_X1 U15491 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18078) );
  NAND2_X1 U15492 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18077) );
  NOR3_X1 U15493 ( .A1(n17764), .A2(n18078), .A3(n18077), .ZN(n12290) );
  NAND2_X1 U15494 ( .A1(n18105), .A2(n12290), .ZN(n18065) );
  NOR2_X1 U15495 ( .A1(n18065), .A2(n18066), .ZN(n18012) );
  NAND2_X1 U15496 ( .A1(n18012), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17690) );
  NAND2_X1 U15497 ( .A1(n17764), .A2(n17780), .ZN(n17763) );
  NOR2_X1 U15498 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17763), .ZN(
        n12281) );
  INV_X1 U15499 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18088) );
  NAND2_X1 U15500 ( .A1(n12281), .A2(n18088), .ZN(n17725) );
  INV_X1 U15501 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17709) );
  NAND3_X1 U15502 ( .A1(n17712), .A2(n18066), .A3(n17709), .ZN(n12282) );
  INV_X1 U15503 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18125) );
  INV_X1 U15504 ( .A(n12284), .ZN(n12285) );
  INV_X1 U15505 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17692) );
  NAND2_X1 U15506 ( .A1(n17693), .A2(n17692), .ZN(n17691) );
  NAND2_X1 U15507 ( .A1(n12290), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18041) );
  NOR2_X1 U15508 ( .A1(n17765), .A2(n18041), .ZN(n17696) );
  NAND3_X1 U15509 ( .A1(n17691), .A2(n17696), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12292) );
  INV_X1 U15510 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18025) );
  NAND2_X1 U15511 ( .A1(n17780), .A2(n17691), .ZN(n17679) );
  NAND2_X1 U15512 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12470) );
  INV_X1 U15513 ( .A(n16597), .ZN(n17649) );
  INV_X1 U15514 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21268) );
  NAND2_X1 U15515 ( .A1(n10072), .A2(n21268), .ZN(n16596) );
  INV_X1 U15516 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16571) );
  INV_X1 U15517 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16011) );
  OAI21_X1 U15518 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n10072), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12294) );
  OAI221_X1 U15519 ( .B1(n16005), .B2(n16011), .C1(n10072), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n12294), .ZN(n12301) );
  NOR2_X1 U15520 ( .A1(n10072), .A2(n16004), .ZN(n12300) );
  OAI21_X1 U15521 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16011), .A(
        n16005), .ZN(n12298) );
  NAND2_X1 U15522 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10072), .ZN(
        n12296) );
  OAI22_X1 U15523 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10072), .B1(
        n12296), .B2(n16011), .ZN(n12297) );
  OAI21_X1 U15524 ( .B1(n12298), .B2(n12300), .A(n12297), .ZN(n12299) );
  OAI21_X1 U15525 ( .B1(n12301), .B2(n12300), .A(n12299), .ZN(n16595) );
  AOI22_X1 U15526 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15527 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15528 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15529 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15530 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12313) );
  AOI22_X1 U15531 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15532 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14185), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15533 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15534 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U15535 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12312) );
  AOI22_X1 U15536 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15537 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15538 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15539 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12314) );
  NAND4_X1 U15540 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12324) );
  AOI22_X1 U15541 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15542 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17272), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15543 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15544 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15545 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12323) );
  NAND2_X1 U15546 ( .A1(n18335), .A2(n18338), .ZN(n12405) );
  NOR2_X1 U15547 ( .A1(n18338), .A2(n18335), .ZN(n12397) );
  INV_X1 U15548 ( .A(n12397), .ZN(n12325) );
  NAND2_X1 U15549 ( .A1(n12405), .A2(n12325), .ZN(n18969) );
  AOI22_X1 U15550 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15551 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15552 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15553 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U15554 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12335) );
  AOI22_X1 U15555 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15556 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15557 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15558 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12330) );
  NAND4_X1 U15559 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12334) );
  AOI22_X1 U15560 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15561 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15562 ( .A1(n17317), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12336) );
  OAI21_X1 U15563 ( .B1(n12337), .B2(n17344), .A(n12336), .ZN(n12343) );
  AOI22_X1 U15564 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15565 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15566 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15567 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12242), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12338) );
  NAND4_X1 U15568 ( .A1(n12341), .A2(n12340), .A3(n12339), .A4(n12338), .ZN(
        n12342) );
  AOI211_X1 U15569 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n12343), .B(n12342), .ZN(n12344) );
  NAND3_X1 U15570 ( .A1(n12346), .A2(n12345), .A3(n12344), .ZN(n18361) );
  AOI22_X1 U15571 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15572 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15573 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12347) );
  OAI21_X1 U15574 ( .B1(n12348), .B2(n17282), .A(n12347), .ZN(n12354) );
  AOI22_X1 U15575 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15576 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15577 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15578 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12349) );
  NAND4_X1 U15579 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12353) );
  AOI211_X1 U15580 ( .C1(n12247), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12354), .B(n12353), .ZN(n12355) );
  NAND3_X1 U15581 ( .A1(n12357), .A2(n12356), .A3(n12355), .ZN(n18342) );
  AOI22_X1 U15582 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9827), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15583 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15584 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15585 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15586 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12367) );
  AOI22_X1 U15587 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15588 ( .A1(n17317), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15589 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15590 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12362) );
  NAND4_X1 U15591 ( .A1(n12365), .A2(n12364), .A3(n12363), .A4(n12362), .ZN(
        n12366) );
  NAND2_X1 U15592 ( .A1(n18357), .A2(n15945), .ZN(n15944) );
  AOI22_X1 U15593 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12368) );
  OAI21_X1 U15594 ( .B1(n12318), .B2(n21204), .A(n12368), .ZN(n12374) );
  AOI22_X1 U15595 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17178), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15596 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15597 ( .A1(n17303), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15598 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15599 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  AOI211_X2 U15600 ( .C1(n14169), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n12374), .B(n12373), .ZN(n12375) );
  AOI22_X1 U15601 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15602 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15603 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12378) );
  OAI21_X1 U15604 ( .B1(n12379), .B2(n21140), .A(n12378), .ZN(n12385) );
  AOI22_X1 U15605 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15606 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15607 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15608 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15609 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12384) );
  AOI211_X1 U15610 ( .C1(n17178), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12385), .B(n12384), .ZN(n12386) );
  NAND3_X1 U15611 ( .A1(n12388), .A2(n12387), .A3(n12386), .ZN(n18346) );
  INV_X1 U15612 ( .A(n12403), .ZN(n12412) );
  NAND2_X1 U15613 ( .A1(n18335), .A2(n18367), .ZN(n12407) );
  NOR2_X1 U15614 ( .A1(n18346), .A2(n12407), .ZN(n12389) );
  NOR2_X1 U15615 ( .A1(n17377), .A2(n12390), .ZN(n12391) );
  NAND3_X1 U15616 ( .A1(n18354), .A2(n12389), .A3(n12391), .ZN(n12404) );
  NOR2_X1 U15617 ( .A1(n12390), .A2(n18361), .ZN(n18787) );
  NOR2_X1 U15618 ( .A1(n17519), .A2(n12391), .ZN(n12395) );
  NOR2_X1 U15619 ( .A1(n17377), .A2(n18357), .ZN(n12401) );
  INV_X1 U15620 ( .A(n18335), .ZN(n16711) );
  NOR3_X1 U15621 ( .A1(n18774), .A2(n12401), .A3(n16711), .ZN(n12393) );
  AOI21_X1 U15622 ( .B1(n12405), .B2(n15945), .A(n12391), .ZN(n12392) );
  AOI21_X1 U15623 ( .B1(n15945), .B2(n12393), .A(n12392), .ZN(n12394) );
  OAI21_X1 U15624 ( .B1(n12395), .B2(n18354), .A(n12394), .ZN(n12396) );
  AOI21_X1 U15625 ( .B1(n18354), .B2(n18787), .A(n12396), .ZN(n15932) );
  OAI21_X1 U15626 ( .B1(n17519), .B2(n18787), .A(n12397), .ZN(n15931) );
  NAND3_X1 U15627 ( .A1(n18346), .A2(n15931), .A3(n12398), .ZN(n12399) );
  OAI21_X1 U15628 ( .B1(n18346), .B2(n12407), .A(n12399), .ZN(n12400) );
  NAND2_X1 U15629 ( .A1(n15932), .A2(n12400), .ZN(n12409) );
  NAND2_X1 U15630 ( .A1(n18972), .A2(n14103), .ZN(n12406) );
  NOR4_X4 U15631 ( .A1(n18335), .A2(n12403), .A3(n12402), .A4(n18357), .ZN(
        n17581) );
  NOR2_X2 U15632 ( .A1(n15945), .A2(n12404), .ZN(n15934) );
  INV_X2 U15633 ( .A(n12408), .ZN(n15935) );
  NAND2_X1 U15634 ( .A1(n18338), .A2(n18761), .ZN(n12411) );
  INV_X1 U15635 ( .A(n12409), .ZN(n12410) );
  AOI21_X4 U15636 ( .B1(n18773), .B2(n15935), .A(n18772), .ZN(n18197) );
  AOI21_X1 U15637 ( .B1(n12413), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12429), .ZN(n12435) );
  AOI22_X1 U15638 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18793), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12414), .ZN(n12434) );
  AOI22_X1 U15639 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18798), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n12415), .ZN(n12421) );
  NAND2_X1 U15640 ( .A1(n12434), .A2(n12429), .ZN(n12416) );
  OAI21_X1 U15641 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12414), .A(
        n12416), .ZN(n12420) );
  NAND2_X1 U15642 ( .A1(n12421), .A2(n12420), .ZN(n12417) );
  OAI22_X1 U15643 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18802), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12418), .ZN(n12423) );
  NOR2_X1 U15644 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18802), .ZN(
        n12419) );
  NAND2_X1 U15645 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12418), .ZN(
        n12422) );
  AOI22_X1 U15646 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12423), .B1(
        n12419), .B2(n12422), .ZN(n12425) );
  AND2_X1 U15647 ( .A1(n12434), .A2(n12425), .ZN(n12428) );
  XOR2_X1 U15648 ( .A(n12421), .B(n12420), .Z(n12426) );
  AND2_X1 U15649 ( .A1(n12422), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12424) );
  OAI22_X1 U15650 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18767), .B1(
        n12424), .B2(n12423), .ZN(n12430) );
  AOI21_X1 U15651 ( .B1(n12426), .B2(n12425), .A(n12430), .ZN(n12427) );
  INV_X1 U15652 ( .A(n12427), .ZN(n15928) );
  NOR2_X1 U15653 ( .A1(n18972), .A2(n18342), .ZN(n15953) );
  INV_X1 U15654 ( .A(n12429), .ZN(n12433) );
  INV_X1 U15655 ( .A(n12430), .ZN(n12432) );
  NAND2_X1 U15656 ( .A1(n12434), .A2(n12433), .ZN(n12431) );
  OAI211_X1 U15657 ( .C1(n12434), .C2(n12433), .A(n12432), .B(n12431), .ZN(
        n15927) );
  OAI21_X1 U15658 ( .B1(n12435), .B2(n15927), .A(n15928), .ZN(n18962) );
  NAND2_X1 U15659 ( .A1(n15953), .A2(n18962), .ZN(n15951) );
  NAND2_X1 U15660 ( .A1(n18972), .A2(n18035), .ZN(n18057) );
  INV_X1 U15661 ( .A(n17825), .ZN(n17975) );
  NAND2_X1 U15662 ( .A1(n17992), .A2(n17520), .ZN(n12441) );
  NAND2_X1 U15663 ( .A1(n12436), .A2(n12441), .ZN(n12440) );
  NAND2_X1 U15664 ( .A1(n12440), .A2(n12437), .ZN(n12450) );
  NOR2_X1 U15665 ( .A1(n17503), .A2(n12450), .ZN(n12439) );
  NAND2_X1 U15666 ( .A1(n12439), .A2(n12438), .ZN(n12457) );
  NOR2_X1 U15667 ( .A1(n17496), .A2(n12457), .ZN(n12461) );
  NAND2_X1 U15668 ( .A1(n12461), .A2(n15959), .ZN(n12462) );
  XNOR2_X1 U15669 ( .A(n12439), .B(n17500), .ZN(n12454) );
  AND2_X1 U15670 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12454), .ZN(
        n12455) );
  XOR2_X1 U15671 ( .A(n12440), .B(n17507), .Z(n12447) );
  NOR2_X1 U15672 ( .A1(n18280), .A2(n12447), .ZN(n12448) );
  XOR2_X1 U15673 ( .A(n12436), .B(n12441), .Z(n12442) );
  NOR2_X1 U15674 ( .A1(n12442), .A2(n18292), .ZN(n12446) );
  XNOR2_X1 U15675 ( .A(n18292), .B(n12442), .ZN(n17973) );
  INV_X1 U15676 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18944) );
  NOR2_X1 U15677 ( .A1(n12258), .A2(n18944), .ZN(n12445) );
  INV_X1 U15678 ( .A(n17992), .ZN(n12444) );
  NAND3_X1 U15679 ( .A1(n12444), .A2(n12258), .A3(n18944), .ZN(n12443) );
  OAI221_X1 U15680 ( .B1(n12445), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n12444), .C2(n12258), .A(n12443), .ZN(n17972) );
  NOR2_X1 U15681 ( .A1(n17973), .A2(n17972), .ZN(n17971) );
  NOR2_X1 U15682 ( .A1(n12446), .A2(n17971), .ZN(n17961) );
  XNOR2_X1 U15683 ( .A(n18280), .B(n12447), .ZN(n17960) );
  NOR2_X1 U15684 ( .A1(n17961), .A2(n17960), .ZN(n17959) );
  NOR2_X1 U15685 ( .A1(n12448), .A2(n17959), .ZN(n12451) );
  XOR2_X1 U15686 ( .A(n12450), .B(n12449), .Z(n12452) );
  NOR2_X1 U15687 ( .A1(n12451), .A2(n12452), .ZN(n12453) );
  INV_X1 U15688 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18261) );
  XNOR2_X1 U15689 ( .A(n12452), .B(n12451), .ZN(n17950) );
  NOR2_X1 U15690 ( .A1(n18261), .A2(n17950), .ZN(n17949) );
  NOR2_X1 U15691 ( .A1(n12453), .A2(n17949), .ZN(n17938) );
  XNOR2_X1 U15692 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12454), .ZN(
        n17937) );
  NOR2_X1 U15693 ( .A1(n17938), .A2(n17937), .ZN(n17936) );
  NOR2_X1 U15694 ( .A1(n12455), .A2(n17936), .ZN(n12458) );
  XOR2_X1 U15695 ( .A(n12457), .B(n12456), .Z(n12459) );
  NOR2_X1 U15696 ( .A1(n12458), .A2(n12459), .ZN(n12460) );
  XNOR2_X1 U15697 ( .A(n12459), .B(n12458), .ZN(n17925) );
  INV_X1 U15698 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18229) );
  NOR2_X1 U15699 ( .A1(n17925), .A2(n18229), .ZN(n17924) );
  NOR2_X1 U15700 ( .A1(n12460), .A2(n17924), .ZN(n12463) );
  XNOR2_X1 U15701 ( .A(n12461), .B(n15959), .ZN(n12464) );
  NAND2_X1 U15702 ( .A1(n12463), .A2(n12464), .ZN(n17907) );
  NAND2_X1 U15703 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17907), .ZN(
        n12466) );
  NOR2_X1 U15704 ( .A1(n12462), .A2(n12466), .ZN(n12468) );
  INV_X1 U15705 ( .A(n12462), .ZN(n12467) );
  OR2_X1 U15706 ( .A1(n12464), .A2(n12463), .ZN(n17908) );
  OAI21_X1 U15707 ( .B1(n12467), .B2(n12466), .A(n17908), .ZN(n12465) );
  AOI21_X1 U15708 ( .B1(n12467), .B2(n12466), .A(n12465), .ZN(n17900) );
  INV_X1 U15709 ( .A(n18123), .ZN(n18133) );
  NAND2_X1 U15710 ( .A1(n17817), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18056) );
  NOR2_X1 U15711 ( .A1(n17690), .A2(n17692), .ZN(n18020) );
  INV_X1 U15712 ( .A(n18020), .ZN(n18024) );
  NOR2_X1 U15713 ( .A1(n18056), .A2(n18024), .ZN(n17678) );
  INV_X1 U15714 ( .A(n12470), .ZN(n18001) );
  NAND2_X1 U15715 ( .A1(n17678), .A2(n18001), .ZN(n16567) );
  NAND2_X1 U15716 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15958) );
  INV_X1 U15717 ( .A(n15958), .ZN(n16569) );
  NAND2_X1 U15718 ( .A1(n16569), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16583) );
  NOR2_X1 U15719 ( .A1(n16567), .A2(n16583), .ZN(n16568) );
  NAND2_X1 U15720 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16568), .ZN(
        n12469) );
  XNOR2_X1 U15721 ( .A(n12469), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16592) );
  INV_X1 U15722 ( .A(n17986), .ZN(n17997) );
  NOR2_X2 U15723 ( .A1(n15959), .A2(n17997), .ZN(n17861) );
  INV_X1 U15724 ( .A(n18189), .ZN(n17810) );
  NAND2_X1 U15725 ( .A1(n18123), .A2(n17810), .ZN(n17809) );
  INV_X1 U15726 ( .A(n18132), .ZN(n17715) );
  NOR2_X1 U15727 ( .A1(n18024), .A2(n12470), .ZN(n16589) );
  INV_X1 U15728 ( .A(n16589), .ZN(n16561) );
  INV_X1 U15729 ( .A(n18002), .ZN(n12471) );
  NOR2_X1 U15730 ( .A1(n16583), .A2(n12471), .ZN(n16570) );
  NAND2_X1 U15731 ( .A1(n16570), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12472) );
  XNOR2_X1 U15732 ( .A(n12472), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16591) );
  AOI22_X1 U15733 ( .A1(n17983), .A2(n16592), .B1(n17861), .B2(n16591), .ZN(
        n12481) );
  NOR2_X1 U15734 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18943) );
  INV_X1 U15735 ( .A(n18943), .ZN(n18983) );
  INV_X1 U15736 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18920) );
  NAND2_X1 U15737 ( .A1(n18819), .A2(n18920), .ZN(n16692) );
  NAND2_X1 U15738 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17829) );
  NAND2_X1 U15739 ( .A1(n17030), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17939) );
  INV_X1 U15740 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17895) );
  NAND3_X1 U15741 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17856) );
  INV_X1 U15742 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17634) );
  NAND2_X1 U15743 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16575), .ZN(
        n12474) );
  INV_X1 U15744 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21196) );
  NAND3_X2 U15745 ( .A1(n18943), .A2(n18819), .A3(n12475), .ZN(n18317) );
  NOR2_X1 U15746 ( .A1(n21196), .A2(n18317), .ZN(n16586) );
  NOR2_X1 U15747 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18920), .ZN(
        n18941) );
  INV_X1 U15748 ( .A(n18941), .ZN(n18930) );
  OAI221_X1 U15749 ( .B1(n18928), .B2(P3_STATE2_REG_2__SCAN_IN), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n18819), .A(n18930), .ZN(n18333) );
  INV_X1 U15750 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18971) );
  NOR3_X1 U15751 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18971), .ZN(n18394) );
  NAND2_X2 U15752 ( .A1(n18626), .A2(n18394), .ZN(n18364) );
  INV_X1 U15753 ( .A(n17843), .ZN(n17794) );
  OR2_X1 U15754 ( .A1(n12476), .A2(n17794), .ZN(n16558) );
  INV_X1 U15755 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16736) );
  XOR2_X1 U15756 ( .A(n16736), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12478) );
  NOR2_X1 U15757 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17700), .ZN(
        n16576) );
  NAND2_X1 U15758 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16578), .ZN(
        n16717) );
  AOI22_X1 U15759 ( .A1(n18705), .A2(n12476), .B1(n17827), .B2(n16717), .ZN(
        n12477) );
  NAND2_X1 U15760 ( .A1(n12477), .A2(n17993), .ZN(n16577) );
  NOR2_X1 U15761 ( .A1(n16576), .A2(n16577), .ZN(n16557) );
  OAI22_X1 U15762 ( .A1(n16558), .A2(n12478), .B1(n16557), .B2(n16736), .ZN(
        n12479) );
  AOI211_X1 U15763 ( .C1(n17846), .C2(n10080), .A(n16586), .B(n12479), .ZN(
        n12480) );
  XNOR2_X1 U15764 ( .A(n14419), .B(n12484), .ZN(n14620) );
  NAND2_X1 U15765 ( .A1(n13010), .A2(n12496), .ZN(n13179) );
  OAI21_X1 U15766 ( .B1(n16015), .B2(n12485), .A(n13179), .ZN(n12486) );
  INV_X1 U15767 ( .A(n12486), .ZN(n12487) );
  OR2_X1 U15768 ( .A1(n13276), .A2(n12487), .ZN(n12491) );
  INV_X1 U15769 ( .A(n12488), .ZN(n12489) );
  NAND3_X1 U15770 ( .A1(n12489), .A2(n13064), .A3(n20972), .ZN(n12490) );
  AND2_X1 U15771 ( .A1(n10412), .A2(n12492), .ZN(n12495) );
  INV_X1 U15772 ( .A(n13353), .ZN(n20342) );
  NOR2_X1 U15773 ( .A1(n12513), .A2(n20042), .ZN(n12493) );
  NAND2_X1 U15774 ( .A1(n13350), .A2(n12496), .ZN(n12497) );
  NAND2_X1 U15775 ( .A1(n13009), .A2(n13353), .ZN(n13365) );
  INV_X1 U15776 ( .A(n14615), .ZN(n12499) );
  NAND2_X1 U15777 ( .A1(n14620), .A2(n12499), .ZN(n12521) );
  NOR4_X1 U15778 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12503) );
  NOR4_X1 U15779 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12502) );
  NOR4_X1 U15780 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12501) );
  NOR4_X1 U15781 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12500) );
  AND4_X1 U15782 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12509) );
  NOR4_X1 U15783 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12507) );
  NOR4_X1 U15784 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12506) );
  NOR4_X1 U15785 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12505) );
  INV_X1 U15786 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12504) );
  AND4_X1 U15787 ( .A1(n12507), .A2(n12506), .A3(n12505), .A4(n12504), .ZN(
        n12508) );
  NAND2_X1 U15788 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  NOR2_X1 U15789 ( .A1(n13003), .A2(n20271), .ZN(n12511) );
  NAND2_X1 U15790 ( .A1(n14600), .A2(n12511), .ZN(n14602) );
  AOI22_X1 U15791 ( .A1(n14610), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14609), .ZN(n12512) );
  INV_X1 U15792 ( .A(n12512), .ZN(n12519) );
  NOR3_X4 U15793 ( .A1(n14609), .A2(n20342), .A3(n12513), .ZN(n14612) );
  INV_X1 U15794 ( .A(DATAI_14_), .ZN(n12515) );
  NAND2_X1 U15795 ( .A1(n20270), .A2(BUF1_REG_14__SCAN_IN), .ZN(n12514) );
  OAI21_X1 U15796 ( .B1(n20270), .B2(n12515), .A(n12514), .ZN(n20202) );
  NOR3_X1 U15797 ( .A1(n14609), .A2(n20270), .A3(n13003), .ZN(n12516) );
  AOI22_X1 U15798 ( .A1(n14612), .A2(n20202), .B1(n14611), .B2(DATAI_30_), 
        .ZN(n12517) );
  INV_X1 U15799 ( .A(n12517), .ZN(n12518) );
  NAND2_X1 U15800 ( .A1(n12521), .A2(n12520), .ZN(P1_U2874) );
  NAND2_X2 U15801 ( .A1(n12525), .A2(n12524), .ZN(n13369) );
  INV_X1 U15802 ( .A(n16502), .ZN(n12560) );
  INV_X1 U15803 ( .A(n12529), .ZN(n12532) );
  INV_X1 U15804 ( .A(n12530), .ZN(n12531) );
  INV_X1 U15805 ( .A(n12538), .ZN(n12533) );
  NOR2_X1 U15806 ( .A1(n12528), .A2(n12533), .ZN(n12543) );
  INV_X1 U15807 ( .A(n12536), .ZN(n12534) );
  INV_X1 U15808 ( .A(n12619), .ZN(n12535) );
  AOI21_X1 U15809 ( .B1(n12535), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n15191), .ZN(n12550) );
  INV_X1 U15810 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12541) );
  OR2_X1 U15811 ( .A1(n12537), .A2(n19150), .ZN(n12559) );
  INV_X1 U15812 ( .A(n12559), .ZN(n12539) );
  NAND3_X1 U15813 ( .A1(n16502), .A2(n12539), .A3(n12566), .ZN(n12620) );
  INV_X1 U15814 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12540) );
  INV_X1 U15815 ( .A(n12542), .ZN(n12549) );
  INV_X1 U15816 ( .A(n12616), .ZN(n19573) );
  INV_X1 U15817 ( .A(n12544), .ZN(n12545) );
  NAND4_X1 U15818 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        n12558) );
  INV_X1 U15819 ( .A(n16502), .ZN(n12552) );
  INV_X1 U15820 ( .A(n12572), .ZN(n12551) );
  INV_X1 U15821 ( .A(n12537), .ZN(n12555) );
  XNOR2_X2 U15822 ( .A(n12555), .B(n12554), .ZN(n13119) );
  INV_X1 U15823 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15920) );
  NOR2_X1 U15824 ( .A1(n12615), .A2(n15920), .ZN(n12557) );
  NOR2_X1 U15825 ( .A1(n12558), .A2(n12557), .ZN(n12582) );
  INV_X1 U15826 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12564) );
  INV_X1 U15827 ( .A(n12633), .ZN(n12563) );
  NOR2_X2 U15828 ( .A1(n12561), .A2(n16502), .ZN(n19366) );
  NAND2_X1 U15829 ( .A1(n19366), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12562) );
  OAI21_X1 U15830 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n12571) );
  INV_X1 U15831 ( .A(n19150), .ZN(n12565) );
  OR2_X2 U15832 ( .A1(n12566), .A2(n12565), .ZN(n12574) );
  NOR2_X2 U15833 ( .A1(n12574), .A2(n12567), .ZN(n12632) );
  INV_X1 U15834 ( .A(n12632), .ZN(n12569) );
  INV_X1 U15835 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15181) );
  NOR2_X1 U15836 ( .A1(n12571), .A2(n12570), .ZN(n12581) );
  NOR2_X2 U15837 ( .A1(n12574), .A2(n16502), .ZN(n12578) );
  INV_X1 U15838 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12576) );
  NAND2_X1 U15839 ( .A1(n13119), .A2(n16502), .ZN(n12573) );
  NOR2_X2 U15840 ( .A1(n12574), .A2(n12573), .ZN(n12625) );
  NAND2_X1 U15841 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12575) );
  OAI21_X1 U15842 ( .B1(n12576), .B2(n19785), .A(n12575), .ZN(n12577) );
  AOI21_X1 U15843 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n19411), .A(
        n12577), .ZN(n12580) );
  AOI22_X1 U15844 ( .A1(n12630), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12631), .ZN(n12579) );
  NAND4_X1 U15845 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12585) );
  OR2_X1 U15846 ( .A1(n12832), .A2(n15910), .ZN(n13233) );
  NOR2_X1 U15847 ( .A1(n13233), .A2(n12831), .ZN(n12836) );
  INV_X1 U15848 ( .A(n12837), .ZN(n12583) );
  OR2_X1 U15849 ( .A1(n12836), .A2(n12583), .ZN(n12584) );
  NAND2_X1 U15850 ( .A1(n12585), .A2(n12584), .ZN(n12650) );
  INV_X1 U15851 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U15852 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12586) );
  INV_X1 U15853 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12589) );
  INV_X1 U15854 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12588) );
  OAI22_X1 U15855 ( .A1(n12589), .A2(n12619), .B1(n12620), .B2(n12588), .ZN(
        n12590) );
  INV_X1 U15856 ( .A(n12590), .ZN(n12595) );
  INV_X1 U15857 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12592) );
  INV_X1 U15858 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12591) );
  INV_X1 U15859 ( .A(n12593), .ZN(n12594) );
  NOR2_X1 U15860 ( .A1(n12597), .A2(n12596), .ZN(n12607) );
  INV_X1 U15861 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12598) );
  INV_X1 U15862 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U15863 ( .A1(n12630), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n12631), .ZN(n12605) );
  NAND2_X1 U15864 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12603) );
  NAND2_X1 U15865 ( .A1(n19366), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12602) );
  NAND2_X1 U15866 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12601) );
  NAND4_X1 U15867 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12608) );
  NAND2_X1 U15868 ( .A1(n12608), .A2(n15910), .ZN(n12611) );
  NAND2_X1 U15869 ( .A1(n12609), .A2(n15191), .ZN(n12610) );
  INV_X1 U15870 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15276) );
  INV_X1 U15871 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12613) );
  OAI22_X1 U15872 ( .A1(n15276), .A2(n12685), .B1(n19785), .B2(n12613), .ZN(
        n12614) );
  AOI21_X1 U15873 ( .B1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n19411), .A(
        n12614), .ZN(n12642) );
  INV_X1 U15874 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12628) );
  INV_X1 U15875 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12618) );
  INV_X1 U15876 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12617) );
  OAI22_X1 U15877 ( .A1(n12618), .A2(n19442), .B1(n12616), .B2(n12617), .ZN(
        n12624) );
  INV_X1 U15878 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12622) );
  INV_X1 U15879 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12621) );
  OAI22_X1 U15880 ( .A1(n12622), .A2(n12619), .B1(n12620), .B2(n12621), .ZN(
        n12623) );
  NOR2_X1 U15881 ( .A1(n12624), .A2(n12623), .ZN(n12627) );
  NAND2_X1 U15882 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12626) );
  OAI211_X1 U15883 ( .C1(n12615), .C2(n12628), .A(n12627), .B(n12626), .ZN(
        n12629) );
  INV_X1 U15884 ( .A(n12629), .ZN(n12641) );
  AOI22_X1 U15885 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12630), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15886 ( .A1(n19366), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12638) );
  NAND2_X1 U15887 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12637) );
  NAND2_X1 U15888 ( .A1(n12633), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12636) );
  AOI22_X1 U15889 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19636), .B1(
        n12634), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12635) );
  NAND4_X1 U15890 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12645) );
  NAND2_X1 U15891 ( .A1(n15191), .A2(n12643), .ZN(n12644) );
  INV_X1 U15892 ( .A(n12702), .ZN(n12649) );
  NAND2_X1 U15893 ( .A1(n12667), .A2(n12647), .ZN(n12648) );
  NAND2_X1 U15894 ( .A1(n12649), .A2(n12648), .ZN(n19128) );
  NAND2_X1 U15895 ( .A1(n13652), .A2(n14364), .ZN(n12653) );
  INV_X1 U15896 ( .A(n12668), .ZN(n12651) );
  OAI21_X1 U15897 ( .B1(n12659), .B2(n12652), .A(n12651), .ZN(n13701) );
  OAI21_X1 U15898 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20006), .A(
        n12654), .ZN(n12897) );
  MUX2_X1 U15899 ( .A(n12832), .B(n12897), .S(n12929), .Z(n12656) );
  MUX2_X1 U15900 ( .A(n12656), .B(n12655), .S(n12883), .Z(n19144) );
  NOR2_X1 U15901 ( .A1(n19144), .A2(n13217), .ZN(n13231) );
  INV_X1 U15902 ( .A(n13231), .ZN(n13169) );
  NAND3_X1 U15903 ( .A1(n12883), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15904 ( .A1(n12660), .A2(n12657), .ZN(n15056) );
  NOR2_X1 U15905 ( .A1(n13169), .A2(n15056), .ZN(n12658) );
  NAND2_X1 U15906 ( .A1(n13169), .A2(n15056), .ZN(n13168) );
  OAI21_X1 U15907 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12658), .A(
        n13168), .ZN(n13247) );
  INV_X1 U15908 ( .A(n12659), .ZN(n12663) );
  NAND2_X1 U15909 ( .A1(n12661), .A2(n12660), .ZN(n12662) );
  NAND2_X1 U15910 ( .A1(n12663), .A2(n12662), .ZN(n13842) );
  XNOR2_X1 U15911 ( .A(n13842), .B(n21237), .ZN(n13246) );
  OR2_X1 U15912 ( .A1(n13247), .A2(n13246), .ZN(n13249) );
  INV_X1 U15913 ( .A(n13842), .ZN(n12664) );
  NAND2_X1 U15914 ( .A1(n12664), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12665) );
  NAND2_X1 U15915 ( .A1(n13249), .A2(n12665), .ZN(n13656) );
  INV_X1 U15916 ( .A(n13656), .ZN(n12666) );
  OAI21_X1 U15917 ( .B1(n12669), .B2(n12668), .A(n12667), .ZN(n13818) );
  XNOR2_X1 U15918 ( .A(n13818), .B(n13996), .ZN(n13718) );
  NAND2_X1 U15919 ( .A1(n12670), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12671) );
  NAND2_X1 U15920 ( .A1(n12672), .A2(n12671), .ZN(n13968) );
  AOI22_X1 U15921 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12632), .B1(
        n12633), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12679) );
  INV_X1 U15922 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15102) );
  INV_X1 U15923 ( .A(n12634), .ZN(n12674) );
  INV_X1 U15924 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12673) );
  AOI21_X1 U15925 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n19366), .A(
        n12675), .ZN(n12678) );
  INV_X1 U15926 ( .A(n19785), .ZN(n19788) );
  AOI22_X1 U15927 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12625), .B1(
        n19788), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12677) );
  NAND2_X1 U15928 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12676) );
  INV_X1 U15929 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12681) );
  INV_X1 U15930 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12680) );
  OAI22_X1 U15931 ( .A1(n12681), .A2(n19442), .B1(n12616), .B2(n12680), .ZN(
        n12684) );
  INV_X1 U15932 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12682) );
  INV_X1 U15933 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15113) );
  OAI22_X1 U15934 ( .A1(n12682), .A2(n12619), .B1(n12620), .B2(n15113), .ZN(
        n12683) );
  NOR2_X1 U15935 ( .A1(n12684), .A2(n12683), .ZN(n12687) );
  NAND2_X1 U15936 ( .A1(n19721), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12686) );
  OAI211_X1 U15937 ( .C1(n12615), .C2(n15100), .A(n12687), .B(n12686), .ZN(
        n12688) );
  INV_X1 U15938 ( .A(n12688), .ZN(n12693) );
  INV_X1 U15939 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19351) );
  INV_X1 U15940 ( .A(n12630), .ZN(n12690) );
  INV_X1 U15941 ( .A(n19411), .ZN(n19405) );
  OAI22_X1 U15942 ( .A1(n19351), .A2(n12690), .B1(n19405), .B2(n12689), .ZN(
        n12691) );
  INV_X1 U15943 ( .A(n12691), .ZN(n12692) );
  NAND3_X1 U15944 ( .A1(n10297), .A2(n12693), .A3(n12692), .ZN(n12696) );
  NAND2_X1 U15945 ( .A1(n12694), .A2(n15191), .ZN(n12695) );
  NOR2_X2 U15946 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  INV_X1 U15947 ( .A(n12707), .ZN(n12700) );
  OAI21_X1 U15948 ( .B1(n12702), .B2(n12701), .A(n12700), .ZN(n19112) );
  XNOR2_X1 U15949 ( .A(n12703), .B(n13966), .ZN(n13969) );
  NAND2_X1 U15950 ( .A1(n12703), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12704) );
  INV_X1 U15951 ( .A(n12705), .ZN(n12706) );
  XNOR2_X1 U15952 ( .A(n12707), .B(n12706), .ZN(n19103) );
  INV_X1 U15953 ( .A(n19103), .ZN(n12708) );
  NAND2_X1 U15954 ( .A1(n12708), .A2(n14036), .ZN(n14029) );
  NOR2_X1 U15955 ( .A1(n12710), .A2(n12709), .ZN(n12711) );
  NOR2_X1 U15956 ( .A1(n12714), .A2(n12711), .ZN(n13835) );
  NAND2_X1 U15957 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12859) );
  INV_X1 U15958 ( .A(n12859), .ZN(n12712) );
  NAND2_X1 U15959 ( .A1(n13835), .A2(n12712), .ZN(n16403) );
  AOI21_X1 U15960 ( .B1(n13835), .B2(n12646), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16404) );
  AND2_X1 U15961 ( .A1(n12883), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12713) );
  XNOR2_X1 U15962 ( .A(n12714), .B(n12713), .ZN(n19092) );
  NAND2_X1 U15963 ( .A1(n19092), .A2(n12646), .ZN(n12715) );
  NAND2_X1 U15964 ( .A1(n12715), .A2(n21159), .ZN(n15605) );
  NAND3_X1 U15965 ( .A1(n12717), .A2(n12883), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n12716) );
  OAI211_X1 U15966 ( .C1(n12717), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12794), .B(
        n12716), .ZN(n19079) );
  OR2_X1 U15967 ( .A1(n19079), .A2(n14364), .ZN(n12719) );
  NAND2_X1 U15968 ( .A1(n12719), .A2(n12718), .ZN(n15831) );
  INV_X1 U15969 ( .A(n12720), .ZN(n12721) );
  AND3_X1 U15970 ( .A1(n12883), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n12721), .ZN(
        n12722) );
  NOR2_X1 U15971 ( .A1(n12723), .A2(n12722), .ZN(n19071) );
  AOI21_X1 U15972 ( .B1(n19071), .B2(n12646), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15814) );
  INV_X1 U15973 ( .A(n15814), .ZN(n12724) );
  NAND2_X1 U15974 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12725) );
  OR2_X1 U15975 ( .A1(n19079), .A2(n12725), .ZN(n15830) );
  AND2_X1 U15976 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12726) );
  NAND2_X1 U15977 ( .A1(n19092), .A2(n12726), .ZN(n15828) );
  NAND2_X1 U15978 ( .A1(n15830), .A2(n15828), .ZN(n15810) );
  INV_X1 U15979 ( .A(n19071), .ZN(n12728) );
  NAND2_X1 U15980 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12727) );
  NOR2_X1 U15981 ( .A1(n12728), .A2(n12727), .ZN(n15813) );
  NOR2_X1 U15982 ( .A1(n15810), .A2(n15813), .ZN(n12729) );
  INV_X1 U15983 ( .A(n12730), .ZN(n12731) );
  OR2_X1 U15984 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  NAND2_X1 U15985 ( .A1(n12763), .A2(n12733), .ZN(n13805) );
  NOR2_X1 U15986 ( .A1(n12735), .A2(n12734), .ZN(n16374) );
  NAND2_X1 U15987 ( .A1(n12735), .A2(n12734), .ZN(n16373) );
  AND3_X1 U15988 ( .A1(n9895), .A2(n12883), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n12736) );
  OR2_X1 U15989 ( .A1(n12737), .A2(n12736), .ZN(n15006) );
  OAI21_X1 U15990 ( .B1(n15006), .B2(n14364), .A(n10262), .ZN(n15532) );
  NOR2_X1 U15991 ( .A1(n12741), .A2(n12738), .ZN(n12739) );
  OR2_X1 U15992 ( .A1(n12744), .A2(n12739), .ZN(n19018) );
  INV_X1 U15993 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15730) );
  OAI21_X1 U15994 ( .B1(n19018), .B2(n14364), .A(n15730), .ZN(n15559) );
  AND2_X1 U15995 ( .A1(n12751), .A2(n12740), .ZN(n12742) );
  OR2_X1 U15996 ( .A1(n12742), .A2(n12741), .ZN(n15033) );
  OAI21_X1 U15997 ( .B1(n15033), .B2(n14364), .A(n15740), .ZN(n15569) );
  AND2_X1 U15998 ( .A1(n15559), .A2(n15569), .ZN(n15545) );
  NAND2_X1 U15999 ( .A1(n12883), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12743) );
  OAI211_X1 U16000 ( .C1(n12744), .C2(n12743), .A(n12794), .B(n9895), .ZN(
        n15021) );
  OR2_X1 U16001 ( .A1(n15021), .A2(n14364), .ZN(n12767) );
  INV_X1 U16002 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U16003 ( .A1(n12767), .A2(n15718), .ZN(n15547) );
  AND2_X1 U16004 ( .A1(n15545), .A2(n15547), .ZN(n15530) );
  NAND3_X1 U16005 ( .A1(n12745), .A2(n12883), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n12746) );
  OAI211_X1 U16006 ( .C1(n12745), .C2(P2_EBX_REG_16__SCAN_IN), .A(n12794), .B(
        n12746), .ZN(n15046) );
  OR2_X1 U16007 ( .A1(n15046), .A2(n14364), .ZN(n12747) );
  XNOR2_X1 U16008 ( .A(n12747), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15526) );
  NAND2_X1 U16009 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  AND2_X1 U16010 ( .A1(n12751), .A2(n12750), .ZN(n19033) );
  NAND2_X1 U16011 ( .A1(n19033), .A2(n12646), .ZN(n12752) );
  INV_X1 U16012 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15757) );
  NAND2_X1 U16013 ( .A1(n12752), .A2(n15757), .ZN(n15583) );
  NAND2_X1 U16014 ( .A1(n12883), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12753) );
  MUX2_X1 U16015 ( .A(n12753), .B(n12883), .S(n9892), .Z(n12755) );
  INV_X1 U16016 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U16017 ( .A1(n9892), .A2(n12754), .ZN(n12758) );
  NAND2_X1 U16018 ( .A1(n12755), .A2(n12758), .ZN(n13851) );
  OR2_X1 U16019 ( .A1(n13851), .A2(n14364), .ZN(n12756) );
  NAND2_X1 U16020 ( .A1(n12756), .A2(n12774), .ZN(n16363) );
  AND2_X1 U16021 ( .A1(n12883), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U16022 ( .A1(n12758), .A2(n12757), .ZN(n12759) );
  NAND2_X1 U16023 ( .A1(n12759), .A2(n12745), .ZN(n19041) );
  OR2_X1 U16024 ( .A1(n19041), .A2(n14364), .ZN(n12760) );
  NAND2_X1 U16025 ( .A1(n12760), .A2(n15788), .ZN(n15780) );
  INV_X1 U16026 ( .A(n12761), .ZN(n12762) );
  XNOR2_X1 U16027 ( .A(n12763), .B(n12762), .ZN(n19060) );
  NAND2_X1 U16028 ( .A1(n19060), .A2(n12646), .ZN(n12764) );
  NAND2_X1 U16029 ( .A1(n12764), .A2(n15803), .ZN(n15523) );
  AND4_X1 U16030 ( .A1(n15583), .A2(n16363), .A3(n15780), .A4(n15523), .ZN(
        n12765) );
  NAND4_X1 U16031 ( .A1(n15532), .A2(n15530), .A3(n15526), .A4(n12765), .ZN(
        n12778) );
  NAND2_X1 U16032 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12766) );
  NOR2_X1 U16033 ( .A1(n15006), .A2(n12766), .ZN(n15531) );
  INV_X1 U16034 ( .A(n19018), .ZN(n12769) );
  AND2_X1 U16035 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12768) );
  NAND2_X1 U16036 ( .A1(n12769), .A2(n12768), .ZN(n15558) );
  INV_X1 U16037 ( .A(n15033), .ZN(n12771) );
  AND2_X1 U16038 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12770) );
  NAND2_X1 U16039 ( .A1(n12771), .A2(n12770), .ZN(n15568) );
  AND2_X1 U16040 ( .A1(n15558), .A2(n15568), .ZN(n15528) );
  AND2_X1 U16041 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12772) );
  NAND2_X1 U16042 ( .A1(n19033), .A2(n12772), .ZN(n15582) );
  OR3_X1 U16043 ( .A1(n15046), .A2(n14364), .A3(n15573), .ZN(n15584) );
  NAND2_X1 U16044 ( .A1(n15582), .A2(n15584), .ZN(n15527) );
  AND2_X1 U16045 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12773) );
  AND2_X1 U16046 ( .A1(n19060), .A2(n12773), .ZN(n15597) );
  OR3_X1 U16047 ( .A1(n13851), .A2(n14364), .A3(n12774), .ZN(n16362) );
  OR3_X1 U16048 ( .A1(n19041), .A2(n14364), .A3(n15788), .ZN(n15779) );
  NAND2_X1 U16049 ( .A1(n16362), .A2(n15779), .ZN(n15525) );
  NOR3_X1 U16050 ( .A1(n15527), .A2(n15597), .A3(n15525), .ZN(n12775) );
  NAND3_X1 U16051 ( .A1(n15548), .A2(n15528), .A3(n12775), .ZN(n12776) );
  NOR2_X1 U16052 ( .A1(n15531), .A2(n12776), .ZN(n12777) );
  NAND2_X1 U16053 ( .A1(n12779), .A2(n12646), .ZN(n12780) );
  NAND2_X1 U16054 ( .A1(n12780), .A2(n15689), .ZN(n15684) );
  NAND2_X1 U16055 ( .A1(n15683), .A2(n15684), .ZN(n12781) );
  OR2_X1 U16056 ( .A1(n12780), .A2(n15689), .ZN(n15685) );
  INV_X1 U16057 ( .A(n12782), .ZN(n12783) );
  XNOR2_X1 U16058 ( .A(n12779), .B(n12783), .ZN(n16315) );
  NAND2_X1 U16059 ( .A1(n16315), .A2(n12646), .ZN(n12784) );
  XNOR2_X1 U16060 ( .A(n12784), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15514) );
  OR2_X1 U16061 ( .A1(n12784), .A2(n15669), .ZN(n12785) );
  NAND3_X1 U16062 ( .A1(n12786), .A2(n12883), .A3(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n12787) );
  NAND2_X1 U16063 ( .A1(n12787), .A2(n12794), .ZN(n12788) );
  OR2_X1 U16064 ( .A1(n12788), .A2(n12791), .ZN(n14978) );
  NOR2_X1 U16065 ( .A1(n14978), .A2(n14364), .ZN(n12789) );
  AND2_X1 U16066 ( .A1(n12789), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15501) );
  INV_X1 U16067 ( .A(n12789), .ZN(n12790) );
  INV_X1 U16068 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15505) );
  NAND2_X1 U16069 ( .A1(n12790), .A2(n15505), .ZN(n15500) );
  NOR2_X1 U16070 ( .A1(n12791), .A2(n15360), .ZN(n12792) );
  NAND2_X1 U16071 ( .A1(n12883), .A2(n12792), .ZN(n12793) );
  AND2_X1 U16072 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U16073 ( .A1(n16294), .A2(n12795), .ZN(n14964) );
  OR2_X1 U16074 ( .A1(n14964), .A2(n14364), .ZN(n12796) );
  NAND2_X1 U16075 ( .A1(n12796), .A2(n14262), .ZN(n15488) );
  INV_X1 U16076 ( .A(n12797), .ZN(n12799) );
  NAND2_X1 U16077 ( .A1(n12799), .A2(n12798), .ZN(n12800) );
  NAND2_X1 U16078 ( .A1(n12809), .A2(n12800), .ZN(n14944) );
  NAND2_X1 U16079 ( .A1(n14338), .A2(n12806), .ZN(n12804) );
  INV_X1 U16080 ( .A(n12801), .ZN(n12802) );
  NAND2_X1 U16081 ( .A1(n12802), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12803) );
  INV_X1 U16082 ( .A(n14341), .ZN(n12805) );
  NAND2_X1 U16083 ( .A1(n10309), .A2(n12805), .ZN(n15480) );
  NOR2_X1 U16084 ( .A1(n15480), .A2(n15481), .ZN(n15479) );
  AOI21_X1 U16085 ( .B1(n14338), .B2(n14342), .A(n12806), .ZN(n12807) );
  NOR2_X1 U16086 ( .A1(n15479), .A2(n12807), .ZN(n12812) );
  NAND2_X1 U16087 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  NAND2_X1 U16088 ( .A1(n14345), .A2(n12810), .ZN(n14927) );
  XOR2_X1 U16089 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14340), .Z(
        n12811) );
  XNOR2_X1 U16090 ( .A(n12812), .B(n12811), .ZN(n12930) );
  INV_X1 U16091 ( .A(n12897), .ZN(n12900) );
  AOI21_X1 U16092 ( .B1(n12900), .B2(n12813), .A(n16521), .ZN(n12814) );
  INV_X1 U16093 ( .A(n12814), .ZN(n12816) );
  AND2_X1 U16094 ( .A1(n13100), .A2(n12815), .ZN(n16527) );
  AOI21_X1 U16095 ( .B1(n13913), .B2(n16527), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n20000) );
  MUX2_X1 U16096 ( .A(n12816), .B(n20000), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20012) );
  NOR2_X1 U16097 ( .A1(n12818), .A2(n15191), .ZN(n12826) );
  NAND2_X1 U16098 ( .A1(n12819), .A2(n12907), .ZN(n12894) );
  NAND2_X1 U16099 ( .A1(n12900), .A2(n12896), .ZN(n12820) );
  AND2_X1 U16100 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  NOR2_X1 U16101 ( .A1(n12894), .A2(n12822), .ZN(n12823) );
  OR2_X1 U16102 ( .A1(n12918), .A2(n12823), .ZN(n20009) );
  AND2_X1 U16103 ( .A1(n15191), .A2(n11435), .ZN(n12884) );
  INV_X1 U16104 ( .A(n12884), .ZN(n12824) );
  NAND2_X1 U16105 ( .A1(n11435), .A2(n13295), .ZN(n12827) );
  INV_X1 U16106 ( .A(n13052), .ZN(n12828) );
  NAND2_X1 U16107 ( .A1(n12930), .A2(n16414), .ZN(n12876) );
  NAND2_X1 U16108 ( .A1(n13233), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13232) );
  INV_X1 U16109 ( .A(n13232), .ZN(n12833) );
  XOR2_X1 U16110 ( .A(n12832), .B(n12831), .Z(n12834) );
  NAND2_X1 U16111 ( .A1(n12833), .A2(n12834), .ZN(n12835) );
  XNOR2_X1 U16112 ( .A(n12834), .B(n13232), .ZN(n13172) );
  NAND2_X1 U16113 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13172), .ZN(
        n13171) );
  NAND2_X1 U16114 ( .A1(n12835), .A2(n13171), .ZN(n12838) );
  XOR2_X1 U16115 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12838), .Z(
        n13245) );
  XOR2_X1 U16116 ( .A(n12837), .B(n12836), .Z(n13244) );
  NAND2_X1 U16117 ( .A1(n13245), .A2(n13244), .ZN(n13243) );
  NAND2_X1 U16118 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12838), .ZN(
        n12839) );
  NAND2_X1 U16119 ( .A1(n13243), .A2(n12839), .ZN(n12840) );
  XNOR2_X1 U16120 ( .A(n12840), .B(n16479), .ZN(n13653) );
  NAND2_X1 U16121 ( .A1(n13652), .A2(n13653), .ZN(n12842) );
  NAND2_X1 U16122 ( .A1(n12840), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12841) );
  AND2_X1 U16123 ( .A1(n12848), .A2(n13997), .ZN(n14002) );
  INV_X1 U16124 ( .A(n12846), .ZN(n12855) );
  NAND2_X1 U16125 ( .A1(n12847), .A2(n12846), .ZN(n12852) );
  NAND2_X1 U16126 ( .A1(n12853), .A2(n12854), .ZN(n12856) );
  NAND2_X1 U16127 ( .A1(n12856), .A2(n12855), .ZN(n12857) );
  XNOR2_X1 U16128 ( .A(n12860), .B(n14364), .ZN(n14026) );
  OAI21_X1 U16129 ( .B1(n12860), .B2(n14364), .A(n21138), .ZN(n12861) );
  NOR2_X1 U16130 ( .A1(n12734), .A2(n15803), .ZN(n16430) );
  AND2_X1 U16131 ( .A1(n16430), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16431) );
  NOR2_X1 U16132 ( .A1(n12718), .A2(n15818), .ZN(n15817) );
  AND2_X1 U16133 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15817), .ZN(
        n15796) );
  AND3_X1 U16134 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15698) );
  NAND2_X1 U16135 ( .A1(n15698), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15717) );
  INV_X1 U16136 ( .A(n15717), .ZN(n12863) );
  NAND2_X1 U16137 ( .A1(n15503), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14255) );
  INV_X1 U16138 ( .A(n14255), .ZN(n12864) );
  NAND2_X1 U16139 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15643) );
  OAI21_X1 U16140 ( .B1(n12865), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14354), .ZN(n12932) );
  NOR2_X2 U16141 ( .A1(n13052), .A2(n15910), .ZN(n16415) );
  NOR2_X1 U16142 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19969) );
  OR2_X1 U16143 ( .A1(n19971), .A2(n19969), .ZN(n19998) );
  NAND2_X1 U16144 ( .A1(n19998), .A2(n19237), .ZN(n12866) );
  INV_X1 U16145 ( .A(n13376), .ZN(n13072) );
  INV_X1 U16146 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n15893) );
  NAND2_X1 U16147 ( .A1(n15893), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12867) );
  NAND2_X1 U16148 ( .A1(n13072), .A2(n12867), .ZN(n13235) );
  NAND2_X1 U16149 ( .A1(n16460), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16150 ( .B1(n16429), .B2(n12868), .A(n12977), .ZN(n12872) );
  OAI21_X1 U16151 ( .B1(n14936), .B2(n12869), .A(n14912), .ZN(n15339) );
  AND2_X1 U16152 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12870) );
  NOR2_X1 U16153 ( .A1(n15339), .A2(n16393), .ZN(n12871) );
  AOI211_X1 U16154 ( .C1(n16420), .C2(n14930), .A(n12872), .B(n12871), .ZN(
        n12873) );
  NAND2_X1 U16155 ( .A1(n12876), .A2(n12875), .ZN(P2_U2986) );
  INV_X1 U16156 ( .A(n16521), .ZN(n12893) );
  MUX2_X1 U16157 ( .A(n12877), .B(n11458), .S(n15191), .Z(n12878) );
  NOR2_X1 U16158 ( .A1(n12878), .A2(n20023), .ZN(n12892) );
  NAND2_X1 U16159 ( .A1(n12879), .A2(n11458), .ZN(n12880) );
  NAND2_X1 U16160 ( .A1(n11613), .A2(n12880), .ZN(n12889) );
  NOR2_X1 U16161 ( .A1(n19337), .A2(n15910), .ZN(n12933) );
  OAI211_X1 U16162 ( .C1(n12933), .C2(n11435), .A(n13630), .B(n19355), .ZN(
        n12881) );
  NAND2_X1 U16163 ( .A1(n12881), .A2(n11458), .ZN(n12888) );
  INV_X1 U16164 ( .A(n12882), .ZN(n12887) );
  AND2_X1 U16165 ( .A1(n12883), .A2(n19347), .ZN(n12885) );
  OAI21_X1 U16166 ( .B1(n12886), .B2(n12885), .A(n12884), .ZN(n12937) );
  NAND4_X1 U16167 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12937), .ZN(
        n12935) );
  OR2_X1 U16168 ( .A1(n13087), .A2(n16521), .ZN(n12890) );
  NOR2_X1 U16169 ( .A1(n12877), .A2(n12890), .ZN(n12891) );
  OR2_X1 U16170 ( .A1(n12935), .A2(n12891), .ZN(n13090) );
  AOI21_X1 U16171 ( .B1(n12893), .B2(n12892), .A(n13090), .ZN(n12926) );
  NAND2_X1 U16172 ( .A1(n12894), .A2(n12929), .ZN(n12910) );
  NAND2_X1 U16173 ( .A1(n19239), .A2(n15910), .ZN(n12895) );
  MUX2_X1 U16174 ( .A(n12929), .B(n12895), .S(n12903), .Z(n12906) );
  INV_X1 U16175 ( .A(n12896), .ZN(n12898) );
  OAI21_X1 U16176 ( .B1(n12898), .B2(n12897), .A(n12911), .ZN(n12902) );
  OAI211_X1 U16177 ( .C1(n15910), .C2(n12900), .A(n20028), .B(n12899), .ZN(
        n12901) );
  OAI211_X1 U16178 ( .C1(n12904), .C2(n12903), .A(n12902), .B(n12901), .ZN(
        n12905) );
  NAND2_X1 U16179 ( .A1(n12906), .A2(n12905), .ZN(n12908) );
  NAND2_X1 U16180 ( .A1(n12908), .A2(n12907), .ZN(n12909) );
  NAND2_X1 U16181 ( .A1(n12910), .A2(n12909), .ZN(n12914) );
  NAND2_X1 U16182 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  NAND2_X1 U16183 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  MUX2_X1 U16184 ( .A(n12916), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19237), .Z(n12921) );
  INV_X1 U16185 ( .A(n19239), .ZN(n12917) );
  NAND2_X1 U16186 ( .A1(n12918), .A2(n12917), .ZN(n12919) );
  NAND2_X1 U16187 ( .A1(n16523), .A2(n15910), .ZN(n19235) );
  AOI21_X1 U16188 ( .B1(n12921), .B2(n12920), .A(n19337), .ZN(n12922) );
  NAND2_X1 U16189 ( .A1(n19235), .A2(n12922), .ZN(n12925) );
  INV_X1 U16190 ( .A(n19235), .ZN(n13089) );
  INV_X1 U16191 ( .A(n11458), .ZN(n12923) );
  INV_X1 U16192 ( .A(n13087), .ZN(n13050) );
  NAND3_X1 U16193 ( .A1(n13089), .A2(n12923), .A3(n13050), .ZN(n12924) );
  NAND4_X1 U16194 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12928) );
  NOR2_X1 U16195 ( .A1(n12818), .A2(n12929), .ZN(n20011) );
  NAND2_X1 U16196 ( .A1(n12930), .A2(n16475), .ZN(n12985) );
  INV_X1 U16197 ( .A(n12931), .ZN(n20010) );
  OR2_X1 U16198 ( .A1(n12932), .A2(n19318), .ZN(n12983) );
  INV_X1 U16199 ( .A(n12933), .ZN(n12934) );
  NAND2_X1 U16200 ( .A1(n12974), .A2(n16517), .ZN(n15750) );
  OR2_X1 U16201 ( .A1(n12936), .A2(n15191), .ZN(n13868) );
  NAND2_X1 U16202 ( .A1(n13868), .A2(n12937), .ZN(n12938) );
  NAND2_X1 U16203 ( .A1(n12938), .A2(n13630), .ZN(n12953) );
  OAI22_X1 U16204 ( .A1(n12939), .A2(n19337), .B1(n11458), .B2(n20028), .ZN(
        n12940) );
  INV_X1 U16205 ( .A(n12940), .ZN(n12950) );
  INV_X1 U16206 ( .A(n12941), .ZN(n12943) );
  NAND2_X1 U16207 ( .A1(n12943), .A2(n12942), .ZN(n12944) );
  NAND2_X1 U16208 ( .A1(n12944), .A2(n12939), .ZN(n12946) );
  NAND2_X1 U16209 ( .A1(n12946), .A2(n12945), .ZN(n12949) );
  NAND2_X1 U16210 ( .A1(n12948), .A2(n12947), .ZN(n13293) );
  AND4_X1 U16211 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n13293), .ZN(
        n12952) );
  NAND2_X1 U16212 ( .A1(n12953), .A2(n12952), .ZN(n16501) );
  INV_X1 U16213 ( .A(n15883), .ZN(n12954) );
  OR2_X1 U16214 ( .A1(n16501), .A2(n12954), .ZN(n12955) );
  NAND2_X1 U16215 ( .A1(n12974), .A2(n12955), .ZN(n15753) );
  INV_X1 U16216 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16479) );
  NOR3_X1 U16217 ( .A1(n16479), .A2(n13997), .A3(n13996), .ZN(n12956) );
  AND2_X1 U16218 ( .A1(n12956), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12957) );
  OR2_X1 U16219 ( .A1(n15864), .A2(n12957), .ZN(n12959) );
  INV_X1 U16220 ( .A(n15750), .ZN(n13239) );
  NOR2_X1 U16221 ( .A1(n13217), .A2(n13218), .ZN(n13257) );
  NOR2_X1 U16222 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13257), .ZN(
        n13241) );
  NOR2_X1 U16223 ( .A1(n15753), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13256) );
  INV_X1 U16224 ( .A(n12974), .ZN(n12958) );
  NAND2_X1 U16225 ( .A1(n12958), .A2(n19324), .ZN(n15863) );
  OAI21_X1 U16226 ( .B1(n15753), .B2(n13257), .A(n15863), .ZN(n13262) );
  AOI211_X1 U16227 ( .C1(n13239), .C2(n13241), .A(n13256), .B(n13262), .ZN(
        n16478) );
  NAND2_X1 U16228 ( .A1(n12959), .A2(n16478), .ZN(n16454) );
  NAND2_X1 U16229 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16461) );
  INV_X1 U16230 ( .A(n16461), .ZN(n12960) );
  NOR2_X1 U16231 ( .A1(n15864), .A2(n12960), .ZN(n12961) );
  NAND2_X1 U16232 ( .A1(n15851), .A2(n15864), .ZN(n15798) );
  NAND2_X1 U16233 ( .A1(n15798), .A2(n15643), .ZN(n12963) );
  NOR2_X1 U16234 ( .A1(n15669), .A2(n15689), .ZN(n15668) );
  INV_X1 U16235 ( .A(n15864), .ZN(n15736) );
  INV_X1 U16236 ( .A(n15715), .ZN(n12962) );
  NOR4_X1 U16237 ( .A1(n12962), .A2(n15718), .A3(n15730), .A4(n15717), .ZN(
        n12965) );
  OAI21_X1 U16238 ( .B1(n15864), .B2(n12965), .A(n15851), .ZN(n15707) );
  AOI21_X1 U16239 ( .B1(n10262), .B2(n15736), .A(n15707), .ZN(n15688) );
  OAI211_X1 U16240 ( .C1(n15864), .C2(n15668), .A(n15688), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15656) );
  NAND2_X1 U16241 ( .A1(n15656), .A2(n15798), .ZN(n15647) );
  NAND2_X1 U16242 ( .A1(n12963), .A2(n15647), .ZN(n15638) );
  INV_X1 U16243 ( .A(n15643), .ZN(n12966) );
  NAND2_X1 U16244 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13257), .ZN(
        n13238) );
  NAND4_X1 U16245 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(n16467), .ZN(n13957) );
  INV_X1 U16246 ( .A(n16462), .ZN(n12964) );
  NAND3_X1 U16247 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n12965), .A3(
        n15855), .ZN(n15690) );
  INV_X1 U16248 ( .A(n15690), .ZN(n15676) );
  NAND2_X1 U16249 ( .A1(n12966), .A2(n15644), .ZN(n15632) );
  NOR2_X1 U16250 ( .A1(n12967), .A2(n15481), .ZN(n15616) );
  NOR2_X1 U16251 ( .A1(n15632), .A2(n15616), .ZN(n12968) );
  OR2_X1 U16252 ( .A1(n15638), .A2(n12968), .ZN(n15622) );
  NAND2_X1 U16253 ( .A1(n16495), .A2(n15191), .ZN(n12969) );
  NAND2_X1 U16254 ( .A1(n12969), .A2(n15884), .ZN(n12970) );
  AND2_X1 U16255 ( .A1(n12972), .A2(n12971), .ZN(n16522) );
  INV_X1 U16256 ( .A(n16522), .ZN(n15878) );
  OAI21_X1 U16257 ( .B1(n15191), .B2(n16519), .A(n15878), .ZN(n12973) );
  AND2_X1 U16258 ( .A1(n14942), .A2(n12975), .ZN(n12976) );
  NOR2_X1 U16259 ( .A1(n9878), .A2(n12976), .ZN(n15417) );
  INV_X1 U16260 ( .A(n12977), .ZN(n12979) );
  NOR3_X1 U16261 ( .A1(n15632), .A2(n15616), .A3(n15481), .ZN(n12978) );
  AOI211_X1 U16262 ( .C1(n19310), .C2(n15417), .A(n12979), .B(n12978), .ZN(
        n12980) );
  OAI21_X1 U16263 ( .B1(n15339), .B2(n19312), .A(n12980), .ZN(n12981) );
  AOI21_X1 U16264 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15622), .A(
        n12981), .ZN(n12982) );
  NAND2_X1 U16265 ( .A1(n12985), .A2(n12984), .ZN(P2_U3018) );
  NOR2_X1 U16266 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .ZN(n12987) );
  NOR4_X1 U16267 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_BE_N_REG_3__SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12986) );
  NAND4_X1 U16268 ( .A1(n12987), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n12986), .ZN(n13000) );
  INV_X1 U16269 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20962) );
  NOR3_X1 U16270 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20962), .ZN(n12989) );
  NOR4_X1 U16271 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12988) );
  NAND4_X1 U16272 ( .A1(n20270), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12989), .A4(
        n12988), .ZN(U214) );
  NOR4_X1 U16273 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12993) );
  NOR4_X1 U16274 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12992) );
  NOR4_X1 U16275 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12991) );
  NOR4_X1 U16276 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12990) );
  NAND4_X1 U16277 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n12990), .ZN(
        n12998) );
  NOR4_X1 U16278 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12996) );
  NOR4_X1 U16279 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12995) );
  NOR4_X1 U16280 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12994) );
  NAND4_X1 U16281 ( .A1(n12996), .A2(n12995), .A3(n12994), .A4(n19911), .ZN(
        n12997) );
  NOR2_X1 U16282 ( .A1(n15399), .A2(n13000), .ZN(n16613) );
  NAND2_X1 U16283 ( .A1(n16613), .A2(U214), .ZN(U212) );
  AOI21_X1 U16284 ( .B1(n13309), .B2(n16016), .A(n16015), .ZN(n13001) );
  NAND2_X1 U16285 ( .A1(n13064), .A2(n13001), .ZN(n13008) );
  INV_X1 U16286 ( .A(n13002), .ZN(n13005) );
  NAND2_X1 U16287 ( .A1(n13003), .A2(n13280), .ZN(n13004) );
  AOI21_X1 U16288 ( .B1(n13190), .B2(n13005), .A(n13004), .ZN(n13006) );
  OR2_X1 U16289 ( .A1(n13276), .A2(n13006), .ZN(n13007) );
  MUX2_X1 U16290 ( .A(n13008), .B(n13007), .S(n20298), .Z(n13016) );
  OR2_X1 U16291 ( .A1(n13009), .A2(n20287), .ZN(n13030) );
  INV_X1 U16292 ( .A(n13030), .ZN(n13014) );
  AND2_X1 U16293 ( .A1(n13010), .A2(n13018), .ZN(n13013) );
  AND2_X1 U16294 ( .A1(n13030), .A2(n13280), .ZN(n13011) );
  NAND2_X1 U16295 ( .A1(n13012), .A2(n13011), .ZN(n13023) );
  OAI21_X1 U16296 ( .B1(n13065), .B2(n13013), .A(n13023), .ZN(n13195) );
  AOI21_X1 U16297 ( .B1(n13276), .B2(n13014), .A(n13195), .ZN(n13015) );
  NAND2_X1 U16298 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  INV_X1 U16299 ( .A(n13018), .ZN(n13022) );
  NAND2_X1 U16300 ( .A1(n13193), .A2(n13019), .ZN(n13020) );
  OAI211_X1 U16301 ( .C1(n11162), .C2(n13668), .A(n13020), .B(n12049), .ZN(
        n13021) );
  AOI21_X1 U16302 ( .B1(n13022), .B2(n10456), .A(n13021), .ZN(n13025) );
  NAND3_X1 U16303 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(n13177) );
  INV_X1 U16304 ( .A(n13026), .ZN(n13027) );
  NOR2_X1 U16305 ( .A1(n13177), .A2(n13027), .ZN(n13028) );
  NOR2_X1 U16306 ( .A1(n13041), .A2(n13028), .ZN(n13038) );
  INV_X1 U16307 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20245) );
  NAND2_X1 U16308 ( .A1(n13038), .A2(n20245), .ZN(n13338) );
  NAND2_X1 U16309 ( .A1(n20252), .A2(n13041), .ZN(n13330) );
  NAND2_X1 U16310 ( .A1(n13338), .A2(n13330), .ZN(n20246) );
  INV_X1 U16311 ( .A(n20246), .ZN(n14212) );
  INV_X1 U16312 ( .A(n13189), .ZN(n13061) );
  NAND2_X1 U16313 ( .A1(n14878), .A2(n20245), .ZN(n13340) );
  AOI21_X1 U16314 ( .B1(n14212), .B2(n13340), .A(n20249), .ZN(n13048) );
  NOR2_X1 U16315 ( .A1(n13031), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13392) );
  INV_X1 U16316 ( .A(n13032), .ZN(n13391) );
  INV_X1 U16317 ( .A(n13039), .ZN(n13035) );
  AND2_X1 U16318 ( .A1(n13033), .A2(n13179), .ZN(n13062) );
  OAI211_X1 U16319 ( .C1(n10412), .C2(n13035), .A(n13034), .B(n13062), .ZN(
        n13036) );
  INV_X1 U16320 ( .A(n13036), .ZN(n13037) );
  NOR3_X1 U16321 ( .A1(n13392), .A2(n13391), .A3(n20250), .ZN(n13047) );
  NAND2_X1 U16322 ( .A1(n13065), .A2(n13309), .ZN(n15965) );
  NOR2_X1 U16323 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13332), .ZN(
        n13600) );
  NOR3_X1 U16324 ( .A1(n14856), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13600), .ZN(n13046) );
  AOI22_X1 U16325 ( .A1(n12020), .A2(n20287), .B1(n13039), .B2(n10412), .ZN(
        n13040) );
  OAI21_X1 U16326 ( .B1(n13043), .B2(n13349), .A(n13042), .ZN(n13671) );
  INV_X1 U16327 ( .A(n13671), .ZN(n13044) );
  NAND2_X1 U16328 ( .A1(n20221), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13390) );
  OAI21_X1 U16329 ( .B1(n20254), .B2(n13044), .A(n13390), .ZN(n13045) );
  OR4_X1 U16330 ( .A1(n13048), .A2(n13047), .A3(n13046), .A4(n13045), .ZN(
        P1_U3030) );
  OR2_X1 U16331 ( .A1(n11613), .A2(n16553), .ZN(n19234) );
  OR2_X1 U16332 ( .A1(n16521), .A2(n19234), .ZN(n15060) );
  INV_X1 U16333 ( .A(n15060), .ZN(n19157) );
  INV_X1 U16334 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20038) );
  OAI211_X1 U16335 ( .C1(n19157), .C2(n20038), .A(n18992), .B(n13079), .ZN(
        P2_U2814) );
  NOR2_X1 U16336 ( .A1(n20019), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13049)
         );
  INV_X1 U16337 ( .A(n12939), .ZN(n20030) );
  AOI22_X1 U16338 ( .A1(n13049), .A2(n18992), .B1(n20019), .B2(n20030), .ZN(
        P2_U3612) );
  INV_X1 U16339 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n16020) );
  AND2_X1 U16340 ( .A1(n12939), .A2(n20026), .ZN(n13091) );
  NOR2_X1 U16341 ( .A1(n13091), .A2(n13050), .ZN(n13051) );
  AND2_X1 U16342 ( .A1(n13092), .A2(n13051), .ZN(n16531) );
  NOR2_X1 U16343 ( .A1(n16531), .A2(n16553), .ZN(n20015) );
  OAI21_X1 U16344 ( .B1(n16020), .B2(n20015), .A(n13052), .ZN(P2_U2819) );
  INV_X1 U16345 ( .A(n20970), .ZN(n13054) );
  NAND2_X1 U16346 ( .A1(n20680), .A2(n20857), .ZN(n20045) );
  INV_X1 U16347 ( .A(n20045), .ZN(n14013) );
  OAI21_X1 U16348 ( .B1(n14013), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13054), 
        .ZN(n13053) );
  OAI21_X1 U16349 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(P1_U3487) );
  INV_X1 U16350 ( .A(n13308), .ZN(n13278) );
  AOI211_X1 U16351 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13056), .A(n14013), 
        .B(n13278), .ZN(n13057) );
  INV_X1 U16352 ( .A(n13057), .ZN(P1_U2801) );
  AOI21_X1 U16353 ( .B1(n13064), .B2(n13065), .A(n12020), .ZN(n13058) );
  AOI21_X1 U16354 ( .B1(n13276), .B2(n13663), .A(n13058), .ZN(n20041) );
  NAND3_X1 U16355 ( .A1(n13663), .A2(n13059), .A3(n16016), .ZN(n13060) );
  NAND2_X1 U16356 ( .A1(n13060), .A2(n20972), .ZN(n20963) );
  AND2_X1 U16357 ( .A1(n20041), .A2(n20963), .ZN(n15986) );
  NOR2_X1 U16358 ( .A1(n15986), .A2(n20042), .ZN(n20050) );
  INV_X1 U16359 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21227) );
  OR2_X1 U16360 ( .A1(n13276), .A2(n13061), .ZN(n13070) );
  NAND2_X1 U16361 ( .A1(n13276), .A2(n12020), .ZN(n13069) );
  INV_X1 U16362 ( .A(n13062), .ZN(n13063) );
  NAND2_X1 U16363 ( .A1(n13276), .A2(n13063), .ZN(n13068) );
  INV_X1 U16364 ( .A(n13064), .ZN(n13066) );
  NAND2_X1 U16365 ( .A1(n13066), .A2(n13065), .ZN(n13067) );
  NAND4_X1 U16366 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n15983) );
  NAND2_X1 U16367 ( .A1(n20050), .A2(n15983), .ZN(n13071) );
  OAI21_X1 U16368 ( .B1(n20050), .B2(n21227), .A(n13071), .ZN(P1_U3484) );
  NAND2_X1 U16369 ( .A1(n19347), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U16370 ( .A1(n13373), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19971), .B2(n20006), .ZN(n13073) );
  NAND2_X1 U16371 ( .A1(n15910), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13075) );
  AND4_X1 U16372 ( .A1(n11429), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13075), 
        .A4(n19825), .ZN(n13076) );
  INV_X1 U16373 ( .A(n16523), .ZN(n16518) );
  NAND2_X1 U16374 ( .A1(n16518), .A2(n16522), .ZN(n13093) );
  NAND2_X1 U16375 ( .A1(n13093), .A2(n15883), .ZN(n13077) );
  MUX2_X1 U16376 ( .A(n12655), .B(n19150), .S(n15395), .Z(n13078) );
  OAI21_X1 U16377 ( .B1(n20002), .B2(n15397), .A(n13078), .ZN(P2_U2887) );
  INV_X1 U16378 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13082) );
  NOR2_X1 U16379 ( .A1(n13079), .A2(n20023), .ZN(n13080) );
  AND2_X1 U16380 ( .A1(n13080), .A2(n15910), .ZN(n19303) );
  INV_X1 U16381 ( .A(n19303), .ZN(n13085) );
  AOI22_X1 U16382 ( .A1(n13789), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15399), .ZN(n19176) );
  INV_X1 U16383 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13081) );
  OAI222_X1 U16384 ( .A1(n13082), .A2(n13101), .B1(n13085), .B2(n19176), .C1(
        n13081), .C2(n19233), .ZN(P2_U2982) );
  INV_X1 U16385 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13084) );
  INV_X1 U16386 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16653) );
  INV_X1 U16387 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U16388 ( .A1(n13789), .A2(n16653), .B1(n18330), .B2(n15399), .ZN(
        n19166) );
  INV_X1 U16389 ( .A(n19166), .ZN(n19325) );
  INV_X1 U16390 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13083) );
  OAI222_X1 U16391 ( .A1(n13084), .A2(n13101), .B1(n13085), .B2(n19325), .C1(
        n19233), .C2(n13083), .ZN(P2_U2967) );
  INV_X1 U16392 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13086) );
  INV_X1 U16393 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19269) );
  OAI222_X1 U16394 ( .A1(n13086), .A2(n13101), .B1(n19233), .B2(n19269), .C1(
        n19325), .C2(n13085), .ZN(P2_U2952) );
  NOR2_X1 U16395 ( .A1(n11613), .A2(n13087), .ZN(n13088) );
  NAND2_X1 U16396 ( .A1(n13089), .A2(n13088), .ZN(n13095) );
  INV_X1 U16397 ( .A(n13090), .ZN(n13094) );
  AOI22_X1 U16398 ( .A1(n16523), .A2(n16517), .B1(n13092), .B2(n13091), .ZN(
        n13294) );
  NAND4_X1 U16399 ( .A1(n13095), .A2(n13094), .A3(n13294), .A4(n13093), .ZN(
        n16533) );
  NAND2_X1 U16400 ( .A1(n16533), .A2(n13295), .ZN(n13097) );
  INV_X1 U16401 ( .A(n19238), .ZN(n19999) );
  NOR2_X1 U16402 ( .A1(n19237), .A2(n19999), .ZN(n16538) );
  AOI22_X1 U16403 ( .A1(n19237), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(
        P2_FLUSH_REG_SCAN_IN), .B2(n16538), .ZN(n13096) );
  INV_X1 U16404 ( .A(n19966), .ZN(n13099) );
  INV_X1 U16405 ( .A(n19969), .ZN(n19963) );
  OR2_X1 U16406 ( .A1(n11613), .A2(n15910), .ZN(n16528) );
  OR4_X1 U16407 ( .A1(n19966), .A2(n16527), .A3(n19963), .A4(n16528), .ZN(
        n13098) );
  OAI21_X1 U16408 ( .B1(n13100), .B2(n13099), .A(n13098), .ZN(P2_U3595) );
  INV_X1 U16409 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19276) );
  NAND2_X1 U16410 ( .A1(n19306), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13104) );
  NAND2_X1 U16411 ( .A1(n15399), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13103) );
  INV_X1 U16412 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16633) );
  OR2_X1 U16413 ( .A1(n15399), .A2(n16633), .ZN(n13102) );
  NAND2_X1 U16414 ( .A1(n13103), .A2(n13102), .ZN(n19183) );
  NAND2_X1 U16415 ( .A1(n19303), .A2(n19183), .ZN(n13113) );
  OAI211_X1 U16416 ( .C1(n19276), .C2(n19233), .A(n13104), .B(n13113), .ZN(
        P2_U2979) );
  INV_X1 U16417 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19280) );
  NAND2_X1 U16418 ( .A1(n19306), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U16419 ( .A1(n15399), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13106) );
  INV_X1 U16420 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16635) );
  OR2_X1 U16421 ( .A1(n15399), .A2(n16635), .ZN(n13105) );
  NAND2_X1 U16422 ( .A1(n13106), .A2(n13105), .ZN(n19188) );
  NAND2_X1 U16423 ( .A1(n19303), .A2(n19188), .ZN(n13108) );
  OAI211_X1 U16424 ( .C1(n19280), .C2(n19233), .A(n13107), .B(n13108), .ZN(
        P2_U2977) );
  INV_X1 U16425 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19247) );
  NAND2_X1 U16426 ( .A1(n19306), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13109) );
  OAI211_X1 U16427 ( .C1(n19247), .C2(n19233), .A(n13109), .B(n13108), .ZN(
        P2_U2962) );
  INV_X1 U16428 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19284) );
  NAND2_X1 U16429 ( .A1(n19306), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U16430 ( .A1(n15399), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13111) );
  INV_X1 U16431 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16638) );
  OR2_X1 U16432 ( .A1(n15399), .A2(n16638), .ZN(n13110) );
  NAND2_X1 U16433 ( .A1(n13111), .A2(n13110), .ZN(n19193) );
  NAND2_X1 U16434 ( .A1(n19303), .A2(n19193), .ZN(n13115) );
  OAI211_X1 U16435 ( .C1(n19284), .C2(n19233), .A(n13112), .B(n13115), .ZN(
        P2_U2975) );
  INV_X1 U16436 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19244) );
  NAND2_X1 U16437 ( .A1(n19306), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13114) );
  OAI211_X1 U16438 ( .C1(n19244), .C2(n19233), .A(n13114), .B(n13113), .ZN(
        P2_U2964) );
  INV_X1 U16439 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19251) );
  NAND2_X1 U16440 ( .A1(n19306), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13116) );
  OAI211_X1 U16441 ( .C1(n19251), .C2(n19233), .A(n13116), .B(n13115), .ZN(
        P2_U2960) );
  NAND2_X1 U16442 ( .A1(n15216), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13272) );
  NAND2_X1 U16443 ( .A1(n13373), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13117) );
  XNOR2_X1 U16444 ( .A(n20006), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19469) );
  NAND2_X1 U16445 ( .A1(n19469), .A2(n19971), .ZN(n19406) );
  NAND2_X1 U16446 ( .A1(n13117), .A2(n19406), .ZN(n13118) );
  MUX2_X1 U16447 ( .A(n13121), .B(n13228), .S(n15395), .Z(n13122) );
  OAI21_X1 U16448 ( .B1(n19990), .B2(n15397), .A(n13122), .ZN(P2_U2886) );
  AOI22_X1 U16449 ( .A1(n19306), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13127) );
  INV_X1 U16450 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13123) );
  OR2_X1 U16451 ( .A1(n15399), .A2(n13123), .ZN(n13125) );
  NAND2_X1 U16452 ( .A1(n15399), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13124) );
  AND2_X1 U16453 ( .A1(n13125), .A2(n13124), .ZN(n19191) );
  INV_X1 U16454 ( .A(n19191), .ZN(n13126) );
  NAND2_X1 U16455 ( .A1(n19303), .A2(n13126), .ZN(n13166) );
  NAND2_X1 U16456 ( .A1(n13127), .A2(n13166), .ZN(P2_U2976) );
  AOI22_X1 U16457 ( .A1(n19306), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16458 ( .A1(n13789), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15399), .ZN(n19232) );
  INV_X1 U16459 ( .A(n19232), .ZN(n13128) );
  NAND2_X1 U16460 ( .A1(n19303), .A2(n13128), .ZN(n13142) );
  NAND2_X1 U16461 ( .A1(n13129), .A2(n13142), .ZN(P2_U2953) );
  AOI22_X1 U16462 ( .A1(n19306), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16463 ( .A1(n13789), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15399), .ZN(n19221) );
  INV_X1 U16464 ( .A(n19221), .ZN(n13130) );
  NAND2_X1 U16465 ( .A1(n19303), .A2(n13130), .ZN(n13139) );
  NAND2_X1 U16466 ( .A1(n13131), .A2(n13139), .ZN(P2_U2955) );
  AOI22_X1 U16467 ( .A1(n19306), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13136) );
  INV_X1 U16468 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13132) );
  OR2_X1 U16469 ( .A1(n15399), .A2(n13132), .ZN(n13134) );
  NAND2_X1 U16470 ( .A1(n15399), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13133) );
  AND2_X1 U16471 ( .A1(n13134), .A2(n13133), .ZN(n19186) );
  INV_X1 U16472 ( .A(n19186), .ZN(n13135) );
  NAND2_X1 U16473 ( .A1(n19303), .A2(n13135), .ZN(n13156) );
  NAND2_X1 U16474 ( .A1(n13136), .A2(n13156), .ZN(P2_U2978) );
  AOI22_X1 U16475 ( .A1(n19306), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16476 ( .A1(n13789), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15399), .ZN(n19343) );
  INV_X1 U16477 ( .A(n19343), .ZN(n19201) );
  NAND2_X1 U16478 ( .A1(n19303), .A2(n19201), .ZN(n13147) );
  NAND2_X1 U16479 ( .A1(n13137), .A2(n13147), .ZN(P2_U2957) );
  AOI22_X1 U16480 ( .A1(n19306), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13138) );
  OAI22_X1 U16481 ( .A1(n15399), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13789), .ZN(n19338) );
  INV_X1 U16482 ( .A(n19338), .ZN(n16325) );
  NAND2_X1 U16483 ( .A1(n19303), .A2(n16325), .ZN(n13160) );
  NAND2_X1 U16484 ( .A1(n13138), .A2(n13160), .ZN(P2_U2971) );
  AOI22_X1 U16485 ( .A1(n19306), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U16486 ( .A1(n13140), .A2(n13139), .ZN(P2_U2970) );
  AOI22_X1 U16487 ( .A1(n19306), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13141) );
  INV_X1 U16488 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16646) );
  INV_X1 U16489 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U16490 ( .A1(n13789), .A2(n16646), .B1(n21142), .B2(n15399), .ZN(
        n16332) );
  NAND2_X1 U16491 ( .A1(n19303), .A2(n16332), .ZN(n13162) );
  NAND2_X1 U16492 ( .A1(n13141), .A2(n13162), .ZN(P2_U2969) );
  AOI22_X1 U16493 ( .A1(n19306), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13143) );
  NAND2_X1 U16494 ( .A1(n13143), .A2(n13142), .ZN(P2_U2968) );
  AOI22_X1 U16495 ( .A1(n19306), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U16496 ( .A1(n13789), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15399), .ZN(n19357) );
  INV_X1 U16497 ( .A(n19357), .ZN(n13144) );
  NAND2_X1 U16498 ( .A1(n19303), .A2(n13144), .ZN(n13154) );
  NAND2_X1 U16499 ( .A1(n13145), .A2(n13154), .ZN(P2_U2974) );
  AOI22_X1 U16500 ( .A1(n19306), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13146) );
  INV_X1 U16501 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16641) );
  INV_X1 U16502 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18362) );
  AOI22_X1 U16503 ( .A1(n13789), .A2(n16641), .B1(n18362), .B2(n15399), .ZN(
        n19197) );
  NAND2_X1 U16504 ( .A1(n19303), .A2(n19197), .ZN(n13158) );
  NAND2_X1 U16505 ( .A1(n13146), .A2(n13158), .ZN(P2_U2973) );
  AOI22_X1 U16506 ( .A1(n19306), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13148) );
  NAND2_X1 U16507 ( .A1(n13148), .A2(n13147), .ZN(P2_U2972) );
  AOI22_X1 U16508 ( .A1(n19306), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13153) );
  INV_X1 U16509 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13149) );
  OR2_X1 U16510 ( .A1(n15399), .A2(n13149), .ZN(n13151) );
  NAND2_X1 U16511 ( .A1(n15399), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13150) );
  AND2_X1 U16512 ( .A1(n13151), .A2(n13150), .ZN(n19181) );
  INV_X1 U16513 ( .A(n19181), .ZN(n13152) );
  NAND2_X1 U16514 ( .A1(n19303), .A2(n13152), .ZN(n13164) );
  NAND2_X1 U16515 ( .A1(n13153), .A2(n13164), .ZN(P2_U2980) );
  AOI22_X1 U16516 ( .A1(n19306), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16517 ( .A1(n13155), .A2(n13154), .ZN(P2_U2959) );
  AOI22_X1 U16518 ( .A1(n19306), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19305), .ZN(n13157) );
  NAND2_X1 U16519 ( .A1(n13157), .A2(n13156), .ZN(P2_U2963) );
  AOI22_X1 U16520 ( .A1(n19306), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19305), .ZN(n13159) );
  NAND2_X1 U16521 ( .A1(n13159), .A2(n13158), .ZN(P2_U2958) );
  AOI22_X1 U16522 ( .A1(n19306), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19305), .ZN(n13161) );
  NAND2_X1 U16523 ( .A1(n13161), .A2(n13160), .ZN(P2_U2956) );
  AOI22_X1 U16524 ( .A1(n19306), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19305), .ZN(n13163) );
  NAND2_X1 U16525 ( .A1(n13163), .A2(n13162), .ZN(P2_U2954) );
  AOI22_X1 U16526 ( .A1(n19306), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19305), .ZN(n13165) );
  NAND2_X1 U16527 ( .A1(n13165), .A2(n13164), .ZN(P2_U2965) );
  AOI22_X1 U16528 ( .A1(n19306), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19305), .ZN(n13167) );
  NAND2_X1 U16529 ( .A1(n13167), .A2(n13166), .ZN(P2_U2961) );
  OAI21_X1 U16530 ( .B1(n15056), .B2(n13169), .A(n13168), .ZN(n13170) );
  XNOR2_X1 U16531 ( .A(n13170), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13225) );
  OAI21_X1 U16532 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13172), .A(
        n13171), .ZN(n13215) );
  OR2_X1 U16533 ( .A1(n19124), .A2(n11471), .ZN(n13216) );
  OAI21_X1 U16534 ( .B1(n16424), .B2(n13215), .A(n13216), .ZN(n13173) );
  AOI21_X1 U16535 ( .B1(n16414), .B2(n13225), .A(n13173), .ZN(n13175) );
  MUX2_X1 U16536 ( .A(n16419), .B(n16429), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13174) );
  OAI211_X1 U16537 ( .C1(n16393), .C2(n13228), .A(n13175), .B(n13174), .ZN(
        P2_U3013) );
  NOR2_X1 U16538 ( .A1(n13177), .A2(n20323), .ZN(n13178) );
  AND2_X1 U16539 ( .A1(n13178), .A2(n12488), .ZN(n13209) );
  OR2_X1 U16540 ( .A1(n20684), .A2(n13209), .ZN(n13186) );
  INV_X1 U16541 ( .A(n13179), .ZN(n13180) );
  OR2_X1 U16542 ( .A1(n13189), .A2(n13180), .ZN(n13499) );
  XNOR2_X1 U16543 ( .A(n14894), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13187) );
  XNOR2_X1 U16544 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13183) );
  INV_X1 U16545 ( .A(n10416), .ZN(n13182) );
  NAND2_X1 U16546 ( .A1(n13182), .A2(n13181), .ZN(n13495) );
  OAI22_X1 U16547 ( .A1(n15965), .A2(n13183), .B1(n13187), .B2(n13495), .ZN(
        n13184) );
  AOI21_X1 U16548 ( .B1(n13499), .B2(n13187), .A(n13184), .ZN(n13185) );
  NAND2_X1 U16549 ( .A1(n13186), .A2(n13185), .ZN(n13485) );
  NOR2_X1 U16550 ( .A1(n20857), .A2(n20245), .ZN(n14902) );
  AOI22_X1 U16551 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20249), .B2(n11269), .ZN(
        n14900) );
  INV_X1 U16552 ( .A(n13187), .ZN(n13188) );
  AOI222_X1 U16553 ( .A1(n13485), .A2(n13205), .B1(n14902), .B2(n14900), .C1(
        n13188), .C2(n15999), .ZN(n13202) );
  NAND2_X1 U16554 ( .A1(n13276), .A2(n13189), .ZN(n13348) );
  INV_X1 U16555 ( .A(n13348), .ZN(n13199) );
  INV_X1 U16556 ( .A(n13190), .ZN(n13191) );
  NAND2_X1 U16557 ( .A1(n15965), .A2(n13191), .ZN(n13192) );
  NAND3_X1 U16558 ( .A1(n13192), .A2(n15991), .A3(n20972), .ZN(n13197) );
  NOR2_X1 U16559 ( .A1(n13668), .A2(n13193), .ZN(n13194) );
  NOR2_X1 U16560 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  OAI21_X1 U16561 ( .B1(n13276), .B2(n13197), .A(n13196), .ZN(n13198) );
  NOR2_X1 U16562 ( .A1(n20968), .A2(n16289), .ZN(n13513) );
  AOI22_X1 U16563 ( .A1(n13507), .A2(n13201), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13513), .ZN(n13206) );
  OAI21_X1 U16564 ( .B1(n20694), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13206), 
        .ZN(n14909) );
  MUX2_X1 U16565 ( .A(n10314), .B(n13202), .S(n14909), .Z(n13203) );
  INV_X1 U16566 ( .A(n13203), .ZN(P1_U3472) );
  INV_X1 U16567 ( .A(n20448), .ZN(n20683) );
  OR2_X1 U16568 ( .A1(n10581), .A2(n20683), .ZN(n13204) );
  XNOR2_X1 U16569 ( .A(n13204), .B(n13208), .ZN(n20113) );
  INV_X1 U16570 ( .A(n13205), .ZN(n14908) );
  OR4_X1 U16571 ( .A1(n20113), .A2(n13206), .A3(n14908), .A4(n12488), .ZN(
        n13207) );
  OAI21_X1 U16572 ( .B1(n13208), .B2(n14909), .A(n13207), .ZN(P1_U3468) );
  INV_X1 U16573 ( .A(n13209), .ZN(n14898) );
  NOR2_X1 U16574 ( .A1(n10416), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13210) );
  AOI21_X1 U16575 ( .B1(n10573), .B2(n14898), .A(n13210), .ZN(n15968) );
  AOI22_X1 U16576 ( .A1(n15999), .A2(n10321), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(n20245), .ZN(n13211) );
  OAI21_X1 U16577 ( .B1(n15968), .B2(n14908), .A(n13211), .ZN(n13213) );
  OAI21_X1 U16578 ( .B1(n15965), .B2(n14908), .A(n14909), .ZN(n13212) );
  AOI22_X1 U16579 ( .A1(n13213), .A2(n14909), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13212), .ZN(n13214) );
  INV_X1 U16580 ( .A(n13214), .ZN(P1_U3474) );
  INV_X1 U16581 ( .A(n13215), .ZN(n13221) );
  OAI21_X1 U16582 ( .B1(n15863), .B2(n13218), .A(n13216), .ZN(n13220) );
  AOI211_X1 U16583 ( .C1(n13218), .C2(n13217), .A(n13257), .B(n15864), .ZN(
        n13219) );
  AOI211_X1 U16584 ( .C1(n15847), .C2(n13221), .A(n13220), .B(n13219), .ZN(
        n13227) );
  OAI21_X1 U16585 ( .B1(n13224), .B2(n13223), .A(n13222), .ZN(n19994) );
  AOI22_X1 U16586 ( .A1(n16475), .A2(n13225), .B1(n19310), .B2(n19994), .ZN(
        n13226) );
  OAI211_X1 U16587 ( .C1(n13228), .C2(n19312), .A(n13227), .B(n13226), .ZN(
        P2_U3045) );
  INV_X1 U16588 ( .A(n19144), .ZN(n13229) );
  NOR2_X1 U16589 ( .A1(n13229), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13230) );
  NOR2_X1 U16590 ( .A1(n13231), .A2(n13230), .ZN(n15862) );
  NOR2_X1 U16591 ( .A1(n19124), .A2(n19007), .ZN(n15861) );
  OAI21_X1 U16592 ( .B1(n13233), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13232), .ZN(n15859) );
  NOR2_X1 U16593 ( .A1(n16424), .A2(n15859), .ZN(n13234) );
  AOI211_X1 U16594 ( .C1(n15862), .C2(n16414), .A(n15861), .B(n13234), .ZN(
        n13237) );
  OAI21_X1 U16595 ( .B1(n16411), .B2(n13235), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13236) );
  OAI211_X1 U16596 ( .C1(n16393), .C2(n19150), .A(n13237), .B(n13236), .ZN(
        P2_U3014) );
  INV_X1 U16597 ( .A(n13238), .ZN(n13240) );
  OAI21_X1 U16598 ( .B1(n13241), .B2(n13240), .A(n13239), .ZN(n13242) );
  OAI21_X1 U16599 ( .B1(n12552), .B2(n19312), .A(n13242), .ZN(n13261) );
  OAI21_X1 U16600 ( .B1(n13245), .B2(n13244), .A(n13243), .ZN(n14248) );
  NAND2_X1 U16601 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  NAND2_X1 U16602 ( .A1(n13249), .A2(n13248), .ZN(n14247) );
  INV_X1 U16603 ( .A(n14247), .ZN(n13255) );
  NAND2_X1 U16604 ( .A1(n13251), .A2(n13250), .ZN(n13254) );
  INV_X1 U16605 ( .A(n13252), .ZN(n13253) );
  AND2_X1 U16606 ( .A1(n13254), .A2(n13253), .ZN(n19983) );
  INV_X1 U16607 ( .A(n19983), .ZN(n13460) );
  AOI22_X1 U16608 ( .A1(n16475), .A2(n13255), .B1(n19310), .B2(n13460), .ZN(
        n13259) );
  AOI22_X1 U16609 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n16460), .B1(n13257), 
        .B2(n13256), .ZN(n13258) );
  OAI211_X1 U16610 ( .C1(n19318), .C2(n14248), .A(n13259), .B(n13258), .ZN(
        n13260) );
  AOI211_X1 U16611 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13262), .A(
        n13261), .B(n13260), .ZN(n13263) );
  INV_X1 U16612 ( .A(n13263), .ZN(P2_U3044) );
  NAND2_X1 U16613 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19688) );
  NAND2_X1 U16614 ( .A1(n19688), .A2(n16505), .ZN(n13264) );
  NOR2_X1 U16615 ( .A1(n16505), .A2(n19996), .ZN(n19781) );
  NAND2_X1 U16616 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19781), .ZN(
        n15895) );
  AOI22_X1 U16617 ( .A1(n13373), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19971), .B2(n19468), .ZN(n13265) );
  INV_X1 U16618 ( .A(n13265), .ZN(n13266) );
  NAND2_X1 U16619 ( .A1(n13270), .A2(n13269), .ZN(n13274) );
  INV_X1 U16620 ( .A(n13271), .ZN(n13872) );
  NAND2_X1 U16621 ( .A1(n13872), .A2(n13272), .ZN(n13273) );
  INV_X1 U16622 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13841) );
  MUX2_X1 U16623 ( .A(n12552), .B(n13841), .S(n15368), .Z(n13275) );
  OAI21_X1 U16624 ( .B1(n19981), .B2(n15397), .A(n13275), .ZN(P2_U2885) );
  INV_X1 U16625 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13282) );
  NOR3_X1 U16626 ( .A1(n13276), .A2(n20042), .A3(n15965), .ZN(n13277) );
  NAND2_X1 U16627 ( .A1(n20170), .A2(n13280), .ZN(n13483) );
  NOR2_X1 U16628 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16289), .ZN(n20186) );
  NOR2_X4 U16629 ( .A1(n20170), .A2(n20973), .ZN(n20175) );
  AOI22_X1 U16630 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13281) );
  OAI21_X1 U16631 ( .B1(n13282), .B2(n13483), .A(n13281), .ZN(P1_U2907) );
  INV_X1 U16632 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14575) );
  AOI22_X1 U16633 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13283) );
  OAI21_X1 U16634 ( .B1(n14575), .B2(n13483), .A(n13283), .ZN(P1_U2911) );
  INV_X1 U16635 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U16636 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13284) );
  OAI21_X1 U16637 ( .B1(n13285), .B2(n13483), .A(n13284), .ZN(P1_U2909) );
  AOI22_X1 U16638 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13286) );
  OAI21_X1 U16639 ( .B1(n11092), .B2(n13483), .A(n13286), .ZN(P1_U2906) );
  INV_X1 U16640 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U16641 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13287) );
  OAI21_X1 U16642 ( .B1(n13288), .B2(n13483), .A(n13287), .ZN(P1_U2912) );
  INV_X1 U16643 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13290) );
  AOI22_X1 U16644 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13289) );
  OAI21_X1 U16645 ( .B1(n13290), .B2(n13483), .A(n13289), .ZN(P1_U2908) );
  INV_X1 U16646 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13292) );
  AOI22_X1 U16647 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13291) );
  OAI21_X1 U16648 ( .B1(n13292), .B2(n13483), .A(n13291), .ZN(P1_U2910) );
  NAND2_X1 U16649 ( .A1(n13294), .A2(n13293), .ZN(n13296) );
  NOR2_X1 U16650 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NOR2_X1 U16651 ( .A1(n13300), .A2(n13299), .ZN(n19141) );
  AND2_X1 U16652 ( .A1(n19158), .A2(n19141), .ZN(n19226) );
  INV_X1 U16653 ( .A(n19226), .ZN(n13302) );
  OAI211_X1 U16654 ( .C1(n19158), .C2(n19141), .A(n13302), .B(n19210), .ZN(
        n13305) );
  AOI22_X1 U16655 ( .A1(n19223), .A2(n19141), .B1(n19222), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13304) );
  OAI211_X1 U16656 ( .C1(n19231), .C2(n19325), .A(n13305), .B(n13304), .ZN(
        P2_U2919) );
  INV_X1 U16657 ( .A(n13521), .ZN(n20195) );
  INV_X1 U16658 ( .A(n13521), .ZN(n20215) );
  AOI22_X1 U16659 ( .A1(n20192), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20215), .ZN(n13312) );
  NAND2_X1 U16660 ( .A1(n13521), .A2(n13309), .ZN(n13345) );
  INV_X1 U16661 ( .A(DATAI_5_), .ZN(n13311) );
  NAND2_X1 U16662 ( .A1(n20270), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13310) );
  OAI21_X1 U16663 ( .B1(n20270), .B2(n13311), .A(n13310), .ZN(n20324) );
  NAND2_X1 U16664 ( .A1(n20203), .A2(n20324), .ZN(n13527) );
  NAND2_X1 U16665 ( .A1(n13312), .A2(n13527), .ZN(P1_U2957) );
  AOI22_X1 U16666 ( .A1(n20192), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20215), .ZN(n13315) );
  INV_X1 U16667 ( .A(DATAI_6_), .ZN(n13314) );
  NAND2_X1 U16668 ( .A1(n20270), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13313) );
  OAI21_X1 U16669 ( .B1(n20270), .B2(n13314), .A(n13313), .ZN(n20333) );
  NAND2_X1 U16670 ( .A1(n20203), .A2(n20333), .ZN(n13537) );
  NAND2_X1 U16671 ( .A1(n13315), .A2(n13537), .ZN(P1_U2958) );
  AOI22_X1 U16672 ( .A1(n20192), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20215), .ZN(n13318) );
  INV_X1 U16673 ( .A(DATAI_2_), .ZN(n13317) );
  NAND2_X1 U16674 ( .A1(n20270), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13316) );
  OAI21_X1 U16675 ( .B1(n20270), .B2(n13317), .A(n13316), .ZN(n20300) );
  NAND2_X1 U16676 ( .A1(n20203), .A2(n20300), .ZN(n13522) );
  NAND2_X1 U16677 ( .A1(n13318), .A2(n13522), .ZN(P1_U2954) );
  AOI22_X1 U16678 ( .A1(n20192), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20215), .ZN(n13321) );
  INV_X1 U16679 ( .A(DATAI_7_), .ZN(n13320) );
  NAND2_X1 U16680 ( .A1(n20270), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13319) );
  OAI21_X1 U16681 ( .B1(n20270), .B2(n13320), .A(n13319), .ZN(n20345) );
  NAND2_X1 U16682 ( .A1(n20203), .A2(n20345), .ZN(n13529) );
  NAND2_X1 U16683 ( .A1(n13321), .A2(n13529), .ZN(P1_U2959) );
  AOI22_X1 U16684 ( .A1(n20192), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20215), .ZN(n13324) );
  INV_X1 U16685 ( .A(DATAI_4_), .ZN(n13323) );
  NAND2_X1 U16686 ( .A1(n20270), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13322) );
  OAI21_X1 U16687 ( .B1(n20270), .B2(n13323), .A(n13322), .ZN(n20317) );
  NAND2_X1 U16688 ( .A1(n20203), .A2(n20317), .ZN(n13541) );
  NAND2_X1 U16689 ( .A1(n13324), .A2(n13541), .ZN(P1_U2956) );
  AOI22_X1 U16690 ( .A1(n20192), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20215), .ZN(n13327) );
  INV_X1 U16691 ( .A(DATAI_3_), .ZN(n13326) );
  NAND2_X1 U16692 ( .A1(n20270), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13325) );
  OAI21_X1 U16693 ( .B1(n20270), .B2(n13326), .A(n13325), .ZN(n20309) );
  NAND2_X1 U16694 ( .A1(n20203), .A2(n20309), .ZN(n13535) );
  NAND2_X1 U16695 ( .A1(n13327), .A2(n13535), .ZN(P1_U2955) );
  OAI21_X1 U16696 ( .B1(n13329), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13328), .ZN(n13360) );
  INV_X1 U16697 ( .A(n13330), .ZN(n13331) );
  OAI21_X1 U16698 ( .B1(n13332), .B2(n13331), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13341) );
  OR2_X1 U16699 ( .A1(n13333), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13335) );
  NAND2_X1 U16700 ( .A1(n13335), .A2(n13334), .ZN(n13679) );
  INV_X1 U16701 ( .A(n13679), .ZN(n13337) );
  INV_X1 U16702 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13336) );
  NOR2_X1 U16703 ( .A1(n20252), .A2(n13336), .ZN(n13362) );
  AOI21_X1 U16704 ( .B1(n20234), .B2(n13337), .A(n13362), .ZN(n13339) );
  AND4_X1 U16705 ( .A1(n13341), .A2(n13340), .A3(n13339), .A4(n13338), .ZN(
        n13342) );
  OAI21_X1 U16706 ( .B1(n13360), .B2(n20250), .A(n13342), .ZN(P1_U3031) );
  INV_X1 U16707 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14070) );
  INV_X1 U16708 ( .A(DATAI_15_), .ZN(n13344) );
  INV_X1 U16709 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13343) );
  MUX2_X1 U16710 ( .A(n13344), .B(n13343), .S(n20270), .Z(n14071) );
  INV_X1 U16711 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20159) );
  OAI222_X1 U16712 ( .A1(n13520), .A2(n14070), .B1(n13345), .B2(n14071), .C1(
        n13521), .C2(n20159), .ZN(P1_U2967) );
  OAI21_X1 U16713 ( .B1(n13347), .B2(n13346), .A(n13414), .ZN(n13678) );
  NAND2_X1 U16714 ( .A1(n13350), .A2(n13349), .ZN(n13351) );
  INV_X1 U16715 ( .A(n20157), .ZN(n14552) );
  AOI22_X1 U16716 ( .A1(n20152), .A2(n13671), .B1(n14552), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13354) );
  OAI21_X1 U16717 ( .B1(n13678), .B2(n14564), .A(n13354), .ZN(P1_U2871) );
  INV_X1 U16718 ( .A(n13355), .ZN(n13358) );
  OAI21_X1 U16719 ( .B1(n13358), .B2(n13357), .A(n13356), .ZN(n13684) );
  NAND2_X1 U16720 ( .A1(n13359), .A2(n14693), .ZN(n13363) );
  NOR2_X1 U16721 ( .A1(n13360), .A2(n20048), .ZN(n13361) );
  AOI211_X1 U16722 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13363), .A(
        n13362), .B(n13361), .ZN(n13364) );
  OAI21_X1 U16723 ( .B1(n14699), .B2(n13684), .A(n13364), .ZN(P1_U2999) );
  INV_X1 U16724 ( .A(DATAI_1_), .ZN(n13367) );
  NAND2_X1 U16725 ( .A1(n20270), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13366) );
  OAI21_X1 U16726 ( .B1(n20270), .B2(n13367), .A(n13366), .ZN(n20291) );
  INV_X1 U16727 ( .A(n20291), .ZN(n13368) );
  INV_X1 U16728 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20185) );
  OAI222_X1 U16729 ( .A1(n13678), .A2(n14615), .B1(n14082), .B2(n13368), .C1(
        n14600), .C2(n20185), .ZN(P1_U2903) );
  NAND2_X1 U16731 ( .A1(n19781), .A2(n19980), .ZN(n19578) );
  INV_X1 U16732 ( .A(n19578), .ZN(n13370) );
  INV_X1 U16733 ( .A(n19609), .ZN(n19606) );
  NAND2_X1 U16734 ( .A1(n15895), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13371) );
  NAND2_X1 U16735 ( .A1(n19606), .A2(n13371), .ZN(n13372) );
  AOI21_X1 U16736 ( .B1(n13373), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19722), .ZN(n13375) );
  INV_X1 U16737 ( .A(n13375), .ZN(n13377) );
  NAND2_X1 U16738 ( .A1(n13381), .A2(n13380), .ZN(n13399) );
  NOR2_X1 U16739 ( .A1(n15395), .A2(n12004), .ZN(n13387) );
  AOI21_X1 U16740 ( .B1(n12566), .B2(n15395), .A(n13387), .ZN(n13388) );
  OAI21_X1 U16741 ( .B1(n19972), .B2(n15397), .A(n13388), .ZN(P2_U2884) );
  OAI222_X1 U16742 ( .A1(n13679), .A2(n20146), .B1(n20157), .B2(n13389), .C1(
        n13684), .C2(n14564), .ZN(P1_U2872) );
  INV_X1 U16743 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13676) );
  OAI21_X1 U16744 ( .B1(n14693), .B2(n13676), .A(n13390), .ZN(n13394) );
  NOR3_X1 U16745 ( .A1(n13392), .A2(n13391), .A3(n20048), .ZN(n13393) );
  AOI211_X1 U16746 ( .C1(n16169), .C2(n13676), .A(n13394), .B(n13393), .ZN(
        n13395) );
  OAI21_X1 U16747 ( .B1(n14699), .B2(n13678), .A(n13395), .ZN(P1_U2998) );
  INV_X1 U16748 ( .A(n13396), .ZN(n13397) );
  NAND2_X1 U16749 ( .A1(n13397), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13398) );
  INV_X1 U16750 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19341) );
  NOR2_X1 U16751 ( .A1(n15261), .A2(n19341), .ZN(n13438) );
  NAND2_X1 U16752 ( .A1(n13591), .A2(n13438), .ZN(n13424) );
  XOR2_X1 U16753 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13424), .Z(n13408)
         );
  NAND2_X1 U16754 ( .A1(n13403), .A2(n13402), .ZN(n13405) );
  INV_X1 U16755 ( .A(n13426), .ZN(n13404) );
  AND2_X1 U16756 ( .A1(n13405), .A2(n13404), .ZN(n19134) );
  INV_X1 U16757 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19125) );
  NOR2_X1 U16758 ( .A1(n15395), .A2(n19125), .ZN(n13406) );
  AOI21_X1 U16759 ( .B1(n19134), .B2(n15395), .A(n13406), .ZN(n13407) );
  OAI21_X1 U16760 ( .B1(n13408), .B2(n15397), .A(n13407), .ZN(P2_U2882) );
  OR2_X1 U16761 ( .A1(n13591), .A2(n13438), .ZN(n13409) );
  NAND2_X1 U16762 ( .A1(n13409), .A2(n13424), .ZN(n19209) );
  OAI21_X1 U16763 ( .B1(n13411), .B2(n13410), .A(n13402), .ZN(n19313) );
  NOR2_X1 U16764 ( .A1(n19313), .A2(n15368), .ZN(n13412) );
  AOI21_X1 U16765 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n15370), .A(n13412), .ZN(
        n13413) );
  OAI21_X1 U16766 ( .B1(n19209), .B2(n15397), .A(n13413), .ZN(P2_U2883) );
  NAND2_X1 U16767 ( .A1(n13415), .A2(n13414), .ZN(n13416) );
  NAND2_X1 U16768 ( .A1(n13417), .A2(n13416), .ZN(n20133) );
  NAND2_X1 U16769 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  NAND2_X1 U16770 ( .A1(n13548), .A2(n13420), .ZN(n20253) );
  INV_X1 U16771 ( .A(n20253), .ZN(n13421) );
  AOI22_X1 U16772 ( .A1(n20152), .A2(n13421), .B1(n14552), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16773 ( .B1(n20133), .B2(n14564), .A(n13422), .ZN(P1_U2870) );
  INV_X1 U16774 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13423) );
  NOR2_X1 U16775 ( .A1(n13424), .A2(n13423), .ZN(n13425) );
  NAND2_X1 U16776 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13435) );
  OR2_X1 U16777 ( .A1(n13424), .A2(n13435), .ZN(n13464) );
  OAI211_X1 U16778 ( .C1(n13425), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15383), .B(n13464), .ZN(n13430) );
  NOR2_X1 U16779 ( .A1(n13427), .A2(n13426), .ZN(n13428) );
  NOR2_X1 U16780 ( .A1(n13467), .A2(n13428), .ZN(n19120) );
  NAND2_X1 U16781 ( .A1(n15395), .A2(n19120), .ZN(n13429) );
  OAI211_X1 U16782 ( .C1(n15395), .C2(n19111), .A(n13430), .B(n13429), .ZN(
        P2_U2881) );
  NOR2_X1 U16783 ( .A1(n13432), .A2(n13433), .ZN(n13434) );
  NOR2_X1 U16784 ( .A1(n13431), .A2(n13434), .ZN(n16455) );
  INV_X1 U16785 ( .A(n16455), .ZN(n13832) );
  AND2_X1 U16786 ( .A1(n13591), .A2(n13438), .ZN(n13436) );
  NOR2_X1 U16787 ( .A1(n19363), .A2(n13435), .ZN(n13437) );
  AND2_X1 U16788 ( .A1(n13436), .A2(n13437), .ZN(n13441) );
  AND2_X1 U16789 ( .A1(n13440), .A2(n13437), .ZN(n13439) );
  AND2_X1 U16790 ( .A1(n13439), .A2(n13438), .ZN(n13561) );
  NAND2_X1 U16791 ( .A1(n13591), .A2(n13561), .ZN(n13558) );
  OAI211_X1 U16792 ( .C1(n13441), .C2(n13440), .A(n13558), .B(n15383), .ZN(
        n13443) );
  NAND2_X1 U16793 ( .A1(n15370), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U16794 ( .C1(n13832), .C2(n15370), .A(n13443), .B(n13442), .ZN(
        P2_U2879) );
  NOR2_X1 U16795 ( .A1(n13445), .A2(n13444), .ZN(n20251) );
  INV_X1 U16796 ( .A(n20251), .ZN(n13446) );
  NAND3_X1 U16797 ( .A1(n13446), .A2(n20225), .A3(n20257), .ZN(n13450) );
  INV_X1 U16798 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20121) );
  OAI22_X1 U16799 ( .A1(n14693), .A2(n13447), .B1(n20252), .B2(n20121), .ZN(
        n13448) );
  AOI21_X1 U16800 ( .B1(n20137), .B2(n16169), .A(n13448), .ZN(n13449) );
  OAI211_X1 U16801 ( .C1(n14699), .C2(n20133), .A(n13450), .B(n13449), .ZN(
        P1_U2997) );
  INV_X1 U16802 ( .A(n20300), .ZN(n13451) );
  INV_X1 U16803 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20183) );
  OAI222_X1 U16804 ( .A1(n20133), .A2(n14615), .B1(n14082), .B2(n13451), .C1(
        n14600), .C2(n20183), .ZN(P1_U2902) );
  INV_X1 U16805 ( .A(DATAI_0_), .ZN(n13453) );
  NAND2_X1 U16806 ( .A1(n20270), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13452) );
  OAI21_X1 U16807 ( .B1(n20270), .B2(n13453), .A(n13452), .ZN(n20276) );
  INV_X1 U16808 ( .A(n20276), .ZN(n13454) );
  INV_X1 U16809 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20189) );
  OAI222_X1 U16810 ( .A1(n13684), .A2(n14615), .B1(n14082), .B2(n13454), .C1(
        n14600), .C2(n20189), .ZN(P1_U2904) );
  XNOR2_X1 U16811 ( .A(n19981), .B(n19983), .ZN(n13459) );
  INV_X1 U16812 ( .A(n19994), .ZN(n13455) );
  NAND2_X1 U16813 ( .A1(n19990), .A2(n13455), .ZN(n13456) );
  OAI21_X1 U16814 ( .B1(n19990), .B2(n13455), .A(n13456), .ZN(n19225) );
  NOR2_X1 U16815 ( .A1(n19225), .A2(n19226), .ZN(n19224) );
  INV_X1 U16816 ( .A(n13456), .ZN(n13457) );
  NOR2_X1 U16817 ( .A1(n19224), .A2(n13457), .ZN(n13458) );
  NOR2_X1 U16818 ( .A1(n13458), .A2(n13459), .ZN(n19202) );
  AOI21_X1 U16819 ( .B1(n13459), .B2(n13458), .A(n19202), .ZN(n13463) );
  AOI22_X1 U16820 ( .A1(n19223), .A2(n13460), .B1(n19222), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U16821 ( .A1(n19200), .A2(n16332), .ZN(n13461) );
  OAI211_X1 U16822 ( .C1(n13463), .C2(n19227), .A(n13462), .B(n13461), .ZN(
        P2_U2917) );
  XOR2_X1 U16823 ( .A(n13464), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13469)
         );
  INV_X1 U16824 ( .A(n13432), .ZN(n13465) );
  OAI21_X1 U16825 ( .B1(n13467), .B2(n13466), .A(n13465), .ZN(n19105) );
  MUX2_X1 U16826 ( .A(n12007), .B(n19105), .S(n15395), .Z(n13468) );
  OAI21_X1 U16827 ( .B1(n13469), .B2(n15397), .A(n13468), .ZN(P2_U2880) );
  INV_X1 U16828 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U16829 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13470) );
  OAI21_X1 U16830 ( .B1(n13471), .B2(n13483), .A(n13470), .ZN(P1_U2918) );
  INV_X1 U16831 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U16832 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13472) );
  OAI21_X1 U16833 ( .B1(n13473), .B2(n13483), .A(n13472), .ZN(P1_U2920) );
  INV_X1 U16834 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14601) );
  AOI22_X1 U16835 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13474) );
  OAI21_X1 U16836 ( .B1(n14601), .B2(n13483), .A(n13474), .ZN(P1_U2917) );
  AOI22_X1 U16837 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13475) );
  OAI21_X1 U16838 ( .B1(n14593), .B2(n13483), .A(n13475), .ZN(P1_U2916) );
  INV_X1 U16839 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U16840 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13476) );
  OAI21_X1 U16841 ( .B1(n13477), .B2(n13483), .A(n13476), .ZN(P1_U2915) );
  INV_X1 U16842 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13479) );
  AOI22_X1 U16843 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13478) );
  OAI21_X1 U16844 ( .B1(n13479), .B2(n13483), .A(n13478), .ZN(P1_U2919) );
  INV_X1 U16845 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U16846 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13480) );
  OAI21_X1 U16847 ( .B1(n13481), .B2(n13483), .A(n13480), .ZN(P1_U2913) );
  INV_X1 U16848 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U16849 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13482) );
  OAI21_X1 U16850 ( .B1(n13484), .B2(n13483), .A(n13482), .ZN(P1_U2914) );
  MUX2_X1 U16851 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13485), .S(
        n13507), .Z(n15975) );
  NOR2_X1 U16852 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20857), .ZN(n13510) );
  AND2_X1 U16853 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13510), .ZN(
        n13486) );
  AOI21_X1 U16854 ( .B1(n15975), .B2(n20857), .A(n13486), .ZN(n13506) );
  NAND2_X1 U16855 ( .A1(n13507), .A2(n20857), .ZN(n13487) );
  NAND2_X1 U16856 ( .A1(n13487), .A2(n10315), .ZN(n13504) );
  NAND2_X1 U16857 ( .A1(n20558), .A2(n14898), .ZN(n13501) );
  INV_X1 U16858 ( .A(n13491), .ZN(n13493) );
  MUX2_X1 U16859 ( .A(n13493), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14894), .Z(n13489) );
  INV_X1 U16860 ( .A(n13490), .ZN(n13488) );
  NAND2_X1 U16861 ( .A1(n13489), .A2(n13488), .ZN(n13498) );
  MUX2_X1 U16862 ( .A(n13490), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n10316), .Z(n13492) );
  NOR2_X1 U16863 ( .A1(n13492), .A2(n13491), .ZN(n13496) );
  OAI21_X1 U16864 ( .B1(n14894), .B2(n10315), .A(n13493), .ZN(n13494) );
  NOR2_X1 U16865 ( .A1(n13494), .A2(n10910), .ZN(n14907) );
  OAI22_X1 U16866 ( .A1(n15965), .A2(n13496), .B1(n14907), .B2(n13495), .ZN(
        n13497) );
  AOI21_X1 U16867 ( .B1(n13499), .B2(n13498), .A(n13497), .ZN(n13500) );
  INV_X1 U16868 ( .A(n13510), .ZN(n13502) );
  NAND3_X1 U16869 ( .A1(n10312), .A2(n13502), .A3(n13507), .ZN(n13503) );
  NAND2_X1 U16870 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  OR2_X1 U16871 ( .A1(n13506), .A2(n13505), .ZN(n15989) );
  OAI21_X1 U16872 ( .B1(n20113), .B2(n12488), .A(n13507), .ZN(n13509) );
  INV_X1 U16873 ( .A(n13507), .ZN(n15970) );
  NAND2_X1 U16874 ( .A1(n15970), .A2(n13208), .ZN(n13508) );
  NAND3_X1 U16875 ( .A1(n13509), .A2(n20857), .A3(n13508), .ZN(n13512) );
  NAND2_X1 U16876 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13510), .ZN(
        n13511) );
  AND2_X1 U16877 ( .A1(n13512), .A2(n13511), .ZN(n15988) );
  OAI21_X1 U16878 ( .B1(n15989), .B2(n10333), .A(n15988), .ZN(n15990) );
  OAI21_X1 U16879 ( .B1(n15990), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13513), .ZN(
        n13514) );
  NAND2_X1 U16880 ( .A1(n13514), .A2(n20454), .ZN(n20953) );
  NAND2_X1 U16881 ( .A1(n20680), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20934) );
  NOR2_X1 U16882 ( .A1(n9846), .A2(n20934), .ZN(n20733) );
  INV_X1 U16883 ( .A(n9846), .ZN(n13517) );
  NAND2_X1 U16884 ( .A1(n20680), .A2(n20965), .ZN(n20936) );
  NOR2_X1 U16885 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20857), .ZN(n20947) );
  OAI22_X1 U16886 ( .A1(n13517), .A2(n20936), .B1(n20947), .B2(n20559), .ZN(
        n13518) );
  OAI21_X1 U16887 ( .B1(n20733), .B2(n13518), .A(n20953), .ZN(n13519) );
  OAI21_X1 U16888 ( .B1(n20953), .B2(n20687), .A(n13519), .ZN(P1_U3477) );
  AOI22_X1 U16889 ( .A1(n20218), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20195), .ZN(n13523) );
  NAND2_X1 U16890 ( .A1(n13523), .A2(n13522), .ZN(P1_U2939) );
  AOI22_X1 U16891 ( .A1(n20218), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20195), .ZN(n13524) );
  NAND2_X1 U16892 ( .A1(n20203), .A2(n20276), .ZN(n13525) );
  NAND2_X1 U16893 ( .A1(n13524), .A2(n13525), .ZN(P1_U2937) );
  AOI22_X1 U16894 ( .A1(n20218), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20215), .ZN(n13526) );
  NAND2_X1 U16895 ( .A1(n13526), .A2(n13525), .ZN(P1_U2952) );
  AOI22_X1 U16896 ( .A1(n20218), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20195), .ZN(n13528) );
  NAND2_X1 U16897 ( .A1(n13528), .A2(n13527), .ZN(P1_U2942) );
  AOI22_X1 U16898 ( .A1(n20218), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20215), .ZN(n13530) );
  NAND2_X1 U16899 ( .A1(n13530), .A2(n13529), .ZN(P1_U2944) );
  AOI22_X1 U16900 ( .A1(n20218), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20215), .ZN(n13533) );
  INV_X1 U16901 ( .A(DATAI_9_), .ZN(n13532) );
  NAND2_X1 U16902 ( .A1(n20270), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13531) );
  OAI21_X1 U16903 ( .B1(n20270), .B2(n13532), .A(n13531), .ZN(n14577) );
  NAND2_X1 U16904 ( .A1(n20203), .A2(n14577), .ZN(n20207) );
  NAND2_X1 U16905 ( .A1(n13533), .A2(n20207), .ZN(P1_U2946) );
  AOI22_X1 U16906 ( .A1(n20218), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20215), .ZN(n13534) );
  NAND2_X1 U16907 ( .A1(n20203), .A2(n20291), .ZN(n13539) );
  NAND2_X1 U16908 ( .A1(n13534), .A2(n13539), .ZN(P1_U2953) );
  AOI22_X1 U16909 ( .A1(n20218), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20215), .ZN(n13536) );
  NAND2_X1 U16910 ( .A1(n13536), .A2(n13535), .ZN(P1_U2940) );
  AOI22_X1 U16911 ( .A1(n20218), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20215), .ZN(n13538) );
  NAND2_X1 U16912 ( .A1(n13538), .A2(n13537), .ZN(P1_U2943) );
  AOI22_X1 U16913 ( .A1(n20218), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20215), .ZN(n13540) );
  NAND2_X1 U16914 ( .A1(n13540), .A2(n13539), .ZN(P1_U2938) );
  AOI22_X1 U16915 ( .A1(n20218), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20215), .ZN(n13542) );
  NAND2_X1 U16916 ( .A1(n13542), .A2(n13541), .ZN(P1_U2941) );
  OAI21_X1 U16917 ( .B1(n13545), .B2(n13544), .A(n13543), .ZN(n13571) );
  INV_X1 U16918 ( .A(n20309), .ZN(n13546) );
  INV_X1 U16919 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20181) );
  OAI222_X1 U16920 ( .A1(n13571), .A2(n14615), .B1(n14082), .B2(n13546), .C1(
        n14600), .C2(n20181), .ZN(P1_U2901) );
  AND2_X1 U16921 ( .A1(n13548), .A2(n13547), .ZN(n13549) );
  OR2_X1 U16922 ( .A1(n13549), .A2(n13579), .ZN(n20231) );
  INV_X1 U16923 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13550) );
  OAI222_X1 U16924 ( .A1(n20231), .A2(n20146), .B1(n20157), .B2(n13550), .C1(
        n14564), .C2(n13571), .ZN(P1_U2869) );
  XOR2_X1 U16925 ( .A(n13559), .B(n13558), .Z(n13555) );
  NOR2_X1 U16926 ( .A1(n13431), .A2(n13552), .ZN(n13553) );
  NOR2_X1 U16927 ( .A1(n13551), .A2(n13553), .ZN(n15849) );
  INV_X1 U16928 ( .A(n15849), .ZN(n19094) );
  MUX2_X1 U16929 ( .A(n12008), .B(n19094), .S(n15395), .Z(n13554) );
  OAI21_X1 U16930 ( .B1(n13555), .B2(n15397), .A(n13554), .ZN(P2_U2878) );
  INV_X1 U16931 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19078) );
  INV_X1 U16932 ( .A(n13559), .ZN(n13557) );
  OAI21_X1 U16933 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(n13563) );
  AND2_X1 U16934 ( .A1(n13560), .A2(n13559), .ZN(n13562) );
  NAND2_X1 U16935 ( .A1(n13591), .A2(n13588), .ZN(n13615) );
  NAND3_X1 U16936 ( .A1(n13563), .A2(n15383), .A3(n13615), .ZN(n13567) );
  INV_X1 U16937 ( .A(n13617), .ZN(n13564) );
  OAI21_X1 U16938 ( .B1(n13551), .B2(n13565), .A(n13564), .ZN(n16392) );
  INV_X1 U16939 ( .A(n16392), .ZN(n19085) );
  NAND2_X1 U16940 ( .A1(n19085), .A2(n15395), .ZN(n13566) );
  OAI211_X1 U16941 ( .C1(n15395), .C2(n19078), .A(n13567), .B(n13566), .ZN(
        P2_U2877) );
  OAI21_X1 U16942 ( .B1(n13570), .B2(n13569), .A(n13568), .ZN(n20235) );
  INV_X1 U16943 ( .A(n13571), .ZN(n13690) );
  INV_X1 U16944 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13572) );
  NOR2_X1 U16945 ( .A1(n20252), .A2(n13572), .ZN(n20232) );
  AOI21_X1 U16946 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20232), .ZN(n13573) );
  OAI21_X1 U16947 ( .B1(n20230), .B2(n13693), .A(n13573), .ZN(n13574) );
  AOI21_X1 U16948 ( .B1(n13690), .B2(n16192), .A(n13574), .ZN(n13575) );
  OAI21_X1 U16949 ( .B1(n20235), .B2(n20048), .A(n13575), .ZN(P1_U2996) );
  XOR2_X1 U16950 ( .A(n13543), .B(n13576), .Z(n20224) );
  INV_X1 U16951 ( .A(n20224), .ZN(n13582) );
  AOI22_X1 U16952 ( .A1(n14314), .A2(n20317), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n14609), .ZN(n13577) );
  OAI21_X1 U16953 ( .B1(n13582), .B2(n14615), .A(n13577), .ZN(P1_U2900) );
  OR2_X1 U16954 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  NAND2_X1 U16955 ( .A1(n16274), .A2(n13580), .ZN(n20120) );
  INV_X1 U16956 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13581) );
  OAI222_X1 U16957 ( .A1(n20120), .A2(n20146), .B1(n14564), .B2(n13582), .C1(
        n20157), .C2(n13581), .ZN(P1_U2868) );
  NOR2_X1 U16958 ( .A1(n13583), .A2(n13584), .ZN(n13585) );
  NOR2_X1 U16959 ( .A1(n13646), .A2(n13585), .ZN(n16448) );
  INV_X1 U16960 ( .A(n16448), .ZN(n13596) );
  AND2_X1 U16961 ( .A1(n13587), .A2(n13586), .ZN(n13589) );
  OAI21_X1 U16962 ( .B1(n13615), .B2(n13614), .A(n13592), .ZN(n13593) );
  NAND3_X1 U16963 ( .A1(n10212), .A2(n15383), .A3(n13593), .ZN(n13595) );
  NAND2_X1 U16964 ( .A1(n15370), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13594) );
  OAI211_X1 U16965 ( .C1(n13596), .C2(n15370), .A(n13595), .B(n13594), .ZN(
        P2_U2875) );
  OAI21_X1 U16966 ( .B1(n13599), .B2(n13598), .A(n13597), .ZN(n20223) );
  NOR2_X1 U16967 ( .A1(n20254), .A2(n20120), .ZN(n13606) );
  NOR2_X1 U16968 ( .A1(n13603), .A2(n20241), .ZN(n16280) );
  OAI21_X1 U16969 ( .B1(n20245), .B2(n20249), .A(n20261), .ZN(n14206) );
  NOR2_X1 U16970 ( .A1(n20261), .A2(n20249), .ZN(n14204) );
  AOI22_X1 U16971 ( .A1(n14878), .A2(n14206), .B1(n20243), .B2(n14204), .ZN(
        n13601) );
  OAI21_X1 U16972 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20236), .ZN(n13604) );
  INV_X1 U16973 ( .A(n14204), .ZN(n13602) );
  NOR2_X1 U16974 ( .A1(n20244), .A2(n14206), .ZN(n20256) );
  AOI211_X1 U16975 ( .C1(n20248), .C2(n13602), .A(n20256), .B(n20246), .ZN(
        n20242) );
  OAI22_X1 U16976 ( .A1(n16280), .A2(n13604), .B1(n20242), .B2(n13603), .ZN(
        n13605) );
  AOI211_X1 U16977 ( .C1(n20221), .C2(P1_REIP_REG_4__SCAN_IN), .A(n13606), .B(
        n13605), .ZN(n13607) );
  OAI21_X1 U16978 ( .B1(n20223), .B2(n20250), .A(n13607), .ZN(P1_U3027) );
  NAND2_X1 U16979 ( .A1(n13610), .A2(n13609), .ZN(n13611) );
  AND2_X1 U16980 ( .A1(n13608), .A2(n13611), .ZN(n20154) );
  INV_X1 U16981 ( .A(n20154), .ZN(n13613) );
  INV_X1 U16982 ( .A(n20324), .ZN(n13612) );
  OAI222_X1 U16983 ( .A1(n13613), .A2(n14615), .B1(n14082), .B2(n13612), .C1(
        n14600), .C2(n10657), .ZN(P1_U2899) );
  XNOR2_X1 U16984 ( .A(n13615), .B(n13614), .ZN(n13621) );
  NOR2_X1 U16985 ( .A1(n13617), .A2(n13616), .ZN(n13618) );
  NOR2_X1 U16986 ( .A1(n13583), .A2(n13618), .ZN(n16386) );
  INV_X1 U16987 ( .A(n16386), .ZN(n19073) );
  MUX2_X1 U16988 ( .A(n13619), .B(n19073), .S(n15395), .Z(n13620) );
  OAI21_X1 U16989 ( .B1(n13621), .B2(n15397), .A(n13620), .ZN(P2_U2876) );
  AND2_X1 U16990 ( .A1(n19972), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19575) );
  INV_X1 U16991 ( .A(n19971), .ZN(n19974) );
  AOI21_X1 U16992 ( .B1(n19575), .B2(n19758), .A(n19974), .ZN(n13626) );
  NAND3_X1 U16993 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19980), .A3(
        n19996), .ZN(n19471) );
  NAND2_X1 U16994 ( .A1(n13626), .A2(n19471), .ZN(n13625) );
  NAND2_X1 U16995 ( .A1(n12633), .A2(n19825), .ZN(n13623) );
  NOR2_X1 U16996 ( .A1(n20006), .A2(n19471), .ZN(n19544) );
  NOR2_X1 U16997 ( .A1(n19971), .A2(n19544), .ZN(n13622) );
  AOI21_X1 U16998 ( .B1(n13623), .B2(n13622), .A(n19576), .ZN(n13624) );
  NAND2_X1 U16999 ( .A1(n13625), .A2(n13624), .ZN(n19541) );
  INV_X1 U17000 ( .A(n19541), .ZN(n19527) );
  INV_X1 U17001 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13634) );
  NOR2_X2 U17002 ( .A1(n19221), .A2(n19576), .ZN(n19851) );
  INV_X1 U17003 ( .A(n13626), .ZN(n13628) );
  OAI21_X1 U17004 ( .B1(n12633), .B2(n19544), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13627) );
  AOI22_X1 U17005 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19352), .ZN(n19855) );
  INV_X1 U17006 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20304) );
  INV_X1 U17007 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18348) );
  OAI22_X2 U17008 ( .A1(n20304), .A2(n19359), .B1(n18348), .B2(n19358), .ZN(
        n19852) );
  NOR2_X2 U17009 ( .A1(n19581), .A2(n19755), .ZN(n19569) );
  NAND2_X1 U17010 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19833), .ZN(n19342) );
  AOI22_X1 U17011 ( .A1(n19852), .A2(n19569), .B1(n19850), .B2(n19544), .ZN(
        n13631) );
  OAI21_X1 U17012 ( .B1(n19534), .B2(n19855), .A(n13631), .ZN(n13632) );
  AOI21_X1 U17013 ( .B1(n19851), .B2(n19540), .A(n13632), .ZN(n13633) );
  OAI21_X1 U17014 ( .B1(n19527), .B2(n13634), .A(n13633), .ZN(P2_U3091) );
  OAI21_X1 U17015 ( .B1(n13648), .B2(n13636), .A(n13635), .ZN(n16436) );
  INV_X1 U17016 ( .A(n13638), .ZN(n13641) );
  OAI211_X1 U17017 ( .C1(n13641), .C2(n13640), .A(n15383), .B(n13730), .ZN(
        n13643) );
  NAND2_X1 U17018 ( .A1(n15370), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13642) );
  OAI211_X1 U17019 ( .C1(n16436), .C2(n15370), .A(n13643), .B(n13642), .ZN(
        P2_U2873) );
  INV_X1 U17020 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13651) );
  OAI211_X1 U17021 ( .C1(n13637), .C2(n13644), .A(n13638), .B(n15383), .ZN(
        n13650) );
  NOR2_X1 U17022 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  NOR2_X1 U17023 ( .A1(n13648), .A2(n13647), .ZN(n19062) );
  NAND2_X1 U17024 ( .A1(n19062), .A2(n15395), .ZN(n13649) );
  OAI211_X1 U17025 ( .C1(n15395), .C2(n13651), .A(n13650), .B(n13649), .ZN(
        P2_U2874) );
  XNOR2_X1 U17026 ( .A(n13652), .B(n13653), .ZN(n16473) );
  NAND2_X1 U17027 ( .A1(n13655), .A2(n13654), .ZN(n13657) );
  XNOR2_X1 U17028 ( .A(n13657), .B(n13656), .ZN(n16476) );
  NAND2_X1 U17029 ( .A1(n16476), .A2(n16414), .ZN(n13662) );
  NAND2_X1 U17030 ( .A1(n16420), .A2(n13696), .ZN(n13658) );
  NAND2_X1 U17031 ( .A1(n16460), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16468) );
  OAI211_X1 U17032 ( .C1(n13659), .C2(n16429), .A(n13658), .B(n16468), .ZN(
        n13660) );
  AOI21_X1 U17033 ( .B1(n16426), .B2(n12566), .A(n13660), .ZN(n13661) );
  OAI211_X1 U17034 ( .C1(n16473), .C2(n16424), .A(n13662), .B(n13661), .ZN(
        P2_U3011) );
  OAI21_X1 U17035 ( .B1(n13667), .B2(n13663), .A(n16104), .ZN(n20117) );
  INV_X1 U17036 ( .A(n20117), .ZN(n20134) );
  INV_X1 U17037 ( .A(n13664), .ZN(n13665) );
  OR2_X1 U17038 ( .A1(n13668), .A2(n13667), .ZN(n20130) );
  INV_X1 U17039 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20954) );
  INV_X1 U17040 ( .A(n20125), .ZN(n20064) );
  NAND2_X1 U17041 ( .A1(n20127), .A2(n20954), .ZN(n20122) );
  OAI21_X1 U17042 ( .B1(n20064), .B2(n13669), .A(n20122), .ZN(n13670) );
  AOI21_X1 U17043 ( .B1(n13671), .B2(n20097), .A(n13670), .ZN(n13672) );
  OAI21_X1 U17044 ( .B1(n20123), .B2(n20954), .A(n13672), .ZN(n13673) );
  AOI21_X1 U17045 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20126), .A(
        n13673), .ZN(n13674) );
  OAI21_X1 U17046 ( .B1(n20559), .B2(n20130), .A(n13674), .ZN(n13675) );
  AOI21_X1 U17047 ( .B1(n20136), .B2(n13676), .A(n13675), .ZN(n13677) );
  OAI21_X1 U17048 ( .B1(n20134), .B2(n13678), .A(n13677), .ZN(P1_U2839) );
  INV_X1 U17049 ( .A(n10573), .ZN(n20946) );
  NOR2_X1 U17050 ( .A1(n20946), .A2(n20130), .ZN(n13681) );
  NOR2_X1 U17051 ( .A1(n16045), .A2(n20127), .ZN(n20096) );
  OAI22_X1 U17052 ( .A1(n20096), .A2(n13336), .B1(n20140), .B2(n13679), .ZN(
        n13680) );
  AOI211_X1 U17053 ( .C1(n20125), .C2(P1_EBX_REG_0__SCAN_IN), .A(n13681), .B(
        n13680), .ZN(n13683) );
  OAI21_X1 U17054 ( .B1(n20136), .B2(n20126), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13682) );
  OAI211_X1 U17055 ( .C1(n20134), .C2(n13684), .A(n13683), .B(n13682), .ZN(
        P1_U2840) );
  OAI221_X1 U17056 ( .B1(n20107), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20107), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20123), .ZN(n13685) );
  AOI22_X1 U17057 ( .A1(n20125), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13685), .ZN(n13687) );
  OR4_X1 U17058 ( .A1(n20107), .A2(n20121), .A3(P1_REIP_REG_3__SCAN_IN), .A4(
        n20954), .ZN(n13686) );
  OAI211_X1 U17059 ( .C1(n20231), .C2(n20140), .A(n13687), .B(n13686), .ZN(
        n13689) );
  INV_X1 U17060 ( .A(n20558), .ZN(n20935) );
  NOR2_X1 U17061 ( .A1(n20935), .A2(n20130), .ZN(n13688) );
  AOI211_X1 U17062 ( .C1(n20126), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13689), .B(n13688), .ZN(n13692) );
  NAND2_X1 U17063 ( .A1(n20117), .A2(n13690), .ZN(n13691) );
  OAI211_X1 U17064 ( .C1(n20114), .C2(n13693), .A(n13692), .B(n13691), .ZN(
        P1_U2837) );
  NAND2_X1 U17065 ( .A1(n11321), .A2(n13694), .ZN(n13695) );
  XNOR2_X1 U17066 ( .A(n13696), .B(n13695), .ZN(n13697) );
  NAND2_X1 U17067 ( .A1(n13697), .A2(n19136), .ZN(n13706) );
  OAI21_X1 U17068 ( .B1(n13700), .B2(n13699), .A(n13698), .ZN(n19214) );
  AOI22_X1 U17069 ( .A1(n19102), .A2(n10277), .B1(n19042), .B2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13702) );
  OAI21_X1 U17070 ( .B1(n19143), .B2(n19214), .A(n13702), .ZN(n13704) );
  OAI22_X1 U17071 ( .A1(n19126), .A2(n12004), .B1(n11513), .B2(n19110), .ZN(
        n13703) );
  AOI211_X1 U17072 ( .C1(n19135), .C2(n12566), .A(n13704), .B(n13703), .ZN(
        n13705) );
  OAI211_X1 U17073 ( .C1(n19972), .C2(n15060), .A(n13706), .B(n13705), .ZN(
        P2_U2852) );
  XOR2_X1 U17074 ( .A(n13608), .B(n13707), .Z(n20090) );
  INV_X1 U17075 ( .A(n20090), .ZN(n13715) );
  INV_X1 U17076 ( .A(n20333), .ZN(n13708) );
  OAI222_X1 U17077 ( .A1(n14615), .A2(n13715), .B1(n14082), .B2(n13708), .C1(
        n14600), .C2(n10675), .ZN(P1_U2898) );
  OR2_X1 U17078 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  AND2_X1 U17079 ( .A1(n13709), .A2(n13712), .ZN(n20148) );
  INV_X1 U17080 ( .A(n20148), .ZN(n13714) );
  INV_X1 U17081 ( .A(n20345), .ZN(n13713) );
  INV_X1 U17082 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20174) );
  OAI222_X1 U17083 ( .A1(n13714), .A2(n14615), .B1(n14082), .B2(n13713), .C1(
        n14600), .C2(n20174), .ZN(P1_U2897) );
  INV_X1 U17084 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13716) );
  INV_X1 U17085 ( .A(n16276), .ZN(n16260) );
  XNOR2_X1 U17086 ( .A(n16260), .B(n16259), .ZN(n16268) );
  OAI222_X1 U17087 ( .A1(n13716), .A2(n20157), .B1(n20146), .B2(n16268), .C1(
        n14564), .C2(n13715), .ZN(P1_U2866) );
  XNOR2_X1 U17088 ( .A(n13717), .B(n13718), .ZN(n19317) );
  OAI21_X1 U17089 ( .B1(n13721), .B2(n13996), .A(n13720), .ZN(n19315) );
  OAI22_X1 U17090 ( .A1(n11650), .A2(n19324), .B1(n16419), .B2(n13809), .ZN(
        n13722) );
  AOI21_X1 U17091 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16411), .A(
        n13722), .ZN(n13723) );
  OAI21_X1 U17092 ( .B1(n16393), .B2(n19313), .A(n13723), .ZN(n13724) );
  AOI21_X1 U17093 ( .B1(n19315), .B2(n16415), .A(n13724), .ZN(n13725) );
  OAI21_X1 U17094 ( .B1(n16421), .B2(n19317), .A(n13725), .ZN(P2_U3010) );
  NOR2_X1 U17095 ( .A1(n13727), .A2(n13726), .ZN(n13728) );
  NOR2_X1 U17096 ( .A1(n13742), .A2(n13728), .ZN(n16356) );
  INV_X1 U17097 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13729) );
  NOR2_X1 U17098 ( .A1(n15395), .A2(n13729), .ZN(n13733) );
  NOR2_X2 U17099 ( .A1(n13730), .A2(n13731), .ZN(n13759) );
  AOI211_X1 U17100 ( .C1(n13731), .C2(n13730), .A(n15397), .B(n13759), .ZN(
        n13732) );
  AOI211_X1 U17101 ( .C1(n16356), .C2(n15395), .A(n13733), .B(n13732), .ZN(
        n13734) );
  INV_X1 U17102 ( .A(n13734), .ZN(P2_U2872) );
  INV_X1 U17103 ( .A(n13735), .ZN(n13736) );
  AOI21_X1 U17104 ( .B1(n13737), .B2(n13709), .A(n13736), .ZN(n14494) );
  INV_X1 U17105 ( .A(n14494), .ZN(n13864) );
  INV_X1 U17106 ( .A(DATAI_8_), .ZN(n13739) );
  NAND2_X1 U17107 ( .A1(n20270), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13738) );
  OAI21_X1 U17108 ( .B1(n20270), .B2(n13739), .A(n13738), .ZN(n20190) );
  AOI22_X1 U17109 ( .A1(n14314), .A2(n20190), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14609), .ZN(n13740) );
  OAI21_X1 U17110 ( .B1(n13864), .B2(n14615), .A(n13740), .ZN(P1_U2896) );
  OAI21_X1 U17111 ( .B1(n13742), .B2(n13741), .A(n13876), .ZN(n16346) );
  NAND2_X1 U17112 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13744) );
  AOI22_X1 U17113 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15144), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13743) );
  OAI211_X1 U17114 ( .C1(n19526), .C2(n13745), .A(n13744), .B(n13743), .ZN(
        n13746) );
  INV_X1 U17115 ( .A(n13746), .ZN(n13750) );
  NAND2_X1 U17116 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13749) );
  NAND2_X1 U17117 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13748) );
  NAND2_X1 U17118 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13747) );
  AND4_X1 U17119 ( .A1(n13750), .A2(n13749), .A3(n13748), .A4(n13747), .ZN(
        n13758) );
  AOI22_X1 U17120 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15101), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U17121 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13754) );
  NAND2_X1 U17122 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13753) );
  NAND2_X1 U17123 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13752) );
  NAND2_X1 U17124 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13751) );
  AND4_X1 U17125 ( .A1(n13754), .A2(n13753), .A3(n13752), .A4(n13751), .ZN(
        n13756) );
  AOI22_X1 U17126 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13755) );
  NAND4_X1 U17127 ( .A1(n13758), .A2(n13757), .A3(n13756), .A4(n13755), .ZN(
        n13760) );
  OR2_X1 U17128 ( .A1(n13759), .A2(n13760), .ZN(n13761) );
  AND2_X1 U17129 ( .A1(n13783), .A2(n13761), .ZN(n19172) );
  NAND2_X1 U17130 ( .A1(n19172), .A2(n15383), .ZN(n13763) );
  NAND2_X1 U17131 ( .A1(n15370), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13762) );
  OAI211_X1 U17132 ( .C1(n16346), .C2(n15370), .A(n13763), .B(n13762), .ZN(
        P2_U2871) );
  NAND2_X1 U17133 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13767) );
  NAND2_X1 U17134 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13766) );
  NAND2_X1 U17135 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13765) );
  NAND2_X1 U17136 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13764) );
  NAND4_X1 U17137 ( .A1(n13767), .A2(n13766), .A3(n13765), .A4(n13764), .ZN(
        n13773) );
  AOI22_X1 U17138 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13771) );
  NAND2_X1 U17139 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13770) );
  NAND2_X1 U17140 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13769) );
  NAND2_X1 U17141 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13768) );
  NAND4_X1 U17142 ( .A1(n13771), .A2(n13770), .A3(n13769), .A4(n13768), .ZN(
        n13772) );
  NOR2_X1 U17143 ( .A1(n13773), .A2(n13772), .ZN(n13782) );
  INV_X1 U17144 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19333) );
  INV_X1 U17145 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13774) );
  OAI22_X1 U17146 ( .A1(n19333), .A2(n13913), .B1(n13912), .B2(n13774), .ZN(
        n13780) );
  NAND2_X1 U17147 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13778) );
  AOI22_X1 U17148 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15144), .ZN(n13777) );
  NAND2_X1 U17149 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13776) );
  NAND2_X1 U17150 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13775) );
  NAND4_X1 U17151 ( .A1(n13778), .A2(n13777), .A3(n13776), .A4(n13775), .ZN(
        n13779) );
  NOR2_X1 U17152 ( .A1(n13780), .A2(n13779), .ZN(n13781) );
  INV_X1 U17153 ( .A(n13785), .ZN(n13784) );
  AOI21_X1 U17154 ( .B1(n13785), .B2(n13783), .A(n13923), .ZN(n13878) );
  INV_X1 U17155 ( .A(n13878), .ZN(n13796) );
  OR2_X1 U17156 ( .A1(n15040), .A2(n13787), .ZN(n13788) );
  NAND2_X1 U17157 ( .A1(n13786), .A2(n13788), .ZN(n19040) );
  INV_X1 U17158 ( .A(n19040), .ZN(n15758) );
  INV_X1 U17159 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19266) );
  OAI22_X1 U17160 ( .A1(n16319), .A2(n19232), .B1(n19198), .B2(n19266), .ZN(
        n13794) );
  INV_X1 U17161 ( .A(n19169), .ZN(n15458) );
  INV_X1 U17162 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n13792) );
  INV_X1 U17163 ( .A(n19168), .ZN(n15456) );
  INV_X1 U17164 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13791) );
  OAI22_X1 U17165 ( .A1(n15458), .A2(n13792), .B1(n15456), .B2(n13791), .ZN(
        n13793) );
  AOI211_X1 U17166 ( .C1(n19223), .C2(n15758), .A(n13794), .B(n13793), .ZN(
        n13795) );
  OAI21_X1 U17167 ( .B1(n13796), .B2(n19227), .A(n13795), .ZN(P2_U2902) );
  AOI21_X1 U17168 ( .B1(n13797), .B2(n13798), .A(n15800), .ZN(n16447) );
  INV_X1 U17169 ( .A(n16447), .ZN(n19185) );
  NOR2_X1 U17170 ( .A1(n19117), .A2(n13799), .ZN(n13800) );
  XNOR2_X1 U17171 ( .A(n13800), .B(n16382), .ZN(n13801) );
  NAND2_X1 U17172 ( .A1(n13801), .A2(n19136), .ZN(n13808) );
  AOI22_X1 U17173 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19115), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19147), .ZN(n13802) );
  NAND2_X1 U17174 ( .A1(n19124), .A2(n13802), .ZN(n13803) );
  AOI21_X1 U17175 ( .B1(n16448), .B2(n19135), .A(n13803), .ZN(n13804) );
  OAI21_X1 U17176 ( .B1(n13805), .B2(n19145), .A(n13804), .ZN(n13806) );
  AOI21_X1 U17177 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n9962), .A(n13806), .ZN(
        n13807) );
  OAI211_X1 U17178 ( .C1(n19185), .C2(n19143), .A(n13808), .B(n13807), .ZN(
        P2_U2843) );
  INV_X1 U17179 ( .A(n13809), .ZN(n13813) );
  NOR2_X1 U17180 ( .A1(n19117), .A2(n13810), .ZN(n13812) );
  AOI21_X1 U17181 ( .B1(n13813), .B2(n13812), .A(n19888), .ZN(n13811) );
  OAI21_X1 U17182 ( .B1(n13813), .B2(n13812), .A(n13811), .ZN(n13824) );
  INV_X1 U17183 ( .A(n19313), .ZN(n13822) );
  NAND2_X1 U17184 ( .A1(n13814), .A2(n13698), .ZN(n13816) );
  INV_X1 U17185 ( .A(n13994), .ZN(n13815) );
  AOI22_X1 U17186 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19115), .B1(
        n16306), .B2(n19309), .ZN(n13817) );
  OAI211_X1 U17187 ( .C1(n19145), .C2(n13818), .A(n13817), .B(n19324), .ZN(
        n13819) );
  AOI21_X1 U17188 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n19147), .A(n13819), .ZN(
        n13820) );
  OAI21_X1 U17189 ( .B1(n19110), .B2(n11650), .A(n13820), .ZN(n13821) );
  AOI21_X1 U17190 ( .B1(n19135), .B2(n13822), .A(n13821), .ZN(n13823) );
  OAI211_X1 U17191 ( .C1(n15060), .C2(n19209), .A(n13824), .B(n13823), .ZN(
        P2_U2851) );
  NOR2_X1 U17192 ( .A1(n19117), .A2(n13825), .ZN(n13826) );
  XNOR2_X1 U17193 ( .A(n13826), .B(n16410), .ZN(n13827) );
  NAND2_X1 U17194 ( .A1(n13827), .A2(n19136), .ZN(n13837) );
  AOI21_X1 U17195 ( .B1(n13830), .B2(n13828), .A(n13829), .ZN(n16453) );
  INV_X1 U17196 ( .A(n16453), .ZN(n19195) );
  AOI22_X1 U17197 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19042), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19147), .ZN(n13831) );
  OAI211_X1 U17198 ( .C1(n19143), .C2(n19195), .A(n13831), .B(n19324), .ZN(
        n13834) );
  NOR2_X1 U17199 ( .A1(n13832), .A2(n19149), .ZN(n13833) );
  AOI211_X1 U17200 ( .C1(n19102), .C2(n13835), .A(n13834), .B(n13833), .ZN(
        n13836) );
  OAI211_X1 U17201 ( .C1(n19110), .C2(n13838), .A(n13837), .B(n13836), .ZN(
        P2_U2847) );
  NOR2_X1 U17202 ( .A1(n19117), .A2(n15049), .ZN(n13839) );
  XNOR2_X1 U17203 ( .A(n13839), .B(n14245), .ZN(n13840) );
  NAND2_X1 U17204 ( .A1(n13840), .A2(n19136), .ZN(n13848) );
  OAI22_X1 U17205 ( .A1(n19126), .A2(n13841), .B1(n11500), .B2(n19110), .ZN(
        n13844) );
  NOR2_X1 U17206 ( .A1(n19145), .A2(n13842), .ZN(n13843) );
  AOI211_X1 U17207 ( .C1(n19042), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13844), .B(n13843), .ZN(n13845) );
  OAI21_X1 U17208 ( .B1(n19983), .B2(n19143), .A(n13845), .ZN(n13846) );
  AOI21_X1 U17209 ( .B1(n19135), .B2(n16502), .A(n13846), .ZN(n13847) );
  OAI211_X1 U17210 ( .C1(n19981), .C2(n15060), .A(n13848), .B(n13847), .ZN(
        P2_U2853) );
  NOR2_X1 U17211 ( .A1(n19117), .A2(n13849), .ZN(n13850) );
  XNOR2_X1 U17212 ( .A(n13850), .B(n16371), .ZN(n13860) );
  NOR2_X1 U17213 ( .A1(n13851), .A2(n19145), .ZN(n13859) );
  AOI21_X1 U17214 ( .B1(n13853), .B2(n15799), .A(n13852), .ZN(n19178) );
  AOI22_X1 U17215 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19115), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19147), .ZN(n13854) );
  NAND2_X1 U17216 ( .A1(n19124), .A2(n13854), .ZN(n13855) );
  AOI21_X1 U17217 ( .B1(n16306), .B2(n19178), .A(n13855), .ZN(n13857) );
  NAND2_X1 U17218 ( .A1(n9962), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n13856) );
  OAI211_X1 U17219 ( .C1(n16436), .C2(n19149), .A(n13857), .B(n13856), .ZN(
        n13858) );
  AOI211_X1 U17220 ( .C1(n13860), .C2(n19136), .A(n13859), .B(n13858), .ZN(
        n13861) );
  INV_X1 U17221 ( .A(n13861), .ZN(P2_U2841) );
  NOR2_X1 U17222 ( .A1(n9948), .A2(n13862), .ZN(n13863) );
  OR2_X1 U17223 ( .A1(n16248), .A2(n13863), .ZN(n14501) );
  INV_X1 U17224 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13865) );
  OAI222_X1 U17225 ( .A1(n14501), .A2(n20146), .B1(n20157), .B2(n13865), .C1(
        n14564), .C2(n13864), .ZN(P1_U2864) );
  INV_X1 U17226 ( .A(n16501), .ZN(n13866) );
  OR2_X1 U17227 ( .A1(n19150), .A2(n13866), .ZN(n13871) );
  INV_X1 U17228 ( .A(n12971), .ZN(n13867) );
  NAND2_X1 U17229 ( .A1(n13868), .A2(n13867), .ZN(n15868) );
  MUX2_X1 U17230 ( .A(n16495), .B(n15868), .S(n11328), .Z(n13869) );
  INV_X1 U17231 ( .A(n13869), .ZN(n13870) );
  NAND2_X1 U17232 ( .A1(n13871), .A2(n13870), .ZN(n16481) );
  INV_X1 U17233 ( .A(n19965), .ZN(n16548) );
  OAI22_X1 U17234 ( .A1(n11321), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19140), .B2(n19117), .ZN(n15872) );
  AOI222_X1 U17235 ( .A1(n16481), .A2(n19969), .B1(n13872), .B2(n16548), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15872), .ZN(n13874) );
  NAND2_X1 U17236 ( .A1(n19966), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13873) );
  OAI21_X1 U17237 ( .B1(n13874), .B2(n19966), .A(n13873), .ZN(P2_U3601) );
  AND2_X1 U17238 ( .A1(n13876), .A2(n13875), .ZN(n13877) );
  OR2_X1 U17239 ( .A1(n13877), .A2(n13944), .ZN(n15761) );
  NAND2_X1 U17240 ( .A1(n13878), .A2(n15383), .ZN(n13880) );
  NAND2_X1 U17241 ( .A1(n15370), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13879) );
  OAI211_X1 U17242 ( .C1(n15761), .C2(n15370), .A(n13880), .B(n13879), .ZN(
        P2_U2870) );
  NAND2_X1 U17243 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13884) );
  NAND2_X1 U17244 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13883) );
  NAND2_X1 U17245 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13882) );
  NAND2_X1 U17246 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13881) );
  NAND4_X1 U17247 ( .A1(n13884), .A2(n13883), .A3(n13882), .A4(n13881), .ZN(
        n13890) );
  AOI22_X1 U17248 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13888) );
  NAND2_X1 U17249 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13887) );
  NAND2_X1 U17250 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13886) );
  NAND2_X1 U17251 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13885) );
  NAND4_X1 U17252 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13889) );
  NOR2_X1 U17253 ( .A1(n13890), .A2(n13889), .ZN(n13899) );
  INV_X1 U17254 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13891) );
  OAI22_X1 U17255 ( .A1(n13913), .A2(n19336), .B1(n13912), .B2(n13891), .ZN(
        n13897) );
  NAND2_X1 U17256 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13895) );
  AOI22_X1 U17257 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n15144), .ZN(n13894) );
  NAND2_X1 U17258 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13893) );
  NAND2_X1 U17259 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13892) );
  NAND4_X1 U17260 ( .A1(n13895), .A2(n13894), .A3(n13893), .A4(n13892), .ZN(
        n13896) );
  NOR2_X1 U17261 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  NAND2_X1 U17262 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13904) );
  NAND2_X1 U17263 ( .A1(n15156), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13903) );
  NAND2_X1 U17264 ( .A1(n15101), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13902) );
  NAND2_X1 U17265 ( .A1(n15110), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13901) );
  NAND4_X1 U17266 ( .A1(n13904), .A2(n13903), .A3(n13902), .A4(n13901), .ZN(
        n13910) );
  AOI22_X1 U17267 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13908) );
  NAND2_X1 U17268 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13907) );
  NAND2_X1 U17269 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13906) );
  NAND2_X1 U17270 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13905) );
  NAND4_X1 U17271 ( .A1(n13908), .A2(n13907), .A3(n13906), .A4(n13905), .ZN(
        n13909) );
  NOR2_X1 U17272 ( .A1(n13910), .A2(n13909), .ZN(n13921) );
  INV_X1 U17273 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13911) );
  OAI22_X1 U17274 ( .A1(n13913), .A2(n15903), .B1(n13912), .B2(n13911), .ZN(
        n13919) );
  NAND2_X1 U17275 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13917) );
  AOI22_X1 U17276 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n15144), .ZN(n13916) );
  NAND2_X1 U17277 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13915) );
  NAND2_X1 U17278 ( .A1(n15064), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13914) );
  NAND4_X1 U17279 ( .A1(n13917), .A2(n13916), .A3(n13915), .A4(n13914), .ZN(
        n13918) );
  NOR2_X1 U17280 ( .A1(n13919), .A2(n13918), .ZN(n13920) );
  AND2_X1 U17281 ( .A1(n13921), .A2(n13920), .ZN(n13947) );
  INV_X1 U17282 ( .A(n13947), .ZN(n13922) );
  NAND2_X1 U17283 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  AOI21_X1 U17284 ( .B1(n13925), .B2(n13924), .A(n9856), .ZN(n14022) );
  INV_X1 U17285 ( .A(n14022), .ZN(n13929) );
  XNOR2_X1 U17286 ( .A(n15024), .B(n9955), .ZN(n19021) );
  INV_X1 U17287 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19262) );
  OAI22_X1 U17288 ( .A1(n16319), .A2(n19221), .B1(n19198), .B2(n19262), .ZN(
        n13927) );
  OAI22_X1 U17289 ( .A1(n15458), .A2(n20304), .B1(n15456), .B2(n18348), .ZN(
        n13926) );
  AOI211_X1 U17290 ( .C1(n19223), .C2(n19021), .A(n13927), .B(n13926), .ZN(
        n13928) );
  OAI21_X1 U17291 ( .B1(n13929), .B2(n19227), .A(n13928), .ZN(P2_U2900) );
  XOR2_X1 U17292 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13931), .Z(
        n13932) );
  XNOR2_X1 U17293 ( .A(n13930), .B(n13932), .ZN(n13942) );
  INV_X1 U17294 ( .A(n14501), .ZN(n13936) );
  NOR2_X1 U17295 ( .A1(n20252), .A2(n21118), .ZN(n13938) );
  INV_X1 U17296 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13933) );
  INV_X1 U17297 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16266) );
  NOR2_X1 U17298 ( .A1(n13933), .A2(n16266), .ZN(n16240) );
  AND2_X1 U17299 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16280), .ZN(
        n14205) );
  NAND2_X1 U17300 ( .A1(n14205), .A2(n20236), .ZN(n16272) );
  NOR2_X1 U17301 ( .A1(n16188), .A2(n16272), .ZN(n16262) );
  OAI21_X1 U17302 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16262), .ZN(n13934) );
  OAI21_X1 U17303 ( .B1(n14856), .B2(n14205), .A(n20242), .ZN(n16277) );
  AOI21_X1 U17304 ( .B1(n16188), .B2(n16238), .A(n16277), .ZN(n16267) );
  OAI22_X1 U17305 ( .A1(n16240), .A2(n13934), .B1(n16267), .B2(n13933), .ZN(
        n13935) );
  AOI211_X1 U17306 ( .C1(n20234), .C2(n13936), .A(n13938), .B(n13935), .ZN(
        n13937) );
  OAI21_X1 U17307 ( .B1(n13942), .B2(n20250), .A(n13937), .ZN(P1_U3023) );
  AOI21_X1 U17308 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13938), .ZN(n13939) );
  OAI21_X1 U17309 ( .B1(n20230), .B2(n14497), .A(n13939), .ZN(n13940) );
  AOI21_X1 U17310 ( .B1(n14494), .B2(n16192), .A(n13940), .ZN(n13941) );
  OAI21_X1 U17311 ( .B1(n13942), .B2(n20048), .A(n13941), .ZN(P1_U2991) );
  OR2_X1 U17312 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  NAND2_X1 U17313 ( .A1(n14020), .A2(n13945), .ZN(n15744) );
  INV_X1 U17314 ( .A(n13924), .ZN(n13946) );
  AOI21_X1 U17315 ( .B1(n13947), .B2(n13900), .A(n13946), .ZN(n16334) );
  NAND2_X1 U17316 ( .A1(n16334), .A2(n15383), .ZN(n13949) );
  NAND2_X1 U17317 ( .A1(n15370), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13948) );
  OAI211_X1 U17318 ( .C1(n15744), .C2(n15370), .A(n13949), .B(n13948), .ZN(
        P2_U2869) );
  AND2_X1 U17319 ( .A1(n13735), .A2(n13951), .ZN(n13952) );
  NOR2_X1 U17320 ( .A1(n13950), .A2(n13952), .ZN(n20142) );
  INV_X1 U17321 ( .A(n20142), .ZN(n13954) );
  AOI22_X1 U17322 ( .A1(n14314), .A2(n14577), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14609), .ZN(n13953) );
  OAI21_X1 U17323 ( .B1(n13954), .B2(n14615), .A(n13953), .ZN(P1_U2895) );
  OAI21_X1 U17324 ( .B1(n13956), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13955), .ZN(n16412) );
  INV_X1 U17325 ( .A(n13957), .ZN(n13967) );
  INV_X1 U17326 ( .A(n19120), .ZN(n13964) );
  NAND2_X1 U17327 ( .A1(n16454), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13963) );
  XNOR2_X1 U17328 ( .A(n13959), .B(n13958), .ZN(n19199) );
  INV_X1 U17329 ( .A(n19199), .ZN(n13961) );
  NOR2_X1 U17330 ( .A1(n11529), .A2(n19124), .ZN(n13960) );
  AOI21_X1 U17331 ( .B1(n19310), .B2(n13961), .A(n13960), .ZN(n13962) );
  OAI211_X1 U17332 ( .C1(n13964), .C2(n19312), .A(n13963), .B(n13962), .ZN(
        n13965) );
  AOI21_X1 U17333 ( .B1(n13967), .B2(n13966), .A(n13965), .ZN(n13972) );
  INV_X1 U17334 ( .A(n13969), .ZN(n13970) );
  XNOR2_X1 U17335 ( .A(n13968), .B(n13970), .ZN(n16413) );
  NAND2_X1 U17336 ( .A1(n16413), .A2(n16475), .ZN(n13971) );
  OAI211_X1 U17337 ( .C1(n16412), .C2(n19318), .A(n13972), .B(n13971), .ZN(
        P2_U3040) );
  INV_X1 U17338 ( .A(n13973), .ZN(n13976) );
  INV_X1 U17339 ( .A(n13950), .ZN(n13975) );
  AOI21_X1 U17340 ( .B1(n13976), .B2(n13975), .A(n13974), .ZN(n14734) );
  INV_X1 U17341 ( .A(n14734), .ZN(n13980) );
  INV_X1 U17342 ( .A(DATAI_10_), .ZN(n13978) );
  NAND2_X1 U17343 ( .A1(n20270), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13977) );
  OAI21_X1 U17344 ( .B1(n20270), .B2(n13978), .A(n13977), .ZN(n20193) );
  AOI22_X1 U17345 ( .A1(n14314), .A2(n20193), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14609), .ZN(n13979) );
  OAI21_X1 U17346 ( .B1(n13980), .B2(n14615), .A(n13979), .ZN(P1_U2894) );
  NAND2_X1 U17347 ( .A1(n16250), .A2(n13981), .ZN(n13982) );
  NAND2_X1 U17348 ( .A1(n14061), .A2(n13982), .ZN(n16241) );
  OAI22_X1 U17349 ( .A1(n16241), .A2(n20146), .B1(n13983), .B2(n20157), .ZN(
        n13984) );
  AOI21_X1 U17350 ( .B1(n14734), .B2(n20153), .A(n13984), .ZN(n13985) );
  INV_X1 U17351 ( .A(n13985), .ZN(P1_U2862) );
  XNOR2_X1 U17352 ( .A(n16173), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13987) );
  XNOR2_X1 U17353 ( .A(n13986), .B(n13987), .ZN(n16246) );
  AOI22_X1 U17354 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13988) );
  OAI21_X1 U17355 ( .B1(n20230), .B2(n13989), .A(n13988), .ZN(n13990) );
  AOI21_X1 U17356 ( .B1(n20142), .B2(n16192), .A(n13990), .ZN(n13991) );
  OAI21_X1 U17357 ( .B1(n16246), .B2(n20048), .A(n13991), .ZN(P1_U2990) );
  XNOR2_X1 U17358 ( .A(n13992), .B(n13993), .ZN(n16422) );
  OAI21_X1 U17359 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n16478), .ZN(n19311) );
  XNOR2_X1 U17360 ( .A(n13995), .B(n13994), .ZN(n19206) );
  NAND2_X1 U17361 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16467), .ZN(
        n19314) );
  AOI221_X1 U17362 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13997), .C2(n13996), .A(
        n19314), .ZN(n13998) );
  AOI21_X1 U17363 ( .B1(n16460), .B2(P2_REIP_REG_5__SCAN_IN), .A(n13998), .ZN(
        n14000) );
  NAND2_X1 U17364 ( .A1(n16471), .A2(n19134), .ZN(n13999) );
  OAI211_X1 U17365 ( .C1(n16469), .C2(n19206), .A(n14000), .B(n13999), .ZN(
        n14006) );
  OAI21_X1 U17366 ( .B1(n14004), .B2(n14002), .A(n14001), .ZN(n14003) );
  OAI21_X1 U17367 ( .B1(n14004), .B2(n12853), .A(n14003), .ZN(n16423) );
  NOR2_X1 U17368 ( .A1(n16423), .A2(n19318), .ZN(n14005) );
  AOI211_X1 U17369 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n19311), .A(
        n14006), .B(n14005), .ZN(n14007) );
  OAI21_X1 U17370 ( .B1(n19316), .B2(n16422), .A(n14007), .ZN(P2_U3041) );
  NAND2_X1 U17371 ( .A1(n14734), .A2(n20089), .ZN(n14018) );
  INV_X1 U17372 ( .A(n14499), .ZN(n14008) );
  AND2_X1 U17373 ( .A1(n20127), .A2(n14008), .ZN(n20094) );
  NAND2_X1 U17374 ( .A1(n20094), .A2(n20887), .ZN(n14009) );
  OAI22_X1 U17375 ( .A1(n20140), .A2(n16241), .B1(n14010), .B2(n14009), .ZN(
        n14016) );
  INV_X1 U17376 ( .A(n14326), .ZN(n14011) );
  NAND2_X1 U17377 ( .A1(n20127), .A2(n14011), .ZN(n14012) );
  AND2_X1 U17378 ( .A1(n20123), .A2(n14012), .ZN(n14325) );
  INV_X1 U17379 ( .A(n14325), .ZN(n16129) );
  AOI22_X1 U17380 ( .A1(n20125), .A2(P1_EBX_REG_10__SCAN_IN), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n16129), .ZN(n14014) );
  NAND2_X1 U17381 ( .A1(n14013), .A2(n20123), .ZN(n20098) );
  OAI211_X1 U17382 ( .C1(n20100), .C2(n21212), .A(n14014), .B(n20098), .ZN(
        n14015) );
  NOR2_X1 U17383 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  OAI211_X1 U17384 ( .C1(n20114), .C2(n14732), .A(n14018), .B(n14017), .ZN(
        P1_U2830) );
  NAND2_X1 U17385 ( .A1(n14020), .A2(n14019), .ZN(n14021) );
  NAND2_X1 U17386 ( .A1(n15014), .A2(n14021), .ZN(n19023) );
  NAND2_X1 U17387 ( .A1(n14022), .A2(n15383), .ZN(n14024) );
  NAND2_X1 U17388 ( .A1(n15368), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14023) );
  OAI211_X1 U17389 ( .C1(n19023), .C2(n15370), .A(n14024), .B(n14023), .ZN(
        P2_U2868) );
  XNOR2_X1 U17390 ( .A(n14026), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14027) );
  XNOR2_X1 U17391 ( .A(n14025), .B(n14027), .ZN(n14046) );
  NAND2_X1 U17392 ( .A1(n9947), .A2(n14029), .ZN(n14030) );
  XNOR2_X1 U17393 ( .A(n14028), .B(n14030), .ZN(n14043) );
  OAI22_X1 U17394 ( .A1(n16429), .A2(n14031), .B1(n11535), .B2(n19124), .ZN(
        n14034) );
  INV_X1 U17395 ( .A(n19100), .ZN(n14032) );
  OAI22_X1 U17396 ( .A1(n16393), .A2(n19105), .B1(n16419), .B2(n14032), .ZN(
        n14033) );
  AOI211_X1 U17397 ( .C1(n14043), .C2(n16414), .A(n14034), .B(n14033), .ZN(
        n14035) );
  OAI21_X1 U17398 ( .B1(n14046), .B2(n16424), .A(n14035), .ZN(P2_U3007) );
  AOI22_X1 U17399 ( .A1(n16460), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n14036), 
        .B2(n16462), .ZN(n14037) );
  OAI21_X1 U17400 ( .B1(n19312), .B2(n19105), .A(n14037), .ZN(n14042) );
  OR2_X1 U17401 ( .A1(n14039), .A2(n14038), .ZN(n14040) );
  NAND2_X1 U17402 ( .A1(n14040), .A2(n13828), .ZN(n19196) );
  NOR2_X1 U17403 ( .A1(n16469), .A2(n19196), .ZN(n14041) );
  AOI211_X1 U17404 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16454), .A(
        n14042), .B(n14041), .ZN(n14045) );
  NAND2_X1 U17405 ( .A1(n14043), .A2(n16475), .ZN(n14044) );
  OAI211_X1 U17406 ( .C1(n14046), .C2(n19318), .A(n14045), .B(n14044), .ZN(
        P2_U3039) );
  NAND2_X1 U17407 ( .A1(n14048), .A2(n14047), .ZN(n14298) );
  AOI21_X1 U17408 ( .B1(n14050), .B2(n14298), .A(n10816), .ZN(n14722) );
  INV_X1 U17409 ( .A(n14722), .ZN(n14052) );
  AOI22_X1 U17410 ( .A1(n14314), .A2(n20202), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14609), .ZN(n14051) );
  OAI21_X1 U17411 ( .B1(n14052), .B2(n14615), .A(n14051), .ZN(P1_U2890) );
  NAND2_X1 U17412 ( .A1(n14319), .A2(n14053), .ZN(n14054) );
  NAND2_X1 U17413 ( .A1(n14560), .A2(n14054), .ZN(n14871) );
  OAI22_X1 U17414 ( .A1(n14871), .A2(n20146), .B1(n14055), .B2(n20157), .ZN(
        n14056) );
  AOI21_X1 U17415 ( .B1(n14722), .B2(n20153), .A(n14056), .ZN(n14057) );
  INV_X1 U17416 ( .A(n14057), .ZN(P1_U2858) );
  OR2_X1 U17417 ( .A1(n13974), .A2(n14059), .ZN(n14060) );
  XOR2_X1 U17418 ( .A(n14073), .B(n14074), .Z(n16178) );
  INV_X1 U17419 ( .A(n16178), .ZN(n14068) );
  AOI21_X1 U17420 ( .B1(n14062), .B2(n14061), .A(n14090), .ZN(n16227) );
  AOI22_X1 U17421 ( .A1(n16227), .A2(n20152), .B1(n14552), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14063) );
  OAI21_X1 U17422 ( .B1(n14068), .B2(n14564), .A(n14063), .ZN(P1_U2861) );
  INV_X1 U17423 ( .A(DATAI_11_), .ZN(n14065) );
  NAND2_X1 U17424 ( .A1(n20270), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14064) );
  OAI21_X1 U17425 ( .B1(n20270), .B2(n14065), .A(n14064), .ZN(n20196) );
  INV_X1 U17426 ( .A(n20196), .ZN(n14067) );
  OAI222_X1 U17427 ( .A1(n14068), .A2(n14615), .B1(n14082), .B2(n14067), .C1(
        n14066), .C2(n14600), .ZN(P1_U2893) );
  AOI21_X1 U17428 ( .B1(n14069), .B2(n14049), .A(n10151), .ZN(n16164) );
  INV_X1 U17429 ( .A(n16164), .ZN(n14563) );
  OAI222_X1 U17430 ( .A1(n14563), .A2(n14615), .B1(n14082), .B2(n14071), .C1(
        n14600), .C2(n14070), .ZN(P1_U2889) );
  INV_X1 U17431 ( .A(n14058), .ZN(n14072) );
  AOI21_X1 U17432 ( .B1(n14074), .B2(n14073), .A(n14072), .ZN(n14077) );
  INV_X1 U17433 ( .A(n14075), .ZN(n14076) );
  NOR2_X1 U17434 ( .A1(n14077), .A2(n14076), .ZN(n14300) );
  AOI21_X1 U17435 ( .B1(n14077), .B2(n14076), .A(n14300), .ZN(n16167) );
  INV_X1 U17436 ( .A(n16167), .ZN(n14091) );
  INV_X1 U17437 ( .A(DATAI_12_), .ZN(n14079) );
  NAND2_X1 U17438 ( .A1(n20270), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14078) );
  OAI21_X1 U17439 ( .B1(n20270), .B2(n14079), .A(n14078), .ZN(n20198) );
  INV_X1 U17440 ( .A(n20198), .ZN(n14081) );
  OAI222_X1 U17441 ( .A1(n14091), .A2(n14615), .B1(n14082), .B2(n14081), .C1(
        n14080), .C2(n14600), .ZN(P1_U2892) );
  AND2_X1 U17442 ( .A1(n14084), .A2(n14083), .ZN(n14085) );
  OR2_X1 U17443 ( .A1(n14085), .A2(n14473), .ZN(n16105) );
  AOI22_X1 U17444 ( .A1(n14610), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14609), .ZN(n14087) );
  AOI22_X1 U17445 ( .A1(n14612), .A2(n20276), .B1(n14611), .B2(DATAI_16_), 
        .ZN(n14086) );
  OAI211_X1 U17446 ( .C1(n16105), .C2(n14615), .A(n14087), .B(n14086), .ZN(
        P1_U2888) );
  INV_X1 U17447 ( .A(n14317), .ZN(n14088) );
  OAI21_X1 U17448 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n16119) );
  INV_X1 U17449 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14092) );
  OAI222_X1 U17450 ( .A1(n16119), .A2(n20146), .B1(n14092), .B2(n20157), .C1(
        n14091), .C2(n14564), .ZN(P1_U2860) );
  AOI22_X1 U17451 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17319), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17323), .ZN(n14096) );
  AOI22_X1 U17452 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17453 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17178), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17454 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17320), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17327), .ZN(n14093) );
  NAND4_X1 U17455 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14102) );
  AOI22_X1 U17456 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14100) );
  AOI22_X1 U17457 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12247), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U17458 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17459 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17317), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17310), .ZN(n14097) );
  NAND4_X1 U17460 ( .A1(n14100), .A2(n14099), .A3(n14098), .A4(n14097), .ZN(
        n14101) );
  NOR2_X1 U17461 ( .A1(n14102), .A2(n14101), .ZN(n17451) );
  INV_X1 U17462 ( .A(n17451), .ZN(n14107) );
  INV_X1 U17463 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16906) );
  INV_X1 U17464 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16942) );
  INV_X1 U17465 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16950) );
  INV_X1 U17466 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17360) );
  NAND3_X1 U17467 ( .A1(n18354), .A2(n17519), .A3(n14103), .ZN(n14104) );
  NAND2_X1 U17468 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17073) );
  NAND2_X1 U17469 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17280), .ZN(n17228) );
  AOI21_X1 U17470 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n14108), .A(
        P3_EBX_REG_17__SCAN_IN), .ZN(n14105) );
  INV_X1 U17471 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21127) );
  INV_X1 U17472 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17214) );
  NOR3_X1 U17473 ( .A1(n17211), .A2(n21127), .A3(n17214), .ZN(n17199) );
  NOR2_X1 U17474 ( .A1(n14105), .A2(n17199), .ZN(n14106) );
  MUX2_X1 U17475 ( .A(n14107), .B(n14106), .S(n17365), .Z(P3_U2686) );
  INV_X1 U17476 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16761) );
  INV_X1 U17477 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17120) );
  NOR2_X1 U17478 ( .A1(n16761), .A2(n17120), .ZN(n14193) );
  NAND2_X1 U17479 ( .A1(n17519), .A2(n17367), .ZN(n17373) );
  INV_X1 U17480 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16796) );
  INV_X1 U17481 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16812) );
  INV_X1 U17482 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17091) );
  NAND2_X1 U17483 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17129), .ZN(n17121) );
  AOI22_X1 U17484 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17485 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U17486 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14110) );
  AOI22_X1 U17487 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12242), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14109) );
  NAND4_X1 U17488 ( .A1(n14112), .A2(n14111), .A3(n14110), .A4(n14109), .ZN(
        n14118) );
  AOI22_X1 U17489 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14116) );
  AOI22_X1 U17490 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U17491 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17492 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14113) );
  NAND4_X1 U17493 ( .A1(n14116), .A2(n14115), .A3(n14114), .A4(n14113), .ZN(
        n14117) );
  NOR2_X1 U17494 ( .A1(n14118), .A2(n14117), .ZN(n17117) );
  AOI22_X1 U17495 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17496 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17497 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U17498 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14119) );
  NAND4_X1 U17499 ( .A1(n14122), .A2(n14121), .A3(n14120), .A4(n14119), .ZN(
        n14128) );
  AOI22_X1 U17500 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17501 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17502 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14124) );
  AOI22_X1 U17503 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14123) );
  NAND4_X1 U17504 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        n14127) );
  NOR2_X1 U17505 ( .A1(n14128), .A2(n14127), .ZN(n17127) );
  AOI22_X1 U17506 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17507 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U17508 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U17509 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14129) );
  NAND4_X1 U17510 ( .A1(n14132), .A2(n14131), .A3(n14130), .A4(n14129), .ZN(
        n14138) );
  AOI22_X1 U17511 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17512 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U17513 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14134) );
  AOI22_X1 U17514 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14133) );
  NAND4_X1 U17515 ( .A1(n14136), .A2(n14135), .A3(n14134), .A4(n14133), .ZN(
        n14137) );
  NOR2_X1 U17516 ( .A1(n14138), .A2(n14137), .ZN(n17135) );
  AOI22_X1 U17517 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17518 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17519 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U17520 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14139) );
  NAND4_X1 U17521 ( .A1(n14142), .A2(n14141), .A3(n14140), .A4(n14139), .ZN(
        n14148) );
  AOI22_X1 U17522 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17523 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U17524 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U17525 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14143) );
  NAND4_X1 U17526 ( .A1(n14146), .A2(n14145), .A3(n14144), .A4(n14143), .ZN(
        n14147) );
  NOR2_X1 U17527 ( .A1(n14148), .A2(n14147), .ZN(n17134) );
  NOR2_X1 U17528 ( .A1(n17135), .A2(n17134), .ZN(n17132) );
  AOI22_X1 U17529 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17317), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17323), .ZN(n14158) );
  AOI22_X1 U17530 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12211), .ZN(n14157) );
  AOI22_X1 U17531 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17283), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14149) );
  OAI21_X1 U17532 ( .B1(n17098), .B2(n21243), .A(n14149), .ZN(n14155) );
  AOI22_X1 U17533 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9827), .B1(
        n14185), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17534 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17319), .ZN(n14152) );
  AOI22_X1 U17535 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17301), .ZN(n14151) );
  AOI22_X1 U17536 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17327), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9813), .ZN(n14150) );
  NAND4_X1 U17537 ( .A1(n14153), .A2(n14152), .A3(n14151), .A4(n14150), .ZN(
        n14154) );
  AOI211_X1 U17538 ( .C1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .C2(n12247), .A(
        n14155), .B(n14154), .ZN(n14156) );
  NAND3_X1 U17539 ( .A1(n14158), .A2(n14157), .A3(n14156), .ZN(n17131) );
  NAND2_X1 U17540 ( .A1(n17132), .A2(n17131), .ZN(n17130) );
  NOR2_X1 U17541 ( .A1(n17127), .A2(n17130), .ZN(n17124) );
  AOI22_X1 U17542 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U17543 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U17544 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14159) );
  OAI21_X1 U17545 ( .B1(n17022), .B2(n21140), .A(n14159), .ZN(n14165) );
  AOI22_X1 U17546 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14163) );
  AOI22_X1 U17547 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U17548 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12242), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U17549 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14160) );
  NAND4_X1 U17550 ( .A1(n14163), .A2(n14162), .A3(n14161), .A4(n14160), .ZN(
        n14164) );
  AOI211_X1 U17551 ( .C1(n17301), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n14165), .B(n14164), .ZN(n14166) );
  NAND3_X1 U17552 ( .A1(n14168), .A2(n14167), .A3(n14166), .ZN(n17123) );
  NAND2_X1 U17553 ( .A1(n17124), .A2(n17123), .ZN(n17122) );
  NOR2_X1 U17554 ( .A1(n17117), .A2(n17122), .ZN(n17116) );
  INV_X1 U17555 ( .A(n17116), .ZN(n17110) );
  AOI22_X1 U17556 ( .A1(n14169), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14173) );
  AOI22_X1 U17557 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14172) );
  AOI22_X1 U17558 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U17559 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12242), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14170) );
  NAND4_X1 U17560 ( .A1(n14173), .A2(n14172), .A3(n14171), .A4(n14170), .ZN(
        n14180) );
  AOI22_X1 U17561 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12302), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14178) );
  AOI22_X1 U17562 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14174), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14177) );
  AOI22_X1 U17563 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14176) );
  AOI22_X1 U17564 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14175) );
  NAND4_X1 U17565 ( .A1(n14178), .A2(n14177), .A3(n14176), .A4(n14175), .ZN(
        n14179) );
  NOR2_X1 U17566 ( .A1(n14180), .A2(n14179), .ZN(n17109) );
  NOR2_X1 U17567 ( .A1(n17110), .A2(n17109), .ZN(n14192) );
  AOI22_X1 U17568 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U17569 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U17570 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14182) );
  AOI22_X1 U17571 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14181) );
  NAND4_X1 U17572 ( .A1(n14184), .A2(n14183), .A3(n14182), .A4(n14181), .ZN(
        n14191) );
  AOI22_X1 U17573 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17178), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U17574 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14188) );
  AOI22_X1 U17575 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U17576 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14186) );
  NAND4_X1 U17577 ( .A1(n14189), .A2(n14188), .A3(n14187), .A4(n14186), .ZN(
        n14190) );
  NOR2_X1 U17578 ( .A1(n14191), .A2(n14190), .ZN(n17111) );
  XNOR2_X1 U17579 ( .A(n14192), .B(n17111), .ZN(n17385) );
  AOI22_X1 U17580 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n15921), .B1(n17371), 
        .B2(n17385), .ZN(n14197) );
  INV_X1 U17581 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n14195) );
  NAND3_X1 U17582 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n14193), .ZN(n17090) );
  INV_X1 U17583 ( .A(n17090), .ZN(n14194) );
  NAND3_X1 U17584 ( .A1(n9902), .A2(n14195), .A3(n14194), .ZN(n14196) );
  NAND2_X1 U17585 ( .A1(n14197), .A2(n14196), .ZN(P3_U2674) );
  NAND3_X1 U17586 ( .A1(n15942), .A2(n14198), .A3(n18767), .ZN(n18324) );
  NOR2_X1 U17587 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18324), .ZN(n14199) );
  NAND3_X1 U17588 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(P3_STATE2_REG_0__SCAN_IN), .ZN(n18918)
         );
  OAI21_X1 U17589 ( .B1(n14199), .B2(n18918), .A(n18674), .ZN(n18329) );
  INV_X1 U17590 ( .A(n18329), .ZN(n14200) );
  INV_X1 U17591 ( .A(n17829), .ZN(n17948) );
  NOR2_X1 U17592 ( .A1(n18966), .A2(n17948), .ZN(n15924) );
  AOI21_X1 U17593 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15924), .ZN(n15925) );
  NOR2_X1 U17594 ( .A1(n14200), .A2(n15925), .ZN(n14202) );
  NOR2_X1 U17595 ( .A1(n18920), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18375) );
  OR2_X1 U17596 ( .A1(n18375), .A2(n14200), .ZN(n15923) );
  OR2_X1 U17597 ( .A1(n18394), .A2(n15923), .ZN(n14201) );
  MUX2_X1 U17598 ( .A(n14202), .B(n14201), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U17599 ( .A1(n14508), .A2(n20254), .ZN(n14229) );
  NAND2_X1 U17600 ( .A1(n14204), .A2(n14205), .ZN(n16233) );
  NAND4_X1 U17601 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16240), .ZN(n14867) );
  NOR2_X1 U17602 ( .A1(n16233), .A2(n14867), .ZN(n14213) );
  NAND2_X1 U17603 ( .A1(n14213), .A2(n20243), .ZN(n14879) );
  NOR3_X1 U17604 ( .A1(n11251), .A2(n11245), .A3(n14879), .ZN(n14798) );
  AND2_X1 U17605 ( .A1(n14206), .A2(n14205), .ZN(n16235) );
  NOR2_X1 U17606 ( .A1(n11251), .A2(n14867), .ZN(n14884) );
  NAND2_X1 U17607 ( .A1(n16235), .A2(n14884), .ZN(n14877) );
  NOR2_X1 U17608 ( .A1(n11245), .A2(n14877), .ZN(n14214) );
  INV_X1 U17609 ( .A(n14214), .ZN(n14207) );
  NOR2_X1 U17610 ( .A1(n20244), .A2(n14207), .ZN(n14208) );
  OR2_X1 U17611 ( .A1(n14798), .A2(n14208), .ZN(n16224) );
  INV_X1 U17612 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16152) );
  NAND2_X1 U17613 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14858) );
  NOR3_X1 U17614 ( .A1(n14209), .A2(n16152), .A3(n14858), .ZN(n14848) );
  AND4_X1 U17615 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n14848), .ZN(n14210) );
  NAND2_X1 U17616 ( .A1(n11257), .A2(n14210), .ZN(n14219) );
  INV_X1 U17617 ( .A(n14219), .ZN(n14211) );
  NAND2_X1 U17618 ( .A1(n14849), .A2(n14211), .ZN(n14780) );
  NOR3_X1 U17619 ( .A1(n14780), .A2(n14779), .A3(n14778), .ZN(n14772) );
  NAND3_X1 U17620 ( .A1(n14772), .A2(n14754), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14739) );
  NOR3_X1 U17621 ( .A1(n14739), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n10044), .ZN(n14228) );
  INV_X1 U17622 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14225) );
  OAI21_X1 U17623 ( .B1(n16236), .B2(n14213), .A(n14212), .ZN(n14876) );
  NAND3_X1 U17624 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U17625 ( .A1(n20248), .A2(n14866), .ZN(n14217) );
  NAND2_X1 U17626 ( .A1(n14214), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14215) );
  NAND2_X1 U17627 ( .A1(n14878), .A2(n14215), .ZN(n14216) );
  NAND2_X1 U17628 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  NAND2_X1 U17629 ( .A1(n16238), .A2(n14219), .ZN(n14220) );
  NAND2_X1 U17630 ( .A1(n14868), .A2(n14220), .ZN(n14811) );
  NOR2_X1 U17631 ( .A1(n20244), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14221) );
  NAND2_X1 U17632 ( .A1(n16238), .A2(n14797), .ZN(n14222) );
  OAI21_X1 U17633 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16236), .A(
        n14222), .ZN(n14223) );
  NOR2_X1 U17634 ( .A1(n14800), .A2(n14223), .ZN(n14787) );
  INV_X1 U17635 ( .A(n14754), .ZN(n14745) );
  NAND2_X1 U17636 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14757) );
  NOR2_X1 U17637 ( .A1(n14745), .A2(n14757), .ZN(n14224) );
  NOR2_X1 U17638 ( .A1(n14800), .A2(n16238), .ZN(n14758) );
  AOI21_X1 U17639 ( .B1(n14787), .B2(n14224), .A(n14758), .ZN(n14748) );
  AOI211_X1 U17640 ( .C1(n14225), .C2(n16238), .A(n10044), .B(n14748), .ZN(
        n14738) );
  NOR3_X1 U17641 ( .A1(n14738), .A2(n14758), .A3(n11269), .ZN(n14226) );
  OAI21_X1 U17642 ( .B1(n14203), .B2(n20250), .A(n14230), .ZN(P1_U3000) );
  AOI22_X1 U17643 ( .A1(n14610), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14609), .ZN(n14232) );
  AOI22_X1 U17644 ( .A1(n14612), .A2(n20198), .B1(n14611), .B2(DATAI_28_), 
        .ZN(n14231) );
  OAI211_X1 U17645 ( .C1(n14244), .C2(n14615), .A(n14232), .B(n14231), .ZN(
        P1_U2876) );
  AOI21_X1 U17646 ( .B1(n14233), .B2(n14434), .A(n14418), .ZN(n14764) );
  AOI22_X1 U17647 ( .A1(n14764), .A2(n20152), .B1(n14552), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n14234) );
  OAI21_X1 U17648 ( .B1(n14244), .B2(n14564), .A(n14234), .ZN(P1_U2844) );
  NAND2_X1 U17649 ( .A1(n20136), .A2(n14235), .ZN(n14240) );
  NOR3_X1 U17650 ( .A1(n20107), .A2(n14422), .A3(n14236), .ZN(n14238) );
  NOR2_X1 U17651 ( .A1(n14425), .A2(n20914), .ZN(n14237) );
  AOI211_X1 U17652 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n20125), .A(n14238), .B(
        n14237), .ZN(n14239) );
  OAI211_X1 U17653 ( .C1(n20100), .C2(n14241), .A(n14240), .B(n14239), .ZN(
        n14242) );
  AOI21_X1 U17654 ( .B1(n14764), .B2(n20097), .A(n14242), .ZN(n14243) );
  OAI21_X1 U17655 ( .B1(n14244), .B2(n16104), .A(n14243), .ZN(P1_U2812) );
  INV_X1 U17656 ( .A(n14245), .ZN(n14251) );
  INV_X1 U17657 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14246) );
  OAI22_X1 U17658 ( .A1(n16421), .A2(n14247), .B1(n16429), .B2(n14246), .ZN(
        n14250) );
  OAI22_X1 U17659 ( .A1(n16424), .A2(n14248), .B1(n11500), .B2(n19324), .ZN(
        n14249) );
  AOI211_X1 U17660 ( .C1(n16420), .C2(n14251), .A(n14250), .B(n14249), .ZN(
        n14252) );
  OAI21_X1 U17661 ( .B1(n12552), .B2(n16393), .A(n14252), .ZN(P2_U3012) );
  NAND2_X1 U17662 ( .A1(n15488), .A2(n15490), .ZN(n14254) );
  XNOR2_X1 U17663 ( .A(n14253), .B(n14254), .ZN(n14275) );
  BUF_X1 U17664 ( .A(n14255), .Z(n14256) );
  INV_X1 U17665 ( .A(n14256), .ZN(n15504) );
  NOR2_X1 U17666 ( .A1(n15504), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14271) );
  NOR2_X1 U17667 ( .A1(n14256), .A2(n14262), .ZN(n15495) );
  NOR3_X1 U17668 ( .A1(n14271), .A2(n15495), .A3(n19318), .ZN(n14266) );
  NOR2_X1 U17669 ( .A1(n14969), .A2(n14257), .ZN(n14258) );
  OR2_X1 U17670 ( .A1(n15352), .A2(n14258), .ZN(n15361) );
  NOR2_X1 U17671 ( .A1(n14973), .A2(n14259), .ZN(n14260) );
  OR2_X1 U17672 ( .A1(n15428), .A2(n14260), .ZN(n14959) );
  INV_X1 U17673 ( .A(n14959), .ZN(n15438) );
  OR2_X1 U17674 ( .A1(n19124), .A2(n19939), .ZN(n14268) );
  NAND2_X1 U17675 ( .A1(n15644), .A2(n14262), .ZN(n14261) );
  OAI211_X1 U17676 ( .C1(n15647), .C2(n14262), .A(n14268), .B(n14261), .ZN(
        n14263) );
  AOI21_X1 U17677 ( .B1(n19310), .B2(n15438), .A(n14263), .ZN(n14264) );
  OAI21_X1 U17678 ( .B1(n15361), .B2(n19312), .A(n14264), .ZN(n14265) );
  NOR2_X1 U17679 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  OAI21_X1 U17680 ( .B1(n19316), .B2(n14275), .A(n14267), .ZN(P2_U3021) );
  INV_X1 U17681 ( .A(n15361), .ZN(n14961) );
  NAND2_X1 U17682 ( .A1(n16420), .A2(n14954), .ZN(n14269) );
  OAI211_X1 U17683 ( .C1(n14270), .C2(n16429), .A(n14269), .B(n14268), .ZN(
        n14273) );
  NOR3_X1 U17684 ( .A1(n14271), .A2(n15495), .A3(n16424), .ZN(n14272) );
  AOI211_X1 U17685 ( .C1(n16426), .C2(n14961), .A(n14273), .B(n14272), .ZN(
        n14274) );
  OAI21_X1 U17686 ( .B1(n16421), .B2(n14275), .A(n14274), .ZN(P2_U2989) );
  AOI22_X1 U17687 ( .A1(n14276), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14279) );
  NAND2_X1 U17688 ( .A1(n14277), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14278) );
  OAI211_X1 U17689 ( .C1(n14281), .C2(n14280), .A(n14279), .B(n14278), .ZN(
        n14282) );
  XNOR2_X1 U17690 ( .A(n14283), .B(n14282), .ZN(n15061) );
  NOR2_X1 U17691 ( .A1(n19117), .A2(n19888), .ZN(n15034) );
  NAND2_X1 U17692 ( .A1(n14284), .A2(n15034), .ZN(n14297) );
  AOI222_X1 U17693 ( .A1(n14286), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14285), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11664), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14287) );
  INV_X1 U17694 ( .A(n14287), .ZN(n14288) );
  AOI22_X1 U17695 ( .A1(n14290), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19042), .ZN(n14291) );
  INV_X1 U17696 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14292) );
  MUX2_X1 U17697 ( .A(n16299), .B(n14294), .S(n12883), .Z(n14365) );
  NOR2_X1 U17698 ( .A1(n14365), .A2(n19145), .ZN(n14295) );
  OAI211_X1 U17699 ( .C1(n15061), .C2(n19149), .A(n14297), .B(n14296), .ZN(
        P2_U2824) );
  OAI21_X1 U17700 ( .B1(n14300), .B2(n14299), .A(n14298), .ZN(n14336) );
  INV_X1 U17701 ( .A(n14301), .ZN(n16174) );
  INV_X1 U17702 ( .A(n14302), .ZN(n14303) );
  AOI21_X1 U17703 ( .B1(n16174), .B2(n14304), .A(n14303), .ZN(n14882) );
  AND2_X1 U17704 ( .A1(n14305), .A2(n14306), .ZN(n14881) );
  NAND2_X1 U17705 ( .A1(n14882), .A2(n14881), .ZN(n14880) );
  NAND2_X1 U17706 ( .A1(n14880), .A2(n14306), .ZN(n14307) );
  XOR2_X1 U17707 ( .A(n14308), .B(n14307), .Z(n16222) );
  NAND2_X1 U17708 ( .A1(n16222), .A2(n20225), .ZN(n14311) );
  OAI22_X1 U17709 ( .A1(n14693), .A2(n14323), .B1(n20252), .B2(n20893), .ZN(
        n14309) );
  AOI21_X1 U17710 ( .B1(n16169), .B2(n14333), .A(n14309), .ZN(n14310) );
  OAI211_X1 U17711 ( .C1(n14699), .C2(n14336), .A(n14311), .B(n14310), .ZN(
        P1_U2986) );
  INV_X1 U17712 ( .A(DATAI_13_), .ZN(n14313) );
  NAND2_X1 U17713 ( .A1(n20270), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14312) );
  OAI21_X1 U17714 ( .B1(n20270), .B2(n14313), .A(n14312), .ZN(n20200) );
  AOI22_X1 U17715 ( .A1(n14314), .A2(n20200), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14609), .ZN(n14315) );
  OAI21_X1 U17716 ( .B1(n14336), .B2(n14615), .A(n14315), .ZN(P1_U2891) );
  OR2_X1 U17717 ( .A1(n14317), .A2(n14316), .ZN(n14318) );
  AND2_X1 U17718 ( .A1(n14319), .A2(n14318), .ZN(n16221) );
  NOR2_X1 U17719 ( .A1(n20157), .A2(n14320), .ZN(n14321) );
  AOI21_X1 U17720 ( .B1(n16221), .B2(n20152), .A(n14321), .ZN(n14322) );
  OAI21_X1 U17721 ( .B1(n14336), .B2(n14564), .A(n14322), .ZN(P1_U2859) );
  OAI21_X1 U17722 ( .B1(n20100), .B2(n14323), .A(n20098), .ZN(n14332) );
  NAND2_X1 U17723 ( .A1(n20127), .A2(n14327), .ZN(n14324) );
  AND2_X1 U17724 ( .A1(n14325), .A2(n14324), .ZN(n16127) );
  NAND2_X1 U17725 ( .A1(n16221), .A2(n20097), .ZN(n14330) );
  NAND2_X1 U17726 ( .A1(n20127), .A2(n14326), .ZN(n14484) );
  NOR3_X1 U17727 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14327), .A3(n14484), 
        .ZN(n14328) );
  AOI21_X1 U17728 ( .B1(n20125), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14328), .ZN(
        n14329) );
  OAI211_X1 U17729 ( .C1(n20893), .C2(n16127), .A(n14330), .B(n14329), .ZN(
        n14331) );
  NOR2_X1 U17730 ( .A1(n14332), .A2(n14331), .ZN(n14335) );
  NAND2_X1 U17731 ( .A1(n20136), .A2(n14333), .ZN(n14334) );
  OAI211_X1 U17732 ( .C1(n14336), .C2(n16104), .A(n14335), .B(n14334), .ZN(
        P1_U2827) );
  INV_X1 U17733 ( .A(n14340), .ZN(n14337) );
  OAI21_X1 U17734 ( .B1(n14338), .B2(n15481), .A(n14337), .ZN(n14339) );
  NAND2_X1 U17735 ( .A1(n14339), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14344) );
  OAI21_X1 U17736 ( .B1(n14341), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14340), .ZN(n14343) );
  NAND3_X1 U17737 ( .A1(n14344), .A2(n14343), .A3(n14342), .ZN(n15466) );
  INV_X1 U17738 ( .A(n14345), .ZN(n14347) );
  XNOR2_X1 U17739 ( .A(n14347), .B(n14346), .ZN(n14348) );
  INV_X1 U17740 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15615) );
  OAI21_X1 U17741 ( .B1(n14348), .B2(n14364), .A(n15615), .ZN(n15464) );
  INV_X1 U17742 ( .A(n14348), .ZN(n14917) );
  NAND3_X1 U17743 ( .A1(n14917), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12646), .ZN(n15465) );
  AOI21_X1 U17744 ( .B1(n14350), .B2(n12646), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14363) );
  AND2_X1 U17745 ( .A1(n12646), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14349) );
  NAND2_X1 U17746 ( .A1(n14350), .A2(n14349), .ZN(n14362) );
  INV_X1 U17747 ( .A(n14362), .ZN(n14351) );
  NOR2_X1 U17748 ( .A1(n14363), .A2(n14351), .ZN(n14352) );
  XNOR2_X1 U17749 ( .A(n14353), .B(n14352), .ZN(n14401) );
  XNOR2_X1 U17750 ( .A(n15468), .B(n14355), .ZN(n14399) );
  NOR2_X1 U17751 ( .A1(n19124), .A2(n14356), .ZN(n14391) );
  AOI21_X1 U17752 ( .B1(n16411), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14391), .ZN(n14359) );
  NAND2_X1 U17753 ( .A1(n16420), .A2(n14357), .ZN(n14358) );
  OAI211_X1 U17754 ( .C1(n14397), .C2(n16393), .A(n14359), .B(n14358), .ZN(
        n14360) );
  AOI21_X1 U17755 ( .B1(n14399), .B2(n16415), .A(n14360), .ZN(n14361) );
  OAI21_X1 U17756 ( .B1(n14401), .B2(n16421), .A(n14361), .ZN(P2_U2984) );
  XOR2_X1 U17757 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14366), .Z(
        n14367) );
  XNOR2_X1 U17758 ( .A(n14368), .B(n14367), .ZN(n14385) );
  XNOR2_X1 U17759 ( .A(n14369), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14383) );
  NAND2_X1 U17760 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15616), .ZN(
        n14390) );
  NOR4_X1 U17761 ( .A1(n15632), .A2(n14355), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n14390), .ZN(n14371) );
  INV_X1 U17762 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14370) );
  NOR2_X1 U17763 ( .A1(n19124), .A2(n14370), .ZN(n14380) );
  AOI21_X1 U17764 ( .B1(n14390), .B2(n15798), .A(n15638), .ZN(n14393) );
  OAI21_X1 U17765 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14393), .ZN(n14373) );
  NAND2_X1 U17766 ( .A1(n14373), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14374) );
  OAI211_X1 U17767 ( .C1(n15061), .C2(n19312), .A(n14375), .B(n14374), .ZN(
        n14376) );
  AOI21_X1 U17768 ( .B1(n14383), .B2(n15847), .A(n14376), .ZN(n14377) );
  OAI21_X1 U17769 ( .B1(n14385), .B2(n19316), .A(n14377), .ZN(P2_U3015) );
  NOR2_X1 U17770 ( .A1(n16419), .A2(n14378), .ZN(n14379) );
  AOI211_X1 U17771 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n16411), .A(
        n14380), .B(n14379), .ZN(n14381) );
  OAI21_X1 U17772 ( .B1(n15061), .B2(n16393), .A(n14381), .ZN(n14382) );
  AOI21_X1 U17773 ( .B1(n14383), .B2(n16415), .A(n14382), .ZN(n14384) );
  OAI21_X1 U17774 ( .B1(n14385), .B2(n16421), .A(n14384), .ZN(P2_U2983) );
  INV_X1 U17775 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20339) );
  AND2_X1 U17776 ( .A1(n14600), .A2(n20342), .ZN(n14386) );
  NAND2_X1 U17777 ( .A1(n14387), .A2(n14386), .ZN(n14389) );
  AOI22_X1 U17778 ( .A1(n14611), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14609), .ZN(n14388) );
  OAI211_X1 U17779 ( .C1(n14602), .C2(n20339), .A(n14389), .B(n14388), .ZN(
        P1_U2873) );
  NOR3_X1 U17780 ( .A1(n15632), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14390), .ZN(n14392) );
  OR2_X1 U17781 ( .A1(n14393), .A2(n14355), .ZN(n14394) );
  OAI21_X1 U17782 ( .B1(n14397), .B2(n19312), .A(n10293), .ZN(n14398) );
  OAI21_X1 U17783 ( .B1(n14401), .B2(n19316), .A(n14400), .ZN(P2_U3016) );
  INV_X1 U17784 ( .A(n14620), .ZN(n14510) );
  NAND2_X1 U17785 ( .A1(n14416), .A2(n10456), .ZN(n14405) );
  INV_X1 U17786 ( .A(n14402), .ZN(n14403) );
  NAND2_X1 U17787 ( .A1(n14418), .A2(n14403), .ZN(n14404) );
  NAND2_X1 U17788 ( .A1(n14405), .A2(n14404), .ZN(n14407) );
  XNOR2_X1 U17789 ( .A(n14407), .B(n14406), .ZN(n14742) );
  INV_X1 U17790 ( .A(n14616), .ZN(n14413) );
  AOI22_X1 U17791 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n20125), .ZN(n14412) );
  INV_X1 U17792 ( .A(n14408), .ZN(n14410) );
  OAI21_X1 U17793 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14410), .A(n14409), 
        .ZN(n14411) );
  OAI211_X1 U17794 ( .C1(n20114), .C2(n14413), .A(n14412), .B(n14411), .ZN(
        n14414) );
  AOI21_X1 U17795 ( .B1(n14742), .B2(n20097), .A(n14414), .ZN(n14415) );
  OAI21_X1 U17796 ( .B1(n14510), .B2(n16104), .A(n14415), .ZN(P1_U2810) );
  OAI21_X1 U17797 ( .B1(n14418), .B2(n14417), .A(n14416), .ZN(n14749) );
  NAND2_X1 U17798 ( .A1(n14627), .A2(n20089), .ZN(n14429) );
  NAND3_X1 U17799 ( .A1(n20127), .A2(n14422), .A3(n20916), .ZN(n14424) );
  NAND2_X1 U17800 ( .A1(n20125), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14423) );
  OAI211_X1 U17801 ( .C1(n14425), .C2(n20916), .A(n14424), .B(n14423), .ZN(
        n14427) );
  NOR2_X1 U17802 ( .A1(n20114), .A2(n14625), .ZN(n14426) );
  AOI211_X1 U17803 ( .C1(n20126), .C2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14427), .B(n14426), .ZN(n14428) );
  OAI211_X1 U17804 ( .C1(n20140), .C2(n14749), .A(n14429), .B(n14428), .ZN(
        P1_U2811) );
  AOI21_X1 U17805 ( .B1(n14431), .B2(n14430), .A(n11272), .ZN(n14635) );
  INV_X1 U17806 ( .A(n14635), .ZN(n14572) );
  NAND2_X1 U17807 ( .A1(n14453), .A2(n14432), .ZN(n14433) );
  NAND2_X1 U17808 ( .A1(n14434), .A2(n14433), .ZN(n14767) );
  INV_X1 U17809 ( .A(n14767), .ZN(n14441) );
  INV_X1 U17810 ( .A(n14435), .ZN(n14436) );
  NOR3_X1 U17811 ( .A1(n20107), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14436), 
        .ZN(n14438) );
  INV_X1 U17812 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U17813 ( .A1(n20127), .A2(n14436), .ZN(n14450) );
  AND2_X1 U17814 ( .A1(n20123), .A2(n14450), .ZN(n14445) );
  INV_X1 U17815 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21202) );
  OAI22_X1 U17816 ( .A1(n20064), .A2(n14512), .B1(n14445), .B2(n21202), .ZN(
        n14437) );
  AOI211_X1 U17817 ( .C1(n20126), .C2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14438), .B(n14437), .ZN(n14439) );
  OAI21_X1 U17818 ( .B1(n20114), .B2(n14633), .A(n14439), .ZN(n14440) );
  AOI21_X1 U17819 ( .B1(n14441), .B2(n20097), .A(n14440), .ZN(n14442) );
  OAI21_X1 U17820 ( .B1(n14572), .B2(n16104), .A(n14442), .ZN(P1_U2813) );
  OAI21_X1 U17821 ( .B1(n14443), .B2(n14444), .A(n14430), .ZN(n14641) );
  NAND2_X1 U17822 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14448) );
  INV_X1 U17823 ( .A(n14445), .ZN(n14446) );
  AOI22_X1 U17824 ( .A1(n20125), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(n14446), .ZN(n14447) );
  OAI211_X1 U17825 ( .C1(n14450), .C2(n14449), .A(n14448), .B(n14447), .ZN(
        n14455) );
  NAND2_X1 U17826 ( .A1(n14461), .A2(n14451), .ZN(n14452) );
  NAND2_X1 U17827 ( .A1(n14453), .A2(n14452), .ZN(n14777) );
  NOR2_X1 U17828 ( .A1(n14777), .A2(n20140), .ZN(n14454) );
  AOI211_X1 U17829 ( .C1(n20136), .C2(n14644), .A(n14455), .B(n14454), .ZN(
        n14456) );
  OAI21_X1 U17830 ( .B1(n14641), .B2(n16104), .A(n14456), .ZN(P1_U2814) );
  AOI21_X1 U17831 ( .B1(n14458), .B2(n14516), .A(n14443), .ZN(n14654) );
  NAND2_X1 U17832 ( .A1(n14654), .A2(n20089), .ZN(n14470) );
  OR2_X1 U17833 ( .A1(n14520), .A2(n14459), .ZN(n14460) );
  AND2_X1 U17834 ( .A1(n14461), .A2(n14460), .ZN(n14790) );
  NAND2_X1 U17835 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14467) );
  NAND2_X1 U17836 ( .A1(n20127), .A2(n16026), .ZN(n14462) );
  NAND2_X1 U17837 ( .A1(n20123), .A2(n14462), .ZN(n16040) );
  NAND2_X1 U17838 ( .A1(n16040), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U17839 ( .A1(n20125), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14465) );
  OAI21_X1 U17840 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n16026), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14463) );
  OAI211_X1 U17841 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n20127), .B(n14463), .ZN(n14464) );
  NAND4_X1 U17842 ( .A1(n14467), .A2(n14466), .A3(n14465), .A4(n14464), .ZN(
        n14468) );
  AOI21_X1 U17843 ( .B1(n14790), .B2(n20097), .A(n14468), .ZN(n14469) );
  OAI211_X1 U17844 ( .C1(n20114), .C2(n14652), .A(n14470), .B(n14469), .ZN(
        P1_U2815) );
  OAI21_X1 U17845 ( .B1(n14473), .B2(n14472), .A(n14471), .ZN(n16154) );
  INV_X1 U17846 ( .A(n16076), .ZN(n14474) );
  NOR2_X1 U17847 ( .A1(n16045), .A2(n16097), .ZN(n14485) );
  AOI21_X1 U17848 ( .B1(n14474), .B2(n14485), .A(n20096), .ZN(n16087) );
  INV_X1 U17849 ( .A(n16087), .ZN(n14481) );
  INV_X1 U17850 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20895) );
  NOR3_X1 U17851 ( .A1(n20107), .A2(n16097), .A3(n20895), .ZN(n16096) );
  AOI21_X1 U17852 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n16096), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14480) );
  AOI21_X1 U17853 ( .B1(n14475), .B2(n14556), .A(n10121), .ZN(n16208) );
  AOI21_X1 U17854 ( .B1(n20125), .B2(P1_EBX_REG_17__SCAN_IN), .A(n20110), .ZN(
        n14476) );
  OAI21_X1 U17855 ( .B1(n20100), .B2(n14477), .A(n14476), .ZN(n14478) );
  AOI21_X1 U17856 ( .B1(n16208), .B2(n20097), .A(n14478), .ZN(n14479) );
  OAI21_X1 U17857 ( .B1(n14481), .B2(n14480), .A(n14479), .ZN(n14482) );
  AOI21_X1 U17858 ( .B1(n20136), .B2(n16155), .A(n14482), .ZN(n14483) );
  OAI21_X1 U17859 ( .B1(n16154), .B2(n16104), .A(n14483), .ZN(P1_U2823) );
  NAND2_X1 U17860 ( .A1(n14722), .A2(n20089), .ZN(n14493) );
  INV_X1 U17861 ( .A(n14484), .ZN(n16128) );
  NOR2_X1 U17862 ( .A1(n20096), .A2(n14485), .ZN(n16110) );
  OAI221_X1 U17863 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14486), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(n16128), .A(n16110), .ZN(n14492) );
  INV_X1 U17864 ( .A(n14720), .ZN(n14487) );
  NAND2_X1 U17865 ( .A1(n20136), .A2(n14487), .ZN(n14491) );
  AOI22_X1 U17866 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20126), .B1(
        n20125), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n14488) );
  OAI211_X1 U17867 ( .C1(n14871), .C2(n20140), .A(n14488), .B(n20098), .ZN(
        n14489) );
  INV_X1 U17868 ( .A(n14489), .ZN(n14490) );
  NAND4_X1 U17869 ( .A1(n14493), .A2(n14492), .A3(n14491), .A4(n14490), .ZN(
        P1_U2826) );
  NAND2_X1 U17870 ( .A1(n14494), .A2(n20089), .ZN(n14506) );
  NOR2_X1 U17871 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14495), .ZN(n14496) );
  AOI22_X1 U17872 ( .A1(n20094), .A2(n14496), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n20125), .ZN(n14505) );
  INV_X1 U17873 ( .A(n14497), .ZN(n14498) );
  NAND2_X1 U17874 ( .A1(n20136), .A2(n14498), .ZN(n14504) );
  NOR2_X1 U17875 ( .A1(n16045), .A2(n14499), .ZN(n20095) );
  AOI21_X1 U17876 ( .B1(n20069), .B2(n20095), .A(n20096), .ZN(n20067) );
  AOI22_X1 U17877 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20126), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20067), .ZN(n14500) );
  OAI211_X1 U17878 ( .C1(n20140), .C2(n14501), .A(n14500), .B(n20098), .ZN(
        n14502) );
  INV_X1 U17879 ( .A(n14502), .ZN(n14503) );
  NAND4_X1 U17880 ( .A1(n14506), .A2(n14505), .A3(n14504), .A4(n14503), .ZN(
        P1_U2832) );
  INV_X1 U17881 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14507) );
  OAI22_X1 U17882 ( .A1(n14508), .A2(n20146), .B1(n14507), .B2(n20157), .ZN(
        P1_U2841) );
  AOI22_X1 U17883 ( .A1(n14742), .A2(n20152), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14552), .ZN(n14509) );
  OAI21_X1 U17884 ( .B1(n14510), .B2(n14564), .A(n14509), .ZN(P1_U2842) );
  INV_X1 U17885 ( .A(n14627), .ZN(n14568) );
  OAI222_X1 U17886 ( .A1(n14511), .A2(n20157), .B1(n20146), .B2(n14749), .C1(
        n14568), .C2(n14564), .ZN(P1_U2843) );
  OAI222_X1 U17887 ( .A1(n14512), .A2(n20157), .B1(n20146), .B2(n14767), .C1(
        n14572), .C2(n14564), .ZN(P1_U2845) );
  OAI222_X1 U17888 ( .A1(n14513), .A2(n20157), .B1(n20146), .B2(n14777), .C1(
        n14641), .C2(n14564), .ZN(P1_U2846) );
  INV_X1 U17889 ( .A(n14654), .ZN(n14580) );
  AOI22_X1 U17890 ( .A1(n14790), .A2(n20152), .B1(n14552), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14514) );
  OAI21_X1 U17891 ( .B1(n14580), .B2(n14564), .A(n14514), .ZN(P1_U2847) );
  OAI21_X1 U17892 ( .B1(n14515), .B2(n14517), .A(n14516), .ZN(n16031) );
  NOR2_X1 U17893 ( .A1(n14807), .A2(n14518), .ZN(n14519) );
  OR2_X1 U17894 ( .A1(n14520), .A2(n14519), .ZN(n16035) );
  OAI22_X1 U17895 ( .A1(n16035), .A2(n20146), .B1(n14521), .B2(n20157), .ZN(
        n14522) );
  INV_X1 U17896 ( .A(n14522), .ZN(n14523) );
  OAI21_X1 U17897 ( .B1(n16031), .B2(n14564), .A(n14523), .ZN(P1_U2848) );
  NAND2_X1 U17898 ( .A1(n14524), .A2(n14525), .ZN(n14526) );
  NAND2_X1 U17899 ( .A1(n14533), .A2(n14527), .ZN(n14528) );
  NAND2_X1 U17900 ( .A1(n14806), .A2(n14528), .ZN(n16054) );
  OAI22_X1 U17901 ( .A1(n16054), .A2(n20146), .B1(n16046), .B2(n20157), .ZN(
        n14529) );
  INV_X1 U17902 ( .A(n14529), .ZN(n14530) );
  OAI21_X1 U17903 ( .B1(n14590), .B2(n14564), .A(n14530), .ZN(P1_U2850) );
  INV_X1 U17904 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14537) );
  OR2_X1 U17905 ( .A1(n14540), .A2(n14531), .ZN(n14532) );
  NAND2_X1 U17906 ( .A1(n14533), .A2(n14532), .ZN(n16061) );
  OAI21_X1 U17908 ( .B1(n14535), .B2(n14536), .A(n14524), .ZN(n16060) );
  OAI222_X1 U17909 ( .A1(n14537), .A2(n20157), .B1(n20146), .B2(n16061), .C1(
        n16060), .C2(n14564), .ZN(P1_U2851) );
  NOR2_X1 U17910 ( .A1(n16082), .A2(n14538), .ZN(n14539) );
  OR2_X1 U17911 ( .A1(n14540), .A2(n14539), .ZN(n16068) );
  INV_X1 U17912 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14544) );
  INV_X1 U17913 ( .A(n14535), .ZN(n14542) );
  OAI21_X1 U17914 ( .B1(n14543), .B2(n14541), .A(n14542), .ZN(n16069) );
  OAI222_X1 U17915 ( .A1(n16068), .A2(n20146), .B1(n20157), .B2(n14544), .C1(
        n14564), .C2(n16069), .ZN(P1_U2852) );
  NAND2_X1 U17916 ( .A1(n14546), .A2(n14545), .ZN(n14547) );
  NAND2_X1 U17917 ( .A1(n16083), .A2(n14547), .ZN(n16095) );
  INV_X1 U17918 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U17919 ( .A1(n14471), .A2(n14549), .ZN(n14550) );
  AND2_X1 U17920 ( .A1(n14598), .A2(n14550), .ZN(n16092) );
  OAI222_X1 U17921 ( .A1(n16095), .A2(n20146), .B1(n20157), .B2(n14551), .C1(
        n14564), .C2(n14700), .ZN(P1_U2854) );
  AOI22_X1 U17922 ( .A1(n16208), .A2(n20152), .B1(n14552), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14553) );
  OAI21_X1 U17923 ( .B1(n16154), .B2(n14564), .A(n14553), .ZN(P1_U2855) );
  INV_X1 U17924 ( .A(n16105), .ZN(n14711) );
  OR2_X1 U17925 ( .A1(n14562), .A2(n14554), .ZN(n14555) );
  NAND2_X1 U17926 ( .A1(n14556), .A2(n14555), .ZN(n16109) );
  OAI22_X1 U17927 ( .A1(n16109), .A2(n20146), .B1(n16101), .B2(n20157), .ZN(
        n14557) );
  AOI21_X1 U17928 ( .B1(n14711), .B2(n20153), .A(n14557), .ZN(n14558) );
  INV_X1 U17929 ( .A(n14558), .ZN(P1_U2856) );
  AND2_X1 U17930 ( .A1(n14560), .A2(n14559), .ZN(n14561) );
  OR2_X1 U17931 ( .A1(n14562), .A2(n14561), .ZN(n16215) );
  INV_X1 U17932 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14565) );
  OAI222_X1 U17933 ( .A1(n16215), .A2(n20146), .B1(n14565), .B2(n20157), .C1(
        n14564), .C2(n14563), .ZN(P1_U2857) );
  AOI22_X1 U17934 ( .A1(n14610), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14609), .ZN(n14567) );
  AOI22_X1 U17935 ( .A1(n14612), .A2(n20200), .B1(n14611), .B2(DATAI_29_), 
        .ZN(n14566) );
  OAI211_X1 U17936 ( .C1(n14568), .C2(n14615), .A(n14567), .B(n14566), .ZN(
        P1_U2875) );
  OAI22_X1 U17937 ( .A1(n14602), .A2(n20306), .B1(n13285), .B2(n14600), .ZN(
        n14569) );
  INV_X1 U17938 ( .A(n14569), .ZN(n14571) );
  AOI22_X1 U17939 ( .A1(n14612), .A2(n20196), .B1(n14611), .B2(DATAI_27_), 
        .ZN(n14570) );
  OAI211_X1 U17940 ( .C1(n14572), .C2(n14615), .A(n14571), .B(n14570), .ZN(
        P1_U2877) );
  AOI22_X1 U17941 ( .A1(n14610), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14609), .ZN(n14574) );
  AOI22_X1 U17942 ( .A1(n14612), .A2(n20193), .B1(n14611), .B2(DATAI_26_), 
        .ZN(n14573) );
  OAI211_X1 U17943 ( .C1(n14641), .C2(n14615), .A(n14574), .B(n14573), .ZN(
        P1_U2878) );
  INV_X1 U17944 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20286) );
  OAI22_X1 U17945 ( .A1(n14602), .A2(n20286), .B1(n14575), .B2(n14600), .ZN(
        n14576) );
  INV_X1 U17946 ( .A(n14576), .ZN(n14579) );
  AOI22_X1 U17947 ( .A1(n14612), .A2(n14577), .B1(n14611), .B2(DATAI_25_), 
        .ZN(n14578) );
  OAI211_X1 U17948 ( .C1(n14580), .C2(n14615), .A(n14579), .B(n14578), .ZN(
        P1_U2879) );
  AOI22_X1 U17949 ( .A1(n14610), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14609), .ZN(n14582) );
  AOI22_X1 U17950 ( .A1(n14612), .A2(n20190), .B1(n14611), .B2(DATAI_24_), 
        .ZN(n14581) );
  OAI211_X1 U17951 ( .C1(n16031), .C2(n14615), .A(n14582), .B(n14581), .ZN(
        P1_U2880) );
  AND2_X1 U17952 ( .A1(n9880), .A2(n14583), .ZN(n14584) );
  OR2_X1 U17953 ( .A1(n14584), .A2(n14515), .ZN(n16135) );
  INV_X1 U17954 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20336) );
  OAI22_X1 U17955 ( .A1(n14602), .A2(n20336), .B1(n13481), .B2(n14600), .ZN(
        n14585) );
  INV_X1 U17956 ( .A(n14585), .ZN(n14587) );
  AOI22_X1 U17957 ( .A1(n14612), .A2(n20345), .B1(n14611), .B2(DATAI_23_), 
        .ZN(n14586) );
  OAI211_X1 U17958 ( .C1(n16135), .C2(n14615), .A(n14587), .B(n14586), .ZN(
        P1_U2881) );
  AOI22_X1 U17959 ( .A1(n14610), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14609), .ZN(n14589) );
  AOI22_X1 U17960 ( .A1(n14612), .A2(n20333), .B1(n14611), .B2(DATAI_22_), 
        .ZN(n14588) );
  OAI211_X1 U17961 ( .C1(n14590), .C2(n14615), .A(n14589), .B(n14588), .ZN(
        P1_U2882) );
  AOI22_X1 U17962 ( .A1(n14610), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14609), .ZN(n14592) );
  AOI22_X1 U17963 ( .A1(n14612), .A2(n20324), .B1(n14611), .B2(DATAI_21_), 
        .ZN(n14591) );
  OAI211_X1 U17964 ( .C1(n16060), .C2(n14615), .A(n14592), .B(n14591), .ZN(
        P1_U2883) );
  INV_X1 U17965 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14594) );
  OAI22_X1 U17966 ( .A1(n14602), .A2(n14594), .B1(n14593), .B2(n14600), .ZN(
        n14595) );
  INV_X1 U17967 ( .A(n14595), .ZN(n14597) );
  AOI22_X1 U17968 ( .A1(n14612), .A2(n20317), .B1(n14611), .B2(DATAI_20_), 
        .ZN(n14596) );
  OAI211_X1 U17969 ( .C1(n16069), .C2(n14615), .A(n14597), .B(n14596), .ZN(
        P1_U2884) );
  AOI21_X1 U17970 ( .B1(n14599), .B2(n14598), .A(n14541), .ZN(n16144) );
  INV_X1 U17971 ( .A(n16144), .ZN(n14606) );
  OAI22_X1 U17972 ( .A1(n14602), .A2(n20304), .B1(n14601), .B2(n14600), .ZN(
        n14603) );
  INV_X1 U17973 ( .A(n14603), .ZN(n14605) );
  AOI22_X1 U17974 ( .A1(n14612), .A2(n20309), .B1(n14611), .B2(DATAI_19_), 
        .ZN(n14604) );
  OAI211_X1 U17975 ( .C1(n14606), .C2(n14615), .A(n14605), .B(n14604), .ZN(
        P1_U2885) );
  AOI22_X1 U17976 ( .A1(n14610), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14609), .ZN(n14608) );
  AOI22_X1 U17977 ( .A1(n14612), .A2(n20300), .B1(n14611), .B2(DATAI_18_), 
        .ZN(n14607) );
  OAI211_X1 U17978 ( .C1(n14700), .C2(n14615), .A(n14608), .B(n14607), .ZN(
        P1_U2886) );
  AOI22_X1 U17979 ( .A1(n14610), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14609), .ZN(n14614) );
  AOI22_X1 U17980 ( .A1(n14612), .A2(n20291), .B1(n14611), .B2(DATAI_17_), 
        .ZN(n14613) );
  OAI211_X1 U17981 ( .C1(n16154), .C2(n14615), .A(n14614), .B(n14613), .ZN(
        P1_U2887) );
  NAND2_X1 U17982 ( .A1(n14616), .A2(n16169), .ZN(n14617) );
  NAND2_X1 U17983 ( .A1(n20221), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14737) );
  OAI211_X1 U17984 ( .C1(n14618), .C2(n14693), .A(n14617), .B(n14737), .ZN(
        n14619) );
  AOI21_X1 U17985 ( .B1(n14620), .B2(n16192), .A(n14619), .ZN(n14621) );
  OAI21_X1 U17986 ( .B1(n14744), .B2(n20048), .A(n14621), .ZN(P1_U2969) );
  NOR2_X1 U17987 ( .A1(n20252), .A2(n20916), .ZN(n14747) );
  AOI21_X1 U17988 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14747), .ZN(n14624) );
  OAI21_X1 U17989 ( .B1(n14625), .B2(n20230), .A(n14624), .ZN(n14626) );
  AOI21_X1 U17990 ( .B1(n14627), .B2(n16192), .A(n14626), .ZN(n14628) );
  OAI21_X1 U17991 ( .B1(n20048), .B2(n14753), .A(n14628), .ZN(P1_U2970) );
  MUX2_X1 U17992 ( .A(n14630), .B(n14629), .S(n14728), .Z(n14631) );
  XNOR2_X1 U17993 ( .A(n14631), .B(n14771), .ZN(n14775) );
  NOR2_X1 U17994 ( .A1(n20252), .A2(n21202), .ZN(n14769) );
  AOI21_X1 U17995 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14769), .ZN(n14632) );
  OAI21_X1 U17996 ( .B1(n14633), .B2(n20230), .A(n14632), .ZN(n14634) );
  AOI21_X1 U17997 ( .B1(n14635), .B2(n16192), .A(n14634), .ZN(n14636) );
  OAI21_X1 U17998 ( .B1(n20048), .B2(n14775), .A(n14636), .ZN(P1_U2972) );
  OAI211_X1 U17999 ( .C1(n14728), .C2(n11275), .A(n14638), .B(n14637), .ZN(
        n14639) );
  XNOR2_X1 U18000 ( .A(n14639), .B(n14778), .ZN(n14785) );
  NAND2_X1 U18001 ( .A1(n20221), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14776) );
  OAI21_X1 U18002 ( .B1(n14693), .B2(n14640), .A(n14776), .ZN(n14643) );
  NOR2_X1 U18003 ( .A1(n14641), .A2(n14699), .ZN(n14642) );
  AOI211_X1 U18004 ( .C1(n16169), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        n14645) );
  OAI21_X1 U18005 ( .B1(n20048), .B2(n14785), .A(n14645), .ZN(P1_U2973) );
  NAND2_X1 U18006 ( .A1(n14658), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14649) );
  INV_X1 U18007 ( .A(n11275), .ZN(n14647) );
  NAND3_X1 U18008 ( .A1(n14647), .A2(n14797), .A3(n14812), .ZN(n14648) );
  MUX2_X1 U18009 ( .A(n14649), .B(n14648), .S(n14728), .Z(n14650) );
  XNOR2_X1 U18010 ( .A(n14650), .B(n14786), .ZN(n14793) );
  INV_X1 U18011 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20909) );
  NOR2_X1 U18012 ( .A1(n20252), .A2(n20909), .ZN(n14789) );
  AOI21_X1 U18013 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14789), .ZN(n14651) );
  OAI21_X1 U18014 ( .B1(n14652), .B2(n20230), .A(n14651), .ZN(n14653) );
  AOI21_X1 U18015 ( .B1(n14654), .B2(n16192), .A(n14653), .ZN(n14655) );
  OAI21_X1 U18016 ( .B1(n20048), .B2(n14793), .A(n14655), .ZN(P1_U2974) );
  INV_X1 U18017 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21260) );
  NOR2_X1 U18018 ( .A1(n20252), .A2(n21260), .ZN(n14795) );
  NOR2_X1 U18019 ( .A1(n14693), .A2(n14656), .ZN(n14657) );
  AOI211_X1 U18020 ( .C1(n16033), .C2(n16169), .A(n14795), .B(n14657), .ZN(
        n14662) );
  NOR2_X1 U18021 ( .A1(n14658), .A2(n11275), .ZN(n14659) );
  MUX2_X1 U18022 ( .A(n14659), .B(n14658), .S(n16173), .Z(n14660) );
  XNOR2_X1 U18023 ( .A(n14660), .B(n14797), .ZN(n14794) );
  NAND2_X1 U18024 ( .A1(n14794), .A2(n20225), .ZN(n14661) );
  OAI211_X1 U18025 ( .C1(n16031), .C2(n14699), .A(n14662), .B(n14661), .ZN(
        P1_U2975) );
  XNOR2_X1 U18026 ( .A(n16173), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14663) );
  XNOR2_X1 U18027 ( .A(n11275), .B(n14663), .ZN(n14816) );
  INV_X1 U18028 ( .A(n16135), .ZN(n14667) );
  INV_X1 U18029 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14664) );
  NOR2_X1 U18030 ( .A1(n20252), .A2(n14664), .ZN(n14810) );
  AOI21_X1 U18031 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14810), .ZN(n14665) );
  OAI21_X1 U18032 ( .B1(n16044), .B2(n20230), .A(n14665), .ZN(n14666) );
  AOI21_X1 U18033 ( .B1(n14667), .B2(n16192), .A(n14666), .ZN(n14668) );
  OAI21_X1 U18034 ( .B1(n14816), .B2(n20048), .A(n14668), .ZN(P1_U2976) );
  NAND2_X1 U18035 ( .A1(n14670), .A2(n14669), .ZN(n14671) );
  XNOR2_X1 U18036 ( .A(n14671), .B(n14823), .ZN(n14828) );
  NAND2_X1 U18037 ( .A1(n16051), .A2(n16192), .ZN(n14675) );
  NOR2_X1 U18038 ( .A1(n20252), .A2(n21166), .ZN(n14820) );
  NOR2_X1 U18039 ( .A1(n14693), .A2(n14672), .ZN(n14673) );
  AOI211_X1 U18040 ( .C1(n16050), .C2(n16169), .A(n14820), .B(n14673), .ZN(
        n14674) );
  OAI211_X1 U18041 ( .C1(n14828), .C2(n20048), .A(n14675), .B(n14674), .ZN(
        P1_U2977) );
  OAI21_X1 U18042 ( .B1(n16173), .B2(n11260), .A(n14676), .ZN(n16142) );
  OR2_X1 U18043 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16141) );
  NAND2_X1 U18044 ( .A1(n16173), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16140) );
  OAI22_X1 U18045 ( .A1(n16142), .A2(n16141), .B1(n14676), .B2(n16140), .ZN(
        n14688) );
  NAND2_X1 U18046 ( .A1(n14688), .A2(n14687), .ZN(n14686) );
  INV_X1 U18047 ( .A(n16140), .ZN(n14677) );
  NAND2_X1 U18048 ( .A1(n14677), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14678) );
  OAI22_X1 U18049 ( .A1(n14686), .A2(n16173), .B1(n14676), .B2(n14678), .ZN(
        n14679) );
  XOR2_X1 U18050 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14679), .Z(
        n14829) );
  NAND2_X1 U18051 ( .A1(n14829), .A2(n20225), .ZN(n14683) );
  INV_X1 U18052 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14680) );
  NOR2_X1 U18053 ( .A1(n20252), .A2(n14680), .ZN(n14831) );
  NOR2_X1 U18054 ( .A1(n16066), .A2(n20230), .ZN(n14681) );
  AOI211_X1 U18055 ( .C1(n20222), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14831), .B(n14681), .ZN(n14682) );
  OAI211_X1 U18056 ( .C1(n14699), .C2(n16060), .A(n14683), .B(n14682), .ZN(
        P1_U2978) );
  NAND2_X1 U18057 ( .A1(n20221), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14838) );
  OAI21_X1 U18058 ( .B1(n14693), .B2(n14684), .A(n14838), .ZN(n14685) );
  AOI21_X1 U18059 ( .B1(n16071), .B2(n16169), .A(n14685), .ZN(n14690) );
  OAI21_X1 U18060 ( .B1(n14688), .B2(n14687), .A(n14686), .ZN(n14837) );
  NAND2_X1 U18061 ( .A1(n14837), .A2(n20225), .ZN(n14689) );
  OAI211_X1 U18062 ( .C1(n16069), .C2(n14699), .A(n14690), .B(n14689), .ZN(
        P1_U2979) );
  INV_X1 U18063 ( .A(n14691), .ZN(n16091) );
  NAND2_X1 U18064 ( .A1(n20221), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14852) );
  OAI21_X1 U18065 ( .B1(n14693), .B2(n14692), .A(n14852), .ZN(n14694) );
  AOI21_X1 U18066 ( .B1(n16169), .B2(n16091), .A(n14694), .ZN(n14698) );
  OR2_X1 U18067 ( .A1(n14696), .A2(n14695), .ZN(n14847) );
  NAND3_X1 U18068 ( .A1(n14847), .A2(n14676), .A3(n20225), .ZN(n14697) );
  OAI211_X1 U18069 ( .C1(n14700), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        P1_U2981) );
  AND2_X1 U18070 ( .A1(n14301), .A2(n14701), .ZN(n14716) );
  OAI21_X1 U18071 ( .B1(n14716), .B2(n14703), .A(n14702), .ZN(n16161) );
  INV_X1 U18072 ( .A(n16160), .ZN(n14704) );
  NOR2_X1 U18073 ( .A1(n16161), .A2(n14704), .ZN(n16149) );
  NOR2_X1 U18074 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14857) );
  NOR2_X1 U18075 ( .A1(n16149), .A2(n14857), .ZN(n14707) );
  INV_X1 U18076 ( .A(n16148), .ZN(n14706) );
  AOI22_X1 U18077 ( .A1(n14707), .A2(n14706), .B1(n16149), .B2(n14705), .ZN(
        n14865) );
  INV_X1 U18078 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14708) );
  NOR2_X1 U18079 ( .A1(n20252), .A2(n14708), .ZN(n14860) );
  AOI21_X1 U18080 ( .B1(n20222), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14860), .ZN(n14709) );
  OAI21_X1 U18081 ( .B1(n20230), .B2(n16103), .A(n14709), .ZN(n14710) );
  AOI21_X1 U18082 ( .B1(n14711), .B2(n16192), .A(n14710), .ZN(n14712) );
  OAI21_X1 U18083 ( .B1(n14865), .B2(n20048), .A(n14712), .ZN(P1_U2983) );
  INV_X1 U18084 ( .A(n14713), .ZN(n14715) );
  OAI21_X1 U18085 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14718) );
  XNOR2_X1 U18086 ( .A(n16173), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14717) );
  XNOR2_X1 U18087 ( .A(n14718), .B(n14717), .ZN(n14875) );
  NAND2_X1 U18088 ( .A1(n20221), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14869) );
  NAND2_X1 U18089 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14719) );
  OAI211_X1 U18090 ( .C1(n20230), .C2(n14720), .A(n14869), .B(n14719), .ZN(
        n14721) );
  AOI21_X1 U18091 ( .B1(n14722), .B2(n16192), .A(n14721), .ZN(n14723) );
  OAI21_X1 U18092 ( .B1(n14875), .B2(n20048), .A(n14723), .ZN(P1_U2985) );
  NAND2_X1 U18093 ( .A1(n14724), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14726) );
  XNOR2_X1 U18094 ( .A(n14301), .B(n14727), .ZN(n14725) );
  MUX2_X1 U18095 ( .A(n14726), .B(n14725), .S(n16173), .Z(n14730) );
  INV_X1 U18096 ( .A(n14724), .ZN(n14729) );
  NAND3_X1 U18097 ( .A1(n14729), .A2(n14728), .A3(n14727), .ZN(n16175) );
  NAND2_X1 U18098 ( .A1(n14730), .A2(n16175), .ZN(n16244) );
  INV_X1 U18099 ( .A(n16244), .ZN(n14736) );
  AOI22_X1 U18100 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14731) );
  OAI21_X1 U18101 ( .B1(n20230), .B2(n14732), .A(n14731), .ZN(n14733) );
  AOI21_X1 U18102 ( .B1(n14734), .B2(n16192), .A(n14733), .ZN(n14735) );
  OAI21_X1 U18103 ( .B1(n14736), .B2(n20048), .A(n14735), .ZN(P1_U2989) );
  INV_X1 U18104 ( .A(n14737), .ZN(n14741) );
  AOI21_X1 U18105 ( .B1(n10044), .B2(n14739), .A(n14738), .ZN(n14740) );
  AOI211_X1 U18106 ( .C1(n14742), .C2(n20234), .A(n14741), .B(n14740), .ZN(
        n14743) );
  OAI21_X1 U18107 ( .B1(n14744), .B2(n20250), .A(n14743), .ZN(P1_U3001) );
  INV_X1 U18108 ( .A(n14772), .ZN(n14756) );
  NOR3_X1 U18109 ( .A1(n14756), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14745), .ZN(n14746) );
  AOI211_X1 U18110 ( .C1(n14748), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14747), .B(n14746), .ZN(n14752) );
  INV_X1 U18111 ( .A(n14749), .ZN(n14750) );
  NAND2_X1 U18112 ( .A1(n14750), .A2(n20234), .ZN(n14751) );
  OAI211_X1 U18113 ( .C1(n14753), .C2(n20250), .A(n14752), .B(n14751), .ZN(
        P1_U3002) );
  NOR3_X1 U18114 ( .A1(n14756), .A2(n14755), .A3(n14754), .ZN(n14763) );
  INV_X1 U18115 ( .A(n14757), .ZN(n14759) );
  AOI21_X1 U18116 ( .B1(n14787), .B2(n14759), .A(n14758), .ZN(n14770) );
  NAND2_X1 U18117 ( .A1(n14770), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14761) );
  NAND2_X1 U18118 ( .A1(n14761), .A2(n14760), .ZN(n14762) );
  AOI211_X1 U18119 ( .C1(n14764), .C2(n20234), .A(n14763), .B(n14762), .ZN(
        n14765) );
  OAI21_X1 U18120 ( .B1(n14766), .B2(n20250), .A(n14765), .ZN(P1_U3003) );
  NOR2_X1 U18121 ( .A1(n14767), .A2(n20254), .ZN(n14768) );
  AOI211_X1 U18122 ( .C1(n14770), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14769), .B(n14768), .ZN(n14774) );
  NAND2_X1 U18123 ( .A1(n14772), .A2(n14771), .ZN(n14773) );
  OAI211_X1 U18124 ( .C1(n14775), .C2(n20250), .A(n14774), .B(n14773), .ZN(
        P1_U3004) );
  OAI21_X1 U18125 ( .B1(n14777), .B2(n20254), .A(n14776), .ZN(n14783) );
  INV_X1 U18126 ( .A(n14780), .ZN(n14813) );
  NAND4_X1 U18127 ( .A1(n14813), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n14786), .ZN(n14791) );
  AOI21_X1 U18128 ( .B1(n14791), .B2(n14787), .A(n14778), .ZN(n14782) );
  NOR3_X1 U18129 ( .A1(n14780), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14779), .ZN(n14781) );
  NOR3_X1 U18130 ( .A1(n14783), .A2(n14782), .A3(n14781), .ZN(n14784) );
  OAI21_X1 U18131 ( .B1(n14785), .B2(n20250), .A(n14784), .ZN(P1_U3005) );
  NOR2_X1 U18132 ( .A1(n14787), .A2(n14786), .ZN(n14788) );
  AOI211_X1 U18133 ( .C1(n14790), .C2(n20234), .A(n14789), .B(n14788), .ZN(
        n14792) );
  OAI211_X1 U18134 ( .C1(n14793), .C2(n20250), .A(n14792), .B(n14791), .ZN(
        P1_U3006) );
  NAND2_X1 U18135 ( .A1(n14794), .A2(n20237), .ZN(n14804) );
  INV_X1 U18136 ( .A(n16035), .ZN(n14796) );
  AOI21_X1 U18137 ( .B1(n14796), .B2(n20234), .A(n14795), .ZN(n14803) );
  NAND3_X1 U18138 ( .A1(n14813), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14797), .ZN(n14802) );
  AND2_X1 U18139 ( .A1(n14798), .A2(n14812), .ZN(n14799) );
  OAI21_X1 U18140 ( .B1(n14800), .B2(n14799), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14801) );
  NAND4_X1 U18141 ( .A1(n14804), .A2(n14803), .A3(n14802), .A4(n14801), .ZN(
        P1_U3007) );
  AND2_X1 U18142 ( .A1(n14806), .A2(n14805), .ZN(n14808) );
  OR2_X1 U18143 ( .A1(n14808), .A2(n14807), .ZN(n16134) );
  NOR2_X1 U18144 ( .A1(n16134), .A2(n20254), .ZN(n14809) );
  AOI211_X1 U18145 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14811), .A(
        n14810), .B(n14809), .ZN(n14815) );
  NAND2_X1 U18146 ( .A1(n14813), .A2(n14812), .ZN(n14814) );
  OAI211_X1 U18147 ( .C1(n14816), .C2(n20250), .A(n14815), .B(n14814), .ZN(
        P1_U3008) );
  AND2_X1 U18148 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14848), .ZN(
        n14822) );
  INV_X1 U18149 ( .A(n14822), .ZN(n14817) );
  NAND2_X1 U18150 ( .A1(n16238), .A2(n14817), .ZN(n14818) );
  AND2_X1 U18151 ( .A1(n14868), .A2(n14818), .ZN(n16201) );
  NAND2_X1 U18152 ( .A1(n16238), .A2(n14841), .ZN(n14819) );
  NAND2_X1 U18153 ( .A1(n16201), .A2(n14819), .ZN(n14832) );
  INV_X1 U18154 ( .A(n14820), .ZN(n14821) );
  OAI21_X1 U18155 ( .B1(n16054), .B2(n20254), .A(n14821), .ZN(n14826) );
  NAND2_X1 U18156 ( .A1(n14849), .A2(n14822), .ZN(n16207) );
  INV_X1 U18157 ( .A(n16207), .ZN(n14843) );
  AOI22_X1 U18158 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(n14823), .B2(n14833), .ZN(
        n14824) );
  AND3_X1 U18159 ( .A1(n14843), .A2(n11257), .A3(n14824), .ZN(n14825) );
  AOI211_X1 U18160 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n14832), .A(
        n14826), .B(n14825), .ZN(n14827) );
  OAI21_X1 U18161 ( .B1(n14828), .B2(n20250), .A(n14827), .ZN(P1_U3009) );
  INV_X1 U18162 ( .A(n14829), .ZN(n14836) );
  NOR2_X1 U18163 ( .A1(n16061), .A2(n20254), .ZN(n14830) );
  AOI211_X1 U18164 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n14832), .A(
        n14831), .B(n14830), .ZN(n14835) );
  NAND3_X1 U18165 ( .A1(n14843), .A2(n11257), .A3(n14833), .ZN(n14834) );
  OAI211_X1 U18166 ( .C1(n14836), .C2(n20250), .A(n14835), .B(n14834), .ZN(
        P1_U3010) );
  INV_X1 U18167 ( .A(n14837), .ZN(n14846) );
  INV_X1 U18168 ( .A(n16201), .ZN(n14840) );
  OAI21_X1 U18169 ( .B1(n16068), .B2(n20254), .A(n14838), .ZN(n14839) );
  AOI21_X1 U18170 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14840), .A(
        n14839), .ZN(n14845) );
  NAND3_X1 U18171 ( .A1(n14843), .A2(n14842), .A3(n14841), .ZN(n14844) );
  OAI211_X1 U18172 ( .C1(n14846), .C2(n20250), .A(n14845), .B(n14844), .ZN(
        P1_U3011) );
  NAND3_X1 U18173 ( .A1(n14847), .A2(n14676), .A3(n20237), .ZN(n14855) );
  OAI21_X1 U18174 ( .B1(n14856), .B2(n14848), .A(n14868), .ZN(n16209) );
  NOR2_X1 U18175 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16152), .ZN(
        n14850) );
  NAND2_X1 U18176 ( .A1(n14849), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16216) );
  NOR2_X1 U18177 ( .A1(n14858), .A2(n16216), .ZN(n16210) );
  AOI22_X1 U18178 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16209), .B1(
        n14850), .B2(n16210), .ZN(n14854) );
  INV_X1 U18179 ( .A(n16095), .ZN(n14851) );
  NAND2_X1 U18180 ( .A1(n14851), .A2(n20234), .ZN(n14853) );
  NAND4_X1 U18181 ( .A1(n14855), .A2(n14854), .A3(n14853), .A4(n14852), .ZN(
        P1_U3013) );
  OAI21_X1 U18182 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14856), .A(
        n14868), .ZN(n16214) );
  NOR2_X1 U18183 ( .A1(n14857), .A2(n16216), .ZN(n14859) );
  AOI22_X1 U18184 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16214), .B1(
        n14859), .B2(n14858), .ZN(n14862) );
  INV_X1 U18185 ( .A(n14860), .ZN(n14861) );
  OAI211_X1 U18186 ( .C1(n16109), .C2(n20254), .A(n14862), .B(n14861), .ZN(
        n14863) );
  INV_X1 U18187 ( .A(n14863), .ZN(n14864) );
  OAI21_X1 U18188 ( .B1(n14865), .B2(n20250), .A(n14864), .ZN(P1_U3015) );
  NOR2_X1 U18189 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14866), .ZN(
        n14873) );
  NOR2_X1 U18190 ( .A1(n14867), .A2(n16272), .ZN(n16228) );
  INV_X1 U18191 ( .A(n14868), .ZN(n16223) );
  NAND2_X1 U18192 ( .A1(n16223), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14870) );
  OAI211_X1 U18193 ( .C1(n20254), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        n14872) );
  AOI21_X1 U18194 ( .B1(n14873), .B2(n16228), .A(n14872), .ZN(n14874) );
  OAI21_X1 U18195 ( .B1(n14875), .B2(n20250), .A(n14874), .ZN(P1_U3017) );
  AOI21_X1 U18196 ( .B1(n14878), .B2(n14877), .A(n14876), .ZN(n16232) );
  OAI21_X1 U18197 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14879), .A(
        n16232), .ZN(n14887) );
  OAI21_X1 U18198 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14883) );
  INV_X1 U18199 ( .A(n14883), .ZN(n16172) );
  NAND2_X1 U18200 ( .A1(n14884), .A2(n11245), .ZN(n14885) );
  OAI22_X1 U18201 ( .A1(n16172), .A2(n20250), .B1(n16272), .B2(n14885), .ZN(
        n14886) );
  AOI21_X1 U18202 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14887), .A(
        n14886), .ZN(n14889) );
  NAND2_X1 U18203 ( .A1(n20221), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14888) );
  OAI211_X1 U18204 ( .C1(n20254), .C2(n16119), .A(n14889), .B(n14888), .ZN(
        P1_U3019) );
  NAND2_X1 U18205 ( .A1(n9846), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20417) );
  NAND2_X1 U18206 ( .A1(n20417), .A2(n20680), .ZN(n14891) );
  MUX2_X1 U18207 ( .A(n14891), .B(n20799), .S(n14890), .Z(n14892) );
  OAI21_X1 U18208 ( .B1(n20947), .B2(n20684), .A(n14892), .ZN(n14893) );
  MUX2_X1 U18209 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14893), .S(
        n20953), .Z(P1_U3476) );
  INV_X1 U18210 ( .A(n10333), .ZN(n14896) );
  INV_X1 U18211 ( .A(n14894), .ZN(n14895) );
  NAND2_X1 U18212 ( .A1(n14896), .A2(n14895), .ZN(n14899) );
  OAI22_X1 U18213 ( .A1(n15965), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14899), .B2(n10416), .ZN(n14897) );
  AOI21_X1 U18214 ( .B1(n10546), .B2(n14898), .A(n14897), .ZN(n15969) );
  INV_X1 U18215 ( .A(n14899), .ZN(n14903) );
  INV_X1 U18216 ( .A(n14900), .ZN(n14901) );
  AOI22_X1 U18217 ( .A1(n15999), .A2(n14903), .B1(n14902), .B2(n14901), .ZN(
        n14904) );
  OAI21_X1 U18218 ( .B1(n15969), .B2(n14908), .A(n14904), .ZN(n14905) );
  MUX2_X1 U18219 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14905), .S(
        n14909), .Z(P1_U3473) );
  OAI22_X1 U18220 ( .A1(n10312), .A2(n14908), .B1(n14907), .B2(n14906), .ZN(
        n14910) );
  MUX2_X1 U18221 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14910), .S(
        n14909), .Z(P1_U3469) );
  NAND2_X1 U18222 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  NAND2_X1 U18223 ( .A1(n14914), .A2(n14913), .ZN(n15625) );
  OR2_X1 U18224 ( .A1(n9878), .A2(n14915), .ZN(n14916) );
  NAND2_X1 U18225 ( .A1(n11983), .A2(n14916), .ZN(n15410) );
  AOI22_X1 U18226 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n9962), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19115), .ZN(n14919) );
  AOI22_X1 U18227 ( .A1(n14917), .A2(n19102), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19147), .ZN(n14918) );
  OAI211_X1 U18228 ( .C1(n15410), .C2(n19143), .A(n14919), .B(n14918), .ZN(
        n14921) );
  OAI21_X1 U18229 ( .B1(n15625), .B2(n19149), .A(n14922), .ZN(P2_U2826) );
  INV_X1 U18230 ( .A(n15339), .ZN(n14933) );
  NAND2_X1 U18231 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19147), .ZN(n14924) );
  AOI22_X1 U18232 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n9962), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19115), .ZN(n14923) );
  NAND2_X1 U18233 ( .A1(n14924), .A2(n14923), .ZN(n14925) );
  AOI21_X1 U18234 ( .B1(n15417), .B2(n16306), .A(n14925), .ZN(n14926) );
  OAI21_X1 U18235 ( .B1(n14927), .B2(n19145), .A(n14926), .ZN(n14932) );
  AOI211_X1 U18236 ( .C1(n14930), .C2(n14929), .A(n14928), .B(n19888), .ZN(
        n14931) );
  AOI211_X1 U18237 ( .C1(n19135), .C2(n14933), .A(n14932), .B(n14931), .ZN(
        n14934) );
  INV_X1 U18238 ( .A(n14934), .ZN(P2_U2827) );
  INV_X1 U18239 ( .A(n14936), .ZN(n14937) );
  OAI21_X1 U18240 ( .B1(n14935), .B2(n14938), .A(n14937), .ZN(n15636) );
  NAND2_X1 U18241 ( .A1(n14939), .A2(n14940), .ZN(n14941) );
  NAND2_X1 U18242 ( .A1(n14942), .A2(n14941), .ZN(n15421) );
  AOI22_X1 U18243 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n9962), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19115), .ZN(n14947) );
  OAI22_X1 U18244 ( .A1(n14944), .A2(n19145), .B1(n19126), .B2(n14943), .ZN(
        n14945) );
  INV_X1 U18245 ( .A(n14945), .ZN(n14946) );
  OAI211_X1 U18246 ( .C1(n15421), .C2(n19143), .A(n14947), .B(n14946), .ZN(
        n14951) );
  AOI211_X1 U18247 ( .C1(n15485), .C2(n14949), .A(n14948), .B(n19888), .ZN(
        n14950) );
  NOR2_X1 U18248 ( .A1(n14951), .A2(n14950), .ZN(n14952) );
  OAI21_X1 U18249 ( .B1(n15636), .B2(n19149), .A(n14952), .ZN(P2_U2828) );
  AOI211_X1 U18250 ( .C1(n14955), .C2(n14954), .A(n19888), .B(n14953), .ZN(
        n14956) );
  INV_X1 U18251 ( .A(n14956), .ZN(n14963) );
  NAND2_X1 U18252 ( .A1(n19147), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U18253 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19042), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n9962), .ZN(n14957) );
  OAI211_X1 U18254 ( .C1(n19143), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n14960) );
  AOI21_X1 U18255 ( .B1(n14961), .B2(n19135), .A(n14960), .ZN(n14962) );
  OAI211_X1 U18256 ( .C1(n19145), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        P2_U2830) );
  AOI211_X1 U18257 ( .C1(n15507), .C2(n10133), .A(n14965), .B(n19888), .ZN(
        n14967) );
  OAI22_X1 U18258 ( .A1(n10142), .A2(n19155), .B1(n19937), .B2(n19110), .ZN(
        n14966) );
  AOI211_X1 U18259 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n19147), .A(n14967), .B(
        n14966), .ZN(n14977) );
  AND2_X1 U18260 ( .A1(n15379), .A2(n14968), .ZN(n14970) );
  OR2_X1 U18261 ( .A1(n14970), .A2(n14969), .ZN(n15663) );
  AND2_X1 U18262 ( .A1(n15449), .A2(n14971), .ZN(n14972) );
  NOR2_X1 U18263 ( .A1(n14973), .A2(n14972), .ZN(n15660) );
  INV_X1 U18264 ( .A(n15660), .ZN(n14974) );
  OAI22_X1 U18265 ( .A1(n15663), .A2(n19149), .B1(n14974), .B2(n19143), .ZN(
        n14975) );
  INV_X1 U18266 ( .A(n14975), .ZN(n14976) );
  OAI211_X1 U18267 ( .C1(n14978), .C2(n19145), .A(n14977), .B(n14976), .ZN(
        P2_U2831) );
  OAI21_X1 U18268 ( .B1(n16344), .B2(n14979), .A(n19136), .ZN(n14981) );
  AOI22_X1 U18269 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19042), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n9962), .ZN(n14980) );
  OAI21_X1 U18270 ( .B1(n14982), .B2(n14981), .A(n14980), .ZN(n14983) );
  AOI21_X1 U18271 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n19147), .A(n14983), .ZN(
        n14990) );
  OR2_X1 U18272 ( .A1(n14998), .A2(n14984), .ZN(n14985) );
  NAND2_X1 U18273 ( .A1(n15377), .A2(n14985), .ZN(n15692) );
  OAI21_X1 U18274 ( .B1(n14986), .B2(n15001), .A(n15447), .ZN(n15691) );
  INV_X1 U18275 ( .A(n15691), .ZN(n16320) );
  AOI22_X1 U18276 ( .A1(n16340), .A2(n19135), .B1(n16320), .B2(n16306), .ZN(
        n14989) );
  INV_X1 U18277 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15386) );
  OAI211_X1 U18278 ( .C1(n10246), .C2(n15386), .A(n12779), .B(n19102), .ZN(
        n14988) );
  NAND3_X1 U18279 ( .A1(n14990), .A2(n14989), .A3(n14988), .ZN(P2_U2833) );
  INV_X1 U18280 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14991) );
  OAI22_X1 U18281 ( .A1(n19126), .A2(n14991), .B1(n19932), .B2(n19110), .ZN(
        n14995) );
  AND2_X1 U18282 ( .A1(n11321), .A2(n14992), .ZN(n15007) );
  OAI21_X1 U18283 ( .B1(n15536), .B2(n15007), .A(n19136), .ZN(n14993) );
  AOI21_X1 U18284 ( .B1(n15536), .B2(n15007), .A(n14993), .ZN(n14994) );
  AOI211_X1 U18285 ( .C1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n19115), .A(
        n14995), .B(n14994), .ZN(n15005) );
  AND2_X1 U18286 ( .A1(n15012), .A2(n14996), .ZN(n14997) );
  NOR2_X1 U18287 ( .A1(n14998), .A2(n14997), .ZN(n15701) );
  OR2_X1 U18288 ( .A1(n14999), .A2(n15000), .ZN(n15003) );
  INV_X1 U18289 ( .A(n15001), .ZN(n15002) );
  NAND2_X1 U18290 ( .A1(n15003), .A2(n15002), .ZN(n15703) );
  INV_X1 U18291 ( .A(n15703), .ZN(n15461) );
  AOI22_X1 U18292 ( .A1(n15701), .A2(n19135), .B1(n15461), .B2(n16306), .ZN(
        n15004) );
  OAI211_X1 U18293 ( .C1(n15006), .C2(n19145), .A(n15005), .B(n15004), .ZN(
        P2_U2834) );
  NAND2_X1 U18294 ( .A1(n19117), .A2(n19136), .ZN(n19154) );
  AOI22_X1 U18295 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n9962), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19147), .ZN(n15010) );
  OAI211_X1 U18296 ( .C1(n15008), .C2(n15552), .A(n19136), .B(n15007), .ZN(
        n15009) );
  OAI211_X1 U18297 ( .C1(n15552), .C2(n19154), .A(n15010), .B(n15009), .ZN(
        n15011) );
  AOI21_X1 U18298 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19115), .A(
        n15011), .ZN(n15020) );
  INV_X1 U18299 ( .A(n15012), .ZN(n15013) );
  AOI21_X1 U18300 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15721) );
  NOR2_X1 U18301 ( .A1(n15017), .A2(n15016), .ZN(n15018) );
  OR2_X1 U18302 ( .A1(n14999), .A2(n15018), .ZN(n15714) );
  INV_X1 U18303 ( .A(n15714), .ZN(n16327) );
  AOI22_X1 U18304 ( .A1(n15721), .A2(n19135), .B1(n16327), .B2(n16306), .ZN(
        n15019) );
  OAI211_X1 U18305 ( .C1(n15021), .C2(n19145), .A(n15020), .B(n15019), .ZN(
        P2_U2835) );
  NOR2_X1 U18306 ( .A1(n19117), .A2(n15022), .ZN(n19035) );
  XNOR2_X1 U18307 ( .A(n19035), .B(n15577), .ZN(n15023) );
  NAND2_X1 U18308 ( .A1(n15023), .A2(n19136), .ZN(n15032) );
  NOR2_X1 U18309 ( .A1(n15744), .A2(n19149), .ZN(n15030) );
  INV_X1 U18310 ( .A(n15024), .ZN(n15025) );
  AOI21_X1 U18311 ( .B1(n15026), .B2(n13786), .A(n15025), .ZN(n16333) );
  INV_X1 U18312 ( .A(n16333), .ZN(n15028) );
  AOI22_X1 U18313 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19042), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19147), .ZN(n15027) );
  OAI211_X1 U18314 ( .C1(n19143), .C2(n15028), .A(n15027), .B(n19324), .ZN(
        n15029) );
  OAI211_X1 U18315 ( .C1(n19145), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        P2_U2837) );
  INV_X1 U18316 ( .A(n15034), .ZN(n19161) );
  NOR2_X1 U18317 ( .A1(n15036), .A2(n19161), .ZN(n19052) );
  INV_X1 U18318 ( .A(n16352), .ZN(n15035) );
  OAI211_X1 U18319 ( .C1(n19117), .C2(n15036), .A(n15035), .B(n19136), .ZN(
        n15045) );
  NOR2_X1 U18320 ( .A1(n19149), .A2(n16346), .ZN(n15043) );
  NOR2_X1 U18321 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  OR2_X1 U18322 ( .A1(n15040), .A2(n15039), .ZN(n19170) );
  AOI22_X1 U18323 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n9962), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19115), .ZN(n15041) );
  OAI211_X1 U18324 ( .C1(n19143), .C2(n19170), .A(n15041), .B(n19324), .ZN(
        n15042) );
  AOI211_X1 U18325 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19147), .A(n15043), .B(
        n15042), .ZN(n15044) );
  OAI211_X1 U18326 ( .C1(n15046), .C2(n19145), .A(n15045), .B(n15044), .ZN(
        n15047) );
  AOI21_X1 U18327 ( .B1(n19052), .B2(n16352), .A(n15047), .ZN(n15048) );
  INV_X1 U18328 ( .A(n15048), .ZN(P2_U2839) );
  AOI211_X1 U18329 ( .C1(n19140), .C2(n15050), .A(n19117), .B(n15049), .ZN(
        n15873) );
  NAND2_X1 U18330 ( .A1(n15873), .A2(n19136), .ZN(n15059) );
  INV_X1 U18331 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15053) );
  INV_X1 U18332 ( .A(n19154), .ZN(n19046) );
  AOI22_X1 U18333 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n9962), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n19147), .ZN(n15051) );
  OAI21_X1 U18334 ( .B1(n19155), .B2(n15053), .A(n15051), .ZN(n15052) );
  AOI21_X1 U18335 ( .B1(n15053), .B2(n19046), .A(n15052), .ZN(n15055) );
  NAND2_X1 U18336 ( .A1(n16306), .A2(n19994), .ZN(n15054) );
  OAI211_X1 U18337 ( .C1(n19145), .C2(n15056), .A(n15055), .B(n15054), .ZN(
        n15057) );
  AOI21_X1 U18338 ( .B1(n13119), .B2(n19135), .A(n15057), .ZN(n15058) );
  OAI211_X1 U18339 ( .C1(n19990), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        P2_U2854) );
  INV_X1 U18340 ( .A(n15061), .ZN(n15062) );
  NAND2_X1 U18341 ( .A1(n15062), .A2(n15395), .ZN(n15063) );
  OAI21_X1 U18342 ( .B1(n15395), .B2(n11990), .A(n15063), .ZN(P2_U2856) );
  INV_X1 U18343 ( .A(n15064), .ZN(n15148) );
  NAND2_X1 U18344 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n15066) );
  AOI22_X1 U18345 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n15144), .ZN(n15065) );
  OAI211_X1 U18346 ( .C1(n15148), .C2(n15245), .A(n15066), .B(n15065), .ZN(
        n15067) );
  INV_X1 U18347 ( .A(n15067), .ZN(n15071) );
  NAND2_X1 U18348 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n15070) );
  NAND2_X1 U18349 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n15069) );
  NAND2_X1 U18350 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n15068) );
  AND4_X1 U18351 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15079) );
  AOI22_X1 U18352 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n15101), .B1(
        n15156), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15078) );
  AOI22_X1 U18353 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15075) );
  NAND2_X1 U18354 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15074) );
  NAND2_X1 U18355 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n15073) );
  NAND2_X1 U18356 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n15072) );
  AND4_X1 U18357 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        n15077) );
  AOI22_X1 U18358 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15076) );
  NAND4_X1 U18359 ( .A1(n15079), .A2(n15078), .A3(n15077), .A4(n15076), .ZN(
        n15392) );
  NAND2_X1 U18360 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n15081) );
  AOI22_X1 U18361 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n15144), .ZN(n15080) );
  OAI211_X1 U18362 ( .C1(n15148), .C2(n15269), .A(n15081), .B(n15080), .ZN(
        n15082) );
  INV_X1 U18363 ( .A(n15082), .ZN(n15086) );
  NAND2_X1 U18364 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n15085) );
  NAND2_X1 U18365 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15084) );
  NAND2_X1 U18366 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n15083) );
  AND4_X1 U18367 ( .A1(n15086), .A2(n15085), .A3(n15084), .A4(n15083), .ZN(
        n15094) );
  AOI22_X1 U18368 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n15101), .B1(
        n15156), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U18369 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U18370 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15089) );
  NAND2_X1 U18371 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n15088) );
  NAND2_X1 U18372 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n15087) );
  AND4_X1 U18373 ( .A1(n15090), .A2(n15089), .A3(n15088), .A4(n15087), .ZN(
        n15092) );
  AOI22_X1 U18374 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15091) );
  NAND4_X1 U18375 ( .A1(n15094), .A2(n15093), .A3(n15092), .A4(n15091), .ZN(
        n15388) );
  INV_X1 U18376 ( .A(n15151), .ZN(n15099) );
  AOI22_X1 U18377 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15150), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15098) );
  INV_X1 U18378 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15287) );
  AOI22_X1 U18379 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n15144), .ZN(n15095) );
  OAI21_X1 U18380 ( .B1(n15148), .B2(n15287), .A(n15095), .ZN(n15096) );
  AOI21_X1 U18381 ( .B1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n15143), .A(
        n15096), .ZN(n15097) );
  OAI211_X1 U18382 ( .C1(n15100), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        n15118) );
  INV_X1 U18383 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15295) );
  INV_X1 U18384 ( .A(n15101), .ZN(n15104) );
  INV_X1 U18385 ( .A(n15156), .ZN(n15103) );
  OAI22_X1 U18386 ( .A1(n15295), .A2(n15104), .B1(n15103), .B2(n15102), .ZN(
        n15117) );
  AOI22_X1 U18387 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15108) );
  NAND2_X1 U18388 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n15107) );
  NAND2_X1 U18389 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n15106) );
  NAND2_X1 U18390 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n15105) );
  NAND4_X1 U18391 ( .A1(n15108), .A2(n15107), .A3(n15106), .A4(n15105), .ZN(
        n15116) );
  INV_X1 U18392 ( .A(n15109), .ZN(n15114) );
  INV_X1 U18393 ( .A(n15110), .ZN(n15112) );
  OAI22_X1 U18394 ( .A1(n15114), .A2(n15113), .B1(n15112), .B2(n15111), .ZN(
        n15115) );
  NOR4_X1 U18395 ( .A1(n15118), .A2(n15117), .A3(n15116), .A4(n15115), .ZN(
        n15382) );
  INV_X1 U18396 ( .A(n15120), .ZN(n15318) );
  AOI22_X1 U18397 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15132) );
  NAND2_X1 U18398 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15122) );
  NAND2_X1 U18399 ( .A1(n15123), .A2(n15122), .ZN(n15311) );
  INV_X1 U18400 ( .A(n15308), .ZN(n15313) );
  INV_X1 U18401 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15124) );
  OR2_X1 U18402 ( .A1(n15313), .A2(n15124), .ZN(n15125) );
  OAI211_X1 U18403 ( .C1(n15121), .C2(n19526), .A(n15311), .B(n15125), .ZN(
        n15126) );
  INV_X1 U18404 ( .A(n15126), .ZN(n15131) );
  AOI22_X1 U18405 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15130) );
  AOI22_X1 U18406 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15128), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15129) );
  NAND4_X1 U18407 ( .A1(n15132), .A2(n15131), .A3(n15130), .A4(n15129), .ZN(
        n15142) );
  AOI22_X1 U18408 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15308), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15140) );
  INV_X1 U18409 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15135) );
  INV_X1 U18410 ( .A(n15311), .ZN(n15293) );
  INV_X1 U18411 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15133) );
  OR2_X1 U18412 ( .A1(n15120), .A2(n15133), .ZN(n15134) );
  OAI211_X1 U18413 ( .C1(n15127), .C2(n15135), .A(n15293), .B(n15134), .ZN(
        n15136) );
  INV_X1 U18414 ( .A(n15136), .ZN(n15139) );
  AOI22_X1 U18415 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U18416 ( .A1(n11627), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15128), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15137) );
  NAND4_X1 U18417 ( .A1(n15140), .A2(n15139), .A3(n15138), .A4(n15137), .ZN(
        n15141) );
  NAND2_X1 U18418 ( .A1(n15910), .A2(n15192), .ZN(n15169) );
  INV_X1 U18419 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U18420 ( .A1(n15143), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n15147) );
  AOI22_X1 U18421 ( .A1(n15145), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n15144), .ZN(n15146) );
  OAI211_X1 U18422 ( .C1(n15148), .C2(n15312), .A(n15147), .B(n15146), .ZN(
        n15149) );
  INV_X1 U18423 ( .A(n15149), .ZN(n15155) );
  NAND2_X1 U18424 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n15154) );
  NAND2_X1 U18425 ( .A1(n15150), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n15153) );
  NAND2_X1 U18426 ( .A1(n15151), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n15152) );
  AND4_X1 U18427 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15168) );
  AOI22_X1 U18428 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n15101), .B1(
        n15156), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U18429 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n15158), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15164) );
  NAND2_X1 U18430 ( .A1(n11916), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n15163) );
  NAND2_X1 U18431 ( .A1(n15159), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n15162) );
  NAND2_X1 U18432 ( .A1(n15160), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n15161) );
  AND4_X1 U18433 ( .A1(n15164), .A2(n15163), .A3(n15162), .A4(n15161), .ZN(
        n15166) );
  AOI22_X1 U18434 ( .A1(n15109), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15165) );
  NAND4_X1 U18435 ( .A1(n15168), .A2(n15167), .A3(n15166), .A4(n15165), .ZN(
        n15172) );
  XNOR2_X1 U18436 ( .A(n15169), .B(n15172), .ZN(n15195) );
  NAND2_X1 U18437 ( .A1(n15191), .A2(n15192), .ZN(n15373) );
  NOR2_X2 U18438 ( .A1(n15372), .A2(n15171), .ZN(n15365) );
  AND2_X1 U18439 ( .A1(n15172), .A2(n15192), .ZN(n15189) );
  AOI22_X1 U18440 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15179) );
  AOI22_X1 U18441 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U18442 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U18443 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n15173) );
  OAI211_X1 U18444 ( .C1(n15313), .C2(n15174), .A(n15173), .B(n15311), .ZN(
        n15175) );
  INV_X1 U18445 ( .A(n15175), .ZN(n15176) );
  NAND4_X1 U18446 ( .A1(n15179), .A2(n15178), .A3(n15177), .A4(n15176), .ZN(
        n15188) );
  AOI22_X1 U18447 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U18448 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15185) );
  AOI22_X1 U18449 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15184) );
  NAND2_X1 U18450 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15180) );
  OAI211_X1 U18451 ( .C1(n15313), .C2(n15181), .A(n15180), .B(n15293), .ZN(
        n15182) );
  INV_X1 U18452 ( .A(n15182), .ZN(n15183) );
  NAND4_X1 U18453 ( .A1(n15186), .A2(n15185), .A3(n15184), .A4(n15183), .ZN(
        n15187) );
  AND2_X1 U18454 ( .A1(n15188), .A2(n15187), .ZN(n15190) );
  NAND2_X1 U18455 ( .A1(n15189), .A2(n15190), .ZN(n15214) );
  OAI211_X1 U18456 ( .C1(n15189), .C2(n15190), .A(n15216), .B(n15214), .ZN(
        n15364) );
  NOR2_X1 U18457 ( .A1(n15365), .A2(n15364), .ZN(n15363) );
  NAND2_X1 U18458 ( .A1(n15191), .A2(n15190), .ZN(n15367) );
  INV_X1 U18459 ( .A(n15192), .ZN(n15193) );
  NOR2_X1 U18460 ( .A1(n15367), .A2(n15193), .ZN(n15194) );
  AOI22_X1 U18461 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15320), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15203) );
  AOI22_X1 U18462 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15202) );
  AOI22_X1 U18463 ( .A1(n11627), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15201) );
  INV_X1 U18464 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U18465 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15197) );
  OAI211_X1 U18466 ( .C1(n15313), .C2(n15198), .A(n15197), .B(n15293), .ZN(
        n15199) );
  INV_X1 U18467 ( .A(n15199), .ZN(n15200) );
  NAND4_X1 U18468 ( .A1(n15203), .A2(n15202), .A3(n15201), .A4(n15200), .ZN(
        n15213) );
  AOI22_X1 U18469 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15211) );
  INV_X1 U18470 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15206) );
  OR2_X1 U18471 ( .A1(n15313), .A2(n15204), .ZN(n15205) );
  OAI211_X1 U18472 ( .C1(n15127), .C2(n15206), .A(n15311), .B(n15205), .ZN(
        n15207) );
  INV_X1 U18473 ( .A(n15207), .ZN(n15210) );
  AOI22_X1 U18474 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15209) );
  AOI22_X1 U18475 ( .A1(n11627), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15128), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15208) );
  NAND4_X1 U18476 ( .A1(n15211), .A2(n15210), .A3(n15209), .A4(n15208), .ZN(
        n15212) );
  NAND2_X1 U18477 ( .A1(n15213), .A2(n15212), .ZN(n15218) );
  NAND2_X1 U18478 ( .A1(n15214), .A2(n15218), .ZN(n15215) );
  NAND3_X1 U18479 ( .A1(n15240), .A2(n15216), .A3(n15215), .ZN(n15219) );
  INV_X1 U18480 ( .A(n15219), .ZN(n15217) );
  NOR2_X1 U18481 ( .A1(n15910), .A2(n15218), .ZN(n15358) );
  INV_X1 U18482 ( .A(n15240), .ZN(n15238) );
  AOI22_X1 U18483 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U18484 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U18485 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15226) );
  NAND2_X1 U18486 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n15222) );
  OAI211_X1 U18487 ( .C1(n15313), .C2(n15223), .A(n15222), .B(n15311), .ZN(
        n15224) );
  INV_X1 U18488 ( .A(n15224), .ZN(n15225) );
  NAND4_X1 U18489 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15237) );
  AOI22_X1 U18490 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U18491 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U18492 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15233) );
  NAND2_X1 U18493 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n15229) );
  OAI211_X1 U18494 ( .C1(n15313), .C2(n15230), .A(n15229), .B(n15293), .ZN(
        n15231) );
  INV_X1 U18495 ( .A(n15231), .ZN(n15232) );
  NAND4_X1 U18496 ( .A1(n15235), .A2(n15234), .A3(n15233), .A4(n15232), .ZN(
        n15236) );
  AND2_X1 U18497 ( .A1(n15237), .A2(n15236), .ZN(n15239) );
  NAND2_X1 U18498 ( .A1(n15238), .A2(n15239), .ZN(n15262) );
  INV_X1 U18499 ( .A(n15239), .ZN(n15242) );
  AOI21_X1 U18500 ( .B1(n15240), .B2(n15242), .A(n15261), .ZN(n15241) );
  NAND2_X1 U18501 ( .A1(n15262), .A2(n15241), .ZN(n15243) );
  NOR2_X1 U18502 ( .A1(n15910), .A2(n15242), .ZN(n15350) );
  AOI22_X1 U18503 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U18504 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15249) );
  AOI22_X1 U18505 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15248) );
  NAND2_X1 U18506 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n15244) );
  OAI211_X1 U18507 ( .C1(n15313), .C2(n15245), .A(n15244), .B(n15311), .ZN(
        n15246) );
  INV_X1 U18508 ( .A(n15246), .ZN(n15247) );
  NAND4_X1 U18509 ( .A1(n15250), .A2(n15249), .A3(n15248), .A4(n15247), .ZN(
        n15259) );
  AOI22_X1 U18510 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U18511 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U18512 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15255) );
  INV_X1 U18513 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U18514 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15251) );
  OAI211_X1 U18515 ( .C1(n15313), .C2(n15252), .A(n15251), .B(n15293), .ZN(
        n15253) );
  INV_X1 U18516 ( .A(n15253), .ZN(n15254) );
  NAND4_X1 U18517 ( .A1(n15257), .A2(n15256), .A3(n15255), .A4(n15254), .ZN(
        n15258) );
  AND2_X1 U18518 ( .A1(n15259), .A2(n15258), .ZN(n15266) );
  INV_X1 U18519 ( .A(n15266), .ZN(n15263) );
  INV_X1 U18520 ( .A(n15262), .ZN(n15260) );
  AOI211_X1 U18521 ( .C1(n15263), .C2(n15262), .A(n15261), .B(n15284), .ZN(
        n15264) );
  NAND2_X1 U18522 ( .A1(n15265), .A2(n15264), .ZN(n15267) );
  OAI21_X1 U18523 ( .B1(n15265), .B2(n15264), .A(n15267), .ZN(n15344) );
  NAND2_X1 U18524 ( .A1(n15191), .A2(n15266), .ZN(n15343) );
  AOI22_X1 U18525 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U18526 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U18527 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15272) );
  NAND2_X1 U18528 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n15268) );
  OAI211_X1 U18529 ( .C1(n15313), .C2(n15269), .A(n15268), .B(n15311), .ZN(
        n15270) );
  INV_X1 U18530 ( .A(n15270), .ZN(n15271) );
  NAND4_X1 U18531 ( .A1(n15274), .A2(n15273), .A3(n15272), .A4(n15271), .ZN(
        n15283) );
  AOI22_X1 U18532 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15281) );
  AOI22_X1 U18533 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U18534 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U18535 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15275) );
  OAI211_X1 U18536 ( .C1(n15313), .C2(n15276), .A(n15275), .B(n15293), .ZN(
        n15277) );
  INV_X1 U18537 ( .A(n15277), .ZN(n15278) );
  NAND4_X1 U18538 ( .A1(n15281), .A2(n15280), .A3(n15279), .A4(n15278), .ZN(
        n15282) );
  AND2_X1 U18539 ( .A1(n15283), .A2(n15282), .ZN(n15337) );
  INV_X1 U18540 ( .A(n15284), .ZN(n15336) );
  NAND2_X1 U18541 ( .A1(n15910), .A2(n15337), .ZN(n15285) );
  NOR2_X1 U18542 ( .A1(n15336), .A2(n15285), .ZN(n15304) );
  AOI22_X1 U18543 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11627), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U18544 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15291) );
  AOI22_X1 U18545 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15128), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U18546 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n15286) );
  OAI211_X1 U18547 ( .C1(n15313), .C2(n15287), .A(n15286), .B(n15311), .ZN(
        n15288) );
  INV_X1 U18548 ( .A(n15288), .ZN(n15289) );
  NAND4_X1 U18549 ( .A1(n15292), .A2(n15291), .A3(n15290), .A4(n15289), .ZN(
        n15302) );
  AOI22_X1 U18550 ( .A1(n11643), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15320), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U18551 ( .A1(n11627), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15318), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U18552 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15298) );
  NAND2_X1 U18553 ( .A1(n15128), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n15294) );
  OAI211_X1 U18554 ( .C1(n15313), .C2(n15295), .A(n15294), .B(n15293), .ZN(
        n15296) );
  INV_X1 U18555 ( .A(n15296), .ZN(n15297) );
  NAND4_X1 U18556 ( .A1(n15300), .A2(n15299), .A3(n15298), .A4(n15297), .ZN(
        n15301) );
  AND2_X1 U18557 ( .A1(n15302), .A2(n15301), .ZN(n15303) );
  NAND2_X1 U18558 ( .A1(n15304), .A2(n15303), .ZN(n15305) );
  OAI21_X1 U18559 ( .B1(n15304), .B2(n15303), .A(n15305), .ZN(n15333) );
  AOI22_X1 U18560 ( .A1(n11635), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15307) );
  AOI22_X1 U18561 ( .A1(n15318), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15128), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15306) );
  NAND2_X1 U18562 ( .A1(n15307), .A2(n15306), .ZN(n15326) );
  AOI22_X1 U18563 ( .A1(n11627), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15320), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15310) );
  AOI21_X1 U18564 ( .B1(n15308), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15311), .ZN(n15309) );
  OAI211_X1 U18565 ( .C1(n15127), .C2(n21090), .A(n15310), .B(n15309), .ZN(
        n15325) );
  OAI21_X1 U18566 ( .B1(n15313), .B2(n15312), .A(n15311), .ZN(n15317) );
  INV_X1 U18567 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15315) );
  INV_X1 U18568 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15314) );
  OAI22_X1 U18569 ( .A1(n15119), .A2(n15315), .B1(n15121), .B2(n15314), .ZN(
        n15316) );
  AOI211_X1 U18570 ( .C1(n11643), .C2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15317), .B(n15316), .ZN(n15323) );
  AOI22_X1 U18571 ( .A1(n15318), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15128), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U18572 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15319), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15321) );
  NAND3_X1 U18573 ( .A1(n15323), .A2(n15322), .A3(n15321), .ZN(n15324) );
  OAI21_X1 U18574 ( .B1(n15326), .B2(n15325), .A(n15324), .ZN(n15327) );
  XNOR2_X1 U18575 ( .A(n15328), .B(n15327), .ZN(n15408) );
  NAND2_X1 U18576 ( .A1(n15329), .A2(n15395), .ZN(n15331) );
  NAND2_X1 U18577 ( .A1(n15370), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15330) );
  OAI211_X1 U18578 ( .C1(n15408), .C2(n15397), .A(n15331), .B(n15330), .ZN(
        P2_U2857) );
  NAND2_X1 U18579 ( .A1(n15332), .A2(n15333), .ZN(n15409) );
  NAND3_X1 U18580 ( .A1(n9851), .A2(n15383), .A3(n15409), .ZN(n15335) );
  NAND2_X1 U18581 ( .A1(n15368), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15334) );
  OAI211_X1 U18582 ( .C1(n15625), .C2(n15370), .A(n15335), .B(n15334), .ZN(
        P2_U2858) );
  NAND2_X1 U18583 ( .A1(n15267), .A2(n15336), .ZN(n15338) );
  XNOR2_X1 U18584 ( .A(n15338), .B(n15337), .ZN(n15420) );
  NOR2_X1 U18585 ( .A1(n15339), .A2(n15368), .ZN(n15340) );
  AOI21_X1 U18586 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15370), .A(n15340), .ZN(
        n15341) );
  OAI21_X1 U18587 ( .B1(n15420), .B2(n15397), .A(n15341), .ZN(P2_U2859) );
  AOI21_X1 U18588 ( .B1(n15344), .B2(n15343), .A(n15342), .ZN(n15345) );
  INV_X1 U18589 ( .A(n15345), .ZN(n15426) );
  NOR2_X1 U18590 ( .A1(n15636), .A2(n15368), .ZN(n15346) );
  AOI21_X1 U18591 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15370), .A(n15346), .ZN(
        n15347) );
  OAI21_X1 U18592 ( .B1(n15426), .B2(n15397), .A(n15347), .ZN(P2_U2860) );
  OAI21_X1 U18593 ( .B1(n15348), .B2(n15350), .A(n15349), .ZN(n15434) );
  INV_X1 U18594 ( .A(n15351), .ZN(n15354) );
  INV_X1 U18595 ( .A(n15352), .ZN(n15353) );
  AOI21_X1 U18596 ( .B1(n15354), .B2(n15353), .A(n14935), .ZN(n16301) );
  INV_X1 U18597 ( .A(n16301), .ZN(n15651) );
  NOR2_X1 U18598 ( .A1(n15651), .A2(n15368), .ZN(n15355) );
  AOI21_X1 U18599 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15370), .A(n15355), .ZN(
        n15356) );
  OAI21_X1 U18600 ( .B1(n15434), .B2(n15397), .A(n15356), .ZN(P2_U2861) );
  OAI21_X1 U18601 ( .B1(n15359), .B2(n15358), .A(n15357), .ZN(n15440) );
  MUX2_X1 U18602 ( .A(n15361), .B(n15360), .S(n15368), .Z(n15362) );
  OAI21_X1 U18603 ( .B1(n15440), .B2(n15397), .A(n15362), .ZN(P2_U2862) );
  AOI21_X1 U18604 ( .B1(n15365), .B2(n15364), .A(n15363), .ZN(n15366) );
  XOR2_X1 U18605 ( .A(n15367), .B(n15366), .Z(n15445) );
  NOR2_X1 U18606 ( .A1(n15663), .A2(n15368), .ZN(n15369) );
  AOI21_X1 U18607 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15370), .A(n15369), .ZN(
        n15371) );
  OAI21_X1 U18608 ( .B1(n15445), .B2(n15397), .A(n15371), .ZN(P2_U2863) );
  AOI21_X1 U18609 ( .B1(n15374), .B2(n15373), .A(n15372), .ZN(n15375) );
  INV_X1 U18610 ( .A(n15375), .ZN(n15454) );
  NAND2_X1 U18611 ( .A1(n15377), .A2(n15376), .ZN(n15378) );
  NAND2_X1 U18612 ( .A1(n15379), .A2(n15378), .ZN(n16313) );
  INV_X1 U18613 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15380) );
  MUX2_X1 U18614 ( .A(n16313), .B(n15380), .S(n15368), .Z(n15381) );
  OAI21_X1 U18615 ( .B1(n15454), .B2(n15397), .A(n15381), .ZN(P2_U2864) );
  AOI21_X1 U18616 ( .B1(n15382), .B2(n15387), .A(n15170), .ZN(n16321) );
  NAND2_X1 U18617 ( .A1(n16321), .A2(n15383), .ZN(n15385) );
  NAND2_X1 U18618 ( .A1(n16340), .A2(n15395), .ZN(n15384) );
  OAI211_X1 U18619 ( .C1(n15395), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        P2_U2865) );
  OAI21_X1 U18620 ( .B1(n15391), .B2(n15388), .A(n15387), .ZN(n15463) );
  NAND2_X1 U18621 ( .A1(n15368), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15390) );
  NAND2_X1 U18622 ( .A1(n15701), .A2(n15395), .ZN(n15389) );
  OAI211_X1 U18623 ( .C1(n15463), .C2(n15397), .A(n15390), .B(n15389), .ZN(
        P2_U2866) );
  OAI21_X1 U18624 ( .B1(n9856), .B2(n15392), .A(n10207), .ZN(n16326) );
  NOR2_X1 U18625 ( .A1(n15395), .A2(n15393), .ZN(n15394) );
  AOI21_X1 U18626 ( .B1(n15721), .B2(n15395), .A(n15394), .ZN(n15396) );
  OAI21_X1 U18627 ( .B1(n16326), .B2(n15397), .A(n15396), .ZN(P2_U2867) );
  NAND2_X1 U18628 ( .A1(n15399), .A2(BUF2_REG_14__SCAN_IN), .ZN(n15401) );
  INV_X1 U18629 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n15398) );
  OR2_X1 U18630 ( .A1(n15399), .A2(n15398), .ZN(n15400) );
  NAND2_X1 U18631 ( .A1(n15401), .A2(n15400), .ZN(n19302) );
  INV_X1 U18632 ( .A(n19302), .ZN(n15403) );
  INV_X1 U18633 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n15402) );
  OAI22_X1 U18634 ( .A1(n16319), .A2(n15403), .B1(n19198), .B2(n15402), .ZN(
        n15404) );
  AOI21_X1 U18635 ( .B1(n15405), .B2(n19223), .A(n15404), .ZN(n15407) );
  AOI22_X1 U18636 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19169), .B1(n19168), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n15406) );
  OAI211_X1 U18637 ( .C1(n15408), .C2(n19227), .A(n15407), .B(n15406), .ZN(
        P2_U2889) );
  NAND3_X1 U18638 ( .A1(n9851), .A2(n19210), .A3(n15409), .ZN(n15414) );
  INV_X1 U18639 ( .A(n15410), .ZN(n15621) );
  INV_X1 U18640 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19242) );
  OAI22_X1 U18641 ( .A1(n16319), .A2(n19181), .B1(n19198), .B2(n19242), .ZN(
        n15411) );
  AOI21_X1 U18642 ( .B1(n19223), .B2(n15621), .A(n15411), .ZN(n15413) );
  AOI22_X1 U18643 ( .A1(n19169), .A2(BUF1_REG_29__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15412) );
  NAND3_X1 U18644 ( .A1(n15414), .A2(n15413), .A3(n15412), .ZN(P2_U2890) );
  INV_X1 U18645 ( .A(n19183), .ZN(n15415) );
  OAI22_X1 U18646 ( .A1(n16319), .A2(n15415), .B1(n19198), .B2(n19244), .ZN(
        n15416) );
  AOI21_X1 U18647 ( .B1(n15417), .B2(n19223), .A(n15416), .ZN(n15419) );
  AOI22_X1 U18648 ( .A1(n19169), .A2(BUF1_REG_28__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15418) );
  OAI211_X1 U18649 ( .C1(n15420), .C2(n19227), .A(n15419), .B(n15418), .ZN(
        P2_U2891) );
  INV_X1 U18650 ( .A(n15421), .ZN(n15634) );
  INV_X1 U18651 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n21193) );
  OAI22_X1 U18652 ( .A1(n16319), .A2(n19186), .B1(n19198), .B2(n21193), .ZN(
        n15424) );
  INV_X1 U18653 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15422) );
  OAI22_X1 U18654 ( .A1(n15458), .A2(n20306), .B1(n15456), .B2(n15422), .ZN(
        n15423) );
  AOI211_X1 U18655 ( .C1(n19223), .C2(n15634), .A(n15424), .B(n15423), .ZN(
        n15425) );
  OAI21_X1 U18656 ( .B1(n15426), .B2(n19227), .A(n15425), .ZN(P2_U2892) );
  OR2_X1 U18657 ( .A1(n15428), .A2(n15427), .ZN(n15429) );
  AND2_X1 U18658 ( .A1(n14939), .A2(n15429), .ZN(n16305) );
  INV_X1 U18659 ( .A(n19188), .ZN(n15430) );
  OAI22_X1 U18660 ( .A1(n16319), .A2(n15430), .B1(n19198), .B2(n19247), .ZN(
        n15431) );
  AOI21_X1 U18661 ( .B1(n19223), .B2(n16305), .A(n15431), .ZN(n15433) );
  AOI22_X1 U18662 ( .A1(n19169), .A2(BUF1_REG_26__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15432) );
  OAI211_X1 U18663 ( .C1(n15434), .C2(n19227), .A(n15433), .B(n15432), .ZN(
        P2_U2893) );
  INV_X1 U18664 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19249) );
  OAI22_X1 U18665 ( .A1(n16319), .A2(n19191), .B1(n19198), .B2(n19249), .ZN(
        n15437) );
  INV_X1 U18666 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15435) );
  OAI22_X1 U18667 ( .A1(n15458), .A2(n20286), .B1(n15456), .B2(n15435), .ZN(
        n15436) );
  AOI211_X1 U18668 ( .C1(n19223), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        n15439) );
  OAI21_X1 U18669 ( .B1(n15440), .B2(n19227), .A(n15439), .ZN(P2_U2894) );
  INV_X1 U18670 ( .A(n19193), .ZN(n15441) );
  OAI22_X1 U18671 ( .A1(n16319), .A2(n15441), .B1(n19198), .B2(n19251), .ZN(
        n15442) );
  AOI21_X1 U18672 ( .B1(n19223), .B2(n15660), .A(n15442), .ZN(n15444) );
  AOI22_X1 U18673 ( .A1(n19169), .A2(BUF1_REG_24__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15443) );
  OAI211_X1 U18674 ( .C1(n15445), .C2(n19227), .A(n15444), .B(n15443), .ZN(
        P2_U2895) );
  NAND2_X1 U18675 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  NAND2_X1 U18676 ( .A1(n15449), .A2(n15448), .ZN(n16318) );
  INV_X1 U18677 ( .A(n16318), .ZN(n15671) );
  INV_X1 U18678 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19253) );
  OAI22_X1 U18679 ( .A1(n16319), .A2(n19357), .B1(n19253), .B2(n19198), .ZN(
        n15452) );
  INV_X1 U18680 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15450) );
  OAI22_X1 U18681 ( .A1(n15458), .A2(n20336), .B1(n15456), .B2(n15450), .ZN(
        n15451) );
  AOI211_X1 U18682 ( .C1(n19223), .C2(n15671), .A(n15452), .B(n15451), .ZN(
        n15453) );
  OAI21_X1 U18683 ( .B1(n15454), .B2(n19227), .A(n15453), .ZN(P2_U2896) );
  INV_X1 U18684 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19258) );
  OAI22_X1 U18685 ( .A1(n16319), .A2(n19343), .B1(n19198), .B2(n19258), .ZN(
        n15460) );
  INV_X1 U18686 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15457) );
  INV_X1 U18687 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15455) );
  OAI22_X1 U18688 ( .A1(n15458), .A2(n15457), .B1(n15456), .B2(n15455), .ZN(
        n15459) );
  AOI211_X1 U18689 ( .C1(n19223), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15462) );
  OAI21_X1 U18690 ( .B1(n15463), .B2(n19227), .A(n15462), .ZN(P2_U2898) );
  NAND2_X1 U18691 ( .A1(n15465), .A2(n15464), .ZN(n15467) );
  AOI21_X1 U18692 ( .B1(n14354), .B2(n15615), .A(n15468), .ZN(n15627) );
  OR2_X1 U18693 ( .A1(n19124), .A2(n19945), .ZN(n15619) );
  OAI21_X1 U18694 ( .B1(n16429), .B2(n15469), .A(n15619), .ZN(n15470) );
  AOI21_X1 U18695 ( .B1(n16420), .B2(n15471), .A(n15470), .ZN(n15472) );
  OAI21_X1 U18696 ( .B1(n15625), .B2(n16393), .A(n15472), .ZN(n15473) );
  AOI21_X1 U18697 ( .B1(n15627), .B2(n16415), .A(n15473), .ZN(n15474) );
  OAI21_X1 U18698 ( .B1(n9876), .B2(n16421), .A(n15474), .ZN(P2_U2985) );
  INV_X1 U18699 ( .A(n15475), .ZN(n15478) );
  INV_X1 U18700 ( .A(n12865), .ZN(n15477) );
  OAI21_X1 U18701 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15478), .A(
        n15477), .ZN(n15641) );
  INV_X1 U18702 ( .A(n15479), .ZN(n15630) );
  NAND2_X1 U18703 ( .A1(n15480), .A2(n15481), .ZN(n15629) );
  NAND3_X1 U18704 ( .A1(n15630), .A2(n16414), .A3(n15629), .ZN(n15487) );
  NAND2_X1 U18705 ( .A1(n16460), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15631) );
  OAI21_X1 U18706 ( .B1(n16429), .B2(n15482), .A(n15631), .ZN(n15484) );
  NOR2_X1 U18707 ( .A1(n15636), .A2(n16393), .ZN(n15483) );
  AOI211_X1 U18708 ( .C1(n16420), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15486) );
  OAI211_X1 U18709 ( .C1(n16424), .C2(n15641), .A(n15487), .B(n15486), .ZN(
        P2_U2987) );
  INV_X1 U18710 ( .A(n15488), .ZN(n15489) );
  AOI21_X1 U18711 ( .B1(n14253), .B2(n15490), .A(n15489), .ZN(n15492) );
  XNOR2_X1 U18712 ( .A(n15492), .B(n15491), .ZN(n15655) );
  NOR2_X1 U18713 ( .A1(n19124), .A2(n19941), .ZN(n15649) );
  AOI21_X1 U18714 ( .B1(n16411), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15649), .ZN(n15493) );
  OAI21_X1 U18715 ( .B1(n16419), .B2(n15494), .A(n15493), .ZN(n15497) );
  OAI21_X1 U18716 ( .B1(n15495), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15475), .ZN(n15642) );
  NOR2_X1 U18717 ( .A1(n15642), .A2(n16424), .ZN(n15496) );
  OAI21_X1 U18718 ( .B1(n16421), .B2(n15655), .A(n15498), .ZN(P2_U2988) );
  NOR2_X1 U18719 ( .A1(n10287), .A2(n15501), .ZN(n15502) );
  XNOR2_X1 U18720 ( .A(n15499), .B(n15502), .ZN(n15667) );
  INV_X1 U18721 ( .A(n15503), .ZN(n15512) );
  AOI21_X1 U18722 ( .B1(n15505), .B2(n15512), .A(n15504), .ZN(n15665) );
  OR2_X1 U18723 ( .A1(n19124), .A2(n19937), .ZN(n15658) );
  OAI21_X1 U18724 ( .B1(n16429), .B2(n10142), .A(n15658), .ZN(n15506) );
  AOI21_X1 U18725 ( .B1(n16420), .B2(n15507), .A(n15506), .ZN(n15508) );
  OAI21_X1 U18726 ( .B1(n15663), .B2(n16393), .A(n15508), .ZN(n15509) );
  AOI21_X1 U18727 ( .B1(n15665), .B2(n16415), .A(n15509), .ZN(n15510) );
  OAI21_X1 U18728 ( .B1(n15667), .B2(n16421), .A(n15510), .ZN(P2_U2990) );
  OAI21_X1 U18729 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15511), .A(
        n15512), .ZN(n15681) );
  NOR2_X1 U18730 ( .A1(n15513), .A2(n15514), .ZN(n15677) );
  NOR2_X1 U18731 ( .A1(n15677), .A2(n16421), .ZN(n15519) );
  OAI22_X1 U18732 ( .A1(n16429), .A2(n11285), .B1(n19935), .B2(n19124), .ZN(
        n15516) );
  AOI21_X1 U18733 ( .B1(n16420), .B2(n16310), .A(n15516), .ZN(n15517) );
  OAI21_X1 U18734 ( .B1(n16313), .B2(n16393), .A(n15517), .ZN(n15518) );
  AOI21_X1 U18735 ( .B1(n15519), .B2(n15515), .A(n15518), .ZN(n15520) );
  OAI21_X1 U18736 ( .B1(n15681), .B2(n16424), .A(n15520), .ZN(P2_U2991) );
  INV_X1 U18737 ( .A(n15597), .ZN(n15521) );
  AND2_X1 U18738 ( .A1(n15521), .A2(n15523), .ZN(n15522) );
  NAND2_X1 U18739 ( .A1(n15595), .A2(n15523), .ZN(n16365) );
  INV_X1 U18740 ( .A(n16363), .ZN(n15524) );
  NOR2_X1 U18741 ( .A1(n16365), .A2(n15524), .ZN(n15778) );
  INV_X1 U18742 ( .A(n15526), .ZN(n15768) );
  INV_X1 U18743 ( .A(n15548), .ZN(n15529) );
  AOI21_X1 U18744 ( .B1(n15546), .B2(n15530), .A(n15529), .ZN(n15535) );
  INV_X1 U18745 ( .A(n15531), .ZN(n15533) );
  NAND2_X1 U18746 ( .A1(n15533), .A2(n15532), .ZN(n15534) );
  XNOR2_X1 U18747 ( .A(n15535), .B(n15534), .ZN(n15709) );
  NAND2_X1 U18748 ( .A1(n16420), .A2(n15536), .ZN(n15537) );
  NAND2_X1 U18749 ( .A1(n16460), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15696) );
  OAI211_X1 U18750 ( .C1(n15538), .C2(n16429), .A(n15537), .B(n15696), .ZN(
        n15543) );
  INV_X1 U18751 ( .A(n15539), .ZN(n15541) );
  OAI21_X1 U18752 ( .B1(n15541), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15540), .ZN(n15704) );
  NOR2_X1 U18753 ( .A1(n15704), .A2(n16424), .ZN(n15542) );
  AOI211_X1 U18754 ( .C1(n16426), .C2(n15701), .A(n15543), .B(n15542), .ZN(
        n15544) );
  OAI21_X1 U18755 ( .B1(n15709), .B2(n16421), .A(n15544), .ZN(P2_U2993) );
  NAND2_X1 U18756 ( .A1(n15546), .A2(n15545), .ZN(n15550) );
  NAND2_X1 U18757 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  XNOR2_X1 U18758 ( .A(n15550), .B(n15549), .ZN(n15725) );
  NOR2_X1 U18759 ( .A1(n19124), .A2(n19930), .ZN(n15711) );
  AOI21_X1 U18760 ( .B1(n16411), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15711), .ZN(n15551) );
  OAI21_X1 U18761 ( .B1(n16419), .B2(n15552), .A(n15551), .ZN(n15556) );
  OAI21_X1 U18762 ( .B1(n15554), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15539), .ZN(n15722) );
  NOR2_X1 U18763 ( .A1(n15722), .A2(n16424), .ZN(n15555) );
  AOI211_X1 U18764 ( .C1(n16426), .C2(n15721), .A(n15556), .B(n15555), .ZN(
        n15557) );
  OAI21_X1 U18765 ( .B1(n15725), .B2(n16421), .A(n15557), .ZN(P2_U2994) );
  NAND2_X1 U18766 ( .A1(n15559), .A2(n15558), .ZN(n15562) );
  INV_X1 U18767 ( .A(n15569), .ZN(n15560) );
  AOI21_X1 U18768 ( .B1(n15571), .B2(n15568), .A(n15560), .ZN(n15561) );
  XOR2_X1 U18769 ( .A(n15562), .B(n15561), .Z(n15735) );
  AOI21_X1 U18770 ( .B1(n15730), .B2(n15563), .A(n15554), .ZN(n15733) );
  NAND2_X1 U18771 ( .A1(n16460), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15726) );
  OAI21_X1 U18772 ( .B1(n16429), .B2(n19017), .A(n15726), .ZN(n15564) );
  AOI21_X1 U18773 ( .B1(n19016), .B2(n16420), .A(n15564), .ZN(n15565) );
  OAI21_X1 U18774 ( .B1(n16393), .B2(n19023), .A(n15565), .ZN(n15566) );
  AOI21_X1 U18775 ( .B1(n15733), .B2(n16415), .A(n15566), .ZN(n15567) );
  OAI21_X1 U18776 ( .B1(n15735), .B2(n16421), .A(n15567), .ZN(P2_U2995) );
  NAND2_X1 U18777 ( .A1(n15569), .A2(n15568), .ZN(n15570) );
  XNOR2_X1 U18778 ( .A(n15571), .B(n15570), .ZN(n15749) );
  NOR2_X1 U18779 ( .A1(n16345), .A2(n15573), .ZN(n15752) );
  AOI21_X1 U18780 ( .B1(n15752), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15575) );
  INV_X1 U18781 ( .A(n15563), .ZN(n15574) );
  NOR2_X1 U18782 ( .A1(n15575), .A2(n15574), .ZN(n15747) );
  NOR2_X1 U18783 ( .A1(n19124), .A2(n15576), .ZN(n15739) );
  NOR2_X1 U18784 ( .A1(n16419), .A2(n15577), .ZN(n15578) );
  AOI211_X1 U18785 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n16411), .A(
        n15739), .B(n15578), .ZN(n15579) );
  OAI21_X1 U18786 ( .B1(n16393), .B2(n15744), .A(n15579), .ZN(n15580) );
  AOI21_X1 U18787 ( .B1(n15747), .B2(n16415), .A(n15580), .ZN(n15581) );
  OAI21_X1 U18788 ( .B1(n15749), .B2(n16421), .A(n15581), .ZN(P2_U2996) );
  NAND2_X1 U18789 ( .A1(n15583), .A2(n15582), .ZN(n15587) );
  INV_X1 U18790 ( .A(n15766), .ZN(n15585) );
  NAND2_X1 U18791 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  XOR2_X1 U18792 ( .A(n15587), .B(n15586), .Z(n15765) );
  INV_X1 U18793 ( .A(n15761), .ZN(n19030) );
  NOR2_X1 U18794 ( .A1(n19925), .A2(n19124), .ZN(n15590) );
  OAI22_X1 U18795 ( .A1(n16429), .A2(n15588), .B1(n16419), .B2(n19036), .ZN(
        n15589) );
  AOI211_X1 U18796 ( .C1(n16426), .C2(n19030), .A(n15590), .B(n15589), .ZN(
        n15594) );
  INV_X1 U18797 ( .A(n15752), .ZN(n15592) );
  OAI21_X1 U18798 ( .B1(n16345), .B2(n15573), .A(n15757), .ZN(n15591) );
  OAI211_X1 U18799 ( .C1(n15592), .C2(n15757), .A(n16415), .B(n15591), .ZN(
        n15593) );
  OAI211_X1 U18800 ( .C1(n15765), .C2(n16421), .A(n15594), .B(n15593), .ZN(
        P2_U2997) );
  INV_X1 U18801 ( .A(n15595), .ZN(n15596) );
  OAI22_X1 U18802 ( .A1(n15597), .A2(n16365), .B1(n15596), .B2(n9918), .ZN(
        n15808) );
  OAI22_X1 U18803 ( .A1(n16429), .A2(n15598), .B1(n11903), .B2(n19324), .ZN(
        n15603) );
  NAND2_X1 U18804 ( .A1(n16420), .A2(n19058), .ZN(n15601) );
  NAND2_X1 U18805 ( .A1(n16415), .A2(n15802), .ZN(n15600) );
  NAND2_X1 U18806 ( .A1(n15601), .A2(n15600), .ZN(n15602) );
  AOI211_X1 U18807 ( .C1(n19062), .C2(n16426), .A(n15603), .B(n15602), .ZN(
        n15604) );
  OAI21_X1 U18808 ( .B1(n15808), .B2(n16421), .A(n15604), .ZN(P2_U3001) );
  NAND2_X1 U18809 ( .A1(n15605), .A2(n15828), .ZN(n15606) );
  XOR2_X1 U18810 ( .A(n15606), .B(n9849), .Z(n15858) );
  INV_X1 U18811 ( .A(n15599), .ZN(n15607) );
  NAND2_X1 U18812 ( .A1(n15607), .A2(n21159), .ZN(n15846) );
  NAND3_X1 U18813 ( .A1(n15848), .A2(n16415), .A3(n15846), .ZN(n15614) );
  NOR2_X1 U18814 ( .A1(n19124), .A2(n15608), .ZN(n15612) );
  INV_X1 U18815 ( .A(n19090), .ZN(n15609) );
  OAI22_X1 U18816 ( .A1(n16429), .A2(n15610), .B1(n16419), .B2(n15609), .ZN(
        n15611) );
  AOI211_X1 U18817 ( .C1(n16426), .C2(n15849), .A(n15612), .B(n15611), .ZN(
        n15613) );
  OAI211_X1 U18818 ( .C1(n16421), .C2(n15858), .A(n15614), .B(n15613), .ZN(
        P2_U3005) );
  INV_X1 U18819 ( .A(n15632), .ZN(n15617) );
  NAND3_X1 U18820 ( .A1(n15617), .A2(n15616), .A3(n15615), .ZN(n15618) );
  NAND2_X1 U18821 ( .A1(n15619), .A2(n15618), .ZN(n15620) );
  AOI21_X1 U18822 ( .B1(n19310), .B2(n15621), .A(n15620), .ZN(n15624) );
  NAND2_X1 U18823 ( .A1(n15622), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15623) );
  OAI211_X1 U18824 ( .C1(n15625), .C2(n19312), .A(n15624), .B(n15623), .ZN(
        n15626) );
  AOI21_X1 U18825 ( .B1(n15627), .B2(n15847), .A(n15626), .ZN(n15628) );
  OAI21_X1 U18826 ( .B1(n9876), .B2(n19316), .A(n15628), .ZN(P2_U3017) );
  NAND3_X1 U18827 ( .A1(n15630), .A2(n16475), .A3(n15629), .ZN(n15640) );
  OAI21_X1 U18828 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15632), .A(
        n15631), .ZN(n15633) );
  AOI21_X1 U18829 ( .B1(n19310), .B2(n15634), .A(n15633), .ZN(n15635) );
  OAI21_X1 U18830 ( .B1(n15636), .B2(n19312), .A(n15635), .ZN(n15637) );
  AOI21_X1 U18831 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15638), .A(
        n15637), .ZN(n15639) );
  OAI211_X1 U18832 ( .C1(n15641), .C2(n19318), .A(n15640), .B(n15639), .ZN(
        P2_U3019) );
  INV_X1 U18833 ( .A(n15642), .ZN(n15653) );
  OAI211_X1 U18834 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n15644), .B(n15643), .ZN(
        n15645) );
  OAI21_X1 U18835 ( .B1(n15647), .B2(n15646), .A(n15645), .ZN(n15648) );
  AOI211_X1 U18836 ( .C1(n19310), .C2(n16305), .A(n15649), .B(n15648), .ZN(
        n15650) );
  OAI21_X1 U18837 ( .B1(n15651), .B2(n19312), .A(n15650), .ZN(n15652) );
  AOI21_X1 U18838 ( .B1(n15653), .B2(n15847), .A(n15652), .ZN(n15654) );
  OAI21_X1 U18839 ( .B1(n19316), .B2(n15655), .A(n15654), .ZN(P2_U3020) );
  OAI21_X1 U18840 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15657), .A(
        n15656), .ZN(n15662) );
  INV_X1 U18841 ( .A(n15658), .ZN(n15659) );
  AOI21_X1 U18842 ( .B1(n19310), .B2(n15660), .A(n15659), .ZN(n15661) );
  OAI211_X1 U18843 ( .C1(n15663), .C2(n19312), .A(n15662), .B(n15661), .ZN(
        n15664) );
  AOI21_X1 U18844 ( .B1(n15665), .B2(n15847), .A(n15664), .ZN(n15666) );
  OAI21_X1 U18845 ( .B1(n15667), .B2(n19316), .A(n15666), .ZN(P2_U3022) );
  AOI21_X1 U18846 ( .B1(n15669), .B2(n15689), .A(n15668), .ZN(n15675) );
  NOR2_X1 U18847 ( .A1(n15688), .A2(n15669), .ZN(n15674) );
  NOR2_X1 U18848 ( .A1(n19935), .A2(n19124), .ZN(n15670) );
  AOI21_X1 U18849 ( .B1(n19310), .B2(n15671), .A(n15670), .ZN(n15672) );
  OAI21_X1 U18850 ( .B1(n16313), .B2(n19312), .A(n15672), .ZN(n15673) );
  AOI211_X1 U18851 ( .C1(n15676), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        n15680) );
  INV_X1 U18852 ( .A(n15677), .ZN(n15678) );
  NAND3_X1 U18853 ( .A1(n15678), .A2(n16475), .A3(n15515), .ZN(n15679) );
  OAI211_X1 U18854 ( .C1(n15681), .C2(n19318), .A(n15680), .B(n15679), .ZN(
        P2_U3023) );
  INV_X1 U18855 ( .A(n15511), .ZN(n15682) );
  NAND2_X1 U18856 ( .A1(n15685), .A2(n15684), .ZN(n15686) );
  XNOR2_X1 U18857 ( .A(n15683), .B(n15686), .ZN(n16341) );
  NAND2_X1 U18858 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n16460), .ZN(n15687) );
  OAI221_X1 U18859 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15690), 
        .C1(n15689), .C2(n15688), .A(n15687), .ZN(n15694) );
  OAI22_X1 U18860 ( .A1(n15692), .A2(n19312), .B1(n16469), .B2(n15691), .ZN(
        n15693) );
  AOI211_X1 U18861 ( .C1(n16341), .C2(n16475), .A(n15694), .B(n15693), .ZN(
        n15695) );
  OAI21_X1 U18862 ( .B1(n16338), .B2(n19318), .A(n15695), .ZN(P2_U3024) );
  INV_X1 U18863 ( .A(n15696), .ZN(n15700) );
  NAND2_X1 U18864 ( .A1(n15796), .A2(n15855), .ZN(n16445) );
  INV_X1 U18865 ( .A(n16445), .ZN(n15697) );
  NAND2_X1 U18866 ( .A1(n16431), .A2(n15697), .ZN(n15786) );
  INV_X1 U18867 ( .A(n15698), .ZN(n15737) );
  NOR2_X1 U18868 ( .A1(n15786), .A2(n15737), .ZN(n15741) );
  NAND3_X1 U18869 ( .A1(n15741), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15710) );
  NOR3_X1 U18870 ( .A1(n15710), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15718), .ZN(n15699) );
  AOI211_X1 U18871 ( .C1(n15701), .C2(n16471), .A(n15700), .B(n15699), .ZN(
        n15702) );
  OAI21_X1 U18872 ( .B1(n16469), .B2(n15703), .A(n15702), .ZN(n15706) );
  NOR2_X1 U18873 ( .A1(n15704), .A2(n19318), .ZN(n15705) );
  AOI211_X1 U18874 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15707), .A(
        n15706), .B(n15705), .ZN(n15708) );
  OAI21_X1 U18875 ( .B1(n15709), .B2(n19316), .A(n15708), .ZN(P2_U3025) );
  INV_X1 U18876 ( .A(n15710), .ZN(n15712) );
  AOI21_X1 U18877 ( .B1(n15712), .B2(n15718), .A(n15711), .ZN(n15713) );
  OAI21_X1 U18878 ( .B1(n16469), .B2(n15714), .A(n15713), .ZN(n15720) );
  OR2_X1 U18879 ( .A1(n15864), .A2(n15715), .ZN(n15716) );
  NAND2_X1 U18880 ( .A1(n15851), .A2(n15716), .ZN(n15793) );
  AOI21_X1 U18881 ( .B1(n15717), .B2(n15736), .A(n15793), .ZN(n15731) );
  NAND3_X1 U18882 ( .A1(n15741), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15730), .ZN(n15727) );
  AOI21_X1 U18883 ( .B1(n15731), .B2(n15727), .A(n15718), .ZN(n15719) );
  AOI211_X1 U18884 ( .C1(n15721), .C2(n16471), .A(n15720), .B(n15719), .ZN(
        n15724) );
  OR2_X1 U18885 ( .A1(n15722), .A2(n19318), .ZN(n15723) );
  OAI211_X1 U18886 ( .C1(n15725), .C2(n19316), .A(n15724), .B(n15723), .ZN(
        P2_U3026) );
  OAI211_X1 U18887 ( .C1(n19312), .C2(n19023), .A(n15727), .B(n15726), .ZN(
        n15728) );
  AOI21_X1 U18888 ( .B1(n19310), .B2(n19021), .A(n15728), .ZN(n15729) );
  OAI21_X1 U18889 ( .B1(n15731), .B2(n15730), .A(n15729), .ZN(n15732) );
  AOI21_X1 U18890 ( .B1(n15733), .B2(n15847), .A(n15732), .ZN(n15734) );
  OAI21_X1 U18891 ( .B1(n15735), .B2(n19316), .A(n15734), .ZN(P2_U3027) );
  AOI21_X1 U18892 ( .B1(n15737), .B2(n15736), .A(n15793), .ZN(n15738) );
  NOR2_X1 U18893 ( .A1(n15738), .A2(n15740), .ZN(n15746) );
  NAND2_X1 U18894 ( .A1(n19310), .A2(n16333), .ZN(n15743) );
  AOI21_X1 U18895 ( .B1(n15741), .B2(n15740), .A(n15739), .ZN(n15742) );
  OAI211_X1 U18896 ( .C1(n15744), .C2(n19312), .A(n15743), .B(n15742), .ZN(
        n15745) );
  AOI211_X1 U18897 ( .C1(n15747), .C2(n15847), .A(n15746), .B(n15745), .ZN(
        n15748) );
  OAI21_X1 U18898 ( .B1(n15749), .B2(n19316), .A(n15748), .ZN(P2_U3028) );
  AND2_X1 U18899 ( .A1(n19318), .A2(n15750), .ZN(n15751) );
  OR2_X1 U18900 ( .A1(n15752), .A2(n15751), .ZN(n15756) );
  NOR2_X1 U18901 ( .A1(n15753), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15754) );
  NOR2_X1 U18902 ( .A1(n15793), .A2(n15754), .ZN(n15755) );
  OAI21_X1 U18903 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15864), .A(
        n15775), .ZN(n15763) );
  OAI22_X1 U18904 ( .A1(n16345), .A2(n19318), .B1(n15788), .B2(n15786), .ZN(
        n15772) );
  NAND3_X1 U18905 ( .A1(n15772), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15757), .ZN(n15760) );
  AOI22_X1 U18906 ( .A1(n19310), .A2(n15758), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n16460), .ZN(n15759) );
  OAI211_X1 U18907 ( .C1(n15761), .C2(n19312), .A(n15760), .B(n15759), .ZN(
        n15762) );
  AOI21_X1 U18908 ( .B1(n15763), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15762), .ZN(n15764) );
  OAI21_X1 U18909 ( .B1(n15765), .B2(n19316), .A(n15764), .ZN(P2_U3029) );
  AOI21_X1 U18910 ( .B1(n15768), .B2(n15767), .A(n15766), .ZN(n16349) );
  NAND2_X1 U18911 ( .A1(n16349), .A2(n16475), .ZN(n15774) );
  NOR2_X1 U18912 ( .A1(n16469), .A2(n19170), .ZN(n15771) );
  OAI22_X1 U18913 ( .A1(n19312), .A2(n16346), .B1(n15769), .B2(n19324), .ZN(
        n15770) );
  AOI211_X1 U18914 ( .C1(n15772), .C2(n15573), .A(n15771), .B(n15770), .ZN(
        n15773) );
  OAI211_X1 U18915 ( .C1(n15573), .C2(n15775), .A(n15774), .B(n15773), .ZN(
        P2_U3030) );
  NAND2_X1 U18916 ( .A1(n15572), .A2(n15788), .ZN(n15776) );
  NAND2_X1 U18917 ( .A1(n16345), .A2(n15776), .ZN(n16353) );
  INV_X1 U18918 ( .A(n16362), .ZN(n15777) );
  NOR2_X1 U18919 ( .A1(n15778), .A2(n15777), .ZN(n15782) );
  NAND2_X1 U18920 ( .A1(n15780), .A2(n15779), .ZN(n15781) );
  XNOR2_X1 U18921 ( .A(n15782), .B(n15781), .ZN(n16354) );
  OR2_X1 U18922 ( .A1(n16354), .A2(n19316), .ZN(n15795) );
  INV_X1 U18923 ( .A(n16356), .ZN(n19044) );
  INV_X1 U18924 ( .A(n15037), .ZN(n15783) );
  OAI21_X1 U18925 ( .B1(n15784), .B2(n13852), .A(n15783), .ZN(n19177) );
  INV_X1 U18926 ( .A(n19177), .ZN(n15785) );
  NAND2_X1 U18927 ( .A1(n19310), .A2(n15785), .ZN(n15791) );
  INV_X1 U18928 ( .A(n15786), .ZN(n15789) );
  NOR2_X1 U18929 ( .A1(n11956), .A2(n19124), .ZN(n15787) );
  AOI21_X1 U18930 ( .B1(n15789), .B2(n15788), .A(n15787), .ZN(n15790) );
  OAI211_X1 U18931 ( .C1(n19044), .C2(n19312), .A(n15791), .B(n15790), .ZN(
        n15792) );
  AOI21_X1 U18932 ( .B1(n15793), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15792), .ZN(n15794) );
  OAI211_X1 U18933 ( .C1(n16353), .C2(n19318), .A(n15795), .B(n15794), .ZN(
        P2_U3031) );
  NAND2_X1 U18934 ( .A1(n15851), .A2(n15796), .ZN(n15797) );
  NAND2_X1 U18935 ( .A1(n15798), .A2(n15797), .ZN(n16444) );
  INV_X1 U18936 ( .A(n16444), .ZN(n15806) );
  OAI21_X1 U18937 ( .B1(n15801), .B2(n15800), .A(n15799), .ZN(n19182) );
  AOI211_X1 U18938 ( .C1(n12734), .C2(n15803), .A(n16430), .B(n16445), .ZN(
        n15804) );
  AOI211_X1 U18939 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15806), .A(
        n15805), .B(n15804), .ZN(n15807) );
  OAI21_X1 U18940 ( .B1(n15808), .B2(n19316), .A(n15807), .ZN(P2_U3033) );
  NOR2_X1 U18941 ( .A1(n15848), .A2(n12718), .ZN(n16391) );
  INV_X1 U18942 ( .A(n16376), .ZN(n15809) );
  OAI21_X1 U18943 ( .B1(n16391), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15809), .ZN(n16384) );
  INV_X1 U18944 ( .A(n15810), .ZN(n15811) );
  NAND2_X1 U18945 ( .A1(n15812), .A2(n15811), .ZN(n15816) );
  NOR2_X1 U18946 ( .A1(n15814), .A2(n15813), .ZN(n15815) );
  XNOR2_X1 U18947 ( .A(n15816), .B(n15815), .ZN(n16383) );
  OAI21_X1 U18948 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15864), .A(
        n15851), .ZN(n15840) );
  NAND2_X1 U18949 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15855), .ZN(
        n15837) );
  AOI211_X1 U18950 ( .C1(n12718), .C2(n15818), .A(n15817), .B(n15837), .ZN(
        n15820) );
  NOR2_X1 U18951 ( .A1(n11862), .A2(n19124), .ZN(n15819) );
  AOI211_X1 U18952 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15840), .A(
        n15820), .B(n15819), .ZN(n15825) );
  OAI21_X1 U18953 ( .B1(n15822), .B2(n15821), .A(n13797), .ZN(n19187) );
  OAI22_X1 U18954 ( .A1(n19187), .A2(n16469), .B1(n19312), .B2(n19073), .ZN(
        n15823) );
  INV_X1 U18955 ( .A(n15823), .ZN(n15824) );
  OAI211_X1 U18956 ( .C1(n16383), .C2(n19316), .A(n15825), .B(n15824), .ZN(
        n15826) );
  INV_X1 U18957 ( .A(n15826), .ZN(n15827) );
  OAI21_X1 U18958 ( .B1(n16384), .B2(n19318), .A(n15827), .ZN(P2_U3035) );
  INV_X1 U18959 ( .A(n15828), .ZN(n15829) );
  NOR2_X1 U18960 ( .A1(n9884), .A2(n15829), .ZN(n15833) );
  NAND2_X1 U18961 ( .A1(n15831), .A2(n15830), .ZN(n15832) );
  XNOR2_X1 U18962 ( .A(n15833), .B(n15832), .ZN(n16394) );
  NOR2_X1 U18963 ( .A1(n15834), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16390) );
  OR3_X1 U18964 ( .A1(n16391), .A2(n16390), .A3(n19318), .ZN(n15845) );
  XNOR2_X1 U18965 ( .A(n15835), .B(n15836), .ZN(n19190) );
  INV_X1 U18966 ( .A(n19190), .ZN(n15843) );
  NOR2_X1 U18967 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15837), .ZN(
        n15839) );
  NOR2_X1 U18968 ( .A1(n11845), .A2(n19124), .ZN(n15838) );
  AOI211_X1 U18969 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n15840), .A(
        n15839), .B(n15838), .ZN(n15841) );
  OAI21_X1 U18970 ( .B1(n16392), .B2(n19312), .A(n15841), .ZN(n15842) );
  AOI21_X1 U18971 ( .B1(n15843), .B2(n19310), .A(n15842), .ZN(n15844) );
  OAI211_X1 U18972 ( .C1(n16394), .C2(n19316), .A(n15845), .B(n15844), .ZN(
        P2_U3036) );
  NAND3_X1 U18973 ( .A1(n15848), .A2(n15847), .A3(n15846), .ZN(n15857) );
  AOI22_X1 U18974 ( .A1(n16471), .A2(n15849), .B1(n16460), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n15850) );
  OAI21_X1 U18975 ( .B1(n15851), .B2(n21159), .A(n15850), .ZN(n15854) );
  OAI21_X1 U18976 ( .B1(n13829), .B2(n15852), .A(n15835), .ZN(n19192) );
  NOR2_X1 U18977 ( .A1(n19192), .A2(n16469), .ZN(n15853) );
  AOI211_X1 U18978 ( .C1(n15855), .C2(n21159), .A(n15854), .B(n15853), .ZN(
        n15856) );
  OAI211_X1 U18979 ( .C1(n15858), .C2(n19316), .A(n15857), .B(n15856), .ZN(
        P2_U3037) );
  NOR2_X1 U18980 ( .A1(n19318), .A2(n15859), .ZN(n15860) );
  AOI211_X1 U18981 ( .C1(n16471), .C2(n12565), .A(n15861), .B(n15860), .ZN(
        n15867) );
  AOI22_X1 U18982 ( .A1(n16475), .A2(n15862), .B1(n19310), .B2(n19141), .ZN(
        n15866) );
  MUX2_X1 U18983 ( .A(n15864), .B(n15863), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n15865) );
  NAND3_X1 U18984 ( .A1(n15867), .A2(n15866), .A3(n15865), .ZN(P2_U3046) );
  NAND2_X1 U18985 ( .A1(n13119), .A2(n16501), .ZN(n15871) );
  OAI21_X1 U18986 ( .B1(n11620), .B2(n11621), .A(n15868), .ZN(n15869) );
  INV_X1 U18987 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15874) );
  NAND2_X1 U18988 ( .A1(n16495), .A2(n15874), .ZN(n16497) );
  AND2_X1 U18989 ( .A1(n15869), .A2(n16497), .ZN(n15870) );
  NAND2_X1 U18990 ( .A1(n15871), .A2(n15870), .ZN(n16485) );
  NOR2_X1 U18991 ( .A1(n16540), .A2(n15872), .ZN(n19960) );
  AOI21_X1 U18992 ( .B1(n19117), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15873), .ZN(n19962) );
  AOI222_X1 U18993 ( .A1(n16485), .A2(n19969), .B1(n19960), .B2(n19962), .C1(
        n15906), .C2(n16548), .ZN(n15876) );
  NAND2_X1 U18994 ( .A1(n19966), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15875) );
  OAI21_X1 U18995 ( .B1(n15876), .B2(n19966), .A(n15875), .ZN(P2_U3600) );
  NAND2_X1 U18996 ( .A1(n15878), .A2(n15877), .ZN(n16488) );
  INV_X1 U18997 ( .A(n11637), .ZN(n15880) );
  NAND2_X1 U18998 ( .A1(n15880), .A2(n15879), .ZN(n16491) );
  NAND2_X1 U18999 ( .A1(n16488), .A2(n16491), .ZN(n15882) );
  INV_X1 U19000 ( .A(n15128), .ZN(n15885) );
  NAND3_X1 U19001 ( .A1(n16495), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15881) );
  NAND3_X1 U19002 ( .A1(n15882), .A2(n15885), .A3(n15881), .ZN(n15889) );
  NAND2_X1 U19003 ( .A1(n15884), .A2(n15883), .ZN(n15886) );
  NAND2_X1 U19004 ( .A1(n15886), .A2(n15885), .ZN(n16492) );
  NAND2_X1 U19005 ( .A1(n16495), .A2(n15879), .ZN(n15887) );
  NAND4_X1 U19006 ( .A1(n16492), .A2(n16497), .A3(n16491), .A4(n15887), .ZN(
        n15888) );
  MUX2_X1 U19007 ( .A(n15889), .B(n15888), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15890) );
  AOI21_X1 U19008 ( .B1(n12566), .B2(n16501), .A(n15890), .ZN(n16514) );
  OAI22_X1 U19009 ( .A1(n19972), .A2(n19965), .B1(n16514), .B2(n19963), .ZN(
        n15891) );
  MUX2_X1 U19010 ( .A(n15891), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n19966), .Z(P2_U3596) );
  INV_X1 U19011 ( .A(n16332), .ZN(n15892) );
  NOR2_X2 U19012 ( .A1(n15892), .A2(n19576), .ZN(n19845) );
  NOR3_X1 U19013 ( .A1(n19879), .A2(n19400), .A3(n19974), .ZN(n15894) );
  AND2_X1 U19014 ( .A1(n19971), .A2(n15893), .ZN(n19970) );
  NOR2_X1 U19015 ( .A1(n15894), .A2(n19970), .ZN(n15897) );
  NOR2_X1 U19016 ( .A1(n19980), .A2(n15895), .ZN(n19874) );
  NOR2_X1 U19017 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19438) );
  NAND2_X1 U19018 ( .A1(n19438), .A2(n19996), .ZN(n19372) );
  NOR2_X1 U19019 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19372), .ZN(
        n19356) );
  NOR2_X1 U19020 ( .A1(n19874), .A2(n19356), .ZN(n15899) );
  OAI21_X1 U19021 ( .B1(n12630), .B2(n19356), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15896) );
  OAI21_X1 U19022 ( .B1(n15897), .B2(n15899), .A(n15896), .ZN(n19360) );
  INV_X1 U19023 ( .A(n15897), .ZN(n15900) );
  AOI211_X1 U19024 ( .C1(n12630), .C2(n19825), .A(n19971), .B(n19356), .ZN(
        n15898) );
  INV_X1 U19025 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20294) );
  INV_X1 U19026 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18343) );
  OAI22_X2 U19027 ( .A1(n20294), .A2(n19359), .B1(n18343), .B2(n19358), .ZN(
        n19846) );
  NOR2_X2 U19028 ( .A1(n11458), .A2(n19342), .ZN(n19844) );
  AOI22_X1 U19029 ( .A1(n19846), .A2(n19400), .B1(n19844), .B2(n19356), .ZN(
        n15902) );
  AOI22_X1 U19030 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19352), .ZN(n19849) );
  INV_X1 U19031 ( .A(n19849), .ZN(n19796) );
  NAND2_X1 U19032 ( .A1(n19796), .A2(n19879), .ZN(n15901) );
  OAI211_X1 U19033 ( .C1(n19364), .C2(n15903), .A(n15902), .B(n15901), .ZN(
        n15904) );
  AOI21_X1 U19034 ( .B1(n19845), .B2(n19360), .A(n15904), .ZN(n15905) );
  INV_X1 U19035 ( .A(n15905), .ZN(P2_U3050) );
  NOR3_X1 U19036 ( .A1(n19682), .A2(n19717), .A3(n19974), .ZN(n15907) );
  NOR2_X1 U19037 ( .A1(n15907), .A2(n19970), .ZN(n15916) );
  INV_X1 U19038 ( .A(n15916), .ZN(n15909) );
  NOR2_X1 U19039 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19980), .ZN(
        n19690) );
  NAND2_X1 U19040 ( .A1(n19469), .A2(n19690), .ZN(n15915) );
  INV_X1 U19041 ( .A(n12615), .ZN(n15913) );
  NOR2_X1 U19042 ( .A1(n19996), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19404) );
  AND2_X1 U19043 ( .A1(n19404), .A2(n19690), .ZN(n19681) );
  AOI211_X1 U19044 ( .C1(n15913), .C2(n19825), .A(n19971), .B(n19681), .ZN(
        n15908) );
  AOI22_X1 U19045 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19352), .ZN(n19843) );
  INV_X1 U19046 ( .A(n19843), .ZN(n19700) );
  NAND2_X1 U19047 ( .A1(n15910), .A2(n19354), .ZN(n19484) );
  INV_X1 U19048 ( .A(n19681), .ZN(n15911) );
  OAI22_X1 U19049 ( .A1(n19703), .A2(n19714), .B1(n19484), .B2(n15911), .ZN(
        n15912) );
  AOI21_X1 U19050 ( .B1(n19682), .B2(n19700), .A(n15912), .ZN(n15919) );
  OAI21_X1 U19051 ( .B1(n15913), .B2(n19681), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15914) );
  NAND2_X1 U19052 ( .A1(n19683), .A2(n15917), .ZN(n15918) );
  OAI211_X1 U19053 ( .C1(n19687), .C2(n15920), .A(n15919), .B(n15918), .ZN(
        P2_U3129) );
  NAND2_X1 U19054 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16761), .ZN(n15922) );
  XNOR2_X1 U19055 ( .A(n17116), .B(n17109), .ZN(n17390) );
  NAND2_X1 U19056 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18554) );
  AOI221_X1 U19057 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18554), .C1(n15924), 
        .C2(n18554), .A(n15923), .ZN(n18328) );
  NOR2_X1 U19058 ( .A1(n15925), .A2(n18793), .ZN(n15926) );
  OAI21_X1 U19059 ( .B1(n15926), .B2(n18394), .A(n18329), .ZN(n18326) );
  AOI22_X1 U19060 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18328), .B1(
        n18326), .B2(n18798), .ZN(P3_U2865) );
  NAND2_X1 U19061 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18973) );
  NOR2_X1 U19062 ( .A1(n18763), .A2(n18836), .ZN(n15937) );
  INV_X1 U19063 ( .A(n15929), .ZN(n15930) );
  NAND2_X1 U19064 ( .A1(n18972), .A2(n17581), .ZN(n18811) );
  NOR2_X2 U19065 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18838), .ZN(n18957) );
  INV_X1 U19066 ( .A(n18981), .ZN(n18980) );
  NAND2_X2 U19067 ( .A1(n18980), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18908) );
  OAI211_X1 U19068 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18845), .B(n18908), .ZN(n18970) );
  OAI211_X1 U19069 ( .C1(n15934), .C2(n15933), .A(n15932), .B(n15931), .ZN(
        n15947) );
  AOI21_X1 U19070 ( .B1(n15937), .B2(n17526), .A(n15947), .ZN(n15939) );
  OAI211_X1 U19071 ( .C1(n18958), .C2(n15940), .A(n15939), .B(n16023), .ZN(
        n18785) );
  NOR2_X1 U19072 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18920), .ZN(n18334) );
  INV_X1 U19073 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21210) );
  NOR2_X1 U19074 ( .A1(n21210), .A2(n18918), .ZN(n15941) );
  AOI21_X1 U19075 ( .B1(n15942), .B2(n18767), .A(n18760), .ZN(n18764) );
  NAND3_X1 U19076 ( .A1(n18945), .A2(n18943), .A3(n18764), .ZN(n15943) );
  OAI21_X1 U19077 ( .B1(n18945), .B2(n18767), .A(n15943), .ZN(P3_U3284) );
  INV_X1 U19078 ( .A(n15944), .ZN(n15949) );
  OAI21_X1 U19079 ( .B1(n15945), .B2(n18338), .A(n18970), .ZN(n15946) );
  OAI21_X1 U19080 ( .B1(n15953), .B2(n15946), .A(n18973), .ZN(n16694) );
  NOR3_X1 U19081 ( .A1(n15949), .A2(n18763), .A3(n16694), .ZN(n15948) );
  AOI211_X1 U19082 ( .C1(n15950), .C2(n15949), .A(n15948), .B(n15947), .ZN(
        n15952) );
  AOI221_X4 U19083 ( .B1(n17377), .B2(n15952), .C1(n15951), .C2(n15952), .A(
        n18817), .ZN(n18315) );
  INV_X1 U19084 ( .A(n18191), .ZN(n17816) );
  INV_X1 U19085 ( .A(n15959), .ZN(n17493) );
  NAND2_X1 U19086 ( .A1(n18035), .A2(n15953), .ZN(n18963) );
  AOI22_X1 U19087 ( .A1(n18959), .A2(n17816), .B1(n17810), .B2(n18190), .ZN(
        n18178) );
  INV_X1 U19088 ( .A(n18197), .ZN(n18786) );
  NAND2_X1 U19089 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18223) );
  NOR2_X1 U19090 ( .A1(n18233), .A2(n18223), .ZN(n18102) );
  INV_X1 U19091 ( .A(n18102), .ZN(n15954) );
  INV_X1 U19092 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18260) );
  NOR3_X1 U19093 ( .A1(n18260), .A2(n18280), .A3(n18261), .ZN(n18250) );
  NOR2_X1 U19094 ( .A1(n18292), .A2(n18927), .ZN(n18268) );
  NAND2_X1 U19095 ( .A1(n18250), .A2(n18268), .ZN(n18225) );
  NOR2_X1 U19096 ( .A1(n15954), .A2(n18225), .ZN(n18149) );
  INV_X1 U19097 ( .A(n18149), .ZN(n18162) );
  NOR2_X1 U19098 ( .A1(n16560), .A2(n18162), .ZN(n18103) );
  NAND2_X1 U19099 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18103), .ZN(
        n18120) );
  INV_X1 U19100 ( .A(n18120), .ZN(n15955) );
  OAI21_X1 U19101 ( .B1(n18944), .B2(n18927), .A(n18292), .ZN(n18296) );
  AND2_X1 U19102 ( .A1(n18296), .A2(n18250), .ZN(n18227) );
  NAND2_X1 U19103 ( .A1(n18227), .A2(n18102), .ZN(n18121) );
  NOR2_X1 U19104 ( .A1(n16560), .A2(n18121), .ZN(n18040) );
  AOI222_X1 U19105 ( .A1(n18786), .A2(n15955), .B1(n18040), .B2(n18784), .C1(
        n18768), .C2(n18103), .ZN(n18026) );
  OAI21_X1 U19106 ( .B1(n18178), .B2(n16560), .A(n18026), .ZN(n18053) );
  NAND2_X1 U19107 ( .A1(n18315), .A2(n18053), .ZN(n18095) );
  NAND2_X1 U19108 ( .A1(n16569), .A2(n18008), .ZN(n15964) );
  NOR2_X1 U19109 ( .A1(n18035), .A2(n18302), .ZN(n18308) );
  NOR2_X2 U19110 ( .A1(n9816), .A2(n18315), .ZN(n18310) );
  INV_X1 U19111 ( .A(n18784), .ZN(n18770) );
  AOI21_X1 U19112 ( .B1(n16589), .B2(n18040), .A(n18770), .ZN(n18006) );
  INV_X1 U19113 ( .A(n18288), .ZN(n18269) );
  AOI21_X1 U19114 ( .B1(n16589), .B2(n18103), .A(n18269), .ZN(n15957) );
  AOI21_X1 U19115 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n18197), .ZN(n15956) );
  NOR4_X1 U19116 ( .A1(n18310), .A2(n18006), .A3(n15957), .A4(n15956), .ZN(
        n16603) );
  NOR2_X1 U19117 ( .A1(n9816), .A2(n16603), .ZN(n16009) );
  NOR2_X1 U19118 ( .A1(n18302), .A2(n18167), .ZN(n16590) );
  INV_X1 U19119 ( .A(n16590), .ZN(n18240) );
  INV_X1 U19120 ( .A(n18307), .ZN(n18322) );
  OAI22_X1 U19121 ( .A1(n18240), .A2(n16570), .B1(n18322), .B2(n16568), .ZN(
        n16010) );
  AOI211_X1 U19122 ( .C1(n18308), .C2(n15958), .A(n16009), .B(n16010), .ZN(
        n15963) );
  AOI21_X1 U19123 ( .B1(n16571), .B2(n15960), .A(n15961), .ZN(n16574) );
  AOI22_X1 U19124 ( .A1(n9816), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18236), 
        .B2(n16574), .ZN(n15962) );
  OAI221_X1 U19125 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15964), 
        .C1(n16571), .C2(n15963), .A(n15962), .ZN(P3_U2833) );
  INV_X1 U19126 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20049) );
  NAND2_X1 U19127 ( .A1(n21227), .A2(n20049), .ZN(n15985) );
  NOR2_X1 U19128 ( .A1(n15970), .A2(n10312), .ZN(n15979) );
  INV_X1 U19129 ( .A(n15975), .ZN(n15977) );
  INV_X1 U19130 ( .A(n15965), .ZN(n15966) );
  AOI21_X1 U19131 ( .B1(n15966), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20952), .ZN(n15967) );
  AND2_X1 U19132 ( .A1(n15968), .A2(n15967), .ZN(n15971) );
  OAI22_X1 U19133 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15971), .B1(
        n15970), .B2(n15969), .ZN(n15973) );
  NAND2_X1 U19134 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15971), .ZN(
        n15972) );
  OAI211_X1 U19135 ( .C1(n15975), .C2(n15974), .A(n15973), .B(n15972), .ZN(
        n15976) );
  OAI21_X1 U19136 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15977), .A(
        n15976), .ZN(n15978) );
  AOI222_X1 U19137 ( .A1(n20945), .A2(n15979), .B1(n20945), .B2(n15978), .C1(
        n15979), .C2(n15978), .ZN(n15981) );
  OAI21_X1 U19138 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n15981), .A(
        n15980), .ZN(n15982) );
  OR2_X1 U19139 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  AOI21_X1 U19140 ( .B1(n15986), .B2(n15985), .A(n15984), .ZN(n15987) );
  NOR2_X1 U19141 ( .A1(n15990), .A2(n16289), .ZN(n20950) );
  INV_X1 U19142 ( .A(n16003), .ZN(n15996) );
  NOR3_X1 U19143 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20964), .A3(n20972), 
        .ZN(n15994) );
  NAND3_X1 U19144 ( .A1(n12020), .A2(n20287), .A3(n15991), .ZN(n15993) );
  NAND2_X1 U19145 ( .A1(n20965), .A2(n20972), .ZN(n15992) );
  OAI22_X1 U19146 ( .A1(n15995), .A2(n15994), .B1(n15993), .B2(n15992), .ZN(
        n16287) );
  AOI221_X1 U19147 ( .B1(n20968), .B2(n20857), .C1(n15996), .C2(n20857), .A(
        n16287), .ZN(n15998) );
  NOR2_X1 U19148 ( .A1(n15998), .A2(n20968), .ZN(n16290) );
  OAI211_X1 U19149 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20972), .A(n16290), 
        .B(n15997), .ZN(n16288) );
  AOI21_X1 U19150 ( .B1(n16000), .B2(n15999), .A(n15998), .ZN(n16001) );
  OAI22_X1 U19151 ( .A1(n20950), .A2(n16288), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16001), .ZN(n16002) );
  OAI21_X1 U19152 ( .B1(n16003), .B2(n20042), .A(n16002), .ZN(P1_U3161) );
  INV_X1 U19153 ( .A(n16004), .ZN(n16006) );
  INV_X1 U19154 ( .A(n16007), .ZN(n16008) );
  XNOR2_X1 U19155 ( .A(n16008), .B(n16011), .ZN(n16566) );
  NOR2_X1 U19156 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16583), .ZN(
        n16562) );
  AOI21_X1 U19157 ( .B1(n18308), .B2(n16583), .A(n16009), .ZN(n16585) );
  INV_X1 U19158 ( .A(n16010), .ZN(n16012) );
  AOI21_X1 U19159 ( .B1(n16585), .B2(n16012), .A(n16011), .ZN(n16013) );
  AOI21_X1 U19160 ( .B1(n18008), .B2(n16562), .A(n16013), .ZN(n16014) );
  NAND2_X1 U19161 ( .A1(n9816), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16556) );
  OAI211_X1 U19162 ( .C1(n16566), .C2(n18221), .A(n16014), .B(n16556), .ZN(
        P3_U2832) );
  INV_X1 U19163 ( .A(HOLD), .ZN(n20866) );
  NOR2_X1 U19164 ( .A1(n20874), .A2(n20866), .ZN(n20861) );
  AOI22_X1 U19165 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n16017) );
  NAND2_X1 U19166 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n16015), .ZN(n20864) );
  OAI211_X1 U19167 ( .C1(n20861), .C2(n16017), .A(n16016), .B(n20864), .ZN(
        P1_U3195) );
  AND2_X1 U19168 ( .A1(n20175), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19169 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16019) );
  NOR2_X1 U19170 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16018) );
  NOR3_X1 U19171 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19237), .A3(n20026), 
        .ZN(n19886) );
  NOR4_X1 U19172 ( .A1(n16019), .A2(n16018), .A3(n19886), .A4(n16538), .ZN(
        P2_U3178) );
  INV_X1 U19173 ( .A(n16538), .ZN(n16555) );
  OAI221_X1 U19174 ( .B1(n16020), .B2(n16555), .C1(n16539), .C2(n16555), .A(
        n19576), .ZN(n20007) );
  NOR2_X1 U19175 ( .A1(n16512), .A2(n20007), .ZN(P2_U3047) );
  NAND3_X1 U19176 ( .A1(n18335), .A2(n18972), .A3(n16021), .ZN(n16022) );
  NAND2_X1 U19177 ( .A1(n17519), .A2(n17517), .ZN(n17491) );
  INV_X1 U19178 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17579) );
  INV_X1 U19179 ( .A(n18787), .ZN(n16024) );
  AOI22_X1 U19180 ( .A1(n17522), .A2(BUF2_REG_0__SCAN_IN), .B1(n17521), .B2(
        n17992), .ZN(n16025) );
  OAI221_X1 U19181 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17491), .C1(n17579), 
        .C2(n17517), .A(n16025), .ZN(P3_U2735) );
  NOR3_X1 U19182 ( .A1(n20107), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n16026), 
        .ZN(n16028) );
  AND2_X1 U19183 ( .A1(n20125), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n16027) );
  AOI211_X1 U19184 ( .C1(n16040), .C2(P1_REIP_REG_24__SCAN_IN), .A(n16028), 
        .B(n16027), .ZN(n16030) );
  NAND2_X1 U19185 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16029) );
  OAI211_X1 U19186 ( .C1(n16031), .C2(n16104), .A(n16030), .B(n16029), .ZN(
        n16032) );
  AOI21_X1 U19187 ( .B1(n16033), .B2(n20136), .A(n16032), .ZN(n16034) );
  OAI21_X1 U19188 ( .B1(n20140), .B2(n16035), .A(n16034), .ZN(P1_U2816) );
  INV_X1 U19189 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21166) );
  NAND3_X1 U19190 ( .A1(n16067), .A2(n20127), .A3(n16036), .ZN(n16047) );
  OAI21_X1 U19191 ( .B1(n21166), .B2(n16047), .A(n14664), .ZN(n16039) );
  INV_X1 U19192 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16037) );
  INV_X1 U19193 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n16138) );
  OAI22_X1 U19194 ( .A1(n20100), .A2(n16037), .B1(n16138), .B2(n20064), .ZN(
        n16038) );
  AOI21_X1 U19195 ( .B1(n16040), .B2(n16039), .A(n16038), .ZN(n16043) );
  OAI22_X1 U19196 ( .A1(n16135), .A2(n16104), .B1(n20140), .B2(n16134), .ZN(
        n16041) );
  INV_X1 U19197 ( .A(n16041), .ZN(n16042) );
  OAI211_X1 U19198 ( .C1(n16044), .C2(n20114), .A(n16043), .B(n16042), .ZN(
        P1_U2817) );
  NAND2_X1 U19199 ( .A1(n16067), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16056) );
  AOI21_X1 U19200 ( .B1(n20127), .B2(n16056), .A(n16045), .ZN(n16075) );
  NAND2_X1 U19201 ( .A1(n20127), .A2(n14680), .ZN(n16057) );
  AOI21_X1 U19202 ( .B1(n16075), .B2(n16057), .A(n21166), .ZN(n16049) );
  OAI22_X1 U19203 ( .A1(n16047), .A2(P1_REIP_REG_22__SCAN_IN), .B1(n16046), 
        .B2(n20064), .ZN(n16048) );
  AOI211_X1 U19204 ( .C1(n20126), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16049), .B(n16048), .ZN(n16053) );
  AOI22_X1 U19205 ( .A1(n16051), .A2(n20089), .B1(n16050), .B2(n20136), .ZN(
        n16052) );
  OAI211_X1 U19206 ( .C1(n20140), .C2(n16054), .A(n16053), .B(n16052), .ZN(
        P1_U2818) );
  NOR2_X1 U19207 ( .A1(n16075), .A2(n14680), .ZN(n16059) );
  AOI22_X1 U19208 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20125), .B2(P1_EBX_REG_21__SCAN_IN), .ZN(n16055) );
  OAI21_X1 U19209 ( .B1(n16057), .B2(n16056), .A(n16055), .ZN(n16058) );
  NOR2_X1 U19210 ( .A1(n16059), .A2(n16058), .ZN(n16065) );
  INV_X1 U19211 ( .A(n16060), .ZN(n16063) );
  INV_X1 U19212 ( .A(n16061), .ZN(n16062) );
  AOI22_X1 U19213 ( .A1(n16063), .A2(n20089), .B1(n16062), .B2(n20097), .ZN(
        n16064) );
  OAI211_X1 U19214 ( .C1(n16066), .C2(n20114), .A(n16065), .B(n16064), .ZN(
        P1_U2819) );
  AOI21_X1 U19215 ( .B1(n16067), .B2(n20127), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n16074) );
  AOI22_X1 U19216 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n20125), .ZN(n16073) );
  OAI22_X1 U19217 ( .A1(n16069), .A2(n16104), .B1(n20140), .B2(n16068), .ZN(
        n16070) );
  AOI21_X1 U19218 ( .B1(n16071), .B2(n20136), .A(n16070), .ZN(n16072) );
  OAI211_X1 U19219 ( .C1(n16075), .C2(n16074), .A(n16073), .B(n16072), .ZN(
        P1_U2820) );
  INV_X1 U19220 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16080) );
  NOR3_X1 U19221 ( .A1(n20107), .A2(n16097), .A3(n16076), .ZN(n16090) );
  XNOR2_X1 U19222 ( .A(P1_REIP_REG_19__SCAN_IN), .B(n20900), .ZN(n16077) );
  AOI22_X1 U19223 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n16087), .B1(n16090), 
        .B2(n16077), .ZN(n16079) );
  AOI21_X1 U19224 ( .B1(n20125), .B2(P1_EBX_REG_19__SCAN_IN), .A(n20110), .ZN(
        n16078) );
  OAI211_X1 U19225 ( .C1(n16080), .C2(n20100), .A(n16079), .B(n16078), .ZN(
        n16081) );
  INV_X1 U19226 ( .A(n16081), .ZN(n16086) );
  AOI21_X1 U19227 ( .B1(n16084), .B2(n16083), .A(n16082), .ZN(n16203) );
  AOI22_X1 U19228 ( .A1(n16144), .A2(n20089), .B1(n20097), .B2(n16203), .ZN(
        n16085) );
  OAI211_X1 U19229 ( .C1(n16147), .C2(n20114), .A(n16086), .B(n16085), .ZN(
        P1_U2821) );
  AOI22_X1 U19230 ( .A1(n16087), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(n20125), .ZN(n16088) );
  OAI211_X1 U19231 ( .C1(n20100), .C2(n14692), .A(n16088), .B(n20098), .ZN(
        n16089) );
  AOI21_X1 U19232 ( .B1(n16090), .B2(n20900), .A(n16089), .ZN(n16094) );
  AOI22_X1 U19233 ( .A1(n16092), .A2(n20089), .B1(n20136), .B2(n16091), .ZN(
        n16093) );
  OAI211_X1 U19234 ( .C1(n20140), .C2(n16095), .A(n16094), .B(n16093), .ZN(
        P1_U2822) );
  INV_X1 U19235 ( .A(n16096), .ZN(n16099) );
  NOR3_X1 U19236 ( .A1(n20107), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n16097), 
        .ZN(n16111) );
  NOR2_X1 U19237 ( .A1(n16110), .A2(n16111), .ZN(n16098) );
  MUX2_X1 U19238 ( .A(n16099), .B(n16098), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n16100) );
  OAI21_X1 U19239 ( .B1(n16101), .B2(n20064), .A(n16100), .ZN(n16102) );
  AOI211_X1 U19240 ( .C1(n20126), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20110), .B(n16102), .ZN(n16108) );
  OAI22_X1 U19241 ( .A1(n16105), .A2(n16104), .B1(n16103), .B2(n20114), .ZN(
        n16106) );
  INV_X1 U19242 ( .A(n16106), .ZN(n16107) );
  OAI211_X1 U19243 ( .C1(n20140), .C2(n16109), .A(n16108), .B(n16107), .ZN(
        P1_U2824) );
  NAND2_X1 U19244 ( .A1(n16110), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16113) );
  AOI211_X1 U19245 ( .C1(n20125), .C2(P1_EBX_REG_15__SCAN_IN), .A(n20110), .B(
        n16111), .ZN(n16112) );
  OAI211_X1 U19246 ( .C1(n16114), .C2(n20100), .A(n16113), .B(n16112), .ZN(
        n16115) );
  AOI21_X1 U19247 ( .B1(n16164), .B2(n20089), .A(n16115), .ZN(n16118) );
  INV_X1 U19248 ( .A(n16215), .ZN(n16116) );
  AOI22_X1 U19249 ( .A1(n16163), .A2(n20136), .B1(n20097), .B2(n16116), .ZN(
        n16117) );
  NAND2_X1 U19250 ( .A1(n16118), .A2(n16117), .ZN(P1_U2825) );
  AOI21_X1 U19251 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16128), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16126) );
  INV_X1 U19252 ( .A(n16119), .ZN(n16123) );
  AOI21_X1 U19253 ( .B1(n20125), .B2(P1_EBX_REG_12__SCAN_IN), .A(n20110), .ZN(
        n16120) );
  OAI21_X1 U19254 ( .B1(n20100), .B2(n16121), .A(n16120), .ZN(n16122) );
  AOI21_X1 U19255 ( .B1(n16123), .B2(n20097), .A(n16122), .ZN(n16125) );
  AOI22_X1 U19256 ( .A1(n16168), .A2(n20136), .B1(n20089), .B2(n16167), .ZN(
        n16124) );
  OAI211_X1 U19257 ( .C1(n16127), .C2(n16126), .A(n16125), .B(n16124), .ZN(
        P1_U2828) );
  INV_X1 U19258 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U19259 ( .A1(n20097), .A2(n16227), .B1(n16128), .B2(n20890), .ZN(
        n16133) );
  INV_X1 U19260 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21272) );
  AOI22_X1 U19261 ( .A1(n16129), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20125), 
        .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n16130) );
  OAI211_X1 U19262 ( .C1(n20100), .C2(n21272), .A(n16130), .B(n20098), .ZN(
        n16131) );
  AOI21_X1 U19263 ( .B1(n20089), .B2(n16178), .A(n16131), .ZN(n16132) );
  OAI211_X1 U19264 ( .C1(n16181), .C2(n20114), .A(n16133), .B(n16132), .ZN(
        P1_U2829) );
  OAI22_X1 U19265 ( .A1(n16135), .A2(n14564), .B1(n16134), .B2(n20146), .ZN(
        n16136) );
  INV_X1 U19266 ( .A(n16136), .ZN(n16137) );
  OAI21_X1 U19267 ( .B1(n20157), .B2(n16138), .A(n16137), .ZN(P1_U2849) );
  AOI22_X1 U19268 ( .A1(n16144), .A2(n20153), .B1(n20152), .B2(n16203), .ZN(
        n16139) );
  OAI21_X1 U19269 ( .B1(n20157), .B2(n21209), .A(n16139), .ZN(P1_U2853) );
  AOI22_X1 U19270 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16146) );
  NAND2_X1 U19271 ( .A1(n16141), .A2(n16140), .ZN(n16143) );
  XOR2_X1 U19272 ( .A(n16143), .B(n16142), .Z(n16204) );
  AOI22_X1 U19273 ( .A1(n16144), .A2(n16192), .B1(n20225), .B2(n16204), .ZN(
        n16145) );
  OAI211_X1 U19274 ( .C1(n20230), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P1_U2980) );
  NAND2_X1 U19275 ( .A1(n16148), .A2(n16150), .ZN(n16151) );
  MUX2_X1 U19276 ( .A(n16151), .B(n16150), .S(n16149), .Z(n16153) );
  XNOR2_X1 U19277 ( .A(n16153), .B(n16152), .ZN(n16213) );
  AOI22_X1 U19278 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16158) );
  INV_X1 U19279 ( .A(n16154), .ZN(n16156) );
  AOI22_X1 U19280 ( .A1(n16156), .A2(n16192), .B1(n16169), .B2(n16155), .ZN(
        n16157) );
  OAI211_X1 U19281 ( .C1(n20048), .C2(n16213), .A(n16158), .B(n16157), .ZN(
        P1_U2982) );
  NAND2_X1 U19282 ( .A1(n16160), .A2(n16159), .ZN(n16162) );
  XOR2_X1 U19283 ( .A(n16162), .B(n16161), .Z(n16220) );
  AOI22_X1 U19284 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16166) );
  AOI22_X1 U19285 ( .A1(n16164), .A2(n16192), .B1(n16163), .B2(n16169), .ZN(
        n16165) );
  OAI211_X1 U19286 ( .C1(n16220), .C2(n20048), .A(n16166), .B(n16165), .ZN(
        P1_U2984) );
  AOI22_X1 U19287 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16171) );
  AOI22_X1 U19288 ( .A1(n16169), .A2(n16168), .B1(n16192), .B2(n16167), .ZN(
        n16170) );
  OAI211_X1 U19289 ( .C1(n16172), .C2(n20048), .A(n16171), .B(n16170), .ZN(
        P1_U2987) );
  AOI22_X1 U19290 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16180) );
  NAND3_X1 U19291 ( .A1(n16174), .A2(n16173), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16176) );
  NAND2_X1 U19292 ( .A1(n16176), .A2(n16175), .ZN(n16177) );
  XNOR2_X1 U19293 ( .A(n16177), .B(n11251), .ZN(n16229) );
  AOI22_X1 U19294 ( .A1(n20225), .A2(n16229), .B1(n16192), .B2(n16178), .ZN(
        n16179) );
  OAI211_X1 U19295 ( .C1(n20230), .C2(n16181), .A(n16180), .B(n16179), .ZN(
        P1_U2988) );
  AOI22_X1 U19296 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16187) );
  NAND2_X1 U19297 ( .A1(n16183), .A2(n16182), .ZN(n16184) );
  XNOR2_X1 U19298 ( .A(n16185), .B(n16184), .ZN(n16263) );
  AOI22_X1 U19299 ( .A1(n16263), .A2(n20225), .B1(n16192), .B2(n20148), .ZN(
        n16186) );
  OAI211_X1 U19300 ( .C1(n20230), .C2(n20083), .A(n16187), .B(n16186), .ZN(
        P1_U2992) );
  AOI22_X1 U19301 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16194) );
  XNOR2_X1 U19302 ( .A(n16189), .B(n16188), .ZN(n16190) );
  XNOR2_X1 U19303 ( .A(n16191), .B(n16190), .ZN(n16269) );
  AOI22_X1 U19304 ( .A1(n16269), .A2(n20225), .B1(n16192), .B2(n20090), .ZN(
        n16193) );
  OAI211_X1 U19305 ( .C1(n20230), .C2(n20093), .A(n16194), .B(n16193), .ZN(
        P1_U2993) );
  AOI22_X1 U19306 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16200) );
  OAI21_X1 U19307 ( .B1(n16197), .B2(n16196), .A(n16195), .ZN(n16198) );
  INV_X1 U19308 ( .A(n16198), .ZN(n16278) );
  AOI22_X1 U19309 ( .A1(n16278), .A2(n20225), .B1(n16192), .B2(n20154), .ZN(
        n16199) );
  OAI211_X1 U19310 ( .C1(n20230), .C2(n20105), .A(n16200), .B(n16199), .ZN(
        P1_U2994) );
  OAI22_X1 U19311 ( .A1(n11258), .A2(n16201), .B1(n20252), .B2(n20898), .ZN(
        n16202) );
  INV_X1 U19312 ( .A(n16202), .ZN(n16206) );
  AOI22_X1 U19313 ( .A1(n16204), .A2(n20237), .B1(n20234), .B2(n16203), .ZN(
        n16205) );
  OAI211_X1 U19314 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16207), .A(
        n16206), .B(n16205), .ZN(P1_U3012) );
  AOI22_X1 U19315 ( .A1(n16208), .A2(n20234), .B1(n20221), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16212) );
  OAI21_X1 U19316 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16210), .A(
        n16209), .ZN(n16211) );
  OAI211_X1 U19317 ( .C1(n16213), .C2(n20250), .A(n16212), .B(n16211), .ZN(
        P1_U3014) );
  AOI22_X1 U19318 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16214), .B1(
        n20221), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16219) );
  OAI22_X1 U19319 ( .A1(n16216), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16215), .B2(n20254), .ZN(n16217) );
  INV_X1 U19320 ( .A(n16217), .ZN(n16218) );
  OAI211_X1 U19321 ( .C1(n16220), .C2(n20250), .A(n16219), .B(n16218), .ZN(
        P1_U3016) );
  AOI22_X1 U19322 ( .A1(n16222), .A2(n20237), .B1(n20234), .B2(n16221), .ZN(
        n16226) );
  OAI21_X1 U19323 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16224), .A(
        n16223), .ZN(n16225) );
  OAI211_X1 U19324 ( .C1(n20893), .C2(n20252), .A(n16226), .B(n16225), .ZN(
        P1_U3018) );
  AOI22_X1 U19325 ( .A1(n16227), .A2(n20234), .B1(n20221), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16231) );
  AOI22_X1 U19326 ( .A1(n16229), .A2(n20237), .B1(n16228), .B2(n11251), .ZN(
        n16230) );
  OAI211_X1 U19327 ( .C1(n16232), .C2(n11251), .A(n16231), .B(n16230), .ZN(
        P1_U3020) );
  INV_X1 U19328 ( .A(n16233), .ZN(n16234) );
  AOI21_X1 U19329 ( .B1(n16236), .B2(n16235), .A(n16234), .ZN(n16239) );
  NAND3_X1 U19330 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16237) );
  AOI221_X1 U19331 ( .B1(n16239), .B2(n16238), .C1(n16237), .C2(n16238), .A(
        n20246), .ZN(n16257) );
  NAND2_X1 U19332 ( .A1(n16240), .A2(n16262), .ZN(n16252) );
  AOI221_X1 U19333 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14727), .C2(n16256), .A(
        n16252), .ZN(n16243) );
  OAI22_X1 U19334 ( .A1(n16241), .A2(n20254), .B1(n20887), .B2(n20252), .ZN(
        n16242) );
  AOI211_X1 U19335 ( .C1(n16244), .C2(n20237), .A(n16243), .B(n16242), .ZN(
        n16245) );
  OAI21_X1 U19336 ( .B1(n16257), .B2(n14727), .A(n16245), .ZN(P1_U3021) );
  INV_X1 U19337 ( .A(n16246), .ZN(n16254) );
  OR2_X1 U19338 ( .A1(n16248), .A2(n16247), .ZN(n16249) );
  AND2_X1 U19339 ( .A1(n16250), .A2(n16249), .ZN(n20141) );
  AOI22_X1 U19340 ( .A1(n20141), .A2(n20234), .B1(n20221), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16251) );
  OAI21_X1 U19341 ( .B1(n16252), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16251), .ZN(n16253) );
  AOI21_X1 U19342 ( .B1(n16254), .B2(n20237), .A(n16253), .ZN(n16255) );
  OAI21_X1 U19343 ( .B1(n16257), .B2(n16256), .A(n16255), .ZN(P1_U3022) );
  AOI21_X1 U19344 ( .B1(n16260), .B2(n16259), .A(n16258), .ZN(n16261) );
  OR2_X1 U19345 ( .A1(n16261), .A2(n9948), .ZN(n20145) );
  INV_X1 U19346 ( .A(n20145), .ZN(n20074) );
  AOI22_X1 U19347 ( .A1(n20234), .A2(n20074), .B1(n20221), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16265) );
  AOI22_X1 U19348 ( .A1(n16263), .A2(n20237), .B1(n16262), .B2(n16266), .ZN(
        n16264) );
  OAI211_X1 U19349 ( .C1(n16267), .C2(n16266), .A(n16265), .B(n16264), .ZN(
        P1_U3024) );
  INV_X1 U19350 ( .A(n16268), .ZN(n20084) );
  AOI22_X1 U19351 ( .A1(n20234), .A2(n20084), .B1(n20221), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16271) );
  AOI22_X1 U19352 ( .A1(n16269), .A2(n20237), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16277), .ZN(n16270) );
  OAI211_X1 U19353 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16272), .A(
        n16271), .B(n16270), .ZN(P1_U3025) );
  NAND2_X1 U19354 ( .A1(n16274), .A2(n16273), .ZN(n16275) );
  AND2_X1 U19355 ( .A1(n16276), .A2(n16275), .ZN(n20151) );
  AOI22_X1 U19356 ( .A1(n20234), .A2(n20151), .B1(n20221), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16283) );
  AOI22_X1 U19357 ( .A1(n16278), .A2(n20237), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16277), .ZN(n16282) );
  NAND3_X1 U19358 ( .A1(n16280), .A2(n16279), .A3(n20236), .ZN(n16281) );
  NAND3_X1 U19359 ( .A1(n16283), .A2(n16282), .A3(n16281), .ZN(P1_U3026) );
  NAND4_X1 U19360 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20964), .A4(n20972), .ZN(n16284) );
  AND2_X1 U19361 ( .A1(n16285), .A2(n16284), .ZN(n20858) );
  NAND2_X1 U19362 ( .A1(n20858), .A2(n16289), .ZN(n16286) );
  AOI22_X1 U19363 ( .A1(n20857), .A2(n16288), .B1(n16287), .B2(n16286), .ZN(
        P1_U3162) );
  OAI22_X1 U19364 ( .A1(n16290), .A2(n20694), .B1(n20968), .B2(n16289), .ZN(
        P1_U3466) );
  AOI211_X1 U19365 ( .C1(n16293), .C2(n16292), .A(n16291), .B(n19888), .ZN(
        n16304) );
  NAND2_X1 U19366 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16294), .ZN(n16295) );
  NAND2_X1 U19367 ( .A1(n19102), .A2(n16295), .ZN(n16298) );
  AOI22_X1 U19368 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19042), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n9962), .ZN(n16297) );
  NAND2_X1 U19369 ( .A1(n19147), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16296) );
  OAI211_X1 U19370 ( .C1(n16299), .C2(n16298), .A(n16297), .B(n16296), .ZN(
        n16300) );
  AOI21_X1 U19371 ( .B1(n16301), .B2(n19135), .A(n16300), .ZN(n16302) );
  INV_X1 U19372 ( .A(n16302), .ZN(n16303) );
  AOI211_X1 U19373 ( .C1(n16306), .C2(n16305), .A(n16304), .B(n16303), .ZN(
        n16307) );
  INV_X1 U19374 ( .A(n16307), .ZN(P2_U2829) );
  AOI211_X1 U19375 ( .C1(n16310), .C2(n16309), .A(n16308), .B(n19888), .ZN(
        n16312) );
  OAI22_X1 U19376 ( .A1(n11285), .A2(n19155), .B1(n19935), .B2(n19110), .ZN(
        n16311) );
  AOI211_X1 U19377 ( .C1(P2_EBX_REG_23__SCAN_IN), .C2(n19147), .A(n16312), .B(
        n16311), .ZN(n16317) );
  INV_X1 U19378 ( .A(n16313), .ZN(n16314) );
  AOI22_X1 U19379 ( .A1(n16315), .A2(n19102), .B1(n19135), .B2(n16314), .ZN(
        n16316) );
  OAI211_X1 U19380 ( .C1(n16318), .C2(n19143), .A(n16317), .B(n16316), .ZN(
        P2_U2832) );
  INV_X1 U19381 ( .A(n16319), .ZN(n19167) );
  AOI22_X1 U19382 ( .A1(n19167), .A2(n19197), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19222), .ZN(n16324) );
  AOI22_X1 U19383 ( .A1(n19169), .A2(BUF1_REG_22__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16323) );
  AOI22_X1 U19384 ( .A1(n16321), .A2(n19210), .B1(n19223), .B2(n16320), .ZN(
        n16322) );
  NAND3_X1 U19385 ( .A1(n16324), .A2(n16323), .A3(n16322), .ZN(P2_U2897) );
  AOI22_X1 U19386 ( .A1(n19167), .A2(n16325), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19222), .ZN(n16331) );
  AOI22_X1 U19387 ( .A1(n19169), .A2(BUF1_REG_20__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16330) );
  INV_X1 U19388 ( .A(n16326), .ZN(n16328) );
  AOI22_X1 U19389 ( .A1(n16328), .A2(n19210), .B1(n19223), .B2(n16327), .ZN(
        n16329) );
  NAND3_X1 U19390 ( .A1(n16331), .A2(n16330), .A3(n16329), .ZN(P2_U2899) );
  AOI22_X1 U19391 ( .A1(n19167), .A2(n16332), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19222), .ZN(n16337) );
  AOI22_X1 U19392 ( .A1(n19169), .A2(BUF1_REG_18__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16336) );
  AOI22_X1 U19393 ( .A1(n16334), .A2(n19210), .B1(n19223), .B2(n16333), .ZN(
        n16335) );
  NAND3_X1 U19394 ( .A1(n16337), .A2(n16336), .A3(n16335), .ZN(P2_U2901) );
  AOI22_X1 U19395 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n16460), .ZN(n16343) );
  INV_X1 U19396 ( .A(n16338), .ZN(n16339) );
  AOI222_X1 U19397 ( .A1(n16341), .A2(n16414), .B1(n16426), .B2(n16340), .C1(
        n16415), .C2(n16339), .ZN(n16342) );
  OAI211_X1 U19398 ( .C1(n16419), .C2(n16344), .A(n16343), .B(n16342), .ZN(
        P2_U2992) );
  AOI22_X1 U19399 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n16460), .ZN(n16351) );
  XNOR2_X1 U19400 ( .A(n16345), .B(n15573), .ZN(n16347) );
  OAI22_X1 U19401 ( .A1(n16347), .A2(n16424), .B1(n16393), .B2(n16346), .ZN(
        n16348) );
  AOI21_X1 U19402 ( .B1(n16349), .B2(n16414), .A(n16348), .ZN(n16350) );
  OAI211_X1 U19403 ( .C1(n16419), .C2(n16352), .A(n16351), .B(n16350), .ZN(
        P2_U2998) );
  AOI22_X1 U19404 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n16460), .B1(n16420), 
        .B2(n19051), .ZN(n16358) );
  OAI22_X1 U19405 ( .A1(n16354), .A2(n16421), .B1(n16424), .B2(n16353), .ZN(
        n16355) );
  AOI21_X1 U19406 ( .B1(n16426), .B2(n16356), .A(n16355), .ZN(n16357) );
  OAI211_X1 U19407 ( .C1(n16429), .C2(n16359), .A(n16358), .B(n16357), .ZN(
        P2_U2999) );
  AOI22_X1 U19408 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n16460), .ZN(n16370) );
  OR2_X1 U19409 ( .A1(n16360), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16361) );
  NAND2_X1 U19410 ( .A1(n16361), .A2(n15572), .ZN(n16439) );
  OR2_X1 U19411 ( .A1(n16436), .A2(n16393), .ZN(n16367) );
  AND2_X1 U19412 ( .A1(n16363), .A2(n16362), .ZN(n16364) );
  XNOR2_X1 U19413 ( .A(n16365), .B(n16364), .ZN(n16435) );
  NAND2_X1 U19414 ( .A1(n16435), .A2(n16414), .ZN(n16366) );
  OAI211_X1 U19415 ( .C1(n16439), .C2(n16424), .A(n16367), .B(n16366), .ZN(
        n16368) );
  INV_X1 U19416 ( .A(n16368), .ZN(n16369) );
  OAI211_X1 U19417 ( .C1(n16419), .C2(n16371), .A(n16370), .B(n16369), .ZN(
        P2_U3000) );
  AOI22_X1 U19418 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n16460), .ZN(n16381) );
  OR2_X1 U19419 ( .A1(n10286), .A2(n16374), .ZN(n16375) );
  XNOR2_X1 U19420 ( .A(n16372), .B(n16375), .ZN(n16449) );
  OR2_X1 U19421 ( .A1(n16376), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16378) );
  NAND2_X1 U19422 ( .A1(n16378), .A2(n16377), .ZN(n16452) );
  INV_X1 U19423 ( .A(n16452), .ZN(n16379) );
  AOI222_X1 U19424 ( .A1(n16449), .A2(n16414), .B1(n16426), .B2(n16448), .C1(
        n16415), .C2(n16379), .ZN(n16380) );
  OAI211_X1 U19425 ( .C1(n16419), .C2(n16382), .A(n16381), .B(n16380), .ZN(
        P2_U3002) );
  AOI22_X1 U19426 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n16460), .B1(n16420), 
        .B2(n19069), .ZN(n16388) );
  OAI22_X1 U19427 ( .A1(n16384), .A2(n16424), .B1(n16383), .B2(n16421), .ZN(
        n16385) );
  AOI21_X1 U19428 ( .B1(n16426), .B2(n16386), .A(n16385), .ZN(n16387) );
  OAI211_X1 U19429 ( .C1(n16429), .C2(n16389), .A(n16388), .B(n16387), .ZN(
        P2_U3003) );
  AOI22_X1 U19430 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n16460), .ZN(n16398) );
  NOR3_X1 U19431 ( .A1(n16391), .A2(n16390), .A3(n16424), .ZN(n16396) );
  OAI22_X1 U19432 ( .A1(n16394), .A2(n16421), .B1(n16393), .B2(n16392), .ZN(
        n16395) );
  NOR2_X1 U19433 ( .A1(n16396), .A2(n16395), .ZN(n16397) );
  OAI211_X1 U19434 ( .C1(n16419), .C2(n19083), .A(n16398), .B(n16397), .ZN(
        P2_U3004) );
  AOI22_X1 U19435 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n16460), .ZN(n16409) );
  OAI21_X1 U19436 ( .B1(n16399), .B2(n16401), .A(n16400), .ZN(n16458) );
  NOR2_X1 U19437 ( .A1(n16404), .A2(n10051), .ZN(n16405) );
  XNOR2_X1 U19438 ( .A(n16402), .B(n16405), .ZN(n16456) );
  AOI22_X1 U19439 ( .A1(n16456), .A2(n16414), .B1(n16426), .B2(n16455), .ZN(
        n16406) );
  OAI21_X1 U19440 ( .B1(n16458), .B2(n16424), .A(n16406), .ZN(n16407) );
  INV_X1 U19441 ( .A(n16407), .ZN(n16408) );
  OAI211_X1 U19442 ( .C1(n16419), .C2(n16410), .A(n16409), .B(n16408), .ZN(
        P2_U3006) );
  AOI22_X1 U19443 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n16460), .ZN(n16418) );
  INV_X1 U19444 ( .A(n16412), .ZN(n16416) );
  AOI222_X1 U19445 ( .A1(n16416), .A2(n16415), .B1(n16414), .B2(n16413), .C1(
        n16426), .C2(n19120), .ZN(n16417) );
  OAI211_X1 U19446 ( .C1(n16419), .C2(n19118), .A(n16418), .B(n16417), .ZN(
        P2_U3008) );
  AOI22_X1 U19447 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n16460), .B1(n16420), 
        .B2(n19133), .ZN(n16428) );
  OAI22_X1 U19448 ( .A1(n16424), .A2(n16423), .B1(n16422), .B2(n16421), .ZN(
        n16425) );
  AOI21_X1 U19449 ( .B1(n16426), .B2(n19134), .A(n16425), .ZN(n16427) );
  OAI211_X1 U19450 ( .C1(n16429), .C2(n19127), .A(n16428), .B(n16427), .ZN(
        P2_U3009) );
  INV_X1 U19451 ( .A(n16430), .ZN(n16432) );
  AOI211_X1 U19452 ( .C1(n16432), .C2(n12774), .A(n16445), .B(n16431), .ZN(
        n16434) );
  NOR2_X1 U19453 ( .A1(n19324), .A2(n11930), .ZN(n16433) );
  AOI211_X1 U19454 ( .C1(n19310), .C2(n19178), .A(n16434), .B(n16433), .ZN(
        n16442) );
  NAND2_X1 U19455 ( .A1(n16435), .A2(n16475), .ZN(n16438) );
  OR2_X1 U19456 ( .A1(n16436), .A2(n19312), .ZN(n16437) );
  OAI211_X1 U19457 ( .C1(n16439), .C2(n19318), .A(n16438), .B(n16437), .ZN(
        n16440) );
  INV_X1 U19458 ( .A(n16440), .ZN(n16441) );
  OAI211_X1 U19459 ( .C1(n16444), .C2(n12774), .A(n16442), .B(n16441), .ZN(
        P2_U3032) );
  NAND2_X1 U19460 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n16460), .ZN(n16443) );
  OAI221_X1 U19461 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16445), 
        .C1(n12734), .C2(n16444), .A(n16443), .ZN(n16446) );
  AOI21_X1 U19462 ( .B1(n19310), .B2(n16447), .A(n16446), .ZN(n16451) );
  AOI22_X1 U19463 ( .A1(n16449), .A2(n16475), .B1(n16471), .B2(n16448), .ZN(
        n16450) );
  OAI211_X1 U19464 ( .C1(n19318), .C2(n16452), .A(n16451), .B(n16450), .ZN(
        P2_U3034) );
  AOI22_X1 U19465 ( .A1(n16454), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19310), .B2(n16453), .ZN(n16466) );
  AOI22_X1 U19466 ( .A1(n16456), .A2(n16475), .B1(n16471), .B2(n16455), .ZN(
        n16457) );
  OAI21_X1 U19467 ( .B1(n16458), .B2(n19318), .A(n16457), .ZN(n16459) );
  INV_X1 U19468 ( .A(n16459), .ZN(n16465) );
  NAND2_X1 U19469 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16460), .ZN(n16464) );
  OAI211_X1 U19470 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16462), .B(n16461), .ZN(n16463) );
  NAND4_X1 U19471 ( .A1(n16466), .A2(n16465), .A3(n16464), .A4(n16463), .ZN(
        P2_U3038) );
  INV_X1 U19472 ( .A(n16467), .ZN(n16480) );
  OAI21_X1 U19473 ( .B1(n16469), .B2(n19214), .A(n16468), .ZN(n16470) );
  AOI21_X1 U19474 ( .B1(n16471), .B2(n12566), .A(n16470), .ZN(n16472) );
  OAI21_X1 U19475 ( .B1(n16473), .B2(n19318), .A(n16472), .ZN(n16474) );
  AOI21_X1 U19476 ( .B1(n16476), .B2(n16475), .A(n16474), .ZN(n16477) );
  OAI221_X1 U19477 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16480), .C1(
        n16479), .C2(n16478), .A(n16477), .ZN(P2_U3043) );
  NAND2_X1 U19478 ( .A1(n16485), .A2(n19996), .ZN(n16483) );
  NOR2_X1 U19479 ( .A1(n16481), .A2(n20006), .ZN(n16482) );
  NAND2_X1 U19480 ( .A1(n16483), .A2(n16482), .ZN(n16484) );
  OAI211_X1 U19481 ( .C1(n19996), .C2(n16485), .A(n16484), .B(n16533), .ZN(
        n16486) );
  AOI21_X1 U19482 ( .B1(n16514), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16486), .ZN(n16506) );
  INV_X1 U19483 ( .A(n16506), .ZN(n16487) );
  NAND2_X1 U19484 ( .A1(n16487), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16504) );
  INV_X1 U19485 ( .A(n16491), .ZN(n16490) );
  INV_X1 U19486 ( .A(n16488), .ZN(n16489) );
  OAI21_X1 U19487 ( .B1(n16490), .B2(n16492), .A(n16489), .ZN(n16494) );
  NAND3_X1 U19488 ( .A1(n16492), .A2(n15885), .A3(n16491), .ZN(n16493) );
  NAND2_X1 U19489 ( .A1(n16494), .A2(n16493), .ZN(n16499) );
  NAND2_X1 U19490 ( .A1(n16495), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16496) );
  MUX2_X1 U19491 ( .A(n16497), .B(n16496), .S(n15879), .Z(n16498) );
  NAND2_X1 U19492 ( .A1(n16499), .A2(n16498), .ZN(n16500) );
  AOI21_X1 U19493 ( .B1(n16502), .B2(n16501), .A(n16500), .ZN(n19964) );
  NOR2_X1 U19494 ( .A1(n16533), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16503) );
  AOI21_X1 U19495 ( .B1(n19964), .B2(n16533), .A(n16503), .ZN(n16509) );
  NAND3_X1 U19496 ( .A1(n16504), .A2(n16509), .A3(n19980), .ZN(n16508) );
  NAND2_X1 U19497 ( .A1(n16506), .A2(n16505), .ZN(n16507) );
  NAND2_X1 U19498 ( .A1(n16508), .A2(n16507), .ZN(n16513) );
  OAI21_X1 U19499 ( .B1(n16513), .B2(n19980), .A(n16512), .ZN(n16511) );
  INV_X1 U19500 ( .A(n16509), .ZN(n16510) );
  NAND2_X1 U19501 ( .A1(n16511), .A2(n16510), .ZN(n16536) );
  NAND2_X1 U19502 ( .A1(n16513), .A2(n16512), .ZN(n16516) );
  MUX2_X1 U19503 ( .A(n11408), .B(n16514), .S(n16533), .Z(n16515) );
  NAND2_X1 U19504 ( .A1(n16516), .A2(n16515), .ZN(n16535) );
  NAND2_X1 U19505 ( .A1(n16518), .A2(n16517), .ZN(n16525) );
  INV_X1 U19506 ( .A(n16519), .ZN(n16520) );
  AOI22_X1 U19507 ( .A1(n16523), .A2(n16522), .B1(n16521), .B2(n16520), .ZN(
        n16524) );
  AND2_X1 U19508 ( .A1(n16525), .A2(n16524), .ZN(n20014) );
  INV_X1 U19509 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n16526) );
  NAND2_X1 U19510 ( .A1(n16020), .A2(n16526), .ZN(n16530) );
  OAI22_X1 U19511 ( .A1(n16528), .A2(n16527), .B1(n20028), .B2(n12818), .ZN(
        n16529) );
  AOI21_X1 U19512 ( .B1(n16531), .B2(n16530), .A(n16529), .ZN(n16532) );
  OAI211_X1 U19513 ( .C1(n16533), .C2(n13100), .A(n20014), .B(n16532), .ZN(
        n16534) );
  AOI21_X1 U19514 ( .B1(n16536), .B2(n16535), .A(n16534), .ZN(n16554) );
  AOI211_X1 U19515 ( .C1(n16539), .C2(n16538), .A(n19886), .B(n16537), .ZN(
        n16552) );
  NAND2_X1 U19516 ( .A1(n16554), .A2(n16540), .ZN(n16541) );
  NAND2_X1 U19517 ( .A1(n16541), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16547) );
  NAND2_X1 U19518 ( .A1(n15191), .A2(n16542), .ZN(n16544) );
  OAI211_X1 U19519 ( .C1(n11612), .C2(n16544), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n16543), .ZN(n16545) );
  INV_X1 U19520 ( .A(n16545), .ZN(n16546) );
  NOR2_X1 U19521 ( .A1(n20026), .A2(n19885), .ZN(n19887) );
  AOI211_X1 U19522 ( .C1(n20024), .C2(n16548), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n19887), .ZN(n16549) );
  AOI21_X1 U19523 ( .B1(n16550), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16549), 
        .ZN(n16551) );
  OAI211_X1 U19524 ( .C1(n16554), .C2(n16553), .A(n16552), .B(n16551), .ZN(
        P2_U3176) );
  OAI221_X1 U19525 ( .B1(n19825), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19825), 
        .C2(n19885), .A(n16555), .ZN(P2_U3593) );
  XOR2_X1 U19526 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16575), .Z(
        n16739) );
  INV_X1 U19527 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16740) );
  OAI221_X1 U19528 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16558), .C1(
        n16740), .C2(n16557), .A(n16556), .ZN(n16559) );
  AOI21_X1 U19529 ( .B1(n17846), .B2(n16739), .A(n16559), .ZN(n16565) );
  OAI22_X1 U19530 ( .A1(n16568), .A2(n17998), .B1(n16570), .B2(n17906), .ZN(
        n16563) );
  OAI22_X2 U19531 ( .A1(n18191), .A2(n17998), .B1(n17906), .B2(n18189), .ZN(
        n17874) );
  NOR2_X1 U19532 ( .A1(n16561), .A2(n17792), .ZN(n17647) );
  AOI22_X1 U19533 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16563), .B1(
        n16562), .B2(n17647), .ZN(n16564) );
  OAI211_X1 U19534 ( .C1(n16566), .C2(n17877), .A(n16565), .B(n16564), .ZN(
        P3_U2800) );
  INV_X1 U19535 ( .A(n16567), .ZN(n18003) );
  NAND2_X1 U19536 ( .A1(n18003), .A2(n16569), .ZN(n16601) );
  AOI211_X1 U19537 ( .C1(n16571), .C2(n16601), .A(n16568), .B(n17998), .ZN(
        n16573) );
  NAND2_X1 U19538 ( .A1(n16569), .A2(n18002), .ZN(n16600) );
  AOI211_X1 U19539 ( .C1(n16571), .C2(n16600), .A(n16570), .B(n17906), .ZN(
        n16572) );
  AOI211_X1 U19540 ( .C1(n16574), .C2(n17903), .A(n16573), .B(n16572), .ZN(
        n16582) );
  NAND2_X1 U19541 ( .A1(n9816), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16581) );
  INV_X1 U19542 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16748) );
  AOI21_X1 U19543 ( .B1(n16748), .B2(n16717), .A(n16575), .ZN(n16747) );
  OAI21_X1 U19544 ( .B1(n16576), .B2(n17846), .A(n16747), .ZN(n16580) );
  OAI221_X1 U19545 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16578), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18705), .A(n16577), .ZN(
        n16579) );
  NAND4_X1 U19546 ( .A1(n16582), .A2(n16581), .A3(n16580), .A4(n16579), .ZN(
        P3_U2801) );
  INV_X1 U19547 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18926) );
  NAND2_X1 U19548 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18926), .ZN(
        n16584) );
  NOR4_X1 U19549 ( .A1(n18026), .A2(n16584), .A3(n16583), .A4(n18302), .ZN(
        n16588) );
  INV_X1 U19550 ( .A(n18308), .ZN(n18273) );
  AOI221_X1 U19551 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16585), 
        .C1(n18273), .C2(n16585), .A(n18926), .ZN(n16587) );
  AOI211_X1 U19552 ( .C1(n16589), .C2(n16588), .A(n16587), .B(n16586), .ZN(
        n16594) );
  AOI22_X1 U19553 ( .A1(n16592), .A2(n18307), .B1(n16591), .B2(n16590), .ZN(
        n16593) );
  OAI211_X1 U19554 ( .C1(n16595), .C2(n18221), .A(n16594), .B(n16593), .ZN(
        P3_U2831) );
  NOR2_X1 U19555 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n9992), .ZN(
        n17643) );
  AOI22_X1 U19556 ( .A1(n9816), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18008), 
        .B2(n17643), .ZN(n16610) );
  INV_X1 U19557 ( .A(n16596), .ZN(n16598) );
  NOR2_X1 U19558 ( .A1(n18302), .A2(n18963), .ZN(n18305) );
  NAND3_X1 U19559 ( .A1(n16598), .A2(n18305), .A3(n17640), .ZN(n16609) );
  AOI21_X1 U19560 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17780), .A(
        n16598), .ZN(n17639) );
  NAND3_X1 U19561 ( .A1(n16597), .A2(n18236), .A3(n17639), .ZN(n16608) );
  NOR2_X1 U19562 ( .A1(n17640), .A2(n17639), .ZN(n17638) );
  NOR3_X1 U19563 ( .A1(n17638), .A2(n16599), .A3(n10301), .ZN(n16606) );
  NOR2_X1 U19564 ( .A1(n18784), .A2(n18768), .ZN(n18205) );
  AOI22_X1 U19565 ( .A1(n18959), .A2(n16601), .B1(n18190), .B2(n16600), .ZN(
        n16602) );
  OAI211_X1 U19566 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18205), .A(
        n16603), .B(n16602), .ZN(n16605) );
  OAI21_X1 U19567 ( .B1(n16606), .B2(n16605), .A(n16604), .ZN(n16607) );
  NAND4_X1 U19568 ( .A1(n16610), .A2(n16609), .A3(n16608), .A4(n16607), .ZN(
        P3_U2834) );
  NOR3_X1 U19569 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16612) );
  NOR4_X1 U19570 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16611) );
  NAND4_X1 U19571 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16612), .A3(n16611), .A4(
        U215), .ZN(U213) );
  INV_X2 U19572 ( .A(U214), .ZN(n16649) );
  NOR2_X1 U19573 ( .A1(n16649), .A2(n16613), .ZN(n16647) );
  INV_X1 U19574 ( .A(U212), .ZN(n16650) );
  AOI222_X1 U19575 ( .A1(n16649), .A2(P1_DATAO_REG_31__SCAN_IN), .B1(n16647), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n16650), .C2(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n16614) );
  INV_X1 U19576 ( .A(n16614), .ZN(U216) );
  INV_X1 U19577 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16686) );
  INV_X1 U19578 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20330) );
  INV_X1 U19579 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n21222) );
  OAI222_X1 U19580 ( .A1(U214), .A2(n16686), .B1(n16652), .B2(n20330), .C1(
        U212), .C2(n21222), .ZN(U217) );
  INV_X1 U19581 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20322) );
  AOI22_X1 U19582 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16649), .ZN(n16615) );
  OAI21_X1 U19583 ( .B1(n20322), .B2(n16652), .A(n16615), .ZN(U218) );
  INV_X1 U19584 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20314) );
  AOI22_X1 U19585 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16649), .ZN(n16616) );
  OAI21_X1 U19586 ( .B1(n20314), .B2(n16652), .A(n16616), .ZN(U219) );
  INV_X1 U19587 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20306) );
  AOI22_X1 U19588 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16649), .ZN(n16617) );
  OAI21_X1 U19589 ( .B1(n20306), .B2(n16652), .A(n16617), .ZN(U220) );
  INV_X1 U19590 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20297) );
  AOI22_X1 U19591 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16649), .ZN(n16618) );
  OAI21_X1 U19592 ( .B1(n20297), .B2(n16652), .A(n16618), .ZN(U221) );
  AOI22_X1 U19593 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16649), .ZN(n16619) );
  OAI21_X1 U19594 ( .B1(n20286), .B2(n16652), .A(n16619), .ZN(U222) );
  INV_X1 U19595 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20272) );
  AOI22_X1 U19596 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16649), .ZN(n16620) );
  OAI21_X1 U19597 ( .B1(n20272), .B2(n16652), .A(n16620), .ZN(U223) );
  AOI22_X1 U19598 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16649), .ZN(n16621) );
  OAI21_X1 U19599 ( .B1(n20336), .B2(n16652), .A(n16621), .ZN(U224) );
  INV_X1 U19600 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n16622) );
  INV_X1 U19601 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20327) );
  INV_X1 U19602 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21180) );
  OAI222_X1 U19603 ( .A1(U214), .A2(n16622), .B1(n16652), .B2(n20327), .C1(
        U212), .C2(n21180), .ZN(U225) );
  AOI22_X1 U19604 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16649), .ZN(n16623) );
  OAI21_X1 U19605 ( .B1(n15457), .B2(n16652), .A(n16623), .ZN(U226) );
  AOI22_X1 U19606 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16649), .ZN(n16624) );
  OAI21_X1 U19607 ( .B1(n14594), .B2(n16652), .A(n16624), .ZN(U227) );
  AOI22_X1 U19608 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16649), .ZN(n16625) );
  OAI21_X1 U19609 ( .B1(n20304), .B2(n16652), .A(n16625), .ZN(U228) );
  AOI22_X1 U19610 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16649), .ZN(n16626) );
  OAI21_X1 U19611 ( .B1(n20294), .B2(n16652), .A(n16626), .ZN(U229) );
  AOI22_X1 U19612 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16649), .ZN(n16627) );
  OAI21_X1 U19613 ( .B1(n13792), .B2(n16652), .A(n16627), .ZN(U230) );
  INV_X1 U19614 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20281) );
  AOI22_X1 U19615 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16649), .ZN(n16628) );
  OAI21_X1 U19616 ( .B1(n20281), .B2(n16652), .A(n16628), .ZN(U231) );
  INV_X1 U19617 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n21137) );
  AOI22_X1 U19618 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16649), .ZN(n16629) );
  OAI21_X1 U19619 ( .B1(n21137), .B2(U212), .A(n16629), .ZN(U232) );
  INV_X1 U19620 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16669) );
  AOI22_X1 U19621 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16649), .ZN(n16630) );
  OAI21_X1 U19622 ( .B1(n16669), .B2(U212), .A(n16630), .ZN(U233) );
  INV_X1 U19623 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n21259) );
  AOI22_X1 U19624 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16649), .ZN(n16631) );
  OAI21_X1 U19625 ( .B1(n21259), .B2(U212), .A(n16631), .ZN(U234) );
  AOI22_X1 U19626 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16649), .ZN(n16632) );
  OAI21_X1 U19627 ( .B1(n16633), .B2(n16652), .A(n16632), .ZN(U235) );
  INV_X1 U19628 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16666) );
  AOI22_X1 U19629 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16649), .ZN(n16634) );
  OAI21_X1 U19630 ( .B1(n16666), .B2(U212), .A(n16634), .ZN(U236) );
  INV_X1 U19631 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n21156) );
  INV_X1 U19632 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16665) );
  OAI222_X1 U19633 ( .A1(U214), .A2(n21156), .B1(n16652), .B2(n16635), .C1(
        U212), .C2(n16665), .ZN(U237) );
  INV_X1 U19634 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16664) );
  AOI22_X1 U19635 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16649), .ZN(n16636) );
  OAI21_X1 U19636 ( .B1(n16664), .B2(U212), .A(n16636), .ZN(U238) );
  AOI22_X1 U19637 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16649), .ZN(n16637) );
  OAI21_X1 U19638 ( .B1(n16638), .B2(n16652), .A(n16637), .ZN(U239) );
  INV_X1 U19639 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16661) );
  AOI22_X1 U19640 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16649), .ZN(n16639) );
  OAI21_X1 U19641 ( .B1(n16661), .B2(U212), .A(n16639), .ZN(U240) );
  AOI22_X1 U19642 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16649), .ZN(n16640) );
  OAI21_X1 U19643 ( .B1(n16641), .B2(n16652), .A(n16640), .ZN(U241) );
  INV_X1 U19644 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16659) );
  AOI22_X1 U19645 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16649), .ZN(n16642) );
  OAI21_X1 U19646 ( .B1(n16659), .B2(U212), .A(n16642), .ZN(U242) );
  INV_X1 U19647 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n21086) );
  AOI22_X1 U19648 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16649), .ZN(n16643) );
  OAI21_X1 U19649 ( .B1(n21086), .B2(n16652), .A(n16643), .ZN(U243) );
  INV_X1 U19650 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16657) );
  AOI22_X1 U19651 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16649), .ZN(n16644) );
  OAI21_X1 U19652 ( .B1(n16657), .B2(U212), .A(n16644), .ZN(U244) );
  AOI22_X1 U19653 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16649), .ZN(n16645) );
  OAI21_X1 U19654 ( .B1(n16646), .B2(n16652), .A(n16645), .ZN(U245) );
  INV_X1 U19655 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16655) );
  AOI22_X1 U19656 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16647), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16649), .ZN(n16648) );
  OAI21_X1 U19657 ( .B1(n16655), .B2(U212), .A(n16648), .ZN(U246) );
  AOI22_X1 U19658 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16650), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16649), .ZN(n16651) );
  OAI21_X1 U19659 ( .B1(n16653), .B2(n16652), .A(n16651), .ZN(U247) );
  INV_X1 U19660 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16654) );
  AOI22_X1 U19661 ( .A1(n16684), .A2(n16654), .B1(n18330), .B2(U215), .ZN(U251) );
  INV_X1 U19662 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U19663 ( .A1(n16670), .A2(n16655), .B1(n18339), .B2(U215), .ZN(U252) );
  INV_X1 U19664 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16656) );
  AOI22_X1 U19665 ( .A1(n16684), .A2(n16656), .B1(n21142), .B2(U215), .ZN(U253) );
  INV_X1 U19666 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18347) );
  AOI22_X1 U19667 ( .A1(n16684), .A2(n16657), .B1(n18347), .B2(U215), .ZN(U254) );
  INV_X1 U19668 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16658) );
  INV_X1 U19669 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U19670 ( .A1(n16670), .A2(n16658), .B1(n18352), .B2(U215), .ZN(U255) );
  INV_X1 U19671 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21246) );
  AOI22_X1 U19672 ( .A1(n16670), .A2(n16659), .B1(n21246), .B2(U215), .ZN(U256) );
  INV_X1 U19673 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16660) );
  AOI22_X1 U19674 ( .A1(n16670), .A2(n16660), .B1(n18362), .B2(U215), .ZN(U257) );
  INV_X1 U19675 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18370) );
  AOI22_X1 U19676 ( .A1(n16670), .A2(n16661), .B1(n18370), .B2(U215), .ZN(U258) );
  INV_X1 U19677 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16662) );
  INV_X1 U19678 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n21192) );
  AOI22_X1 U19679 ( .A1(n16670), .A2(n16662), .B1(n21192), .B2(U215), .ZN(U259) );
  INV_X1 U19680 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n16663) );
  AOI22_X1 U19681 ( .A1(n16684), .A2(n16664), .B1(n16663), .B2(U215), .ZN(U260) );
  INV_X1 U19682 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U19683 ( .A1(n16670), .A2(n16665), .B1(n17614), .B2(U215), .ZN(U261) );
  INV_X1 U19684 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U19685 ( .A1(n16670), .A2(n16666), .B1(n17616), .B2(U215), .ZN(U262) );
  INV_X1 U19686 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16667) );
  INV_X1 U19687 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U19688 ( .A1(n16684), .A2(n16667), .B1(n17618), .B2(U215), .ZN(U263) );
  INV_X1 U19689 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U19690 ( .A1(n16670), .A2(n21259), .B1(n17622), .B2(U215), .ZN(U264) );
  INV_X1 U19691 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16668) );
  AOI22_X1 U19692 ( .A1(n16670), .A2(n16669), .B1(n16668), .B2(U215), .ZN(U265) );
  INV_X1 U19693 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U19694 ( .A1(n16684), .A2(n21137), .B1(n17628), .B2(U215), .ZN(U266) );
  OAI22_X1 U19695 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16684), .ZN(n16671) );
  INV_X1 U19696 ( .A(n16671), .ZN(U267) );
  INV_X1 U19697 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16672) );
  AOI22_X1 U19698 ( .A1(n16684), .A2(n16672), .B1(n13791), .B2(U215), .ZN(U268) );
  INV_X1 U19699 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16673) );
  AOI22_X1 U19700 ( .A1(n16684), .A2(n16673), .B1(n18343), .B2(U215), .ZN(U269) );
  INV_X1 U19701 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16674) );
  AOI22_X1 U19702 ( .A1(n16684), .A2(n16674), .B1(n18348), .B2(U215), .ZN(U270) );
  INV_X1 U19703 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16675) );
  INV_X1 U19704 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U19705 ( .A1(n16684), .A2(n16675), .B1(n18351), .B2(U215), .ZN(U271) );
  INV_X1 U19706 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16676) );
  AOI22_X1 U19707 ( .A1(n16684), .A2(n16676), .B1(n15455), .B2(U215), .ZN(U272) );
  INV_X1 U19708 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U19709 ( .A1(n16684), .A2(n21180), .B1(n18363), .B2(U215), .ZN(U273) );
  INV_X1 U19710 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16677) );
  AOI22_X1 U19711 ( .A1(n16684), .A2(n16677), .B1(n15450), .B2(U215), .ZN(U274) );
  OAI22_X1 U19712 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16684), .ZN(n16678) );
  INV_X1 U19713 ( .A(n16678), .ZN(U275) );
  OAI22_X1 U19714 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16684), .ZN(n16679) );
  INV_X1 U19715 ( .A(n16679), .ZN(U276) );
  OAI22_X1 U19716 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16684), .ZN(n16680) );
  INV_X1 U19717 ( .A(n16680), .ZN(U277) );
  OAI22_X1 U19718 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16684), .ZN(n16681) );
  INV_X1 U19719 ( .A(n16681), .ZN(U278) );
  INV_X1 U19720 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16682) );
  INV_X1 U19721 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21189) );
  AOI22_X1 U19722 ( .A1(n16684), .A2(n16682), .B1(n21189), .B2(U215), .ZN(U279) );
  INV_X1 U19723 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16683) );
  INV_X1 U19724 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18358) );
  AOI22_X1 U19725 ( .A1(n16684), .A2(n16683), .B1(n18358), .B2(U215), .ZN(U280) );
  INV_X1 U19726 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19346) );
  AOI22_X1 U19727 ( .A1(n16684), .A2(n21222), .B1(n19346), .B2(U215), .ZN(U281) );
  INV_X1 U19728 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n21176) );
  INV_X1 U19729 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U19730 ( .A1(n16684), .A2(n21176), .B1(n18369), .B2(U215), .ZN(U282) );
  INV_X1 U19731 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16685) );
  OAI222_X1 U19732 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n21222), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n16686), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16685), .ZN(n16687) );
  INV_X1 U19733 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18867) );
  INV_X1 U19734 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19918) );
  AOI22_X1 U19735 ( .A1(n16689), .A2(n18867), .B1(n19918), .B2(n16688), .ZN(
        U347) );
  INV_X1 U19736 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18865) );
  INV_X1 U19737 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19917) );
  AOI22_X1 U19738 ( .A1(n16689), .A2(n18865), .B1(n19917), .B2(n16688), .ZN(
        U348) );
  INV_X1 U19739 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18862) );
  INV_X1 U19740 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19916) );
  AOI22_X1 U19741 ( .A1(n16689), .A2(n18862), .B1(n19916), .B2(n16688), .ZN(
        U349) );
  INV_X1 U19742 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18861) );
  INV_X1 U19743 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U19744 ( .A1(n16689), .A2(n18861), .B1(n19915), .B2(n16688), .ZN(
        U350) );
  INV_X1 U19745 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18859) );
  INV_X1 U19746 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19747 ( .A1(n16689), .A2(n18859), .B1(n19914), .B2(n16687), .ZN(
        U351) );
  INV_X1 U19748 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18857) );
  INV_X1 U19749 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U19750 ( .A1(n16689), .A2(n18857), .B1(n19913), .B2(n16687), .ZN(
        U352) );
  INV_X2 U19751 ( .A(n16688), .ZN(n16689) );
  INV_X1 U19752 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18855) );
  INV_X1 U19753 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19912) );
  AOI22_X1 U19754 ( .A1(n16689), .A2(n18855), .B1(n19912), .B2(n16687), .ZN(
        U353) );
  INV_X1 U19755 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18853) );
  AOI22_X1 U19756 ( .A1(n16689), .A2(n18853), .B1(n19911), .B2(n16688), .ZN(
        U354) );
  INV_X1 U19757 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18906) );
  INV_X1 U19758 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U19759 ( .A1(n16689), .A2(n18906), .B1(n19949), .B2(n16688), .ZN(
        U355) );
  INV_X1 U19760 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18904) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19946) );
  AOI22_X1 U19762 ( .A1(n16689), .A2(n18904), .B1(n19946), .B2(n16688), .ZN(
        U356) );
  INV_X1 U19763 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18902) );
  INV_X1 U19764 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19944) );
  AOI22_X1 U19765 ( .A1(n16689), .A2(n18902), .B1(n19944), .B2(n16688), .ZN(
        U357) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18900) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19942) );
  AOI22_X1 U19768 ( .A1(n16689), .A2(n18900), .B1(n19942), .B2(n16688), .ZN(
        U358) );
  INV_X1 U19769 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18899) );
  INV_X1 U19770 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21231) );
  AOI22_X1 U19771 ( .A1(n16689), .A2(n18899), .B1(n21231), .B2(n16688), .ZN(
        U359) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18897) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19940) );
  AOI22_X1 U19774 ( .A1(n16689), .A2(n18897), .B1(n19940), .B2(n16687), .ZN(
        U360) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18895) );
  INV_X1 U19776 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19938) );
  AOI22_X1 U19777 ( .A1(n16689), .A2(n18895), .B1(n19938), .B2(n16687), .ZN(
        U361) );
  INV_X1 U19778 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18892) );
  INV_X1 U19779 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19936) );
  AOI22_X1 U19780 ( .A1(n16689), .A2(n18892), .B1(n19936), .B2(n16687), .ZN(
        U362) );
  INV_X1 U19781 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18891) );
  INV_X1 U19782 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19934) );
  AOI22_X1 U19783 ( .A1(n16689), .A2(n18891), .B1(n19934), .B2(n16687), .ZN(
        U363) );
  INV_X1 U19784 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18888) );
  INV_X1 U19785 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19933) );
  AOI22_X1 U19786 ( .A1(n16689), .A2(n18888), .B1(n19933), .B2(n16687), .ZN(
        U364) );
  INV_X1 U19787 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18851) );
  INV_X1 U19788 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19910) );
  AOI22_X1 U19789 ( .A1(n16689), .A2(n18851), .B1(n19910), .B2(n16688), .ZN(
        U365) );
  INV_X1 U19790 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18887) );
  INV_X1 U19791 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U19792 ( .A1(n16689), .A2(n18887), .B1(n19931), .B2(n16688), .ZN(
        U366) );
  INV_X1 U19793 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18885) );
  INV_X1 U19794 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U19795 ( .A1(n16689), .A2(n18885), .B1(n19929), .B2(n16688), .ZN(
        U367) );
  INV_X1 U19796 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18883) );
  INV_X1 U19797 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U19798 ( .A1(n16689), .A2(n18883), .B1(n19927), .B2(n16688), .ZN(
        U368) );
  INV_X1 U19799 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18880) );
  INV_X1 U19800 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19926) );
  AOI22_X1 U19801 ( .A1(n16689), .A2(n18880), .B1(n19926), .B2(n16688), .ZN(
        U369) );
  INV_X1 U19802 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18879) );
  INV_X1 U19803 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19924) );
  AOI22_X1 U19804 ( .A1(n16689), .A2(n18879), .B1(n19924), .B2(n16688), .ZN(
        U370) );
  INV_X1 U19805 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18877) );
  INV_X1 U19806 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U19807 ( .A1(n16689), .A2(n18877), .B1(n19923), .B2(n16688), .ZN(
        U371) );
  INV_X1 U19808 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18874) );
  INV_X1 U19809 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19922) );
  AOI22_X1 U19810 ( .A1(n16689), .A2(n18874), .B1(n19922), .B2(n16688), .ZN(
        U372) );
  INV_X1 U19811 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18873) );
  INV_X1 U19812 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19921) );
  AOI22_X1 U19813 ( .A1(n16689), .A2(n18873), .B1(n19921), .B2(n16688), .ZN(
        U373) );
  INV_X1 U19814 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18871) );
  INV_X1 U19815 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19920) );
  AOI22_X1 U19816 ( .A1(n16689), .A2(n18871), .B1(n19920), .B2(n16688), .ZN(
        U374) );
  INV_X1 U19817 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18869) );
  INV_X1 U19818 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19919) );
  AOI22_X1 U19819 ( .A1(n16689), .A2(n18869), .B1(n19919), .B2(n16688), .ZN(
        U375) );
  INV_X1 U19820 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18848) );
  INV_X1 U19821 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U19822 ( .A1(n16689), .A2(n18848), .B1(n19909), .B2(n16688), .ZN(
        U376) );
  INV_X1 U19823 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16690) );
  INV_X1 U19824 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18847) );
  NAND2_X1 U19825 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18847), .ZN(n18833) );
  AOI22_X1 U19826 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18833), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18845), .ZN(n18917) );
  OAI21_X1 U19827 ( .B1(n18845), .B2(n16690), .A(n18915), .ZN(P3_U2633) );
  INV_X1 U19828 ( .A(n17580), .ZN(n16710) );
  OAI21_X1 U19829 ( .B1(n16696), .B2(n16710), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16691) );
  OAI21_X1 U19830 ( .B1(n16692), .B2(n18822), .A(n16691), .ZN(P3_U2634) );
  AOI21_X1 U19831 ( .B1(n18845), .B2(n18847), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16693) );
  AOI22_X1 U19832 ( .A1(n18980), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16693), 
        .B2(n18981), .ZN(P3_U2635) );
  NOR2_X1 U19833 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18830) );
  OAI21_X1 U19834 ( .B1(n18830), .B2(BS16), .A(n18917), .ZN(n18916) );
  OAI21_X1 U19835 ( .B1(n18917), .B2(n18971), .A(n18916), .ZN(P3_U2636) );
  INV_X1 U19836 ( .A(n16694), .ZN(n16695) );
  NOR3_X1 U19837 ( .A1(n16696), .A2(n18763), .A3(n16695), .ZN(n18765) );
  NOR2_X1 U19838 ( .A1(n18765), .A2(n18817), .ZN(n18964) );
  OAI21_X1 U19839 ( .B1(n18964), .B2(n21210), .A(n16697), .ZN(P3_U2637) );
  NOR4_X1 U19840 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16707) );
  NOR4_X1 U19841 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16706) );
  INV_X1 U19842 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21254) );
  INV_X1 U19843 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21102) );
  NOR4_X1 U19844 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16698) );
  OAI21_X1 U19845 ( .B1(n21254), .B2(n21102), .A(n16698), .ZN(n16704) );
  NOR4_X1 U19846 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16702) );
  NOR4_X1 U19847 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16701) );
  NOR4_X1 U19848 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16700) );
  NOR4_X1 U19849 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16699) );
  NAND4_X1 U19850 ( .A1(n16702), .A2(n16701), .A3(n16700), .A4(n16699), .ZN(
        n16703) );
  NOR4_X1 U19851 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(n16704), .A4(n16703), .ZN(n16705)
         );
  NAND3_X1 U19852 ( .A1(n16707), .A2(n16706), .A3(n16705), .ZN(n18953) );
  NOR2_X1 U19853 ( .A1(n18953), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18955) );
  INV_X1 U19854 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18954) );
  NAND3_X1 U19855 ( .A1(n18954), .A2(n21254), .A3(n21102), .ZN(n16709) );
  INV_X1 U19856 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18912) );
  AOI22_X1 U19857 ( .A1(n18955), .A2(n16709), .B1(n18953), .B2(n18912), .ZN(
        P3_U2638) );
  AOI22_X1 U19858 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18953), .B1(n18955), .B2(n21102), .ZN(n16708) );
  OAI21_X1 U19859 ( .B1(n18953), .B2(n16709), .A(n16708), .ZN(P3_U2639) );
  NOR3_X1 U19860 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18829) );
  NAND2_X1 U19861 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18829), .ZN(n18825) );
  NOR2_X1 U19862 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18920), .ZN(n18820) );
  INV_X1 U19863 ( .A(n18820), .ZN(n18699) );
  OR2_X1 U19864 ( .A1(n18822), .A2(n18699), .ZN(n18815) );
  INV_X1 U19865 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18903) );
  INV_X1 U19866 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18901) );
  INV_X1 U19867 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21163) );
  NOR3_X1 U19868 ( .A1(n18903), .A2(n18901), .A3(n21163), .ZN(n16713) );
  AOI211_X1 U19869 ( .C1(n18972), .C2(n18970), .A(n18836), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16714) );
  INV_X1 U19870 ( .A(n16714), .ZN(n18810) );
  NAND2_X1 U19871 ( .A1(n17021), .A2(n16711), .ZN(n16716) );
  INV_X1 U19872 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18894) );
  INV_X1 U19873 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18872) );
  INV_X1 U19874 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18868) );
  INV_X1 U19875 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18860) );
  INV_X1 U19876 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18856) );
  INV_X1 U19877 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18852) );
  NAND2_X1 U19878 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17055) );
  NOR2_X1 U19879 ( .A1(n18852), .A2(n17055), .ZN(n17033) );
  NAND2_X1 U19880 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17033), .ZN(n17009) );
  NOR2_X1 U19881 ( .A1(n18856), .A2(n17009), .ZN(n16992) );
  NAND2_X1 U19882 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16992), .ZN(n16986) );
  NOR2_X1 U19883 ( .A1(n18860), .A2(n16986), .ZN(n16973) );
  NAND2_X1 U19884 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16973), .ZN(n16945) );
  NAND2_X1 U19885 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16948) );
  NOR3_X1 U19886 ( .A1(n18868), .A2(n16945), .A3(n16948), .ZN(n16927) );
  NAND2_X1 U19887 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16927), .ZN(n16914) );
  NOR2_X1 U19888 ( .A1(n18872), .A2(n16914), .ZN(n16730) );
  INV_X1 U19889 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18881) );
  NAND2_X1 U19890 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16868) );
  NOR2_X1 U19891 ( .A1(n18881), .A2(n16868), .ZN(n16854) );
  AND4_X1 U19892 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(n16854), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16731) );
  NAND2_X1 U19893 ( .A1(n16902), .A2(n16731), .ZN(n16828) );
  INV_X1 U19894 ( .A(n16828), .ZN(n16820) );
  NAND4_X1 U19895 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16820), .A4(P3_REIP_REG_22__SCAN_IN), .ZN(n16802) );
  NOR2_X1 U19896 ( .A1(n18894), .A2(n16802), .ZN(n16792) );
  NAND3_X1 U19897 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16792), .A3(
        P3_REIP_REG_25__SCAN_IN), .ZN(n16712) );
  NAND2_X1 U19898 ( .A1(n17087), .A2(n17076), .ZN(n17085) );
  NAND2_X1 U19899 ( .A1(n16712), .A2(n17085), .ZN(n16786) );
  OAI21_X1 U19900 ( .B1(n16713), .B2(n17076), .A(n16786), .ZN(n16751) );
  AOI211_X4 U19901 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18338), .A(n16714), .B(
        n16716), .ZN(n17028) );
  AOI22_X1 U19902 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n16751), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17028), .ZN(n16735) );
  NAND2_X1 U19903 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18338), .ZN(n16715) );
  AOI211_X4 U19904 ( .C1(n18971), .C2(n18973), .A(n16716), .B(n16715), .ZN(
        n17047) );
  NOR3_X1 U19905 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U19906 ( .A1(n17052), .A2(n17360), .ZN(n17046) );
  NOR2_X1 U19907 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17046), .ZN(n17025) );
  NAND2_X1 U19908 ( .A1(n17025), .A2(n17347), .ZN(n17014) );
  NAND2_X1 U19909 ( .A1(n17001), .A2(n16988), .ZN(n16987) );
  NAND2_X1 U19910 ( .A1(n16964), .A2(n17297), .ZN(n16947) );
  NAND2_X1 U19911 ( .A1(n16946), .A2(n16942), .ZN(n16941) );
  NAND2_X1 U19912 ( .A1(n16924), .A2(n17252), .ZN(n16916) );
  INV_X1 U19913 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21271) );
  NAND2_X1 U19914 ( .A1(n16905), .A2(n21271), .ZN(n16892) );
  NAND2_X1 U19915 ( .A1(n16878), .A2(n21127), .ZN(n16874) );
  INV_X1 U19916 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16852) );
  NAND2_X1 U19917 ( .A1(n16859), .A2(n16852), .ZN(n16850) );
  NAND2_X1 U19918 ( .A1(n16840), .A2(n17091), .ZN(n16831) );
  NAND2_X1 U19919 ( .A1(n16818), .A2(n16812), .ZN(n16810) );
  NAND2_X1 U19920 ( .A1(n16800), .A2(n16796), .ZN(n16795) );
  NAND2_X1 U19921 ( .A1(n16776), .A2(n17120), .ZN(n16772) );
  NOR2_X1 U19922 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16772), .ZN(n16760) );
  NAND2_X1 U19923 ( .A1(n16760), .A2(n14195), .ZN(n16737) );
  NOR2_X1 U19924 ( .A1(n17083), .A2(n16737), .ZN(n16743) );
  INV_X1 U19925 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17096) );
  NOR2_X1 U19926 ( .A1(n17989), .A2(n17635), .ZN(n16720) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16720), .A(
        n16717), .ZN(n17646) );
  INV_X1 U19928 ( .A(n17646), .ZN(n16759) );
  INV_X1 U19929 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17705) );
  INV_X1 U19930 ( .A(n16718), .ZN(n17748) );
  INV_X1 U19931 ( .A(n17747), .ZN(n16719) );
  NAND2_X1 U19932 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16847), .ZN(
        n16728) );
  NAND2_X1 U19933 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16727), .ZN(
        n17671) );
  NOR2_X1 U19934 ( .A1(n17705), .A2(n17671), .ZN(n16725) );
  NAND3_X1 U19935 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n16725), .ZN(n17632) );
  INV_X1 U19936 ( .A(n17632), .ZN(n16722) );
  NAND2_X1 U19937 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16722), .ZN(
        n16721) );
  AOI21_X1 U19938 ( .B1(n10092), .B2(n16721), .A(n16720), .ZN(n17654) );
  OAI21_X1 U19939 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16722), .A(
        n16721), .ZN(n17662) );
  INV_X1 U19940 ( .A(n17662), .ZN(n16779) );
  INV_X1 U19941 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17688) );
  INV_X1 U19942 ( .A(n16725), .ZN(n16724) );
  NOR2_X1 U19943 ( .A1(n17688), .A2(n16724), .ZN(n16723) );
  OAI21_X1 U19944 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16723), .A(
        n17632), .ZN(n17674) );
  INV_X1 U19945 ( .A(n17674), .ZN(n16790) );
  AOI21_X1 U19946 ( .B1(n17688), .B2(n16724), .A(n16723), .ZN(n17685) );
  AOI21_X1 U19947 ( .B1(n17705), .B2(n17671), .A(n16725), .ZN(n17701) );
  OAI21_X1 U19948 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16727), .A(
        n17671), .ZN(n16726) );
  INV_X1 U19949 ( .A(n16726), .ZN(n17718) );
  AOI21_X1 U19950 ( .B1(n10094), .B2(n16728), .A(n16727), .ZN(n17730) );
  OAI21_X1 U19951 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n16847), .A(
        n16728), .ZN(n17736) );
  INV_X1 U19952 ( .A(n17736), .ZN(n16839) );
  NOR3_X1 U19953 ( .A1(n17989), .A2(n17813), .A3(n17812), .ZN(n17784) );
  NAND2_X1 U19954 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17784), .ZN(
        n16890) );
  NOR2_X1 U19955 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16890), .ZN(
        n16901) );
  AOI21_X1 U19956 ( .B1(n16847), .B2(n16901), .A(n16974), .ZN(n16838) );
  NOR2_X1 U19957 ( .A1(n16837), .A2(n16974), .ZN(n16830) );
  NOR2_X1 U19958 ( .A1(n17730), .A2(n16830), .ZN(n16829) );
  NOR2_X1 U19959 ( .A1(n16829), .A2(n16974), .ZN(n16822) );
  NOR2_X1 U19960 ( .A1(n16821), .A2(n16974), .ZN(n16809) );
  NOR2_X1 U19961 ( .A1(n16790), .A2(n16789), .ZN(n16788) );
  NOR2_X1 U19962 ( .A1(n16788), .A2(n16974), .ZN(n16778) );
  NOR2_X1 U19963 ( .A1(n16777), .A2(n16974), .ZN(n16769) );
  NOR2_X1 U19964 ( .A1(n16768), .A2(n16729), .ZN(n16758) );
  NOR2_X1 U19965 ( .A1(n16759), .A2(n16758), .ZN(n16757) );
  NOR2_X1 U19966 ( .A1(n16757), .A2(n16729), .ZN(n16746) );
  NAND2_X1 U19967 ( .A1(n10080), .A2(n17066), .ZN(n16999) );
  NOR3_X1 U19968 ( .A1(n16739), .A2(n16738), .A3(n16999), .ZN(n16733) );
  INV_X1 U19969 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18907) );
  INV_X1 U19970 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18898) );
  INV_X1 U19971 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18889) );
  INV_X1 U19972 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18875) );
  NAND2_X1 U19973 ( .A1(n17054), .A2(n16730), .ZN(n16904) );
  NAND2_X1 U19974 ( .A1(n16731), .A2(n16897), .ZN(n16836) );
  NAND3_X1 U19975 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(n16825), .ZN(n16804) );
  NOR2_X1 U19976 ( .A1(n18894), .A2(n16804), .ZN(n16787) );
  NAND2_X1 U19977 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16787), .ZN(n16785) );
  NAND4_X1 U19978 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16756), .ZN(n16741) );
  AOI221_X1 U19979 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n21196), .C2(n18907), .A(n16741), .ZN(n16732) );
  AOI211_X1 U19980 ( .C1(n16743), .C2(n17096), .A(n16733), .B(n16732), .ZN(
        n16734) );
  OAI211_X1 U19981 ( .C1(n16736), .C2(n17059), .A(n16735), .B(n16734), .ZN(
        P3_U2640) );
  NAND2_X1 U19982 ( .A1(n17047), .A2(n16737), .ZN(n16754) );
  OAI22_X1 U19983 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16741), .B1(n16740), 
        .B2(n17059), .ZN(n16742) );
  OAI21_X1 U19984 ( .B1(n17028), .B2(n16743), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16744) );
  NOR2_X1 U19985 ( .A1(n16760), .A2(n14195), .ZN(n16755) );
  AOI211_X1 U19986 ( .C1(n16747), .C2(n16746), .A(n16745), .B(n18825), .ZN(
        n16750) );
  OAI22_X1 U19987 ( .A1(n16748), .A2(n17059), .B1(n17084), .B2(n14195), .ZN(
        n16749) );
  AOI211_X1 U19988 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16751), .A(n16750), 
        .B(n16749), .ZN(n16753) );
  NAND4_X1 U19989 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16756), .A4(n18903), .ZN(n16752) );
  OAI211_X1 U19990 ( .C1(n16755), .C2(n16754), .A(n16753), .B(n16752), .ZN(
        P3_U2642) );
  NAND2_X1 U19991 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16756), .ZN(n16767) );
  NAND2_X1 U19992 ( .A1(n16756), .A2(n21163), .ZN(n16774) );
  AOI21_X1 U19993 ( .B1(n16786), .B2(n16774), .A(n18901), .ZN(n16765) );
  AOI211_X1 U19994 ( .C1(n16759), .C2(n16758), .A(n16757), .B(n18825), .ZN(
        n16764) );
  AOI211_X1 U19995 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16772), .A(n16760), .B(
        n17083), .ZN(n16763) );
  OAI22_X1 U19996 ( .A1(n17634), .A2(n17059), .B1(n17084), .B2(n16761), .ZN(
        n16762) );
  NOR4_X1 U19997 ( .A1(n16765), .A2(n16764), .A3(n16763), .A4(n16762), .ZN(
        n16766) );
  OAI21_X1 U19998 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n16767), .A(n16766), 
        .ZN(P3_U2643) );
  AOI211_X1 U19999 ( .C1(n17654), .C2(n16769), .A(n16768), .B(n18825), .ZN(
        n16771) );
  OAI22_X1 U20000 ( .A1(n10092), .A2(n17059), .B1(n21163), .B2(n16786), .ZN(
        n16770) );
  AOI211_X1 U20001 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17028), .A(n16771), .B(
        n16770), .ZN(n16775) );
  OAI211_X1 U20002 ( .C1(n16776), .C2(n17120), .A(n17047), .B(n16772), .ZN(
        n16773) );
  NAND3_X1 U20003 ( .A1(n16775), .A2(n16774), .A3(n16773), .ZN(P3_U2644) );
  AOI211_X1 U20004 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16795), .A(n16776), .B(
        n17083), .ZN(n16783) );
  AOI211_X1 U20005 ( .C1(n16779), .C2(n16778), .A(n16777), .B(n18825), .ZN(
        n16782) );
  INV_X1 U20006 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16780) );
  OAI22_X1 U20007 ( .A1(n17660), .A2(n17059), .B1(n17084), .B2(n16780), .ZN(
        n16781) );
  NOR3_X1 U20008 ( .A1(n16783), .A2(n16782), .A3(n16781), .ZN(n16784) );
  OAI221_X1 U20009 ( .B1(n16786), .B2(n18898), .C1(n16786), .C2(n16785), .A(
        n16784), .ZN(P3_U2645) );
  INV_X1 U20010 ( .A(n16787), .ZN(n16799) );
  AOI211_X1 U20011 ( .C1(n16790), .C2(n16789), .A(n16788), .B(n18825), .ZN(
        n16794) );
  NAND2_X1 U20012 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17085), .ZN(n16791) );
  INV_X1 U20013 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17672) );
  OAI22_X1 U20014 ( .A1(n16792), .A2(n16791), .B1(n17672), .B2(n17059), .ZN(
        n16793) );
  AOI211_X1 U20015 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n17028), .A(n16794), .B(
        n16793), .ZN(n16798) );
  OAI211_X1 U20016 ( .C1(n16800), .C2(n16796), .A(n17047), .B(n16795), .ZN(
        n16797) );
  OAI211_X1 U20017 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16799), .A(n16798), 
        .B(n16797), .ZN(P3_U2646) );
  AOI211_X1 U20018 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16810), .A(n16800), .B(
        n17083), .ZN(n16807) );
  AOI211_X1 U20019 ( .C1(n17685), .C2(n9944), .A(n16801), .B(n18825), .ZN(
        n16806) );
  NAND2_X1 U20020 ( .A1(n17085), .A2(n16802), .ZN(n16816) );
  AOI22_X1 U20021 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17071), .B1(
        n17028), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16803) );
  OAI221_X1 U20022 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16804), .C1(n18894), 
        .C2(n16816), .A(n16803), .ZN(n16805) );
  OR3_X1 U20023 ( .A1(n16807), .A2(n16806), .A3(n16805), .ZN(P3_U2647) );
  NAND2_X1 U20024 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16825), .ZN(n16817) );
  INV_X1 U20025 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18893) );
  AOI211_X1 U20026 ( .C1(n17701), .C2(n16809), .A(n16808), .B(n18825), .ZN(
        n16814) );
  OAI211_X1 U20027 ( .C1(n16818), .C2(n16812), .A(n17047), .B(n16810), .ZN(
        n16811) );
  OAI21_X1 U20028 ( .B1(n16812), .B2(n17084), .A(n16811), .ZN(n16813) );
  AOI211_X1 U20029 ( .C1(n17071), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16814), .B(n16813), .ZN(n16815) );
  OAI221_X1 U20030 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n16817), .C1(n18893), 
        .C2(n16816), .A(n16815), .ZN(P3_U2648) );
  AOI211_X1 U20031 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16831), .A(n16818), .B(
        n17083), .ZN(n16819) );
  AOI21_X1 U20032 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17028), .A(n16819), .ZN(
        n16827) );
  INV_X1 U20033 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18890) );
  INV_X1 U20034 ( .A(n17085), .ZN(n16903) );
  OAI22_X1 U20035 ( .A1(n16903), .A2(n16820), .B1(P3_REIP_REG_21__SCAN_IN), 
        .B2(n16836), .ZN(n16824) );
  AOI211_X1 U20036 ( .C1(n17718), .C2(n16822), .A(n16821), .B(n18825), .ZN(
        n16823) );
  AOI221_X1 U20037 ( .B1(n16825), .B2(n18890), .C1(n16824), .C2(
        P3_REIP_REG_22__SCAN_IN), .A(n16823), .ZN(n16826) );
  OAI211_X1 U20038 ( .C1(n10095), .C2(n17059), .A(n16827), .B(n16826), .ZN(
        P3_U2649) );
  NAND2_X1 U20039 ( .A1(n17085), .A2(n16828), .ZN(n16845) );
  AOI211_X1 U20040 ( .C1(n17730), .C2(n16830), .A(n16829), .B(n18825), .ZN(
        n16834) );
  OAI211_X1 U20041 ( .C1(n16840), .C2(n17091), .A(n17047), .B(n16831), .ZN(
        n16832) );
  OAI21_X1 U20042 ( .B1(n17091), .B2(n17084), .A(n16832), .ZN(n16833) );
  AOI211_X1 U20043 ( .C1(n17071), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16834), .B(n16833), .ZN(n16835) );
  OAI221_X1 U20044 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16836), .C1(n18889), 
        .C2(n16845), .A(n16835), .ZN(P3_U2650) );
  INV_X1 U20045 ( .A(n16897), .ZN(n16884) );
  NOR3_X1 U20046 ( .A1(n18881), .A2(n16868), .A3(n16884), .ZN(n16865) );
  NAND3_X1 U20047 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16865), .ZN(n16846) );
  INV_X1 U20048 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18886) );
  AOI211_X1 U20049 ( .C1(n16839), .C2(n16838), .A(n16837), .B(n18825), .ZN(
        n16843) );
  AOI211_X1 U20050 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16850), .A(n16840), .B(
        n17083), .ZN(n16842) );
  OAI22_X1 U20051 ( .A1(n21100), .A2(n17059), .B1(n17084), .B2(n10193), .ZN(
        n16841) );
  NOR3_X1 U20052 ( .A1(n16843), .A2(n16842), .A3(n16841), .ZN(n16844) );
  OAI221_X1 U20053 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16846), .C1(n18886), 
        .C2(n16845), .A(n16844), .ZN(P3_U2651) );
  NAND2_X1 U20054 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17747), .ZN(
        n16861) );
  INV_X1 U20055 ( .A(n16861), .ZN(n16848) );
  INV_X1 U20056 ( .A(n16847), .ZN(n17716) );
  OAI21_X1 U20057 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16848), .A(
        n17716), .ZN(n17752) );
  OAI21_X1 U20058 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16861), .A(
        n10080), .ZN(n16849) );
  XNOR2_X1 U20059 ( .A(n17752), .B(n16849), .ZN(n16858) );
  OAI211_X1 U20060 ( .C1(n16859), .C2(n16852), .A(n17047), .B(n16850), .ZN(
        n16851) );
  OAI211_X1 U20061 ( .C1(n17084), .C2(n16852), .A(n18317), .B(n16851), .ZN(
        n16853) );
  AOI21_X1 U20062 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17071), .A(
        n16853), .ZN(n16857) );
  AOI21_X1 U20063 ( .B1(n16902), .B2(n16854), .A(n16903), .ZN(n16873) );
  INV_X1 U20064 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18882) );
  XNOR2_X1 U20065 ( .A(P3_REIP_REG_19__SCAN_IN), .B(n18882), .ZN(n16855) );
  AOI22_X1 U20066 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16873), .B1(n16865), 
        .B2(n16855), .ZN(n16856) );
  OAI211_X1 U20067 ( .C1(n18825), .C2(n16858), .A(n16857), .B(n16856), .ZN(
        P3_U2652) );
  INV_X1 U20068 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17761) );
  AOI211_X1 U20069 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16874), .A(n16859), .B(
        n17083), .ZN(n16860) );
  AOI211_X1 U20070 ( .C1(n17028), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9816), .B(
        n16860), .ZN(n16867) );
  OAI21_X1 U20071 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17747), .A(
        n16861), .ZN(n17758) );
  INV_X1 U20072 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21228) );
  NAND2_X1 U20073 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21228), .ZN(
        n17064) );
  OAI21_X1 U20074 ( .B1(n17748), .B2(n17064), .A(n10080), .ZN(n16863) );
  OAI21_X1 U20075 ( .B1(n17758), .B2(n16863), .A(n17066), .ZN(n16862) );
  AOI21_X1 U20076 ( .B1(n17758), .B2(n16863), .A(n16862), .ZN(n16864) );
  AOI221_X1 U20077 ( .B1(n16873), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16865), 
        .C2(n18882), .A(n16864), .ZN(n16866) );
  OAI211_X1 U20078 ( .C1(n17761), .C2(n17059), .A(n16867), .B(n16866), .ZN(
        P3_U2653) );
  AOI22_X1 U20079 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17071), .B1(
        n17028), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16877) );
  NOR2_X1 U20080 ( .A1(n16868), .A2(n16884), .ZN(n16872) );
  INV_X1 U20081 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17798) );
  INV_X1 U20082 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16889) );
  NOR2_X1 U20083 ( .A1(n17798), .A2(n16889), .ZN(n17788) );
  NAND2_X1 U20084 ( .A1(n17788), .A2(n17784), .ZN(n16880) );
  AOI21_X1 U20085 ( .B1(n17773), .B2(n16880), .A(n17747), .ZN(n17775) );
  AOI21_X1 U20086 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16901), .A(
        n16729), .ZN(n16870) );
  OAI21_X1 U20087 ( .B1(n17775), .B2(n16870), .A(n17066), .ZN(n16869) );
  AOI21_X1 U20088 ( .B1(n17775), .B2(n16870), .A(n16869), .ZN(n16871) );
  AOI221_X1 U20089 ( .B1(n16873), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16872), 
        .C2(n18881), .A(n16871), .ZN(n16876) );
  OAI211_X1 U20090 ( .C1(n16878), .C2(n21127), .A(n17047), .B(n16874), .ZN(
        n16875) );
  NAND4_X1 U20091 ( .A1(n16877), .A2(n16876), .A3(n18317), .A4(n16875), .ZN(
        P3_U2654) );
  AOI211_X1 U20092 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16892), .A(n16878), .B(
        n17083), .ZN(n16879) );
  AOI211_X1 U20093 ( .C1(n17028), .C2(P3_EBX_REG_16__SCAN_IN), .A(n9816), .B(
        n16879), .ZN(n16888) );
  AOI21_X1 U20094 ( .B1(n16902), .B2(P3_REIP_REG_15__SCAN_IN), .A(n16903), 
        .ZN(n16896) );
  INV_X1 U20095 ( .A(n16880), .ZN(n16881) );
  AOI21_X1 U20096 ( .B1(n16889), .B2(n16890), .A(n16881), .ZN(n17785) );
  NOR2_X1 U20097 ( .A1(n16901), .A2(n16974), .ZN(n16883) );
  OAI21_X1 U20098 ( .B1(n17785), .B2(n16883), .A(n17066), .ZN(n16882) );
  AOI21_X1 U20099 ( .B1(n17785), .B2(n16883), .A(n16882), .ZN(n16886) );
  INV_X1 U20100 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18876) );
  NOR3_X1 U20101 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18876), .A3(n16884), 
        .ZN(n16885) );
  AOI211_X1 U20102 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16896), .A(n16886), 
        .B(n16885), .ZN(n16887) );
  OAI211_X1 U20103 ( .C1(n16889), .C2(n17059), .A(n16888), .B(n16887), .ZN(
        P3_U2655) );
  INV_X1 U20104 ( .A(n16999), .ZN(n17072) );
  OAI21_X1 U20105 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17784), .A(
        n16890), .ZN(n17795) );
  NAND2_X1 U20106 ( .A1(n17072), .A2(n17795), .ZN(n16900) );
  INV_X1 U20107 ( .A(n17784), .ZN(n16891) );
  OAI21_X1 U20108 ( .B1(n16974), .B2(n21228), .A(n17066), .ZN(n17082) );
  AOI211_X1 U20109 ( .C1(n10080), .C2(n16891), .A(n17795), .B(n17082), .ZN(
        n16895) );
  OAI211_X1 U20110 ( .C1(n16905), .C2(n21271), .A(n17047), .B(n16892), .ZN(
        n16893) );
  OAI211_X1 U20111 ( .C1(n17084), .C2(n21271), .A(n18317), .B(n16893), .ZN(
        n16894) );
  AOI211_X1 U20112 ( .C1(n17071), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16895), .B(n16894), .ZN(n16899) );
  OAI21_X1 U20113 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16897), .A(n16896), 
        .ZN(n16898) );
  OAI211_X1 U20114 ( .C1(n16901), .C2(n16900), .A(n16899), .B(n16898), .ZN(
        P3_U2656) );
  OR2_X1 U20115 ( .A1(n17989), .A2(n17813), .ZN(n16913) );
  AOI21_X1 U20116 ( .B1(n17812), .B2(n16913), .A(n17784), .ZN(n17815) );
  NAND2_X1 U20117 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17830) );
  INV_X1 U20118 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17869) );
  NOR2_X1 U20119 ( .A1(n17989), .A2(n17894), .ZN(n16960) );
  NAND3_X1 U20120 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16960), .ZN(n16962) );
  NOR2_X1 U20121 ( .A1(n17869), .A2(n16962), .ZN(n16953) );
  NAND2_X1 U20122 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16953), .ZN(
        n17826) );
  NOR3_X1 U20123 ( .A1(n17830), .A2(n17826), .A3(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16910) );
  OR2_X1 U20124 ( .A1(n16999), .A2(n16910), .ZN(n16922) );
  AOI211_X1 U20125 ( .C1(n18875), .C2(n16904), .A(n16903), .B(n16902), .ZN(
        n16909) );
  AOI211_X1 U20126 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16916), .A(n16905), .B(
        n17083), .ZN(n16908) );
  OAI22_X1 U20127 ( .A1(n17812), .A2(n17059), .B1(n17084), .B2(n16906), .ZN(
        n16907) );
  NOR4_X1 U20128 ( .A1(n9816), .A2(n16909), .A3(n16908), .A4(n16907), .ZN(
        n16912) );
  OAI211_X1 U20129 ( .C1(n16910), .C2(n16729), .A(n17066), .B(n17815), .ZN(
        n16911) );
  OAI211_X1 U20130 ( .C1(n17815), .C2(n16922), .A(n16912), .B(n16911), .ZN(
        P3_U2657) );
  INV_X1 U20131 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16929) );
  NOR2_X1 U20132 ( .A1(n16929), .A2(n17826), .ZN(n16928) );
  OAI21_X1 U20133 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16928), .A(
        n16913), .ZN(n17832) );
  INV_X1 U20134 ( .A(n17832), .ZN(n16923) );
  INV_X1 U20135 ( .A(n17082), .ZN(n16998) );
  OAI21_X1 U20136 ( .B1(n16928), .B2(n16974), .A(n16998), .ZN(n16921) );
  OAI21_X1 U20137 ( .B1(n16927), .B2(n17076), .A(n17087), .ZN(n16936) );
  NOR2_X1 U20138 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17076), .ZN(n16926) );
  NOR3_X1 U20139 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17076), .A3(n16914), 
        .ZN(n16915) );
  AOI211_X1 U20140 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17071), .A(
        n9816), .B(n16915), .ZN(n16918) );
  OAI211_X1 U20141 ( .C1(n16924), .C2(n17252), .A(n17047), .B(n16916), .ZN(
        n16917) );
  OAI211_X1 U20142 ( .C1(n17252), .C2(n17084), .A(n16918), .B(n16917), .ZN(
        n16919) );
  AOI221_X1 U20143 ( .B1(n16936), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16926), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16919), .ZN(n16920) );
  OAI221_X1 U20144 ( .B1(n16923), .B2(n16922), .C1(n17832), .C2(n16921), .A(
        n16920), .ZN(P3_U2658) );
  AOI211_X1 U20145 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16941), .A(n16924), .B(
        n17083), .ZN(n16925) );
  AOI21_X1 U20146 ( .B1(n17071), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16925), .ZN(n16934) );
  AOI22_X1 U20147 ( .A1(n17028), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16927), 
        .B2(n16926), .ZN(n16933) );
  AOI21_X1 U20148 ( .B1(n16929), .B2(n17826), .A(n16928), .ZN(n17845) );
  OAI21_X1 U20149 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17826), .A(
        n10080), .ZN(n16930) );
  XNOR2_X1 U20150 ( .A(n17845), .B(n16930), .ZN(n16931) );
  AOI22_X1 U20151 ( .A1(n17066), .A2(n16931), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16936), .ZN(n16932) );
  NAND4_X1 U20152 ( .A1(n16934), .A2(n16933), .A3(n16932), .A4(n18317), .ZN(
        P3_U2659) );
  INV_X1 U20153 ( .A(n16948), .ZN(n16935) );
  NOR2_X1 U20154 ( .A1(n17076), .A2(n16945), .ZN(n16959) );
  AOI21_X1 U20155 ( .B1(n16935), .B2(n16959), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16939) );
  INV_X1 U20156 ( .A(n16936), .ZN(n16938) );
  AOI21_X1 U20157 ( .B1(n16953), .B2(n21228), .A(n16729), .ZN(n16956) );
  OAI21_X1 U20158 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16953), .A(
        n17826), .ZN(n17857) );
  XOR2_X1 U20159 ( .A(n16956), .B(n17857), .Z(n16937) );
  OAI22_X1 U20160 ( .A1(n16939), .A2(n16938), .B1(n18825), .B2(n16937), .ZN(
        n16940) );
  AOI211_X1 U20161 ( .C1(n17028), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9816), .B(
        n16940), .ZN(n16944) );
  OAI211_X1 U20162 ( .C1(n16946), .C2(n16942), .A(n17047), .B(n16941), .ZN(
        n16943) );
  OAI211_X1 U20163 ( .C1(n17059), .C2(n17859), .A(n16944), .B(n16943), .ZN(
        P3_U2660) );
  INV_X1 U20164 ( .A(n17087), .ZN(n17079) );
  AOI21_X1 U20165 ( .B1(n17054), .B2(n16945), .A(n17079), .ZN(n16979) );
  INV_X1 U20166 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18866) );
  AOI211_X1 U20167 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16947), .A(n16946), .B(
        n17083), .ZN(n16952) );
  OAI211_X1 U20168 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16959), .B(n16948), .ZN(n16949) );
  OAI211_X1 U20169 ( .C1(n17084), .C2(n16950), .A(n18317), .B(n16949), .ZN(
        n16951) );
  AOI211_X1 U20170 ( .C1(n17071), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16952), .B(n16951), .ZN(n16958) );
  AOI21_X1 U20171 ( .B1(n17869), .B2(n16962), .A(n16953), .ZN(n17872) );
  NAND2_X1 U20172 ( .A1(n17066), .A2(n16729), .ZN(n17070) );
  INV_X1 U20173 ( .A(n17070), .ZN(n16955) );
  AOI221_X1 U20174 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17872), .C1(
        n16962), .C2(n17872), .A(n18825), .ZN(n16954) );
  OAI22_X1 U20175 ( .A1(n17872), .A2(n16956), .B1(n16955), .B2(n16954), .ZN(
        n16957) );
  OAI211_X1 U20176 ( .C1(n16979), .C2(n18866), .A(n16958), .B(n16957), .ZN(
        P3_U2661) );
  INV_X1 U20177 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18864) );
  NOR2_X1 U20178 ( .A1(n16964), .A2(n17083), .ZN(n16971) );
  AOI22_X1 U20179 ( .A1(n16959), .A2(n18864), .B1(n16971), .B2(n17297), .ZN(
        n16970) );
  INV_X1 U20180 ( .A(n16960), .ZN(n16997) );
  NOR2_X1 U20181 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16997), .ZN(
        n17000) );
  AOI21_X1 U20182 ( .B1(n17892), .B2(n17000), .A(n16974), .ZN(n16963) );
  INV_X1 U20183 ( .A(n17892), .ZN(n16961) );
  NOR2_X1 U20184 ( .A1(n16961), .A2(n16997), .ZN(n16975) );
  OAI21_X1 U20185 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16975), .A(
        n16962), .ZN(n17883) );
  XNOR2_X1 U20186 ( .A(n16963), .B(n17883), .ZN(n16968) );
  INV_X1 U20187 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16966) );
  AOI21_X1 U20188 ( .B1(n17047), .B2(n16964), .A(n17028), .ZN(n16965) );
  OAI22_X1 U20189 ( .A1(n16966), .A2(n17059), .B1(n17297), .B2(n16965), .ZN(
        n16967) );
  AOI211_X1 U20190 ( .C1(n17066), .C2(n16968), .A(n9816), .B(n16967), .ZN(
        n16969) );
  OAI211_X1 U20191 ( .C1(n18864), .C2(n16979), .A(n16970), .B(n16969), .ZN(
        P3_U2662) );
  INV_X1 U20192 ( .A(n16971), .ZN(n16972) );
  AOI21_X1 U20193 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16987), .A(n16972), .ZN(
        n16982) );
  AOI21_X1 U20194 ( .B1(n17054), .B2(n16973), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16980) );
  NOR3_X1 U20195 ( .A1(n17989), .A2(n17894), .A3(n17912), .ZN(n16984) );
  AOI21_X1 U20196 ( .B1(n16984), .B2(n21228), .A(n16974), .ZN(n16977) );
  INV_X1 U20197 ( .A(n16975), .ZN(n16976) );
  OAI21_X1 U20198 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16984), .A(
        n16976), .ZN(n17896) );
  XOR2_X1 U20199 ( .A(n16977), .B(n17896), .Z(n16978) );
  OAI22_X1 U20200 ( .A1(n16980), .A2(n16979), .B1(n18825), .B2(n16978), .ZN(
        n16981) );
  AOI211_X1 U20201 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17028), .A(n16982), .B(
        n16981), .ZN(n16983) );
  OAI211_X1 U20202 ( .C1(n17895), .C2(n17059), .A(n16983), .B(n18317), .ZN(
        P3_U2663) );
  AOI21_X1 U20203 ( .B1(n17912), .B2(n16997), .A(n16984), .ZN(n17916) );
  NOR2_X1 U20204 ( .A1(n17000), .A2(n16729), .ZN(n16985) );
  XNOR2_X1 U20205 ( .A(n17916), .B(n16985), .ZN(n16995) );
  NOR3_X1 U20206 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17076), .A3(n16986), .ZN(
        n16991) );
  OAI211_X1 U20207 ( .C1(n17001), .C2(n16988), .A(n17047), .B(n16987), .ZN(
        n16989) );
  OAI211_X1 U20208 ( .C1(n17912), .C2(n17059), .A(n18317), .B(n16989), .ZN(
        n16990) );
  AOI211_X1 U20209 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17028), .A(n16991), .B(
        n16990), .ZN(n16994) );
  INV_X1 U20210 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18858) );
  AND3_X1 U20211 ( .A1(n18858), .A2(n17054), .A3(n16992), .ZN(n17002) );
  OAI21_X1 U20212 ( .B1(n16992), .B2(n17076), .A(n17087), .ZN(n17019) );
  OAI21_X1 U20213 ( .B1(n17002), .B2(n17019), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n16993) );
  OAI211_X1 U20214 ( .C1(n16995), .C2(n18825), .A(n16994), .B(n16993), .ZN(
        P3_U2664) );
  INV_X1 U20215 ( .A(n17920), .ZN(n16996) );
  NOR2_X1 U20216 ( .A1(n17989), .A2(n16996), .ZN(n17011) );
  OAI21_X1 U20217 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17011), .A(
        n16997), .ZN(n17931) );
  INV_X1 U20218 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17921) );
  OAI21_X1 U20219 ( .B1(n17921), .B2(n16729), .A(n16998), .ZN(n17008) );
  NOR2_X1 U20220 ( .A1(n17000), .A2(n16999), .ZN(n17004) );
  AOI211_X1 U20221 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17014), .A(n17001), .B(
        n17083), .ZN(n17003) );
  AOI211_X1 U20222 ( .C1(n17004), .C2(n17931), .A(n17003), .B(n17002), .ZN(
        n17007) );
  OAI22_X1 U20223 ( .A1(n17921), .A2(n17059), .B1(n17084), .B2(n17337), .ZN(
        n17005) );
  AOI211_X1 U20224 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n17019), .A(n9816), .B(
        n17005), .ZN(n17006) );
  OAI211_X1 U20225 ( .C1(n17931), .C2(n17008), .A(n17007), .B(n17006), .ZN(
        P3_U2665) );
  OAI21_X1 U20226 ( .B1(n17076), .B2(n17009), .A(n18856), .ZN(n17018) );
  INV_X1 U20227 ( .A(n17939), .ZN(n17010) );
  NAND2_X1 U20228 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17010), .ZN(
        n17024) );
  AOI21_X1 U20229 ( .B1(n17940), .B2(n17024), .A(n17011), .ZN(n17941) );
  OAI21_X1 U20230 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17024), .A(
        n10080), .ZN(n17031) );
  INV_X1 U20231 ( .A(n17031), .ZN(n17013) );
  INV_X1 U20232 ( .A(n17941), .ZN(n17012) );
  OAI221_X1 U20233 ( .B1(n17941), .B2(n17013), .C1(n17012), .C2(n17031), .A(
        n17066), .ZN(n17016) );
  OAI211_X1 U20234 ( .C1(n17025), .C2(n17347), .A(n17047), .B(n17014), .ZN(
        n17015) );
  OAI211_X1 U20235 ( .C1(n17059), .C2(n17940), .A(n17016), .B(n17015), .ZN(
        n17017) );
  AOI21_X1 U20236 ( .B1(n17019), .B2(n17018), .A(n17017), .ZN(n17020) );
  OAI211_X1 U20237 ( .C1(n17084), .C2(n17347), .A(n17020), .B(n18317), .ZN(
        P3_U2666) );
  NAND2_X1 U20238 ( .A1(n18335), .A2(n17021), .ZN(n18987) );
  AOI21_X1 U20239 ( .B1(n17022), .B2(n18767), .A(n18987), .ZN(n17023) );
  AOI211_X1 U20240 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n17071), .A(
        n9816), .B(n17023), .ZN(n17037) );
  INV_X1 U20241 ( .A(n17030), .ZN(n17947) );
  NOR2_X1 U20242 ( .A1(n17989), .A2(n17947), .ZN(n17038) );
  OAI21_X1 U20243 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17038), .A(
        n17024), .ZN(n17029) );
  NOR2_X1 U20244 ( .A1(n17029), .A2(n17070), .ZN(n17027) );
  AOI211_X1 U20245 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17046), .A(n17025), .B(
        n17083), .ZN(n17026) );
  AOI211_X1 U20246 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17028), .A(n17027), .B(
        n17026), .ZN(n17036) );
  INV_X1 U20247 ( .A(n17029), .ZN(n17955) );
  INV_X1 U20248 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17958) );
  NAND2_X1 U20249 ( .A1(n17030), .A2(n17958), .ZN(n17951) );
  OAI22_X1 U20250 ( .A1(n17955), .A2(n17031), .B1(n17064), .B2(n17951), .ZN(
        n17032) );
  OAI21_X1 U20251 ( .B1(n17033), .B2(n17076), .A(n17087), .ZN(n17045) );
  AOI22_X1 U20252 ( .A1(n17066), .A2(n17032), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n17045), .ZN(n17035) );
  INV_X1 U20253 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18854) );
  NAND3_X1 U20254 ( .A1(n17054), .A2(n17033), .A3(n18854), .ZN(n17034) );
  NAND4_X1 U20255 ( .A1(n17037), .A2(n17036), .A3(n17035), .A4(n17034), .ZN(
        P3_U2667) );
  OAI21_X1 U20256 ( .B1(n17076), .B2(n17055), .A(n18852), .ZN(n17044) );
  NAND2_X1 U20257 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17051) );
  AOI21_X1 U20258 ( .B1(n17050), .B2(n17051), .A(n17038), .ZN(n17963) );
  OAI21_X1 U20259 ( .B1(n17051), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n10080), .ZN(n17039) );
  INV_X1 U20260 ( .A(n17039), .ZN(n17065) );
  OAI21_X1 U20261 ( .B1(n17963), .B2(n17065), .A(n17066), .ZN(n17040) );
  AOI21_X1 U20262 ( .B1(n17963), .B2(n17065), .A(n17040), .ZN(n17043) );
  NAND2_X1 U20263 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18769) );
  INV_X1 U20264 ( .A(n18769), .ZN(n18781) );
  NAND2_X1 U20265 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18781), .ZN(
        n17041) );
  AOI21_X1 U20266 ( .B1(n17041), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n9813), .ZN(n18921) );
  OAI22_X1 U20267 ( .A1(n18921), .A2(n18987), .B1(n17084), .B2(n17360), .ZN(
        n17042) );
  AOI211_X1 U20268 ( .C1(n17045), .C2(n17044), .A(n17043), .B(n17042), .ZN(
        n17049) );
  OAI211_X1 U20269 ( .C1(n17052), .C2(n17360), .A(n17047), .B(n17046), .ZN(
        n17048) );
  OAI211_X1 U20270 ( .C1(n17059), .C2(n17050), .A(n17049), .B(n17048), .ZN(
        P3_U2668) );
  OAI21_X1 U20271 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17051), .ZN(n17976) );
  OR2_X1 U20272 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n17053) );
  AOI211_X1 U20273 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17053), .A(n17052), .B(
        n17083), .ZN(n17063) );
  OAI211_X1 U20274 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17055), .B(n17054), .ZN(n17056) );
  INV_X1 U20275 ( .A(n17056), .ZN(n17062) );
  INV_X1 U20276 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17057) );
  INV_X1 U20277 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18850) );
  OAI22_X1 U20278 ( .A1(n17084), .A2(n17057), .B1(n17087), .B2(n18850), .ZN(
        n17061) );
  INV_X1 U20279 ( .A(n17075), .ZN(n18780) );
  NOR2_X1 U20280 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18780), .ZN(
        n18776) );
  AOI21_X1 U20281 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18781), .A(
        n18776), .ZN(n17058) );
  INV_X1 U20282 ( .A(n17058), .ZN(n18929) );
  OAI22_X1 U20283 ( .A1(n17980), .A2(n17059), .B1(n18929), .B2(n18987), .ZN(
        n17060) );
  NOR4_X1 U20284 ( .A1(n17063), .A2(n17062), .A3(n17061), .A4(n17060), .ZN(
        n17069) );
  INV_X1 U20285 ( .A(n17064), .ZN(n17067) );
  OAI211_X1 U20286 ( .C1(n17067), .C2(n17976), .A(n17066), .B(n17065), .ZN(
        n17068) );
  OAI211_X1 U20287 ( .C1(n17976), .C2(n17070), .A(n17069), .B(n17068), .ZN(
        P3_U2669) );
  AOI21_X1 U20288 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17072), .A(
        n17071), .ZN(n17081) );
  INV_X1 U20289 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17368) );
  OAI21_X1 U20290 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17073), .ZN(n17369) );
  OAI22_X1 U20291 ( .A1(n17084), .A2(n17368), .B1(n17083), .B2(n17369), .ZN(
        n17078) );
  NAND2_X1 U20292 ( .A1(n17075), .A2(n17074), .ZN(n18934) );
  OAI22_X1 U20293 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17076), .B1(n18934), 
        .B2(n18987), .ZN(n17077) );
  AOI211_X1 U20294 ( .C1(n17079), .C2(P3_REIP_REG_1__SCAN_IN), .A(n17078), .B(
        n17077), .ZN(n17080) );
  OAI221_X1 U20295 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17082), .C1(
        n17989), .C2(n17081), .A(n17080), .ZN(P3_U2670) );
  NAND2_X1 U20296 ( .A1(n17084), .A2(n17083), .ZN(n17086) );
  AOI22_X1 U20297 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17086), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17085), .ZN(n17089) );
  NAND3_X1 U20298 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18983), .A3(
        n17087), .ZN(n17088) );
  OAI211_X1 U20299 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18987), .A(
        n17089), .B(n17088), .ZN(P3_U2671) );
  NOR2_X1 U20300 ( .A1(n10193), .A2(n17185), .ZN(n17149) );
  NOR4_X1 U20301 ( .A1(n14195), .A2(n10188), .A3(n17091), .A4(n17090), .ZN(
        n17092) );
  NAND4_X1 U20302 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n17149), .A4(n17092), .ZN(n17095) );
  NAND2_X1 U20303 ( .A1(n17365), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17094) );
  NAND2_X1 U20304 ( .A1(n17115), .A2(n17519), .ZN(n17093) );
  OAI22_X1 U20305 ( .A1(n17115), .A2(n17094), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17093), .ZN(P3_U2672) );
  NAND2_X1 U20306 ( .A1(n17096), .A2(n17095), .ZN(n17097) );
  NAND2_X1 U20307 ( .A1(n17097), .A2(n17365), .ZN(n17114) );
  AOI22_X1 U20308 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20309 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12302), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20310 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20311 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17099) );
  NAND4_X1 U20312 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17108) );
  AOI22_X1 U20313 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20314 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20315 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20316 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17103) );
  NAND4_X1 U20317 ( .A1(n17106), .A2(n17105), .A3(n17104), .A4(n17103), .ZN(
        n17107) );
  NOR2_X1 U20318 ( .A1(n17108), .A2(n17107), .ZN(n17113) );
  NOR3_X1 U20319 ( .A1(n17111), .A2(n17110), .A3(n17109), .ZN(n17112) );
  XOR2_X1 U20320 ( .A(n17113), .B(n17112), .Z(n17381) );
  OAI22_X1 U20321 ( .A1(n17115), .A2(n17114), .B1(n17381), .B2(n17365), .ZN(
        P3_U2673) );
  AOI21_X1 U20322 ( .B1(n17117), .B2(n17122), .A(n17116), .ZN(n17394) );
  NAND2_X1 U20323 ( .A1(n17371), .A2(n17394), .ZN(n17118) );
  OAI221_X1 U20324 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17121), .C1(n17120), 
        .C2(n17119), .A(n17118), .ZN(P3_U2676) );
  INV_X1 U20325 ( .A(n17121), .ZN(n17126) );
  AOI21_X1 U20326 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17365), .A(n17129), .ZN(
        n17125) );
  OAI21_X1 U20327 ( .B1(n17124), .B2(n17123), .A(n17122), .ZN(n17403) );
  OAI22_X1 U20328 ( .A1(n17126), .A2(n17125), .B1(n17365), .B2(n17403), .ZN(
        P3_U2677) );
  AOI21_X1 U20329 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17365), .A(n9902), .ZN(
        n17128) );
  XNOR2_X1 U20330 ( .A(n17127), .B(n17130), .ZN(n17408) );
  OAI22_X1 U20331 ( .A1(n17129), .A2(n17128), .B1(n17365), .B2(n17408), .ZN(
        P3_U2678) );
  AOI21_X1 U20332 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17365), .A(n9903), .ZN(
        n17133) );
  OAI21_X1 U20333 ( .B1(n17132), .B2(n17131), .A(n17130), .ZN(n17413) );
  OAI22_X1 U20334 ( .A1(n9902), .A2(n17133), .B1(n17365), .B2(n17413), .ZN(
        P3_U2679) );
  AOI21_X1 U20335 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17365), .A(n9904), .ZN(
        n17136) );
  XNOR2_X1 U20336 ( .A(n17135), .B(n17134), .ZN(n17418) );
  OAI22_X1 U20337 ( .A1(n9903), .A2(n17136), .B1(n17356), .B2(n17418), .ZN(
        P3_U2680) );
  AOI21_X1 U20338 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17365), .A(n17137), .ZN(
        n17148) );
  AOI22_X1 U20339 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20340 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20341 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20342 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17138) );
  NAND4_X1 U20343 ( .A1(n17141), .A2(n17140), .A3(n17139), .A4(n17138), .ZN(
        n17147) );
  AOI22_X1 U20344 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20345 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20346 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20347 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17142) );
  NAND4_X1 U20348 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17146) );
  NOR2_X1 U20349 ( .A1(n17147), .A2(n17146), .ZN(n17420) );
  OAI22_X1 U20350 ( .A1(n9904), .A2(n17148), .B1(n17420), .B2(n17365), .ZN(
        P3_U2681) );
  NOR2_X1 U20351 ( .A1(n17371), .A2(n17149), .ZN(n17172) );
  AOI22_X1 U20352 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20353 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17158) );
  INV_X1 U20354 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21129) );
  AOI22_X1 U20355 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17150) );
  OAI21_X1 U20356 ( .B1(n9874), .B2(n21129), .A(n17150), .ZN(n17156) );
  AOI22_X1 U20357 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20358 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20359 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20360 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17178), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17151) );
  NAND4_X1 U20361 ( .A1(n17154), .A2(n17153), .A3(n17152), .A4(n17151), .ZN(
        n17155) );
  AOI211_X1 U20362 ( .C1(n17320), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n17156), .B(n17155), .ZN(n17157) );
  NAND3_X1 U20363 ( .A1(n17159), .A2(n17158), .A3(n17157), .ZN(n17425) );
  AOI22_X1 U20364 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17172), .B1(n17371), 
        .B2(n17425), .ZN(n17160) );
  OAI21_X1 U20365 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17161), .A(n17160), .ZN(
        P3_U2682) );
  AOI22_X1 U20366 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20367 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20368 ( .A1(n12245), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20369 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17162) );
  NAND4_X1 U20370 ( .A1(n17165), .A2(n17164), .A3(n17163), .A4(n17162), .ZN(
        n17171) );
  AOI22_X1 U20371 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20372 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20373 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20374 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17166) );
  NAND4_X1 U20375 ( .A1(n17169), .A2(n17168), .A3(n17167), .A4(n17166), .ZN(
        n17170) );
  NOR2_X1 U20376 ( .A1(n17171), .A2(n17170), .ZN(n17432) );
  OAI21_X1 U20377 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n9923), .A(n17172), .ZN(
        n17173) );
  OAI21_X1 U20378 ( .B1(n17432), .B2(n17356), .A(n17173), .ZN(P3_U2683) );
  AOI22_X1 U20379 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20380 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20381 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20382 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17174) );
  NAND4_X1 U20383 ( .A1(n17177), .A2(n17176), .A3(n17175), .A4(n17174), .ZN(
        n17184) );
  AOI22_X1 U20384 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20385 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20386 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17178), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20387 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17179) );
  NAND4_X1 U20388 ( .A1(n17182), .A2(n17181), .A3(n17180), .A4(n17179), .ZN(
        n17183) );
  NOR2_X1 U20389 ( .A1(n17184), .A2(n17183), .ZN(n17440) );
  OAI21_X1 U20390 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17197), .A(n17185), .ZN(
        n17186) );
  AOI22_X1 U20391 ( .A1(n17371), .A2(n17440), .B1(n17186), .B2(n17356), .ZN(
        P3_U2684) );
  AOI22_X1 U20392 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20393 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20394 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14185), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20395 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17187) );
  NAND4_X1 U20396 ( .A1(n17190), .A2(n17189), .A3(n17188), .A4(n17187), .ZN(
        n17196) );
  AOI22_X1 U20397 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20398 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20399 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20400 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17191) );
  NAND4_X1 U20401 ( .A1(n17194), .A2(n17193), .A3(n17192), .A4(n17191), .ZN(
        n17195) );
  NOR2_X1 U20402 ( .A1(n17196), .A2(n17195), .ZN(n17444) );
  NOR2_X1 U20403 ( .A1(n17371), .A2(n17197), .ZN(n17198) );
  OAI21_X1 U20404 ( .B1(n17199), .B2(P3_EBX_REG_18__SCAN_IN), .A(n17198), .ZN(
        n17200) );
  OAI21_X1 U20405 ( .B1(n17444), .B2(n17356), .A(n17200), .ZN(P3_U2685) );
  NAND2_X1 U20406 ( .A1(n17356), .A2(n17211), .ZN(n17226) );
  AOI22_X1 U20407 ( .A1(n12211), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20408 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20409 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17201) );
  OAI21_X1 U20410 ( .B1(n12318), .B2(n21178), .A(n17201), .ZN(n17207) );
  AOI22_X1 U20411 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U20412 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20413 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9827), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20414 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17202) );
  NAND4_X1 U20415 ( .A1(n17205), .A2(n17204), .A3(n17203), .A4(n17202), .ZN(
        n17206) );
  AOI211_X1 U20416 ( .C1(n9822), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17207), .B(n17206), .ZN(n17208) );
  NAND3_X1 U20417 ( .A1(n17210), .A2(n17209), .A3(n17208), .ZN(n17452) );
  NOR2_X1 U20418 ( .A1(n18367), .A2(n17211), .ZN(n17212) );
  AOI22_X1 U20419 ( .A1(n17371), .A2(n17452), .B1(n17212), .B2(n17214), .ZN(
        n17213) );
  OAI21_X1 U20420 ( .B1(n17214), .B2(n17226), .A(n17213), .ZN(P3_U2687) );
  AOI22_X1 U20421 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20422 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20423 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20424 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17215) );
  NAND4_X1 U20425 ( .A1(n17218), .A2(n17217), .A3(n17216), .A4(n17215), .ZN(
        n17224) );
  AOI22_X1 U20426 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20427 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20428 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20429 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17302), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17219) );
  NAND4_X1 U20430 ( .A1(n17222), .A2(n17221), .A3(n17220), .A4(n17219), .ZN(
        n17223) );
  NOR2_X1 U20431 ( .A1(n17224), .A2(n17223), .ZN(n17461) );
  NOR2_X1 U20432 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17225), .ZN(n17227) );
  OAI22_X1 U20433 ( .A1(n17461), .A2(n17365), .B1(n17227), .B2(n17226), .ZN(
        P3_U2688) );
  NOR2_X1 U20434 ( .A1(n18367), .A2(n17228), .ZN(n17253) );
  NAND2_X1 U20435 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17253), .ZN(n17240) );
  AOI22_X1 U20436 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20437 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20438 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20439 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17229) );
  NAND4_X1 U20440 ( .A1(n17232), .A2(n17231), .A3(n17230), .A4(n17229), .ZN(
        n17238) );
  AOI22_X1 U20441 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20442 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20443 ( .A1(n17317), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20444 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17233) );
  NAND4_X1 U20445 ( .A1(n17236), .A2(n17235), .A3(n17234), .A4(n17233), .ZN(
        n17237) );
  NOR2_X1 U20446 ( .A1(n17238), .A2(n17237), .ZN(n17467) );
  NAND3_X1 U20447 ( .A1(n17240), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17356), 
        .ZN(n17239) );
  OAI221_X1 U20448 ( .B1(n17240), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17356), 
        .C2(n17467), .A(n17239), .ZN(P3_U2689) );
  AOI22_X1 U20449 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U20450 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20451 ( .A1(n9827), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9813), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20452 ( .A1(n12242), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17241) );
  NAND4_X1 U20453 ( .A1(n17244), .A2(n17243), .A3(n17242), .A4(n17241), .ZN(
        n17251) );
  AOI22_X1 U20454 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U20455 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20456 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20457 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17246) );
  NAND4_X1 U20458 ( .A1(n17249), .A2(n17248), .A3(n17247), .A4(n17246), .ZN(
        n17250) );
  NOR2_X1 U20459 ( .A1(n17251), .A2(n17250), .ZN(n17468) );
  NOR2_X1 U20460 ( .A1(n17371), .A2(n17253), .ZN(n17265) );
  AOI22_X1 U20461 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17265), .B1(n17253), 
        .B2(n17252), .ZN(n17254) );
  OAI21_X1 U20462 ( .B1(n17468), .B2(n17356), .A(n17254), .ZN(P3_U2690) );
  AOI22_X1 U20463 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20464 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U20465 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20466 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17255) );
  NAND4_X1 U20467 ( .A1(n17258), .A2(n17257), .A3(n17256), .A4(n17255), .ZN(
        n17264) );
  AOI22_X1 U20468 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17262) );
  AOI22_X1 U20469 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U20470 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20471 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9827), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17259) );
  NAND4_X1 U20472 ( .A1(n17262), .A2(n17261), .A3(n17260), .A4(n17259), .ZN(
        n17263) );
  NOR2_X1 U20473 ( .A1(n17264), .A2(n17263), .ZN(n17471) );
  OAI21_X1 U20474 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17280), .A(n17265), .ZN(
        n17266) );
  OAI21_X1 U20475 ( .B1(n17471), .B2(n17356), .A(n17266), .ZN(P3_U2691) );
  OAI21_X1 U20476 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17267), .A(n17365), .ZN(
        n17279) );
  AOI22_X1 U20477 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17283), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20478 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20479 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17303), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20480 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12242), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17268) );
  NAND4_X1 U20481 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17278) );
  AOI22_X1 U20482 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20483 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20484 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20485 ( .A1(n17302), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17273) );
  NAND4_X1 U20486 ( .A1(n17276), .A2(n17275), .A3(n17274), .A4(n17273), .ZN(
        n17277) );
  NOR2_X1 U20487 ( .A1(n17278), .A2(n17277), .ZN(n17475) );
  OAI22_X1 U20488 ( .A1(n17280), .A2(n17279), .B1(n17475), .B2(n17365), .ZN(
        P3_U2692) );
  AOI22_X1 U20489 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20490 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20491 ( .A1(n12242), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17281) );
  OAI21_X1 U20492 ( .B1(n17322), .B2(n17282), .A(n17281), .ZN(n17289) );
  AOI22_X1 U20493 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20494 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9827), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20495 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20496 ( .A1(n17283), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17284) );
  NAND4_X1 U20497 ( .A1(n17287), .A2(n17286), .A3(n17285), .A4(n17284), .ZN(
        n17288) );
  AOI211_X1 U20498 ( .C1(n17320), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17289), .B(n17288), .ZN(n17290) );
  NAND3_X1 U20499 ( .A1(n17292), .A2(n17291), .A3(n17290), .ZN(n17480) );
  INV_X1 U20500 ( .A(n17480), .ZN(n17296) );
  OAI21_X1 U20501 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17294), .A(n17293), .ZN(
        n17295) );
  AOI22_X1 U20502 ( .A1(n17371), .A2(n17296), .B1(n17295), .B2(n17356), .ZN(
        P3_U2693) );
  AOI21_X1 U20503 ( .B1(n17297), .B2(n17338), .A(n17371), .ZN(n17314) );
  AOI22_X1 U20504 ( .A1(n17324), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12247), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U20505 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20506 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17298), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20507 ( .B1(n17300), .B2(n21243), .A(n17299), .ZN(n17309) );
  AOI22_X1 U20508 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17323), .ZN(n17307) );
  AOI22_X1 U20509 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12302), .B1(
        n17301), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U20510 ( .A1(n14185), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12211), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U20511 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17303), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17327), .ZN(n17304) );
  NAND4_X1 U20512 ( .A1(n17307), .A2(n17306), .A3(n17305), .A4(n17304), .ZN(
        n17308) );
  AOI211_X1 U20513 ( .C1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .C2(n17310), .A(
        n17309), .B(n17308), .ZN(n17311) );
  NAND3_X1 U20514 ( .A1(n17313), .A2(n17312), .A3(n17311), .ZN(n17484) );
  AOI22_X1 U20515 ( .A1(n17315), .A2(n17314), .B1(n17484), .B2(n17371), .ZN(
        n17316) );
  INV_X1 U20516 ( .A(n17316), .ZN(P3_U2694) );
  AOI22_X1 U20517 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17317), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20518 ( .A1(n17178), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17335) );
  AOI22_X1 U20519 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12302), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17321) );
  OAI21_X1 U20520 ( .B1(n17322), .B2(n21178), .A(n17321), .ZN(n17333) );
  AOI22_X1 U20521 ( .A1(n17301), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17323), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U20522 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17324), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20523 ( .A1(n17326), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20524 ( .A1(n12247), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17328) );
  NAND4_X1 U20525 ( .A1(n17331), .A2(n17330), .A3(n17329), .A4(n17328), .ZN(
        n17332) );
  AOI211_X1 U20526 ( .C1(n9822), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17333), .B(n17332), .ZN(n17334) );
  NAND3_X1 U20527 ( .A1(n17336), .A2(n17335), .A3(n17334), .ZN(n17487) );
  INV_X1 U20528 ( .A(n17487), .ZN(n17340) );
  NOR3_X1 U20529 ( .A1(n17352), .A2(n17337), .A3(n17347), .ZN(n17346) );
  OAI221_X1 U20530 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17346), .A(n17338), .ZN(n17339) );
  AOI22_X1 U20531 ( .A1(n17371), .A2(n17340), .B1(n17339), .B2(n17356), .ZN(
        P3_U2695) );
  OAI21_X1 U20532 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17346), .A(n17356), .ZN(
        n17342) );
  INV_X1 U20533 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17341) );
  OAI22_X1 U20534 ( .A1(n17343), .A2(n17342), .B1(n17341), .B2(n17365), .ZN(
        P3_U2696) );
  NOR3_X1 U20535 ( .A1(n18367), .A2(n17347), .A3(n17352), .ZN(n17351) );
  AOI21_X1 U20536 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17365), .A(n17351), .ZN(
        n17345) );
  OAI22_X1 U20537 ( .A1(n17346), .A2(n17345), .B1(n17344), .B2(n17365), .ZN(
        P3_U2697) );
  AOI21_X1 U20538 ( .B1(n17347), .B2(n17352), .A(n17371), .ZN(n17348) );
  INV_X1 U20539 ( .A(n17348), .ZN(n17350) );
  INV_X1 U20540 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17349) );
  OAI22_X1 U20541 ( .A1(n17351), .A2(n17350), .B1(n17349), .B2(n17365), .ZN(
        P3_U2698) );
  INV_X1 U20542 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17355) );
  OAI21_X1 U20543 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17353), .A(n17352), .ZN(
        n17354) );
  AOI22_X1 U20544 ( .A1(n17371), .A2(n17355), .B1(n17354), .B2(n17356), .ZN(
        P3_U2699) );
  NAND2_X1 U20545 ( .A1(n17356), .A2(n17357), .ZN(n17363) );
  NOR3_X1 U20546 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18367), .A3(n17357), .ZN(
        n17358) );
  AOI21_X1 U20547 ( .B1(n17371), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n17358), .ZN(n17359) );
  OAI21_X1 U20548 ( .B1(n17360), .B2(n17363), .A(n17359), .ZN(P3_U2700) );
  NOR2_X1 U20549 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17361), .ZN(n17364) );
  INV_X1 U20550 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17362) );
  OAI22_X1 U20551 ( .A1(n17364), .A2(n17363), .B1(n17362), .B2(n17365), .ZN(
        P3_U2701) );
  INV_X1 U20552 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17366) );
  OAI222_X1 U20553 ( .A1(n17369), .A2(n17373), .B1(n17368), .B2(n17367), .C1(
        n17366), .C2(n17365), .ZN(P3_U2702) );
  AOI22_X1 U20554 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17371), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17370), .ZN(n17372) );
  OAI21_X1 U20555 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17373), .A(n17372), .ZN(
        P3_U2703) );
  INV_X1 U20556 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17534) );
  INV_X1 U20557 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17630) );
  NAND4_X1 U20558 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n17492) );
  NAND4_X1 U20559 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_7__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17374) );
  NOR2_X1 U20560 ( .A1(n17492), .A2(n17374), .ZN(n17462) );
  NAND2_X1 U20561 ( .A1(n17517), .A2(n17462), .ZN(n17489) );
  NAND2_X1 U20562 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17463) );
  INV_X1 U20563 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17626) );
  INV_X1 U20564 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17552) );
  NAND4_X1 U20565 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(n17375), .ZN(n17464) );
  NOR2_X2 U20566 ( .A1(n17630), .A2(n17464), .ZN(n17458) );
  NAND2_X1 U20567 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17419) );
  NAND4_X1 U20568 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n17376)
         );
  NOR3_X2 U20569 ( .A1(n17454), .A2(n17419), .A3(n17376), .ZN(n17415) );
  NAND2_X1 U20570 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17415), .ZN(n17414) );
  NOR2_X1 U20571 ( .A1(n18367), .A2(n17414), .ZN(n17410) );
  NAND2_X1 U20572 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17410), .ZN(n17409) );
  NOR2_X2 U20573 ( .A1(n17534), .A2(n17404), .ZN(n17399) );
  NAND2_X1 U20574 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17398), .ZN(n17391) );
  NAND2_X1 U20575 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17387), .ZN(n17386) );
  INV_X1 U20576 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17600) );
  OR2_X1 U20577 ( .A1(n17386), .A2(n17600), .ZN(n17380) );
  NOR2_X1 U20578 ( .A1(n17377), .A2(n9811), .ZN(n17453) );
  NAND2_X1 U20579 ( .A1(n9812), .A2(n17386), .ZN(n17384) );
  OAI21_X1 U20580 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17491), .A(n17384), .ZN(
        n17378) );
  AOI22_X1 U20581 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17453), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17378), .ZN(n17379) );
  OAI21_X1 U20582 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17380), .A(n17379), .ZN(
        P3_U2704) );
  INV_X1 U20583 ( .A(n17453), .ZN(n17431) );
  OAI22_X1 U20584 ( .A1(n17381), .A2(n17512), .B1(n19346), .B2(n17431), .ZN(
        n17382) );
  AOI21_X1 U20585 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n9809), .A(n17382), .ZN(
        n17383) );
  OAI221_X1 U20586 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17386), .C1(n17600), 
        .C2(n17384), .A(n17383), .ZN(P3_U2705) );
  AOI22_X1 U20587 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9809), .B1(n17385), .B2(
        n17521), .ZN(n17389) );
  OAI211_X1 U20588 ( .C1(n17387), .C2(P3_EAX_REG_29__SCAN_IN), .A(n9812), .B(
        n17386), .ZN(n17388) );
  OAI211_X1 U20589 ( .C1(n17431), .C2(n18358), .A(n17389), .B(n17388), .ZN(
        P3_U2706) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9809), .B1(n17390), .B2(
        n17521), .ZN(n17393) );
  OAI211_X1 U20591 ( .C1(n17398), .C2(P3_EAX_REG_28__SCAN_IN), .A(n9812), .B(
        n17391), .ZN(n17392) );
  OAI211_X1 U20592 ( .C1(n17431), .C2(n21189), .A(n17393), .B(n17392), .ZN(
        P3_U2707) );
  AOI21_X1 U20593 ( .B1(P3_EAX_REG_27__SCAN_IN), .B2(n9812), .A(n17399), .ZN(
        n17397) );
  AOI22_X1 U20594 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17453), .B1(n17394), .B2(
        n17521), .ZN(n17396) );
  NAND2_X1 U20595 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9809), .ZN(n17395) );
  OAI211_X1 U20596 ( .C1(n17398), .C2(n17397), .A(n17396), .B(n17395), .ZN(
        P3_U2708) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17453), .ZN(n17402) );
  AOI211_X1 U20598 ( .C1(n17534), .C2(n17404), .A(n17399), .B(n17483), .ZN(
        n17400) );
  INV_X1 U20599 ( .A(n17400), .ZN(n17401) );
  OAI211_X1 U20600 ( .C1(n17512), .C2(n17403), .A(n17402), .B(n17401), .ZN(
        P3_U2709) );
  AOI22_X1 U20601 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17453), .ZN(n17407) );
  OAI211_X1 U20602 ( .C1(n17405), .C2(P3_EAX_REG_25__SCAN_IN), .A(n9812), .B(
        n17404), .ZN(n17406) );
  OAI211_X1 U20603 ( .C1(n17512), .C2(n17408), .A(n17407), .B(n17406), .ZN(
        P3_U2710) );
  AOI22_X1 U20604 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17453), .ZN(n17412) );
  OAI211_X1 U20605 ( .C1(n17410), .C2(P3_EAX_REG_24__SCAN_IN), .A(n9812), .B(
        n17409), .ZN(n17411) );
  OAI211_X1 U20606 ( .C1(n17512), .C2(n17413), .A(n17412), .B(n17411), .ZN(
        P3_U2711) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17453), .ZN(n17417) );
  OAI211_X1 U20608 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17415), .A(n9812), .B(
        n17414), .ZN(n17416) );
  OAI211_X1 U20609 ( .C1(n17512), .C2(n17418), .A(n17417), .B(n17416), .ZN(
        P3_U2712) );
  INV_X1 U20611 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17545) );
  OR3_X1 U20612 ( .A1(n18367), .A2(n17454), .A3(n17419), .ZN(n17441) );
  NAND2_X1 U20613 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17436), .ZN(n17426) );
  NAND2_X1 U20614 ( .A1(n9812), .A2(n17426), .ZN(n17430) );
  OAI21_X1 U20615 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17491), .A(n17430), .ZN(
        n17423) );
  INV_X1 U20616 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17542) );
  NOR3_X1 U20617 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17542), .A3(n17426), .ZN(
        n17422) );
  OAI22_X1 U20618 ( .A1(n17420), .A2(n17512), .B1(n18363), .B2(n17431), .ZN(
        n17421) );
  AOI211_X1 U20619 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17423), .A(n17422), .B(
        n17421), .ZN(n17424) );
  OAI21_X1 U20620 ( .B1(n18362), .B2(n17445), .A(n17424), .ZN(P3_U2713) );
  AOI22_X1 U20621 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17453), .B1(n17521), .B2(
        n17425), .ZN(n17429) );
  OAI22_X1 U20622 ( .A1(n21246), .A2(n17445), .B1(n17426), .B2(
        P3_EAX_REG_21__SCAN_IN), .ZN(n17427) );
  INV_X1 U20623 ( .A(n17427), .ZN(n17428) );
  OAI211_X1 U20624 ( .C1(n17542), .C2(n17430), .A(n17429), .B(n17428), .ZN(
        P3_U2714) );
  INV_X1 U20625 ( .A(n17430), .ZN(n17434) );
  INV_X1 U20626 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21083) );
  OAI22_X1 U20627 ( .A1(n17432), .A2(n17512), .B1(n18351), .B2(n17431), .ZN(
        n17433) );
  AOI221_X1 U20628 ( .B1(n17434), .B2(P3_EAX_REG_20__SCAN_IN), .C1(n17436), 
        .C2(n21083), .A(n17433), .ZN(n17435) );
  OAI21_X1 U20629 ( .B1(n18352), .B2(n17445), .A(n17435), .ZN(P3_U2715) );
  AOI22_X1 U20630 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17453), .ZN(n17439) );
  AOI211_X1 U20631 ( .C1(n17545), .C2(n17441), .A(n17436), .B(n17483), .ZN(
        n17437) );
  INV_X1 U20632 ( .A(n17437), .ZN(n17438) );
  OAI211_X1 U20633 ( .C1(n17440), .C2(n17512), .A(n17439), .B(n17438), .ZN(
        P3_U2716) );
  AOI22_X1 U20634 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17453), .ZN(n17443) );
  INV_X1 U20635 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17585) );
  NOR2_X1 U20636 ( .A1(n17454), .A2(n17585), .ZN(n17446) );
  OAI211_X1 U20637 ( .C1(n17446), .C2(P3_EAX_REG_18__SCAN_IN), .A(n9812), .B(
        n17441), .ZN(n17442) );
  OAI211_X1 U20638 ( .C1(n17444), .C2(n17512), .A(n17443), .B(n17442), .ZN(
        P3_U2717) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9809), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17453), .ZN(n17450) );
  INV_X1 U20640 ( .A(n17454), .ZN(n17448) );
  INV_X1 U20641 ( .A(n17446), .ZN(n17447) );
  OAI211_X1 U20642 ( .C1(n17448), .C2(P3_EAX_REG_17__SCAN_IN), .A(n9812), .B(
        n17447), .ZN(n17449) );
  OAI211_X1 U20643 ( .C1(n17451), .C2(n17512), .A(n17450), .B(n17449), .ZN(
        P3_U2718) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17453), .B1(n17521), .B2(
        n17452), .ZN(n17456) );
  OAI211_X1 U20645 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17458), .A(n9812), .B(
        n17454), .ZN(n17455) );
  OAI211_X1 U20646 ( .C1(n17445), .C2(n18330), .A(n17456), .B(n17455), .ZN(
        P3_U2719) );
  AOI211_X1 U20647 ( .C1(n17630), .C2(n17464), .A(n17483), .B(n17458), .ZN(
        n17459) );
  AOI21_X1 U20648 ( .B1(n17522), .B2(BUF2_REG_15__SCAN_IN), .A(n17459), .ZN(
        n17460) );
  OAI21_X1 U20649 ( .B1(n17461), .B2(n17512), .A(n17460), .ZN(P3_U2720) );
  INV_X1 U20650 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n21252) );
  INV_X1 U20651 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17612) );
  INV_X1 U20652 ( .A(n17491), .ZN(n17516) );
  NAND2_X1 U20653 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17495), .ZN(n17486) );
  NOR3_X1 U20654 ( .A1(n21252), .A2(n17612), .A3(n17486), .ZN(n17474) );
  INV_X1 U20655 ( .A(n17474), .ZN(n17478) );
  NOR2_X1 U20656 ( .A1(n17463), .A2(n17478), .ZN(n17473) );
  AND2_X1 U20657 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17473), .ZN(n17470) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17522), .B1(n17470), .B2(
        n17626), .ZN(n17466) );
  NAND3_X1 U20659 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n9812), .A3(n17464), .ZN(
        n17465) );
  OAI211_X1 U20660 ( .C1(n17467), .C2(n17512), .A(n17466), .B(n17465), .ZN(
        P3_U2721) );
  AOI21_X1 U20661 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n9812), .A(n17473), .ZN(
        n17469) );
  OAI222_X1 U20662 ( .A1(n17515), .A2(n17622), .B1(n17470), .B2(n17469), .C1(
        n17512), .C2(n17468), .ZN(P3_U2722) );
  AOI22_X1 U20663 ( .A1(n17474), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n9812), .ZN(n17472) );
  OAI222_X1 U20664 ( .A1(n17515), .A2(n17618), .B1(n17473), .B2(n17472), .C1(
        n17512), .C2(n17471), .ZN(P3_U2723) );
  INV_X1 U20665 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17556) );
  NOR2_X1 U20666 ( .A1(n17556), .A2(n17478), .ZN(n17477) );
  AOI21_X1 U20667 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n9812), .A(n17474), .ZN(
        n17476) );
  OAI222_X1 U20668 ( .A1(n17515), .A2(n17616), .B1(n17477), .B2(n17476), .C1(
        n17512), .C2(n17475), .ZN(P3_U2724) );
  INV_X1 U20669 ( .A(n17486), .ZN(n17479) );
  OAI221_X1 U20670 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(P3_EAX_REG_9__SCAN_IN), 
        .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17479), .A(n17478), .ZN(n17482) );
  AOI22_X1 U20671 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17522), .B1(n17521), .B2(
        n17480), .ZN(n17481) );
  OAI21_X1 U20672 ( .B1(n17483), .B2(n17482), .A(n17481), .ZN(P3_U2725) );
  NAND2_X1 U20673 ( .A1(n9812), .A2(n17486), .ZN(n17490) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17522), .B1(n17521), .B2(
        n17484), .ZN(n17485) );
  OAI221_X1 U20675 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17486), .C1(n17612), 
        .C2(n17490), .A(n17485), .ZN(P3_U2726) );
  INV_X1 U20676 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17560) );
  AOI22_X1 U20677 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17522), .B1(n17521), .B2(
        n17487), .ZN(n17488) );
  OAI221_X1 U20678 ( .B1(n17490), .B2(n17489), .C1(n17490), .C2(n17560), .A(
        n17488), .ZN(P3_U2727) );
  INV_X1 U20679 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17603) );
  NOR3_X1 U20680 ( .A1(n17603), .A2(n17579), .A3(n17491), .ZN(n17510) );
  NAND2_X1 U20681 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17510), .ZN(n17506) );
  NOR2_X1 U20682 ( .A1(n17492), .A2(n17506), .ZN(n17498) );
  AOI21_X1 U20683 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n9812), .A(n17498), .ZN(
        n17494) );
  OAI222_X1 U20684 ( .A1(n18370), .A2(n17515), .B1(n17495), .B2(n17494), .C1(
        n17512), .C2(n17493), .ZN(P3_U2728) );
  INV_X1 U20685 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17567) );
  INV_X1 U20686 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17572) );
  NOR2_X1 U20687 ( .A1(n17572), .A2(n17506), .ZN(n17509) );
  NAND2_X1 U20688 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17509), .ZN(n17499) );
  NOR2_X1 U20689 ( .A1(n17567), .A2(n17499), .ZN(n17502) );
  AOI21_X1 U20690 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n9812), .A(n17502), .ZN(
        n17497) );
  OAI222_X1 U20691 ( .A1(n18362), .A2(n17515), .B1(n17498), .B2(n17497), .C1(
        n17512), .C2(n17496), .ZN(P3_U2729) );
  INV_X1 U20692 ( .A(n17499), .ZN(n17505) );
  AOI21_X1 U20693 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n9812), .A(n17505), .ZN(
        n17501) );
  OAI222_X1 U20694 ( .A1(n21246), .A2(n17515), .B1(n17502), .B2(n17501), .C1(
        n17512), .C2(n17500), .ZN(P3_U2730) );
  AOI21_X1 U20695 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n9812), .A(n17509), .ZN(
        n17504) );
  OAI222_X1 U20696 ( .A1(n18352), .A2(n17515), .B1(n17505), .B2(n17504), .C1(
        n17512), .C2(n17503), .ZN(P3_U2731) );
  INV_X1 U20697 ( .A(n17506), .ZN(n17514) );
  AOI21_X1 U20698 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n9812), .A(n17514), .ZN(
        n17508) );
  OAI222_X1 U20699 ( .A1(n18347), .A2(n17515), .B1(n17509), .B2(n17508), .C1(
        n17512), .C2(n17507), .ZN(P3_U2732) );
  AOI21_X1 U20700 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n9812), .A(n17510), .ZN(
        n17513) );
  OAI222_X1 U20701 ( .A1(n21142), .A2(n17515), .B1(n17514), .B2(n17513), .C1(
        n17512), .C2(n12436), .ZN(P3_U2733) );
  NAND2_X1 U20702 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17516), .ZN(n17525) );
  INV_X1 U20703 ( .A(n17517), .ZN(n17518) );
  AOI21_X1 U20704 ( .B1(n17519), .B2(n17579), .A(n17518), .ZN(n17524) );
  AOI22_X1 U20705 ( .A1(n17522), .A2(BUF2_REG_1__SCAN_IN), .B1(n17521), .B2(
        n17520), .ZN(n17523) );
  OAI221_X1 U20706 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17525), .C1(n17603), 
        .C2(n17524), .A(n17523), .ZN(P3_U2734) );
  INV_X1 U20707 ( .A(n17827), .ZN(n17994) );
  AND2_X1 U20708 ( .A1(n20977), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NOR2_X1 U20709 ( .A1(n18335), .A2(n17578), .ZN(n20978) );
  AOI22_X1 U20710 ( .A1(n17576), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U20711 ( .B1(n17600), .B2(n17548), .A(n17527), .ZN(P3_U2737) );
  INV_X1 U20712 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17529) );
  AOI22_X1 U20713 ( .A1(n17576), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20714 ( .B1(n17529), .B2(n17548), .A(n17528), .ZN(P3_U2738) );
  INV_X1 U20715 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21203) );
  AOI22_X1 U20716 ( .A1(n17576), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17530) );
  OAI21_X1 U20717 ( .B1(n21203), .B2(n17548), .A(n17530), .ZN(P3_U2739) );
  INV_X1 U20718 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U20719 ( .A1(n17576), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20720 ( .B1(n17532), .B2(n17548), .A(n17531), .ZN(P3_U2740) );
  INV_X2 U20721 ( .A(n17570), .ZN(n17576) );
  AOI22_X1 U20722 ( .A1(n17576), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20723 ( .B1(n17534), .B2(n17548), .A(n17533), .ZN(P3_U2741) );
  INV_X1 U20724 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U20725 ( .A1(n17576), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20726 ( .B1(n17594), .B2(n17548), .A(n17535), .ZN(P3_U2742) );
  INV_X1 U20727 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U20728 ( .A1(n17576), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U20729 ( .B1(n17537), .B2(n17548), .A(n17536), .ZN(P3_U2743) );
  INV_X1 U20730 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20731 ( .A1(n17576), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17538) );
  OAI21_X1 U20732 ( .B1(n17539), .B2(n17548), .A(n17538), .ZN(P3_U2744) );
  INV_X1 U20733 ( .A(P3_UWORD_REG_6__SCAN_IN), .ZN(n21088) );
  AOI22_X1 U20734 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20978), .B1(n20977), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17540) );
  OAI21_X1 U20735 ( .B1(n17570), .B2(n21088), .A(n17540), .ZN(P3_U2745) );
  AOI22_X1 U20736 ( .A1(n17576), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17541) );
  OAI21_X1 U20737 ( .B1(n17542), .B2(n17548), .A(n17541), .ZN(P3_U2746) );
  AOI22_X1 U20738 ( .A1(n17576), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17543) );
  OAI21_X1 U20739 ( .B1(n21083), .B2(n17548), .A(n17543), .ZN(P3_U2747) );
  AOI22_X1 U20740 ( .A1(n17576), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17544) );
  OAI21_X1 U20741 ( .B1(n17545), .B2(n17548), .A(n17544), .ZN(P3_U2748) );
  AOI22_X1 U20742 ( .A1(n17576), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17546) );
  OAI21_X1 U20743 ( .B1(n17585), .B2(n17548), .A(n17546), .ZN(P3_U2750) );
  INV_X1 U20744 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U20745 ( .A1(n17576), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17547) );
  OAI21_X1 U20746 ( .B1(n17583), .B2(n17548), .A(n17547), .ZN(P3_U2751) );
  AOI22_X1 U20747 ( .A1(n17576), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17549) );
  OAI21_X1 U20748 ( .B1(n17630), .B2(n17578), .A(n17549), .ZN(P3_U2752) );
  AOI22_X1 U20749 ( .A1(n17576), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17550) );
  OAI21_X1 U20750 ( .B1(n17626), .B2(n17578), .A(n17550), .ZN(P3_U2753) );
  AOI22_X1 U20751 ( .A1(n17576), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17551) );
  OAI21_X1 U20752 ( .B1(n17552), .B2(n17578), .A(n17551), .ZN(P3_U2754) );
  INV_X1 U20753 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20754 ( .A1(n17576), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17553) );
  OAI21_X1 U20755 ( .B1(n17554), .B2(n17578), .A(n17553), .ZN(P3_U2755) );
  AOI22_X1 U20756 ( .A1(n17576), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17555) );
  OAI21_X1 U20757 ( .B1(n17556), .B2(n17578), .A(n17555), .ZN(P3_U2756) );
  AOI22_X1 U20758 ( .A1(n17576), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17557) );
  OAI21_X1 U20759 ( .B1(n21252), .B2(n17578), .A(n17557), .ZN(P3_U2757) );
  AOI22_X1 U20760 ( .A1(n17576), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17558) );
  OAI21_X1 U20761 ( .B1(n17612), .B2(n17578), .A(n17558), .ZN(P3_U2758) );
  AOI22_X1 U20762 ( .A1(n17576), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17559) );
  OAI21_X1 U20763 ( .B1(n17560), .B2(n17578), .A(n17559), .ZN(P3_U2759) );
  INV_X1 U20764 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U20765 ( .A1(n17576), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17561), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17562) );
  OAI21_X1 U20766 ( .B1(n17563), .B2(n17578), .A(n17562), .ZN(P3_U2760) );
  INV_X1 U20767 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17565) );
  AOI22_X1 U20768 ( .A1(n17576), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17564) );
  OAI21_X1 U20769 ( .B1(n17565), .B2(n17578), .A(n17564), .ZN(P3_U2761) );
  AOI22_X1 U20770 ( .A1(n17576), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17566) );
  OAI21_X1 U20771 ( .B1(n17567), .B2(n17578), .A(n17566), .ZN(P3_U2762) );
  INV_X1 U20772 ( .A(P3_LWORD_REG_4__SCAN_IN), .ZN(n21274) );
  AOI22_X1 U20773 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17568), .B1(n20977), .B2(
        P3_DATAO_REG_4__SCAN_IN), .ZN(n17569) );
  OAI21_X1 U20774 ( .B1(n17570), .B2(n21274), .A(n17569), .ZN(P3_U2763) );
  AOI22_X1 U20775 ( .A1(n17576), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17571) );
  OAI21_X1 U20776 ( .B1(n17572), .B2(n17578), .A(n17571), .ZN(P3_U2764) );
  INV_X1 U20777 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U20778 ( .A1(n17576), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17573) );
  OAI21_X1 U20779 ( .B1(n17574), .B2(n17578), .A(n17573), .ZN(P3_U2765) );
  AOI22_X1 U20780 ( .A1(n17576), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U20781 ( .B1(n17603), .B2(n17578), .A(n17575), .ZN(P3_U2766) );
  AOI22_X1 U20782 ( .A1(n17576), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n20977), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17577) );
  OAI21_X1 U20783 ( .B1(n17579), .B2(n17578), .A(n17577), .ZN(P3_U2767) );
  NAND3_X1 U20784 ( .A1(n18972), .A2(n17581), .A3(n17580), .ZN(n17631) );
  AOI22_X1 U20785 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17623), .ZN(n17582) );
  OAI21_X1 U20786 ( .B1(n17583), .B2(n17631), .A(n17582), .ZN(P3_U2768) );
  AOI22_X1 U20787 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17623), .ZN(n17584) );
  OAI21_X1 U20788 ( .B1(n17585), .B2(n17631), .A(n17584), .ZN(P3_U2769) );
  AOI22_X1 U20789 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17623), .ZN(n17586) );
  OAI21_X1 U20790 ( .B1(n21142), .B2(n17627), .A(n17586), .ZN(P3_U2770) );
  AOI22_X1 U20791 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17623), .ZN(n17587) );
  OAI21_X1 U20792 ( .B1(n18347), .B2(n17627), .A(n17587), .ZN(P3_U2771) );
  AOI22_X1 U20793 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17623), .ZN(n17588) );
  OAI21_X1 U20794 ( .B1(n18352), .B2(n17627), .A(n17588), .ZN(P3_U2772) );
  AOI22_X1 U20795 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17623), .ZN(n17589) );
  OAI21_X1 U20796 ( .B1(n21246), .B2(n17627), .A(n17589), .ZN(P3_U2773) );
  AOI22_X1 U20797 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17623), .ZN(n17590) );
  OAI21_X1 U20798 ( .B1(n18362), .B2(n17627), .A(n17590), .ZN(P3_U2774) );
  AOI22_X1 U20799 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17623), .ZN(n17591) );
  OAI21_X1 U20800 ( .B1(n18370), .B2(n17627), .A(n17591), .ZN(P3_U2775) );
  AOI22_X1 U20801 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17623), .ZN(n17592) );
  OAI21_X1 U20802 ( .B1(n21192), .B2(n17627), .A(n17592), .ZN(P3_U2776) );
  AOI22_X1 U20803 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17623), .ZN(n17593) );
  OAI21_X1 U20804 ( .B1(n17594), .B2(n17631), .A(n17593), .ZN(P3_U2777) );
  AOI22_X1 U20805 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17623), .ZN(n17595) );
  OAI21_X1 U20806 ( .B1(n17614), .B2(n17627), .A(n17595), .ZN(P3_U2778) );
  AOI22_X1 U20807 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17619), .ZN(n17596) );
  OAI21_X1 U20808 ( .B1(n17616), .B2(n17627), .A(n17596), .ZN(P3_U2779) );
  AOI22_X1 U20809 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17619), .ZN(n17597) );
  OAI21_X1 U20810 ( .B1(n17618), .B2(n17627), .A(n17597), .ZN(P3_U2780) );
  AOI22_X1 U20811 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17619), .ZN(n17598) );
  OAI21_X1 U20812 ( .B1(n17622), .B2(n17627), .A(n17598), .ZN(P3_U2781) );
  AOI22_X1 U20813 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17624), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17623), .ZN(n17599) );
  OAI21_X1 U20814 ( .B1(n17600), .B2(n17631), .A(n17599), .ZN(P3_U2782) );
  AOI22_X1 U20815 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17619), .ZN(n17601) );
  OAI21_X1 U20816 ( .B1(n18330), .B2(n17627), .A(n17601), .ZN(P3_U2783) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17623), .ZN(n17602) );
  OAI21_X1 U20818 ( .B1(n17603), .B2(n17631), .A(n17602), .ZN(P3_U2784) );
  AOI22_X1 U20819 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17619), .ZN(n17604) );
  OAI21_X1 U20820 ( .B1(n21142), .B2(n17627), .A(n17604), .ZN(P3_U2785) );
  AOI22_X1 U20821 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17619), .ZN(n17605) );
  OAI21_X1 U20822 ( .B1(n18347), .B2(n17627), .A(n17605), .ZN(P3_U2786) );
  AOI22_X1 U20823 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17623), .ZN(n17606) );
  OAI21_X1 U20824 ( .B1(n18352), .B2(n17627), .A(n17606), .ZN(P3_U2787) );
  AOI22_X1 U20825 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17623), .ZN(n17607) );
  OAI21_X1 U20826 ( .B1(n21246), .B2(n17627), .A(n17607), .ZN(P3_U2788) );
  AOI22_X1 U20827 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17623), .ZN(n17608) );
  OAI21_X1 U20828 ( .B1(n18362), .B2(n17627), .A(n17608), .ZN(P3_U2789) );
  AOI22_X1 U20829 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17623), .ZN(n17609) );
  OAI21_X1 U20830 ( .B1(n18370), .B2(n17627), .A(n17609), .ZN(P3_U2790) );
  AOI22_X1 U20831 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17623), .ZN(n17610) );
  OAI21_X1 U20832 ( .B1(n21192), .B2(n17627), .A(n17610), .ZN(P3_U2791) );
  AOI22_X1 U20833 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17623), .ZN(n17611) );
  OAI21_X1 U20834 ( .B1(n17612), .B2(n17631), .A(n17611), .ZN(P3_U2792) );
  AOI22_X1 U20835 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17619), .ZN(n17613) );
  OAI21_X1 U20836 ( .B1(n17614), .B2(n17627), .A(n17613), .ZN(P3_U2793) );
  AOI22_X1 U20837 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17619), .ZN(n17615) );
  OAI21_X1 U20838 ( .B1(n17616), .B2(n17627), .A(n17615), .ZN(P3_U2794) );
  AOI22_X1 U20839 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17619), .ZN(n17617) );
  OAI21_X1 U20840 ( .B1(n17618), .B2(n17627), .A(n17617), .ZN(P3_U2795) );
  AOI22_X1 U20841 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17619), .ZN(n17621) );
  OAI21_X1 U20842 ( .B1(n17622), .B2(n17627), .A(n17621), .ZN(P3_U2796) );
  AOI22_X1 U20843 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17624), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17623), .ZN(n17625) );
  OAI21_X1 U20844 ( .B1(n17626), .B2(n17631), .A(n17625), .ZN(P3_U2797) );
  INV_X1 U20845 ( .A(P3_LWORD_REG_15__SCAN_IN), .ZN(n21062) );
  OAI222_X1 U20846 ( .A1(n17631), .A2(n17630), .B1(n21062), .B2(n17629), .C1(
        n17628), .C2(n17627), .ZN(P3_U2798) );
  INV_X1 U20847 ( .A(n17700), .ZN(n17735) );
  NAND2_X1 U20848 ( .A1(n17827), .A2(n17632), .ZN(n17633) );
  OAI211_X1 U20849 ( .C1(n9951), .C2(n17829), .A(n17993), .B(n17633), .ZN(
        n17665) );
  AOI21_X1 U20850 ( .B1(n17735), .B2(n17660), .A(n17665), .ZN(n17657) );
  NAND3_X1 U20851 ( .A1(n9951), .A2(n17843), .A3(n10092), .ZN(n17655) );
  AOI21_X1 U20852 ( .B1(n17657), .B2(n17655), .A(n17634), .ZN(n17637) );
  NOR3_X1 U20853 ( .A1(n17794), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17635), .ZN(n17636) );
  AOI211_X1 U20854 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n9816), .A(n17637), .B(
        n17636), .ZN(n17645) );
  NOR2_X1 U20855 ( .A1(n17983), .A2(n17861), .ZN(n17740) );
  OAI22_X1 U20856 ( .A1(n18003), .A2(n17998), .B1(n18002), .B2(n17906), .ZN(
        n17667) );
  NOR2_X1 U20857 ( .A1(n9992), .A2(n17667), .ZN(n17652) );
  NOR3_X1 U20858 ( .A1(n17740), .A2(n17652), .A3(n21268), .ZN(n17642) );
  AOI211_X1 U20859 ( .C1(n17640), .C2(n17639), .A(n17638), .B(n17877), .ZN(
        n17641) );
  AOI211_X1 U20860 ( .C1(n17643), .C2(n17647), .A(n17642), .B(n17641), .ZN(
        n17644) );
  OAI211_X1 U20861 ( .C1(n17831), .C2(n17646), .A(n17645), .B(n17644), .ZN(
        P3_U2802) );
  NOR2_X1 U20862 ( .A1(n18317), .A2(n21163), .ZN(n17999) );
  NOR2_X1 U20863 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17647), .ZN(
        n17651) );
  NAND2_X1 U20864 ( .A1(n17649), .A2(n17648), .ZN(n17650) );
  XNOR2_X1 U20865 ( .A(n17650), .B(n10072), .ZN(n18011) );
  OAI22_X1 U20866 ( .A1(n17652), .A2(n17651), .B1(n18011), .B2(n17877), .ZN(
        n17653) );
  AOI211_X1 U20867 ( .C1(n17846), .C2(n17654), .A(n17999), .B(n17653), .ZN(
        n17656) );
  OAI211_X1 U20868 ( .C1(n17657), .C2(n10092), .A(n17656), .B(n17655), .ZN(
        P3_U2803) );
  AOI21_X1 U20869 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17659), .A(
        n17658), .ZN(n18019) );
  OAI21_X1 U20870 ( .B1(n18364), .B2(n17661), .A(n17660), .ZN(n17664) );
  AOI21_X1 U20871 ( .B1(n17831), .B2(n17700), .A(n17662), .ZN(n17663) );
  NOR2_X1 U20872 ( .A1(n18317), .A2(n18898), .ZN(n18016) );
  AOI211_X1 U20873 ( .C1(n17665), .C2(n17664), .A(n17663), .B(n18016), .ZN(
        n17669) );
  NOR2_X1 U20874 ( .A1(n17709), .A2(n17692), .ZN(n18000) );
  NAND3_X1 U20875 ( .A1(n10060), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n18000), .ZN(n18013) );
  INV_X1 U20876 ( .A(n18013), .ZN(n17666) );
  INV_X1 U20877 ( .A(n17792), .ZN(n17776) );
  AND2_X1 U20878 ( .A1(n18012), .A2(n17776), .ZN(n17710) );
  AOI22_X1 U20879 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17667), .B1(
        n17666), .B2(n17710), .ZN(n17668) );
  OAI211_X1 U20880 ( .C1(n18019), .C2(n17877), .A(n17669), .B(n17668), .ZN(
        P3_U2804) );
  NAND2_X1 U20881 ( .A1(n18132), .A2(n18020), .ZN(n17670) );
  XNOR2_X1 U20882 ( .A(n17670), .B(n18025), .ZN(n18033) );
  NOR2_X1 U20883 ( .A1(n17673), .A2(n18364), .ZN(n17702) );
  AOI211_X1 U20884 ( .C1(n17827), .C2(n17671), .A(n17946), .B(n17702), .ZN(
        n17706) );
  OAI21_X1 U20885 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17700), .A(
        n17706), .ZN(n17687) );
  INV_X1 U20886 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18896) );
  NOR2_X1 U20887 ( .A1(n18317), .A2(n18896), .ZN(n18028) );
  NOR2_X1 U20888 ( .A1(n17688), .A2(n17672), .ZN(n17676) );
  OAI211_X1 U20889 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17673), .B(n17843), .ZN(n17675) );
  OAI22_X1 U20890 ( .A1(n17676), .A2(n17675), .B1(n17674), .B2(n17831), .ZN(
        n17677) );
  AOI211_X1 U20891 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17687), .A(
        n18028), .B(n17677), .ZN(n17683) );
  XNOR2_X1 U20892 ( .A(n17678), .B(n18025), .ZN(n18030) );
  OAI21_X1 U20893 ( .B1(n17780), .B2(n17680), .A(n17679), .ZN(n17681) );
  XNOR2_X1 U20894 ( .A(n17681), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18029) );
  AOI22_X1 U20895 ( .A1(n17983), .A2(n18030), .B1(n17903), .B2(n18029), .ZN(
        n17682) );
  OAI211_X1 U20896 ( .C1(n17906), .C2(n18033), .A(n17683), .B(n17682), .ZN(
        P3_U2805) );
  OR2_X1 U20897 ( .A1(n17690), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18046) );
  NOR2_X1 U20898 ( .A1(n17794), .A2(n17684), .ZN(n17689) );
  OAI22_X1 U20899 ( .A1(n18317), .A2(n18894), .B1(n17831), .B2(n10085), .ZN(
        n17686) );
  AOI221_X1 U20900 ( .B1(n17689), .B2(n17688), .C1(n17687), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17686), .ZN(n17695) );
  NOR2_X1 U20901 ( .A1(n17690), .A2(n17715), .ZN(n18036) );
  OAI21_X1 U20902 ( .B1(n18056), .B2(n17690), .A(n18959), .ZN(n18038) );
  OAI22_X1 U20903 ( .A1(n18036), .A2(n17906), .B1(n17975), .B2(n18038), .ZN(
        n17708) );
  OAI21_X1 U20904 ( .B1(n17693), .B2(n17692), .A(n17691), .ZN(n18034) );
  AOI22_X1 U20905 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17708), .B1(
        n17903), .B2(n18034), .ZN(n17694) );
  OAI211_X1 U20906 ( .C1(n17792), .C2(n18046), .A(n17695), .B(n17694), .ZN(
        P3_U2806) );
  OAI22_X1 U20907 ( .A1(n10072), .A2(n18066), .B1(n17712), .B2(n17696), .ZN(
        n17698) );
  NOR2_X1 U20908 ( .A1(n17698), .A2(n17697), .ZN(n17699) );
  XNOR2_X1 U20909 ( .A(n17699), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18052) );
  NAND2_X1 U20910 ( .A1(n17831), .A2(n17700), .ZN(n17985) );
  AOI22_X1 U20911 ( .A1(n17703), .A2(n17702), .B1(n17701), .B2(n17985), .ZN(
        n17704) );
  NAND2_X1 U20912 ( .A1(n9816), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18051) );
  OAI211_X1 U20913 ( .C1(n17706), .C2(n17705), .A(n17704), .B(n18051), .ZN(
        n17707) );
  AOI221_X1 U20914 ( .B1(n17710), .B2(n17709), .C1(n17708), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17707), .ZN(n17711) );
  OAI21_X1 U20915 ( .B1(n17877), .B2(n18052), .A(n17711), .ZN(P3_U2807) );
  INV_X1 U20916 ( .A(n17712), .ZN(n17713) );
  AOI221_X1 U20917 ( .B1(n17781), .B2(n17713), .C1(n18065), .C2(n17713), .A(
        n17697), .ZN(n17714) );
  XNOR2_X1 U20918 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17714), .ZN(
        n18071) );
  INV_X1 U20919 ( .A(n18065), .ZN(n18055) );
  AOI22_X1 U20920 ( .A1(n17983), .A2(n18056), .B1(n17861), .B2(n17715), .ZN(
        n17791) );
  OAI21_X1 U20921 ( .B1(n18055), .B2(n17740), .A(n17791), .ZN(n17731) );
  NAND2_X1 U20922 ( .A1(n9958), .A2(n17843), .ZN(n17728) );
  AOI221_X1 U20923 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n10094), .C2(n10095), .A(
        n17728), .ZN(n17721) );
  AOI21_X1 U20924 ( .B1(n17827), .B2(n17716), .A(n17946), .ZN(n17717) );
  OAI21_X1 U20925 ( .B1(n9958), .B2(n17829), .A(n17717), .ZN(n17739) );
  AOI21_X1 U20926 ( .B1(n17735), .B2(n21100), .A(n17739), .ZN(n17727) );
  AOI22_X1 U20927 ( .A1(n9816), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17846), 
        .B2(n17718), .ZN(n17719) );
  OAI21_X1 U20928 ( .B1(n17727), .B2(n10095), .A(n17719), .ZN(n17720) );
  AOI211_X1 U20929 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17731), .A(
        n17721), .B(n17720), .ZN(n17723) );
  NAND3_X1 U20930 ( .A1(n18055), .A2(n17776), .A3(n18066), .ZN(n17722) );
  OAI211_X1 U20931 ( .C1(n17877), .C2(n18071), .A(n17723), .B(n17722), .ZN(
        P3_U2808) );
  NAND3_X1 U20932 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10072), .A3(
        n17724), .ZN(n17744) );
  INV_X1 U20933 ( .A(n17765), .ZN(n17745) );
  OAI22_X1 U20934 ( .A1(n18077), .A2(n17744), .B1(n17725), .B2(n17745), .ZN(
        n17726) );
  XNOR2_X1 U20935 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17726), .ZN(
        n18084) );
  NAND2_X1 U20936 ( .A1(n9816), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18082) );
  OAI221_X1 U20937 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17728), .C1(
        n10094), .C2(n17727), .A(n18082), .ZN(n17729) );
  AOI21_X1 U20938 ( .B1(n17846), .B2(n17730), .A(n17729), .ZN(n17733) );
  NOR2_X1 U20939 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18077), .ZN(
        n18081) );
  NAND2_X1 U20940 ( .A1(n18105), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18072) );
  NOR2_X1 U20941 ( .A1(n17792), .A2(n18072), .ZN(n17755) );
  AOI22_X1 U20942 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17731), .B1(
        n18081), .B2(n17755), .ZN(n17732) );
  OAI211_X1 U20943 ( .C1(n18084), .C2(n17877), .A(n17733), .B(n17732), .ZN(
        P3_U2809) );
  INV_X1 U20944 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18101) );
  NOR2_X1 U20945 ( .A1(n18101), .A2(n18072), .ZN(n18086) );
  NAND2_X1 U20946 ( .A1(n18086), .A2(n18088), .ZN(n18094) );
  OAI21_X1 U20947 ( .B1(n18364), .B2(n17734), .A(n21100), .ZN(n17738) );
  AOI21_X1 U20948 ( .B1(n17831), .B2(n17700), .A(n17736), .ZN(n17737) );
  NOR2_X1 U20949 ( .A1(n18317), .A2(n18886), .ZN(n18091) );
  AOI211_X1 U20950 ( .C1(n17739), .C2(n17738), .A(n17737), .B(n18091), .ZN(
        n17743) );
  OAI21_X1 U20951 ( .B1(n17740), .B2(n18086), .A(n17791), .ZN(n17754) );
  AOI221_X1 U20952 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17744), 
        .C1(n18101), .C2(n17763), .A(n17697), .ZN(n17741) );
  XNOR2_X1 U20953 ( .A(n17741), .B(n18088), .ZN(n18092) );
  AOI22_X1 U20954 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17754), .B1(
        n17903), .B2(n18092), .ZN(n17742) );
  OAI211_X1 U20955 ( .C1(n17792), .C2(n18094), .A(n17743), .B(n17742), .ZN(
        P3_U2810) );
  OAI21_X1 U20956 ( .B1(n17745), .B2(n17763), .A(n17744), .ZN(n17746) );
  XOR2_X1 U20957 ( .A(n17746), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18097) );
  INV_X1 U20958 ( .A(n18097), .ZN(n17757) );
  OAI21_X1 U20959 ( .B1(n17946), .B2(n17748), .A(n17882), .ZN(n17771) );
  OAI21_X1 U20960 ( .B1(n17747), .B2(n17994), .A(n17771), .ZN(n17760) );
  AOI22_X1 U20961 ( .A1(n9816), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17760), .ZN(n17751) );
  NOR2_X1 U20962 ( .A1(n17794), .A2(n17748), .ZN(n17762) );
  OAI211_X1 U20963 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17762), .B(n17749), .ZN(n17750) );
  OAI211_X1 U20964 ( .C1(n17831), .C2(n17752), .A(n17751), .B(n17750), .ZN(
        n17753) );
  AOI221_X1 U20965 ( .B1(n17755), .B2(n18101), .C1(n17754), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17753), .ZN(n17756) );
  OAI21_X1 U20966 ( .B1(n17757), .B2(n17877), .A(n17756), .ZN(P3_U2811) );
  NAND2_X1 U20967 ( .A1(n18105), .A2(n17764), .ZN(n18112) );
  OAI22_X1 U20968 ( .A1(n18317), .A2(n18882), .B1(n17831), .B2(n17758), .ZN(
        n17759) );
  AOI221_X1 U20969 ( .B1(n17762), .B2(n17761), .C1(n17760), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17759), .ZN(n17768) );
  OAI21_X1 U20970 ( .B1(n18105), .B2(n17792), .A(n17791), .ZN(n17777) );
  OAI21_X1 U20971 ( .B1(n17764), .B2(n17780), .A(n17763), .ZN(n17766) );
  XNOR2_X1 U20972 ( .A(n17766), .B(n17765), .ZN(n18108) );
  AOI22_X1 U20973 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17777), .B1(
        n17903), .B2(n18108), .ZN(n17767) );
  OAI211_X1 U20974 ( .C1(n17792), .C2(n18112), .A(n17768), .B(n17767), .ZN(
        P3_U2812) );
  AOI21_X1 U20975 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17770), .A(
        n17769), .ZN(n18119) );
  NOR2_X1 U20976 ( .A1(n18317), .A2(n18881), .ZN(n18115) );
  AOI221_X1 U20977 ( .B1(n18364), .B2(n17773), .C1(n17772), .C2(n17773), .A(
        n17771), .ZN(n17774) );
  AOI211_X1 U20978 ( .C1(n17775), .C2(n17985), .A(n18115), .B(n17774), .ZN(
        n17779) );
  NOR2_X1 U20979 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18125), .ZN(
        n18117) );
  AOI22_X1 U20980 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17777), .B1(
        n17776), .B2(n18117), .ZN(n17778) );
  OAI211_X1 U20981 ( .C1(n18119), .C2(n17877), .A(n17779), .B(n17778), .ZN(
        P3_U2813) );
  NOR2_X1 U20982 ( .A1(n17780), .A2(n18189), .ZN(n17879) );
  AOI22_X1 U20983 ( .A1(n17879), .A2(n10077), .B1(n17781), .B2(n17780), .ZN(
        n17782) );
  XNOR2_X1 U20984 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17782), .ZN(
        n18128) );
  OAI211_X1 U20985 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17783), .B(n17843), .ZN(n17787) );
  INV_X1 U20986 ( .A(n17783), .ZN(n17793) );
  AOI21_X1 U20987 ( .B1(n17948), .B2(n17793), .A(n17946), .ZN(n17811) );
  OAI21_X1 U20988 ( .B1(n17784), .B2(n17994), .A(n17811), .ZN(n17797) );
  AOI22_X1 U20989 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17797), .B1(
        n17846), .B2(n17785), .ZN(n17786) );
  NAND2_X1 U20990 ( .A1(n9816), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18129) );
  OAI211_X1 U20991 ( .C1(n17788), .C2(n17787), .A(n17786), .B(n18129), .ZN(
        n17789) );
  AOI21_X1 U20992 ( .B1(n17903), .B2(n18128), .A(n17789), .ZN(n17790) );
  OAI221_X1 U20993 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17792), 
        .C1(n18125), .C2(n17791), .A(n17790), .ZN(P3_U2814) );
  NOR2_X1 U20994 ( .A1(n17817), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18138) );
  NAND2_X1 U20995 ( .A1(n17983), .A2(n18056), .ZN(n17808) );
  NOR2_X1 U20996 ( .A1(n17794), .A2(n17793), .ZN(n17799) );
  OAI22_X1 U20997 ( .A1(n18317), .A2(n18876), .B1(n17831), .B2(n17795), .ZN(
        n17796) );
  AOI221_X1 U20998 ( .B1(n17799), .B2(n17798), .C1(n17797), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17796), .ZN(n17807) );
  OAI21_X1 U20999 ( .B1(n17802), .B2(n17800), .A(n17801), .ZN(n17803) );
  OAI221_X1 U21000 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n12276), 
        .C1(n18169), .C2(n10072), .A(n17803), .ZN(n17804) );
  XNOR2_X1 U21001 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17804), .ZN(
        n18140) );
  NOR2_X1 U21002 ( .A1(n18132), .A2(n17906), .ZN(n17805) );
  NAND2_X1 U21003 ( .A1(n12277), .A2(n17809), .ZN(n18136) );
  AOI22_X1 U21004 ( .A1(n17903), .A2(n18140), .B1(n17805), .B2(n18136), .ZN(
        n17806) );
  OAI211_X1 U21005 ( .C1(n18138), .C2(n17808), .A(n17807), .B(n17806), .ZN(
        P3_U2815) );
  NAND2_X1 U21006 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18175), .ZN(
        n18146) );
  NOR2_X1 U21007 ( .A1(n18150), .A2(n18146), .ZN(n18148) );
  OAI221_X1 U21008 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17810), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18148), .A(n17809), .ZN(
        n18161) );
  AOI221_X1 U21009 ( .B1(n17813), .B2(n17812), .C1(n18364), .C2(n17812), .A(
        n17811), .ZN(n17814) );
  NOR2_X1 U21010 ( .A1(n18317), .A2(n18875), .ZN(n18156) );
  AOI211_X1 U21011 ( .C1(n17815), .C2(n17985), .A(n17814), .B(n18156), .ZN(
        n17822) );
  INV_X1 U21012 ( .A(n18146), .ZN(n18145) );
  NAND2_X1 U21013 ( .A1(n18145), .A2(n17816), .ZN(n18165) );
  AOI221_X1 U21014 ( .B1(n18150), .B2(n12276), .C1(n18165), .C2(n12276), .A(
        n17817), .ZN(n18158) );
  INV_X1 U21015 ( .A(n17879), .ZN(n17866) );
  INV_X1 U21016 ( .A(n18148), .ZN(n18152) );
  OAI21_X1 U21017 ( .B1(n17866), .B2(n18152), .A(n17819), .ZN(n17820) );
  XOR2_X1 U21018 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17820), .Z(
        n18157) );
  AOI22_X1 U21019 ( .A1(n17983), .A2(n18158), .B1(n17903), .B2(n18157), .ZN(
        n17821) );
  OAI211_X1 U21020 ( .C1(n17906), .C2(n18161), .A(n17822), .B(n17821), .ZN(
        P3_U2816) );
  AND2_X1 U21021 ( .A1(n18959), .A2(n18165), .ZN(n17824) );
  NOR2_X1 U21022 ( .A1(n18189), .A2(n18146), .ZN(n18168) );
  INV_X1 U21023 ( .A(n18168), .ZN(n17823) );
  AOI22_X1 U21024 ( .A1(n17825), .A2(n17824), .B1(n17861), .B2(n17823), .ZN(
        n17852) );
  AOI21_X1 U21025 ( .B1(n17827), .B2(n17826), .A(n17946), .ZN(n17828) );
  OAI21_X1 U21026 ( .B1(n17844), .B2(n17829), .A(n17828), .ZN(n17847) );
  NOR2_X1 U21027 ( .A1(n18317), .A2(n18872), .ZN(n17836) );
  INV_X1 U21028 ( .A(n17830), .ZN(n17834) );
  OAI211_X1 U21029 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17844), .B(n17843), .ZN(n17833) );
  OAI22_X1 U21030 ( .A1(n17834), .A2(n17833), .B1(n17832), .B2(n17831), .ZN(
        n17835) );
  AOI211_X1 U21031 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17847), .A(
        n17836), .B(n17835), .ZN(n17841) );
  OAI22_X1 U21032 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n10072), .B1(
        n18146), .B2(n17800), .ZN(n17838) );
  OAI21_X1 U21033 ( .B1(n10072), .B2(n17837), .A(n17838), .ZN(n17839) );
  XNOR2_X1 U21034 ( .A(n17839), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18172) );
  NOR2_X1 U21035 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18146), .ZN(
        n18171) );
  AOI22_X1 U21036 ( .A1(n17903), .A2(n18172), .B1(n18171), .B2(n17874), .ZN(
        n17840) );
  OAI211_X1 U21037 ( .C1(n17852), .C2(n18150), .A(n17841), .B(n17840), .ZN(
        P3_U2817) );
  NAND2_X1 U21038 ( .A1(n18175), .A2(n17874), .ZN(n17853) );
  AOI21_X1 U21039 ( .B1(n18175), .B2(n17879), .A(n17837), .ZN(n17842) );
  XNOR2_X1 U21040 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17842), .ZN(
        n18183) );
  NAND2_X1 U21041 ( .A1(n17844), .A2(n17843), .ZN(n17849) );
  AOI22_X1 U21042 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17847), .B1(
        n17846), .B2(n17845), .ZN(n17848) );
  NAND2_X1 U21043 ( .A1(n9816), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18184) );
  OAI211_X1 U21044 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17849), .A(
        n17848), .B(n18184), .ZN(n17850) );
  AOI21_X1 U21045 ( .B1(n17903), .B2(n18183), .A(n17850), .ZN(n17851) );
  OAI221_X1 U21046 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17853), 
        .C1(n18169), .C2(n17852), .A(n17851), .ZN(P3_U2818) );
  INV_X1 U21047 ( .A(n18196), .ZN(n17862) );
  AOI21_X1 U21048 ( .B1(n17879), .B2(n17862), .A(n17854), .ZN(n17855) );
  XNOR2_X1 U21049 ( .A(n17855), .B(n21056), .ZN(n18202) );
  INV_X1 U21050 ( .A(n17894), .ZN(n17891) );
  NAND2_X1 U21051 ( .A1(n18705), .A2(n17891), .ZN(n17923) );
  NOR2_X1 U21052 ( .A1(n17856), .A2(n17923), .ZN(n17868) );
  NOR2_X1 U21053 ( .A1(n17859), .A2(n17868), .ZN(n17860) );
  OAI22_X1 U21054 ( .A1(n17977), .A2(n17857), .B1(n18317), .B2(n18868), .ZN(
        n17858) );
  AOI221_X1 U21055 ( .B1(n17882), .B2(n17860), .C1(n17859), .C2(n17868), .A(
        n17858), .ZN(n17864) );
  INV_X1 U21056 ( .A(n17874), .ZN(n17890) );
  AOI22_X1 U21057 ( .A1(n17983), .A2(n18191), .B1(n17861), .B2(n18189), .ZN(
        n17889) );
  OAI21_X1 U21058 ( .B1(n17862), .B2(n17890), .A(n17889), .ZN(n17873) );
  NOR2_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18196), .ZN(
        n18187) );
  AOI22_X1 U21060 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17873), .B1(
        n18187), .B2(n17874), .ZN(n17863) );
  OAI211_X1 U21061 ( .C1(n18202), .C2(n17877), .A(n17864), .B(n17863), .ZN(
        P3_U2819) );
  OAI21_X1 U21062 ( .B1(n18212), .B2(n17866), .A(n17865), .ZN(n17867) );
  XNOR2_X1 U21063 ( .A(n17867), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18210) );
  INV_X1 U21064 ( .A(n17923), .ZN(n17913) );
  NAND3_X1 U21065 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17913), .ZN(n17881) );
  INV_X1 U21066 ( .A(n17882), .ZN(n17990) );
  AOI211_X1 U21067 ( .C1(n17881), .C2(n17869), .A(n17990), .B(n17868), .ZN(
        n17871) );
  NOR2_X1 U21068 ( .A1(n18317), .A2(n18866), .ZN(n17870) );
  AOI211_X1 U21069 ( .C1(n17872), .C2(n17985), .A(n17871), .B(n17870), .ZN(
        n17876) );
  OAI221_X1 U21070 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17874), .A(n17873), .ZN(
        n17875) );
  OAI211_X1 U21071 ( .C1(n18210), .C2(n17877), .A(n17876), .B(n17875), .ZN(
        P3_U2820) );
  NOR2_X1 U21072 ( .A1(n17879), .A2(n17878), .ZN(n17880) );
  XOR2_X1 U21073 ( .A(n17880), .B(n18212), .Z(n18211) );
  NOR2_X1 U21074 ( .A1(n18317), .A2(n18864), .ZN(n17887) );
  INV_X1 U21075 ( .A(n17881), .ZN(n17885) );
  AOI22_X1 U21076 ( .A1(n17892), .A2(n17913), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17882), .ZN(n17884) );
  OAI22_X1 U21077 ( .A1(n17885), .A2(n17884), .B1(n17977), .B2(n17883), .ZN(
        n17886) );
  AOI211_X1 U21078 ( .C1(n17903), .C2(n18211), .A(n17887), .B(n17886), .ZN(
        n17888) );
  OAI221_X1 U21079 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17890), .C1(
        n18212), .C2(n17889), .A(n17888), .ZN(P3_U2821) );
  NAND2_X1 U21080 ( .A1(n17891), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17893) );
  AOI211_X1 U21081 ( .C1(n17895), .C2(n17893), .A(n17892), .B(n18364), .ZN(
        n17898) );
  AOI21_X1 U21082 ( .B1(n17948), .B2(n17894), .A(n17946), .ZN(n17910) );
  OAI22_X1 U21083 ( .A1(n17977), .A2(n17896), .B1(n17910), .B2(n17895), .ZN(
        n17897) );
  AOI211_X1 U21084 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n9816), .A(n17898), .B(
        n17897), .ZN(n17905) );
  AOI21_X1 U21085 ( .B1(n17900), .B2(n18233), .A(n17899), .ZN(n18237) );
  OAI21_X1 U21086 ( .B1(n10072), .B2(n17902), .A(n17901), .ZN(n18235) );
  AOI22_X1 U21087 ( .A1(n17983), .A2(n18237), .B1(n17903), .B2(n18235), .ZN(
        n17904) );
  OAI211_X1 U21088 ( .C1(n17906), .C2(n18241), .A(n17905), .B(n17904), .ZN(
        P3_U2822) );
  NAND2_X1 U21089 ( .A1(n17908), .A2(n17907), .ZN(n17909) );
  XOR2_X1 U21090 ( .A(n17909), .B(n18228), .Z(n18245) );
  INV_X1 U21091 ( .A(n18245), .ZN(n17919) );
  INV_X1 U21092 ( .A(n17910), .ZN(n17911) );
  NOR2_X1 U21093 ( .A1(n18317), .A2(n18860), .ZN(n18243) );
  AOI221_X1 U21094 ( .B1(n17913), .B2(n17912), .C1(n17911), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18243), .ZN(n17918) );
  AOI21_X1 U21095 ( .B1(n18228), .B2(n17915), .A(n17914), .ZN(n18244) );
  AOI22_X1 U21096 ( .A1(n17986), .A2(n18244), .B1(n17916), .B2(n17985), .ZN(
        n17917) );
  OAI211_X1 U21097 ( .C1(n17998), .C2(n17919), .A(n17918), .B(n17917), .ZN(
        P3_U2823) );
  NAND2_X1 U21098 ( .A1(n18705), .A2(n17920), .ZN(n17942) );
  OAI21_X1 U21099 ( .B1(n17990), .B2(n17921), .A(n17942), .ZN(n17922) );
  AOI22_X1 U21100 ( .A1(n9816), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17923), .B2(
        n17922), .ZN(n17930) );
  AOI21_X1 U21101 ( .B1(n17925), .B2(n18229), .A(n17924), .ZN(n18254) );
  AOI21_X1 U21102 ( .B1(n17926), .B2(n17928), .A(n17927), .ZN(n18253) );
  AOI22_X1 U21103 ( .A1(n17983), .A2(n18254), .B1(n17986), .B2(n18253), .ZN(
        n17929) );
  OAI211_X1 U21104 ( .C1(n17977), .C2(n17931), .A(n17930), .B(n17929), .ZN(
        P3_U2824) );
  OAI21_X1 U21105 ( .B1(n17934), .B2(n17932), .A(n17933), .ZN(n17935) );
  XNOR2_X1 U21106 ( .A(n17935), .B(n18260), .ZN(n18266) );
  AOI21_X1 U21107 ( .B1(n17938), .B2(n17937), .A(n17936), .ZN(n18258) );
  AOI22_X1 U21108 ( .A1(n17983), .A2(n18258), .B1(n9816), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17945) );
  AOI221_X1 U21109 ( .B1(n17946), .B2(n17940), .C1(n17939), .C2(n17940), .A(
        n17990), .ZN(n17943) );
  AOI22_X1 U21110 ( .A1(n17943), .A2(n17942), .B1(n17941), .B2(n17985), .ZN(
        n17944) );
  OAI211_X1 U21111 ( .C1(n17997), .C2(n18266), .A(n17945), .B(n17944), .ZN(
        P3_U2825) );
  AOI21_X1 U21112 ( .B1(n17948), .B2(n17947), .A(n17946), .ZN(n17966) );
  AOI21_X1 U21113 ( .B1(n18261), .B2(n17950), .A(n17949), .ZN(n18274) );
  OAI22_X1 U21114 ( .A1(n18317), .A2(n18854), .B1(n18364), .B2(n17951), .ZN(
        n17952) );
  AOI21_X1 U21115 ( .B1(n17983), .B2(n18274), .A(n17952), .ZN(n17957) );
  AOI21_X1 U21116 ( .B1(n9957), .B2(n17954), .A(n17953), .ZN(n18267) );
  AOI22_X1 U21117 ( .A1(n17986), .A2(n18267), .B1(n17955), .B2(n17985), .ZN(
        n17956) );
  OAI211_X1 U21118 ( .C1(n17958), .C2(n17966), .A(n17957), .B(n17956), .ZN(
        P3_U2826) );
  AOI21_X1 U21119 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17993), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17967) );
  AOI21_X1 U21120 ( .B1(n17961), .B2(n17960), .A(n17959), .ZN(n18285) );
  AOI22_X1 U21121 ( .A1(n17983), .A2(n18285), .B1(n9816), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17965) );
  AOI21_X1 U21122 ( .B1(n18280), .B2(n17962), .A(n9987), .ZN(n18284) );
  AOI22_X1 U21123 ( .A1(n17986), .A2(n18284), .B1(n17963), .B2(n17985), .ZN(
        n17964) );
  OAI211_X1 U21124 ( .C1(n17967), .C2(n17966), .A(n17965), .B(n17964), .ZN(
        P3_U2827) );
  AOI21_X1 U21125 ( .B1(n17970), .B2(n17969), .A(n17968), .ZN(n18299) );
  NOR2_X1 U21126 ( .A1(n18317), .A2(n18850), .ZN(n18300) );
  AOI21_X1 U21127 ( .B1(n17973), .B2(n17972), .A(n17971), .ZN(n17974) );
  NAND2_X1 U21128 ( .A1(n18959), .A2(n17974), .ZN(n18295) );
  OAI22_X1 U21129 ( .A1(n17977), .A2(n17976), .B1(n17975), .B2(n18295), .ZN(
        n17978) );
  AOI211_X1 U21130 ( .C1(n17986), .C2(n18299), .A(n18300), .B(n17978), .ZN(
        n17979) );
  OAI221_X1 U21131 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18364), .C1(
        n17980), .C2(n17993), .A(n17979), .ZN(P3_U2828) );
  NOR2_X1 U21132 ( .A1(n17992), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17982) );
  XNOR2_X1 U21133 ( .A(n17982), .B(n17981), .ZN(n18306) );
  AOI22_X1 U21134 ( .A1(n17983), .A2(n18306), .B1(n9816), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17988) );
  AOI21_X1 U21135 ( .B1(n17981), .B2(n17991), .A(n17984), .ZN(n18304) );
  AOI22_X1 U21136 ( .A1(n17986), .A2(n18304), .B1(n17989), .B2(n17985), .ZN(
        n17987) );
  OAI211_X1 U21137 ( .C1(n17990), .C2(n17989), .A(n17988), .B(n17987), .ZN(
        P3_U2829) );
  OAI21_X1 U21138 ( .B1(n17992), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17991), .ZN(n18321) );
  INV_X1 U21139 ( .A(n18321), .ZN(n18323) );
  NAND3_X1 U21140 ( .A1(n18928), .A2(n17994), .A3(n17993), .ZN(n17995) );
  AOI22_X1 U21141 ( .A1(n9816), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17995), .ZN(n17996) );
  OAI221_X1 U21142 ( .B1(n18323), .B2(n17998), .C1(n18321), .C2(n17997), .A(
        n17996), .ZN(P3_U2830) );
  AOI21_X1 U21143 ( .B1(n18310), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17999), .ZN(n18010) );
  NOR2_X1 U21144 ( .A1(n18197), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18271) );
  INV_X1 U21145 ( .A(n18271), .ZN(n18290) );
  AND3_X1 U21146 ( .A1(n18290), .A2(n18103), .A3(n18012), .ZN(n18054) );
  AOI21_X1 U21147 ( .B1(n18054), .B2(n18000), .A(n18269), .ZN(n18022) );
  OAI22_X1 U21148 ( .A1(n18788), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18197), .B2(n18001), .ZN(n18005) );
  OAI22_X1 U21149 ( .A1(n18003), .A2(n18057), .B1(n18002), .B2(n18167), .ZN(
        n18004) );
  NOR4_X1 U21150 ( .A1(n18006), .A2(n18022), .A3(n18005), .A4(n18004), .ZN(
        n18014) );
  OAI211_X1 U21151 ( .C1(n18788), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18014), .ZN(n18007) );
  OAI211_X1 U21152 ( .C1(n18008), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18315), .B(n18007), .ZN(n18009) );
  OAI211_X1 U21153 ( .C1(n18011), .C2(n18221), .A(n18010), .B(n18009), .ZN(
        P3_U2835) );
  NAND2_X1 U21154 ( .A1(n18012), .A2(n18053), .ZN(n18047) );
  OAI22_X1 U21155 ( .A1(n18014), .A2(n10060), .B1(n18013), .B2(n18047), .ZN(
        n18015) );
  AOI22_X1 U21156 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18310), .B1(
        n18315), .B2(n18015), .ZN(n18018) );
  INV_X1 U21157 ( .A(n18016), .ZN(n18017) );
  OAI211_X1 U21158 ( .C1(n18019), .C2(n18221), .A(n18018), .B(n18017), .ZN(
        P3_U2836) );
  OAI221_X1 U21159 ( .B1(n18770), .B2(n18020), .C1(n18770), .C2(n18040), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18021) );
  OAI21_X1 U21160 ( .B1(n18022), .B2(n18021), .A(n18315), .ZN(n18023) );
  AOI221_X1 U21161 ( .B1(n18026), .B2(n18025), .C1(n18024), .C2(n18025), .A(
        n18023), .ZN(n18027) );
  AOI211_X1 U21162 ( .C1(n18310), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18028), .B(n18027), .ZN(n18032) );
  AOI22_X1 U21163 ( .A1(n18307), .A2(n18030), .B1(n18236), .B2(n18029), .ZN(
        n18031) );
  OAI211_X1 U21164 ( .C1(n18240), .C2(n18033), .A(n18032), .B(n18031), .ZN(
        P3_U2837) );
  AOI22_X1 U21165 ( .A1(n9816), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18236), 
        .B2(n18034), .ZN(n18045) );
  INV_X1 U21166 ( .A(n18035), .ZN(n18230) );
  INV_X1 U21167 ( .A(n18310), .ZN(n18272) );
  OAI21_X1 U21168 ( .B1(n18167), .B2(n18036), .A(n18272), .ZN(n18037) );
  INV_X1 U21169 ( .A(n18037), .ZN(n18039) );
  OAI211_X1 U21170 ( .C1(n18269), .C2(n18054), .A(n18039), .B(n18038), .ZN(
        n18043) );
  AOI21_X1 U21171 ( .B1(n18105), .B2(n18040), .A(n18770), .ZN(n18058) );
  AOI211_X1 U21172 ( .C1(n18784), .C2(n18041), .A(n18058), .B(n18043), .ZN(
        n18042) );
  AOI21_X1 U21173 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18042), .A(
        n9816), .ZN(n18048) );
  OAI211_X1 U21174 ( .C1(n18230), .C2(n18043), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18048), .ZN(n18044) );
  OAI211_X1 U21175 ( .C1(n18046), .C2(n18095), .A(n18045), .B(n18044), .ZN(
        P3_U2838) );
  NOR2_X1 U21176 ( .A1(n18310), .A2(n18047), .ZN(n18049) );
  OAI21_X1 U21177 ( .B1(n18049), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18048), .ZN(n18050) );
  OAI211_X1 U21178 ( .C1(n18052), .C2(n18221), .A(n18051), .B(n18050), .ZN(
        P3_U2839) );
  INV_X1 U21179 ( .A(n18053), .ZN(n18067) );
  AOI21_X1 U21180 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18197), .A(
        n18054), .ZN(n18063) );
  NOR2_X1 U21181 ( .A1(n18959), .A2(n18190), .ZN(n18188) );
  OAI22_X1 U21182 ( .A1(n18788), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18055), .B2(n18188), .ZN(n18076) );
  INV_X1 U21183 ( .A(n18056), .ZN(n18139) );
  OAI22_X1 U21184 ( .A1(n18139), .A2(n18057), .B1(n18132), .B2(n18167), .ZN(
        n18124) );
  NOR2_X1 U21185 ( .A1(n18058), .A2(n18124), .ZN(n18104) );
  AOI21_X1 U21186 ( .B1(n18103), .B2(n18086), .A(n18788), .ZN(n18059) );
  INV_X1 U21187 ( .A(n18059), .ZN(n18060) );
  OAI211_X1 U21188 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n18770), .A(
        n18104), .B(n18060), .ZN(n18074) );
  INV_X1 U21189 ( .A(n18077), .ZN(n18061) );
  OAI22_X1 U21190 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18205), .B1(
        n18061), .B2(n18770), .ZN(n18062) );
  NOR4_X1 U21191 ( .A1(n18063), .A2(n18076), .A3(n18074), .A4(n18062), .ZN(
        n18064) );
  AOI221_X1 U21192 ( .B1(n18067), .B2(n18066), .C1(n18065), .C2(n18066), .A(
        n18064), .ZN(n18068) );
  AOI22_X1 U21193 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18310), .B1(
        n18315), .B2(n18068), .ZN(n18070) );
  NAND2_X1 U21194 ( .A1(n9816), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18069) );
  OAI211_X1 U21195 ( .C1(n18071), .C2(n18221), .A(n18070), .B(n18069), .ZN(
        P3_U2840) );
  NOR2_X1 U21196 ( .A1(n18095), .A2(n18072), .ZN(n18096) );
  OAI21_X1 U21197 ( .B1(n18120), .B2(n18072), .A(n18786), .ZN(n18073) );
  INV_X1 U21198 ( .A(n18073), .ZN(n18075) );
  NOR3_X1 U21199 ( .A1(n18075), .A2(n18074), .A3(n18302), .ZN(n18085) );
  NAND2_X1 U21200 ( .A1(n18197), .A2(n18770), .ZN(n18309) );
  AOI21_X1 U21201 ( .B1(n18077), .B2(n18309), .A(n18076), .ZN(n18079) );
  AOI211_X1 U21202 ( .C1(n18085), .C2(n18079), .A(n9816), .B(n18078), .ZN(
        n18080) );
  AOI21_X1 U21203 ( .B1(n18096), .B2(n18081), .A(n18080), .ZN(n18083) );
  OAI211_X1 U21204 ( .C1(n18084), .C2(n18221), .A(n18083), .B(n18082), .ZN(
        P3_U2841) );
  OAI21_X1 U21205 ( .B1(n18086), .B2(n18188), .A(n18085), .ZN(n18087) );
  NAND2_X1 U21206 ( .A1(n18087), .A2(n18317), .ZN(n18100) );
  NAND3_X1 U21207 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18101), .A3(n18309), 
        .ZN(n18089) );
  AOI21_X1 U21208 ( .B1(n18100), .B2(n18089), .A(n18088), .ZN(n18090) );
  AOI211_X1 U21209 ( .C1(n18092), .C2(n18236), .A(n18091), .B(n18090), .ZN(
        n18093) );
  OAI21_X1 U21210 ( .B1(n18095), .B2(n18094), .A(n18093), .ZN(P3_U2842) );
  AOI22_X1 U21211 ( .A1(n18236), .A2(n18097), .B1(n18096), .B2(n18101), .ZN(
        n18099) );
  NAND2_X1 U21212 ( .A1(n9816), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18098) );
  OAI211_X1 U21213 ( .C1(n18101), .C2(n18100), .A(n18099), .B(n18098), .ZN(
        P3_U2843) );
  OAI21_X1 U21214 ( .B1(n18197), .B2(n18944), .A(n18788), .ZN(n18293) );
  AOI22_X1 U21215 ( .A1(n18784), .A2(n18296), .B1(n18268), .B2(n18293), .ZN(
        n18281) );
  INV_X1 U21216 ( .A(n18250), .ZN(n18224) );
  NOR2_X1 U21217 ( .A1(n18281), .A2(n18224), .ZN(n18242) );
  NAND2_X1 U21218 ( .A1(n18102), .A2(n18242), .ZN(n18177) );
  NAND2_X1 U21219 ( .A1(n10077), .A2(n18213), .ZN(n18131) );
  NAND2_X1 U21220 ( .A1(n18103), .A2(n18290), .ZN(n18107) );
  OAI211_X1 U21221 ( .C1(n18105), .C2(n18188), .A(n18315), .B(n18104), .ZN(
        n18106) );
  AOI221_X1 U21222 ( .B1(n18125), .B2(n18288), .C1(n18107), .C2(n18288), .A(
        n18106), .ZN(n18113) );
  AOI221_X1 U21223 ( .B1(n18269), .B2(n18113), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18113), .A(n9816), .ZN(
        n18109) );
  AOI22_X1 U21224 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18109), .B1(
        n18236), .B2(n18108), .ZN(n18111) );
  NAND2_X1 U21225 ( .A1(n9816), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18110) );
  OAI211_X1 U21226 ( .C1(n18112), .C2(n18131), .A(n18111), .B(n18110), .ZN(
        P3_U2844) );
  INV_X1 U21227 ( .A(n18131), .ZN(n18116) );
  NOR3_X1 U21228 ( .A1(n9816), .A2(n18113), .A3(n10064), .ZN(n18114) );
  AOI211_X1 U21229 ( .C1(n18117), .C2(n18116), .A(n18115), .B(n18114), .ZN(
        n18118) );
  OAI21_X1 U21230 ( .B1(n18119), .B2(n18221), .A(n18118), .ZN(P3_U2845) );
  OAI21_X1 U21231 ( .B1(n18223), .B2(n18225), .A(n18768), .ZN(n18214) );
  OAI21_X1 U21232 ( .B1(n18788), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n18214), .ZN(n18207) );
  AOI211_X1 U21233 ( .C1(n18120), .C2(n18786), .A(n18207), .B(n12277), .ZN(
        n18122) );
  NAND2_X1 U21234 ( .A1(n18784), .A2(n18121), .ZN(n18192) );
  OAI211_X1 U21235 ( .C1(n18123), .C2(n18205), .A(n18122), .B(n18192), .ZN(
        n18135) );
  AOI211_X1 U21236 ( .C1(n18230), .C2(n18135), .A(n18302), .B(n18124), .ZN(
        n18126) );
  NOR3_X1 U21237 ( .A1(n9816), .A2(n18126), .A3(n18125), .ZN(n18127) );
  AOI21_X1 U21238 ( .B1(n18236), .B2(n18128), .A(n18127), .ZN(n18130) );
  OAI211_X1 U21239 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18131), .A(
        n18130), .B(n18129), .ZN(P3_U2846) );
  NOR2_X1 U21240 ( .A1(n18132), .A2(n18167), .ZN(n18137) );
  OAI21_X1 U21241 ( .B1(n18133), .B2(n18177), .A(n12277), .ZN(n18134) );
  AOI22_X1 U21242 ( .A1(n18137), .A2(n18136), .B1(n18135), .B2(n18134), .ZN(
        n18144) );
  AOI22_X1 U21243 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18310), .B1(
        n9816), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18143) );
  NOR2_X1 U21244 ( .A1(n18139), .A2(n18138), .ZN(n18141) );
  AOI22_X1 U21245 ( .A1(n18307), .A2(n18141), .B1(n18236), .B2(n18140), .ZN(
        n18142) );
  OAI211_X1 U21246 ( .C1(n18144), .C2(n18302), .A(n18143), .B(n18142), .ZN(
        P3_U2847) );
  NOR2_X1 U21247 ( .A1(n18944), .A2(n18162), .ZN(n18216) );
  OAI221_X1 U21248 ( .B1(n18197), .B2(n18145), .C1(n18197), .C2(n18216), .A(
        n18192), .ZN(n18164) );
  AOI211_X1 U21249 ( .C1(n18784), .C2(n18146), .A(n12276), .B(n18164), .ZN(
        n18147) );
  OAI221_X1 U21250 ( .B1(n18788), .B2(n18149), .C1(n18788), .C2(n18148), .A(
        n18147), .ZN(n18151) );
  OAI221_X1 U21251 ( .B1(n18151), .B2(n18150), .C1(n18151), .C2(n18309), .A(
        n18315), .ZN(n18154) );
  OR2_X1 U21252 ( .A1(n18177), .A2(n18152), .ZN(n18153) );
  AOI222_X1 U21253 ( .A1(n12276), .A2(n18154), .B1(n12276), .B2(n18153), .C1(
        n18154), .C2(n18272), .ZN(n18155) );
  AOI211_X1 U21254 ( .C1(n18236), .C2(n18157), .A(n18156), .B(n18155), .ZN(
        n18160) );
  NAND2_X1 U21255 ( .A1(n18307), .A2(n18158), .ZN(n18159) );
  OAI211_X1 U21256 ( .C1(n18161), .C2(n18240), .A(n18160), .B(n18159), .ZN(
        P3_U2848) );
  OAI21_X1 U21257 ( .B1(n18196), .B2(n18162), .A(n18768), .ZN(n18163) );
  OAI21_X1 U21258 ( .B1(n18175), .B2(n18770), .A(n18163), .ZN(n18199) );
  AOI211_X1 U21259 ( .C1(n18959), .C2(n18165), .A(n18164), .B(n18199), .ZN(
        n18166) );
  OAI21_X1 U21260 ( .B1(n18168), .B2(n18167), .A(n18166), .ZN(n18180) );
  AOI21_X1 U21261 ( .B1(n18768), .B2(n21056), .A(n18169), .ZN(n18179) );
  OAI21_X1 U21262 ( .B1(n18205), .B2(n18179), .A(n18272), .ZN(n18170) );
  OAI21_X1 U21263 ( .B1(n18180), .B2(n18170), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U21264 ( .A1(n18236), .A2(n18172), .B1(n18213), .B2(n18171), .ZN(
        n18173) );
  OAI221_X1 U21265 ( .B1(n9816), .B2(n18174), .C1(n18317), .C2(n18872), .A(
        n18173), .ZN(P3_U2849) );
  INV_X1 U21266 ( .A(n18175), .ZN(n18176) );
  AOI21_X1 U21267 ( .B1(n18178), .B2(n18177), .A(n18176), .ZN(n18182) );
  INV_X1 U21268 ( .A(n18179), .ZN(n18181) );
  OAI22_X1 U21269 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18182), .B1(
        n18181), .B2(n18180), .ZN(n18186) );
  AOI22_X1 U21270 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18310), .B1(
        n18236), .B2(n18183), .ZN(n18185) );
  OAI211_X1 U21271 ( .C1(n18302), .C2(n18186), .A(n18185), .B(n18184), .ZN(
        P3_U2850) );
  AOI22_X1 U21272 ( .A1(n9816), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18213), 
        .B2(n18187), .ZN(n18201) );
  INV_X1 U21273 ( .A(n18188), .ZN(n18195) );
  AOI21_X1 U21274 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18216), .A(
        n18197), .ZN(n18194) );
  AOI22_X1 U21275 ( .A1(n18959), .A2(n18191), .B1(n18190), .B2(n18189), .ZN(
        n18193) );
  NAND2_X1 U21276 ( .A1(n18193), .A2(n18192), .ZN(n18218) );
  AOI211_X1 U21277 ( .C1(n18196), .C2(n18195), .A(n18194), .B(n18218), .ZN(
        n18204) );
  OAI211_X1 U21278 ( .C1(n18197), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18315), .B(n18204), .ZN(n18198) );
  OAI211_X1 U21279 ( .C1(n18199), .C2(n18198), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18317), .ZN(n18200) );
  OAI211_X1 U21280 ( .C1(n18202), .C2(n18221), .A(n18201), .B(n18200), .ZN(
        P3_U2851) );
  NOR2_X1 U21281 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18212), .ZN(
        n18203) );
  AOI22_X1 U21282 ( .A1(n9816), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18213), 
        .B2(n18203), .ZN(n18209) );
  OAI211_X1 U21283 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18205), .A(
        n18204), .B(n18272), .ZN(n18206) );
  OAI211_X1 U21284 ( .C1(n18207), .C2(n18206), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18317), .ZN(n18208) );
  OAI211_X1 U21285 ( .C1(n18210), .C2(n18221), .A(n18209), .B(n18208), .ZN(
        P3_U2852) );
  INV_X1 U21286 ( .A(n18211), .ZN(n18222) );
  AOI22_X1 U21287 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n9816), .B1(n18213), .B2(
        n18212), .ZN(n18220) );
  AOI21_X1 U21288 ( .B1(n18768), .B2(n18233), .A(n18786), .ZN(n18215) );
  OAI211_X1 U21289 ( .C1(n18216), .C2(n18215), .A(n18315), .B(n18214), .ZN(
        n18217) );
  OAI211_X1 U21290 ( .C1(n18218), .C2(n18217), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18317), .ZN(n18219) );
  OAI211_X1 U21291 ( .C1(n18222), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2853) );
  NOR4_X1 U21292 ( .A1(n18281), .A2(n18224), .A3(n18302), .A4(n18223), .ZN(
        n18234) );
  AOI21_X1 U21293 ( .B1(n18288), .B2(n18225), .A(n18271), .ZN(n18226) );
  OAI21_X1 U21294 ( .B1(n18227), .B2(n18770), .A(n18226), .ZN(n18251) );
  AOI211_X1 U21295 ( .C1(n18230), .C2(n18229), .A(n18228), .B(n18251), .ZN(
        n18249) );
  OAI21_X1 U21296 ( .B1(n18249), .B2(n18273), .A(n18272), .ZN(n18232) );
  INV_X1 U21297 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18863) );
  NOR2_X1 U21298 ( .A1(n18317), .A2(n18863), .ZN(n18231) );
  AOI221_X1 U21299 ( .B1(n18234), .B2(n18233), .C1(n18232), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18231), .ZN(n18239) );
  AOI22_X1 U21300 ( .A1(n18307), .A2(n18237), .B1(n18236), .B2(n18235), .ZN(
        n18238) );
  OAI211_X1 U21301 ( .C1(n18241), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        P3_U2854) );
  OAI221_X1 U21302 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18242), .A(n18315), .ZN(
        n18248) );
  AOI21_X1 U21303 ( .B1(n18310), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18243), .ZN(n18247) );
  AOI22_X1 U21304 ( .A1(n18307), .A2(n18245), .B1(n18305), .B2(n18244), .ZN(
        n18246) );
  OAI211_X1 U21305 ( .C1(n18249), .C2(n18248), .A(n18247), .B(n18246), .ZN(
        P3_U2855) );
  NOR2_X1 U21306 ( .A1(n18281), .A2(n18302), .ZN(n18259) );
  NAND2_X1 U21307 ( .A1(n18250), .A2(n18259), .ZN(n18257) );
  INV_X1 U21308 ( .A(n18251), .ZN(n18252) );
  AOI21_X1 U21309 ( .B1(n18315), .B2(n18252), .A(n9816), .ZN(n18262) );
  AOI22_X1 U21310 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18262), .B1(
        n9816), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U21311 ( .A1(n18307), .A2(n18254), .B1(n18305), .B2(n18253), .ZN(
        n18255) );
  OAI211_X1 U21312 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18257), .A(
        n18256), .B(n18255), .ZN(P3_U2856) );
  INV_X1 U21313 ( .A(n18305), .ZN(n18320) );
  AOI22_X1 U21314 ( .A1(n9816), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18307), .B2(
        n18258), .ZN(n18265) );
  NAND2_X1 U21315 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18259), .ZN(
        n18278) );
  OAI21_X1 U21316 ( .B1(n18261), .B2(n18278), .A(n18260), .ZN(n18263) );
  NAND2_X1 U21317 ( .A1(n18263), .A2(n18262), .ZN(n18264) );
  OAI211_X1 U21318 ( .C1(n18320), .C2(n18266), .A(n18265), .B(n18264), .ZN(
        P3_U2857) );
  AOI22_X1 U21319 ( .A1(n9816), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18305), .B2(
        n18267), .ZN(n18277) );
  OAI22_X1 U21320 ( .A1(n18269), .A2(n18268), .B1(n18770), .B2(n18296), .ZN(
        n18270) );
  NOR3_X1 U21321 ( .A1(n18271), .A2(n18280), .A3(n18270), .ZN(n18279) );
  OAI21_X1 U21322 ( .B1(n18279), .B2(n18273), .A(n18272), .ZN(n18275) );
  AOI22_X1 U21323 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18275), .B1(
        n18307), .B2(n18274), .ZN(n18276) );
  OAI211_X1 U21324 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18278), .A(
        n18277), .B(n18276), .ZN(P3_U2858) );
  NOR2_X1 U21325 ( .A1(n18317), .A2(n18852), .ZN(n18283) );
  AOI211_X1 U21326 ( .C1(n18281), .C2(n18280), .A(n18279), .B(n18302), .ZN(
        n18282) );
  AOI211_X1 U21327 ( .C1(n18310), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18283), .B(n18282), .ZN(n18287) );
  AOI22_X1 U21328 ( .A1(n18307), .A2(n18285), .B1(n18305), .B2(n18284), .ZN(
        n18286) );
  NAND2_X1 U21329 ( .A1(n18287), .A2(n18286), .ZN(P3_U2859) );
  NOR2_X1 U21330 ( .A1(n18944), .A2(n18927), .ZN(n18289) );
  AOI22_X1 U21331 ( .A1(n18784), .A2(n18289), .B1(n18288), .B2(n18927), .ZN(
        n18291) );
  AOI21_X1 U21332 ( .B1(n18291), .B2(n18290), .A(n18292), .ZN(n18298) );
  NAND3_X1 U21333 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18293), .A3(
        n18292), .ZN(n18294) );
  OAI211_X1 U21334 ( .C1(n18296), .C2(n18770), .A(n18295), .B(n18294), .ZN(
        n18297) );
  AOI211_X1 U21335 ( .C1(n18299), .C2(n18808), .A(n18298), .B(n18297), .ZN(
        n18303) );
  AOI21_X1 U21336 ( .B1(n18310), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18300), .ZN(n18301) );
  OAI21_X1 U21337 ( .B1(n18303), .B2(n18302), .A(n18301), .ZN(P3_U2860) );
  AOI22_X1 U21338 ( .A1(n18307), .A2(n18306), .B1(n18305), .B2(n18304), .ZN(
        n18314) );
  NAND2_X1 U21339 ( .A1(n9816), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18313) );
  OAI211_X1 U21340 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18768), .A(
        n18308), .B(n18927), .ZN(n18312) );
  AND3_X1 U21341 ( .A1(n18944), .A2(n18309), .A3(n18315), .ZN(n18316) );
  OAI21_X1 U21342 ( .B1(n18310), .B2(n18316), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18311) );
  NAND4_X1 U21343 ( .A1(n18314), .A2(n18313), .A3(n18312), .A4(n18311), .ZN(
        P3_U2861) );
  AOI21_X1 U21344 ( .B1(n18788), .B2(n18315), .A(n18944), .ZN(n18318) );
  AOI221_X1 U21345 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n9816), .C1(n18318), 
        .C2(n18317), .A(n18316), .ZN(n18319) );
  OAI221_X1 U21346 ( .B1(n18323), .B2(n18322), .C1(n18321), .C2(n18320), .A(
        n18319), .ZN(P3_U2862) );
  INV_X1 U21347 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18791) );
  AOI211_X1 U21348 ( .C1(n21210), .C2(n18324), .A(n18928), .B(n18819), .ZN(
        n18812) );
  OAI21_X1 U21349 ( .B1(n18812), .B2(n18375), .A(n18329), .ZN(n18325) );
  OAI221_X1 U21350 ( .B1(n18791), .B2(n18966), .C1(n18791), .C2(n18329), .A(
        n18325), .ZN(P3_U2863) );
  INV_X1 U21351 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18801) );
  NOR2_X1 U21352 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18798), .ZN(
        n18509) );
  INV_X1 U21353 ( .A(n18509), .ZN(n18485) );
  NAND2_X1 U21354 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18798), .ZN(
        n18602) );
  INV_X1 U21355 ( .A(n18602), .ZN(n18577) );
  NAND2_X1 U21356 ( .A1(n18394), .A2(n18577), .ZN(n18623) );
  AND2_X1 U21357 ( .A1(n18485), .A2(n18623), .ZN(n18327) );
  OAI22_X1 U21358 ( .A1(n18328), .A2(n18801), .B1(n18327), .B2(n18326), .ZN(
        P3_U2866) );
  NOR2_X1 U21359 ( .A1(n18802), .A2(n18329), .ZN(P3_U2867) );
  NAND2_X1 U21360 ( .A1(n18705), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18679) );
  NOR2_X1 U21361 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18793), .ZN(
        n18578) );
  INV_X1 U21362 ( .A(n18578), .ZN(n18486) );
  NAND2_X1 U21363 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18331) );
  NOR2_X2 U21364 ( .A1(n18486), .A2(n18331), .ZN(n18686) );
  INV_X1 U21365 ( .A(n18686), .ZN(n18698) );
  NAND2_X1 U21366 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18705), .ZN(n18710) );
  INV_X1 U21367 ( .A(n18710), .ZN(n18672) );
  NOR2_X1 U21368 ( .A1(n18331), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18704) );
  NAND2_X1 U21369 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18704), .ZN(
        n18735) );
  INV_X1 U21370 ( .A(n18735), .ZN(n18751) );
  NOR2_X2 U21371 ( .A1(n18674), .A2(n18330), .ZN(n18700) );
  NOR2_X1 U21372 ( .A1(n18801), .A2(n18554), .ZN(n18703) );
  NAND2_X1 U21373 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18703), .ZN(
        n18759) );
  INV_X1 U21374 ( .A(n18759), .ZN(n18732) );
  NAND2_X1 U21375 ( .A1(n18793), .A2(n18791), .ZN(n18794) );
  NAND2_X1 U21376 ( .A1(n18798), .A2(n18801), .ZN(n18415) );
  NOR2_X2 U21377 ( .A1(n18794), .A2(n18415), .ZN(n18434) );
  NOR2_X1 U21378 ( .A1(n18732), .A2(n18434), .ZN(n18395) );
  NOR2_X1 U21379 ( .A1(n18820), .A2(n18395), .ZN(n18371) );
  AOI22_X1 U21380 ( .A1(n18672), .A2(n18751), .B1(n18700), .B2(n18371), .ZN(
        n18337) );
  NOR2_X1 U21381 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18791), .ZN(
        n18463) );
  NOR2_X1 U21382 ( .A1(n18578), .A2(n18463), .ZN(n18624) );
  NOR2_X1 U21383 ( .A1(n18624), .A2(n18331), .ZN(n18671) );
  AOI211_X1 U21384 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18395), .B(n18674), .ZN(
        n18332) );
  AOI21_X1 U21385 ( .B1(n18705), .B2(n18671), .A(n18332), .ZN(n18372) );
  NAND2_X1 U21386 ( .A1(n18334), .A2(n18333), .ZN(n18353) );
  NOR2_X2 U21387 ( .A1(n18335), .A2(n18353), .ZN(n18706) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18372), .B1(
        n18434), .B2(n18706), .ZN(n18336) );
  OAI211_X1 U21389 ( .C1(n18679), .C2(n18698), .A(n18337), .B(n18336), .ZN(
        P3_U2868) );
  INV_X1 U21390 ( .A(n18434), .ZN(n18428) );
  INV_X1 U21391 ( .A(n18353), .ZN(n18368) );
  NAND2_X1 U21392 ( .A1(n18368), .A2(n18338), .ZN(n18716) );
  AND2_X1 U21393 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18705), .ZN(n18713) );
  NOR2_X2 U21394 ( .A1(n18674), .A2(n18339), .ZN(n18711) );
  AOI22_X1 U21395 ( .A1(n18713), .A2(n18751), .B1(n18711), .B2(n18371), .ZN(
        n18341) );
  NOR2_X2 U21396 ( .A1(n18364), .A2(n13791), .ZN(n18712) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18372), .B1(
        n18712), .B2(n18686), .ZN(n18340) );
  OAI211_X1 U21398 ( .C1(n18428), .C2(n18716), .A(n18341), .B(n18340), .ZN(
        P3_U2869) );
  NAND2_X1 U21399 ( .A1(n18368), .A2(n18342), .ZN(n18722) );
  NOR2_X2 U21400 ( .A1(n18674), .A2(n21142), .ZN(n18717) );
  AND2_X1 U21401 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18705), .ZN(n18719) );
  AOI22_X1 U21402 ( .A1(n18717), .A2(n18371), .B1(n18719), .B2(n18751), .ZN(
        n18345) );
  NOR2_X2 U21403 ( .A1(n18364), .A2(n18343), .ZN(n18718) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18372), .B1(
        n18718), .B2(n18686), .ZN(n18344) );
  OAI211_X1 U21405 ( .C1(n18428), .C2(n18722), .A(n18345), .B(n18344), .ZN(
        P3_U2870) );
  NAND2_X1 U21406 ( .A1(n18368), .A2(n18346), .ZN(n18728) );
  NOR2_X2 U21407 ( .A1(n18674), .A2(n18347), .ZN(n18723) );
  AND2_X1 U21408 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18705), .ZN(n18725) );
  AOI22_X1 U21409 ( .A1(n18723), .A2(n18371), .B1(n18725), .B2(n18751), .ZN(
        n18350) );
  NOR2_X2 U21410 ( .A1(n18364), .A2(n18348), .ZN(n18724) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18372), .B1(
        n18724), .B2(n18686), .ZN(n18349) );
  OAI211_X1 U21412 ( .C1(n18428), .C2(n18728), .A(n18350), .B(n18349), .ZN(
        P3_U2871) );
  NOR2_X1 U21413 ( .A1(n18364), .A2(n18351), .ZN(n18657) );
  NAND2_X1 U21414 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18705), .ZN(n18661) );
  INV_X1 U21415 ( .A(n18661), .ZN(n18730) );
  NOR2_X2 U21416 ( .A1(n18674), .A2(n18352), .ZN(n18729) );
  AOI22_X1 U21417 ( .A1(n18730), .A2(n18751), .B1(n18729), .B2(n18371), .ZN(
        n18356) );
  NOR2_X2 U21418 ( .A1(n18354), .A2(n18353), .ZN(n18731) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18372), .B1(
        n18434), .B2(n18731), .ZN(n18355) );
  OAI211_X1 U21420 ( .C1(n18736), .C2(n18698), .A(n18356), .B(n18355), .ZN(
        P3_U2872) );
  NAND2_X1 U21421 ( .A1(n18368), .A2(n18357), .ZN(n18742) );
  NOR2_X2 U21422 ( .A1(n18364), .A2(n15455), .ZN(n18739) );
  NOR2_X2 U21423 ( .A1(n18674), .A2(n21246), .ZN(n18737) );
  AOI22_X1 U21424 ( .A1(n18739), .A2(n18686), .B1(n18737), .B2(n18371), .ZN(
        n18360) );
  NOR2_X2 U21425 ( .A1(n18358), .A2(n18364), .ZN(n18738) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18372), .B1(
        n18738), .B2(n18751), .ZN(n18359) );
  OAI211_X1 U21427 ( .C1(n18428), .C2(n18742), .A(n18360), .B(n18359), .ZN(
        P3_U2873) );
  NAND2_X1 U21428 ( .A1(n18368), .A2(n18361), .ZN(n18748) );
  NOR2_X2 U21429 ( .A1(n18674), .A2(n18362), .ZN(n18744) );
  NOR2_X2 U21430 ( .A1(n19346), .A2(n18364), .ZN(n18743) );
  AOI22_X1 U21431 ( .A1(n18744), .A2(n18371), .B1(n18743), .B2(n18751), .ZN(
        n18366) );
  NOR2_X2 U21432 ( .A1(n18364), .A2(n18363), .ZN(n18745) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18372), .B1(
        n18745), .B2(n18686), .ZN(n18365) );
  OAI211_X1 U21434 ( .C1(n18428), .C2(n18748), .A(n18366), .B(n18365), .ZN(
        P3_U2874) );
  NAND2_X1 U21435 ( .A1(n18368), .A2(n18367), .ZN(n18758) );
  NOR2_X2 U21436 ( .A1(n18364), .A2(n18369), .ZN(n18754) );
  NOR2_X2 U21437 ( .A1(n18674), .A2(n18370), .ZN(n18750) );
  AOI22_X1 U21438 ( .A1(n18754), .A2(n18751), .B1(n18750), .B2(n18371), .ZN(
        n18374) );
  NOR2_X2 U21439 ( .A1(n18364), .A2(n15450), .ZN(n18752) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18372), .B1(
        n18752), .B2(n18686), .ZN(n18373) );
  OAI211_X1 U21441 ( .C1(n18428), .C2(n18758), .A(n18374), .B(n18373), .ZN(
        P3_U2875) );
  INV_X1 U21442 ( .A(n18679), .ZN(n18701) );
  NAND2_X1 U21443 ( .A1(n18793), .A2(n18699), .ZN(n18553) );
  NOR2_X1 U21444 ( .A1(n18415), .A2(n18553), .ZN(n18390) );
  AOI22_X1 U21445 ( .A1(n18732), .A2(n18701), .B1(n18700), .B2(n18390), .ZN(
        n18377) );
  INV_X1 U21446 ( .A(n18415), .ZN(n18417) );
  NOR2_X1 U21447 ( .A1(n18674), .A2(n18375), .ZN(n18702) );
  INV_X1 U21448 ( .A(n18702), .ZN(n18416) );
  NOR2_X1 U21449 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18416), .ZN(
        n18461) );
  AOI22_X1 U21450 ( .A1(n18705), .A2(n18703), .B1(n18417), .B2(n18461), .ZN(
        n18391) );
  NAND2_X1 U21451 ( .A1(n18417), .A2(n18463), .ZN(n18451) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18391), .B1(
        n18457), .B2(n18706), .ZN(n18376) );
  OAI211_X1 U21453 ( .C1(n18710), .C2(n18698), .A(n18377), .B(n18376), .ZN(
        P3_U2876) );
  AOI22_X1 U21454 ( .A1(n18713), .A2(n18686), .B1(n18711), .B2(n18390), .ZN(
        n18379) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18391), .B1(
        n18732), .B2(n18712), .ZN(n18378) );
  OAI211_X1 U21456 ( .C1(n18451), .C2(n18716), .A(n18379), .B(n18378), .ZN(
        P3_U2877) );
  AOI22_X1 U21457 ( .A1(n18732), .A2(n18718), .B1(n18717), .B2(n18390), .ZN(
        n18381) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18391), .B1(
        n18719), .B2(n18686), .ZN(n18380) );
  OAI211_X1 U21459 ( .C1(n18451), .C2(n18722), .A(n18381), .B(n18380), .ZN(
        P3_U2878) );
  AOI22_X1 U21460 ( .A1(n18732), .A2(n18724), .B1(n18723), .B2(n18390), .ZN(
        n18383) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18391), .B1(
        n18725), .B2(n18686), .ZN(n18382) );
  OAI211_X1 U21462 ( .C1(n18451), .C2(n18728), .A(n18383), .B(n18382), .ZN(
        P3_U2879) );
  AOI22_X1 U21463 ( .A1(n18730), .A2(n18686), .B1(n18729), .B2(n18390), .ZN(
        n18385) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18391), .B1(
        n18457), .B2(n18731), .ZN(n18384) );
  OAI211_X1 U21465 ( .C1(n18759), .C2(n18736), .A(n18385), .B(n18384), .ZN(
        P3_U2880) );
  AOI22_X1 U21466 ( .A1(n18738), .A2(n18686), .B1(n18737), .B2(n18390), .ZN(
        n18387) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18391), .B1(
        n18732), .B2(n18739), .ZN(n18386) );
  OAI211_X1 U21468 ( .C1(n18451), .C2(n18742), .A(n18387), .B(n18386), .ZN(
        P3_U2881) );
  AOI22_X1 U21469 ( .A1(n18732), .A2(n18745), .B1(n18744), .B2(n18390), .ZN(
        n18389) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18391), .B1(
        n18743), .B2(n18686), .ZN(n18388) );
  OAI211_X1 U21471 ( .C1(n18451), .C2(n18748), .A(n18389), .B(n18388), .ZN(
        P3_U2882) );
  AOI22_X1 U21472 ( .A1(n18754), .A2(n18686), .B1(n18750), .B2(n18390), .ZN(
        n18393) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18391), .B1(
        n18732), .B2(n18752), .ZN(n18392) );
  OAI211_X1 U21474 ( .C1(n18451), .C2(n18758), .A(n18393), .B(n18392), .ZN(
        P3_U2883) );
  NAND2_X1 U21475 ( .A1(n18578), .A2(n18417), .ZN(n18474) );
  AOI21_X1 U21476 ( .B1(n18474), .B2(n18451), .A(n18820), .ZN(n18411) );
  AOI22_X1 U21477 ( .A1(n18434), .A2(n18701), .B1(n18700), .B2(n18411), .ZN(
        n18398) );
  INV_X1 U21478 ( .A(n18394), .ZN(n18579) );
  AOI221_X1 U21479 ( .B1(n18395), .B2(n18451), .C1(n18579), .C2(n18451), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18396) );
  OAI21_X1 U21480 ( .B1(n18480), .B2(n18396), .A(n18626), .ZN(n18412) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18412), .B1(
        n18480), .B2(n18706), .ZN(n18397) );
  OAI211_X1 U21482 ( .C1(n18759), .C2(n18710), .A(n18398), .B(n18397), .ZN(
        P3_U2884) );
  AOI22_X1 U21483 ( .A1(n18732), .A2(n18713), .B1(n18411), .B2(n18711), .ZN(
        n18400) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18712), .ZN(n18399) );
  OAI211_X1 U21485 ( .C1(n18474), .C2(n18716), .A(n18400), .B(n18399), .ZN(
        P3_U2885) );
  AOI22_X1 U21486 ( .A1(n18732), .A2(n18719), .B1(n18411), .B2(n18717), .ZN(
        n18402) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18718), .ZN(n18401) );
  OAI211_X1 U21488 ( .C1(n18474), .C2(n18722), .A(n18402), .B(n18401), .ZN(
        P3_U2886) );
  AOI22_X1 U21489 ( .A1(n18732), .A2(n18725), .B1(n18411), .B2(n18723), .ZN(
        n18404) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18724), .ZN(n18403) );
  OAI211_X1 U21491 ( .C1(n18474), .C2(n18728), .A(n18404), .B(n18403), .ZN(
        P3_U2887) );
  AOI22_X1 U21492 ( .A1(n18434), .A2(n18657), .B1(n18411), .B2(n18729), .ZN(
        n18406) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18412), .B1(
        n18480), .B2(n18731), .ZN(n18405) );
  OAI211_X1 U21494 ( .C1(n18759), .C2(n18661), .A(n18406), .B(n18405), .ZN(
        P3_U2888) );
  AOI22_X1 U21495 ( .A1(n18732), .A2(n18738), .B1(n18411), .B2(n18737), .ZN(
        n18408) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18739), .ZN(n18407) );
  OAI211_X1 U21497 ( .C1(n18474), .C2(n18742), .A(n18408), .B(n18407), .ZN(
        P3_U2889) );
  AOI22_X1 U21498 ( .A1(n18732), .A2(n18743), .B1(n18411), .B2(n18744), .ZN(
        n18410) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18745), .ZN(n18409) );
  OAI211_X1 U21500 ( .C1(n18474), .C2(n18748), .A(n18410), .B(n18409), .ZN(
        P3_U2890) );
  AOI22_X1 U21501 ( .A1(n18732), .A2(n18754), .B1(n18411), .B2(n18750), .ZN(
        n18414) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18752), .ZN(n18413) );
  OAI211_X1 U21503 ( .C1(n18474), .C2(n18758), .A(n18414), .B(n18413), .ZN(
        P3_U2891) );
  NOR2_X1 U21504 ( .A1(n18793), .A2(n18415), .ZN(n18462) );
  AND2_X1 U21505 ( .A1(n18699), .A2(n18462), .ZN(n18433) );
  AOI22_X1 U21506 ( .A1(n18434), .A2(n18672), .B1(n18700), .B2(n18433), .ZN(
        n18419) );
  AOI21_X1 U21507 ( .B1(n18793), .B2(n18579), .A(n18416), .ZN(n18510) );
  NAND2_X1 U21508 ( .A1(n18417), .A2(n18510), .ZN(n18435) );
  NAND2_X1 U21509 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18462), .ZN(
        n18491) );
  INV_X1 U21510 ( .A(n18491), .ZN(n18505) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18435), .B1(
        n18706), .B2(n18505), .ZN(n18418) );
  OAI211_X1 U21512 ( .C1(n18451), .C2(n18679), .A(n18419), .B(n18418), .ZN(
        P3_U2892) );
  AOI22_X1 U21513 ( .A1(n18434), .A2(n18713), .B1(n18711), .B2(n18433), .ZN(
        n18421) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18435), .B1(
        n18457), .B2(n18712), .ZN(n18420) );
  OAI211_X1 U21515 ( .C1(n18716), .C2(n18491), .A(n18421), .B(n18420), .ZN(
        P3_U2893) );
  AOI22_X1 U21516 ( .A1(n18434), .A2(n18719), .B1(n18717), .B2(n18433), .ZN(
        n18423) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18435), .B1(
        n18457), .B2(n18718), .ZN(n18422) );
  OAI211_X1 U21518 ( .C1(n18722), .C2(n18491), .A(n18423), .B(n18422), .ZN(
        P3_U2894) );
  AOI22_X1 U21519 ( .A1(n18457), .A2(n18724), .B1(n18723), .B2(n18433), .ZN(
        n18425) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18725), .ZN(n18424) );
  OAI211_X1 U21521 ( .C1(n18728), .C2(n18491), .A(n18425), .B(n18424), .ZN(
        P3_U2895) );
  AOI22_X1 U21522 ( .A1(n18457), .A2(n18657), .B1(n18729), .B2(n18433), .ZN(
        n18427) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18435), .B1(
        n18731), .B2(n18505), .ZN(n18426) );
  OAI211_X1 U21524 ( .C1(n18428), .C2(n18661), .A(n18427), .B(n18426), .ZN(
        P3_U2896) );
  AOI22_X1 U21525 ( .A1(n18434), .A2(n18738), .B1(n18737), .B2(n18433), .ZN(
        n18430) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18435), .B1(
        n18457), .B2(n18739), .ZN(n18429) );
  OAI211_X1 U21527 ( .C1(n18742), .C2(n18491), .A(n18430), .B(n18429), .ZN(
        P3_U2897) );
  AOI22_X1 U21528 ( .A1(n18434), .A2(n18743), .B1(n18744), .B2(n18433), .ZN(
        n18432) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18435), .B1(
        n18457), .B2(n18745), .ZN(n18431) );
  OAI211_X1 U21530 ( .C1(n18748), .C2(n18491), .A(n18432), .B(n18431), .ZN(
        P3_U2898) );
  AOI22_X1 U21531 ( .A1(n18434), .A2(n18754), .B1(n18750), .B2(n18433), .ZN(
        n18437) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18435), .B1(
        n18457), .B2(n18752), .ZN(n18436) );
  OAI211_X1 U21533 ( .C1(n18758), .C2(n18491), .A(n18437), .B(n18436), .ZN(
        P3_U2899) );
  INV_X1 U21534 ( .A(n18794), .ZN(n18438) );
  NAND2_X1 U21535 ( .A1(n18438), .A2(n18509), .ZN(n18521) );
  AOI21_X1 U21536 ( .B1(n18491), .B2(n18521), .A(n18820), .ZN(n18456) );
  AOI22_X1 U21537 ( .A1(n18480), .A2(n18701), .B1(n18700), .B2(n18456), .ZN(
        n18442) );
  NOR2_X1 U21538 ( .A1(n18480), .A2(n18457), .ZN(n18439) );
  AOI221_X1 U21539 ( .B1(n18439), .B2(n18491), .C1(n18579), .C2(n18491), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18440) );
  OAI21_X1 U21540 ( .B1(n18527), .B2(n18440), .A(n18626), .ZN(n18458) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18458), .B1(
        n18706), .B2(n18527), .ZN(n18441) );
  OAI211_X1 U21542 ( .C1(n18451), .C2(n18710), .A(n18442), .B(n18441), .ZN(
        P3_U2900) );
  AOI22_X1 U21543 ( .A1(n18457), .A2(n18713), .B1(n18711), .B2(n18456), .ZN(
        n18444) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18458), .B1(
        n18480), .B2(n18712), .ZN(n18443) );
  OAI211_X1 U21545 ( .C1(n18716), .C2(n18521), .A(n18444), .B(n18443), .ZN(
        P3_U2901) );
  AOI22_X1 U21546 ( .A1(n18480), .A2(n18718), .B1(n18717), .B2(n18456), .ZN(
        n18446) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18458), .B1(
        n18457), .B2(n18719), .ZN(n18445) );
  OAI211_X1 U21548 ( .C1(n18722), .C2(n18521), .A(n18446), .B(n18445), .ZN(
        P3_U2902) );
  AOI22_X1 U21549 ( .A1(n18457), .A2(n18725), .B1(n18723), .B2(n18456), .ZN(
        n18448) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18458), .B1(
        n18480), .B2(n18724), .ZN(n18447) );
  OAI211_X1 U21551 ( .C1(n18728), .C2(n18521), .A(n18448), .B(n18447), .ZN(
        P3_U2903) );
  AOI22_X1 U21552 ( .A1(n18480), .A2(n18657), .B1(n18729), .B2(n18456), .ZN(
        n18450) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18458), .B1(
        n18731), .B2(n18527), .ZN(n18449) );
  OAI211_X1 U21554 ( .C1(n18451), .C2(n18661), .A(n18450), .B(n18449), .ZN(
        P3_U2904) );
  AOI22_X1 U21555 ( .A1(n18480), .A2(n18739), .B1(n18737), .B2(n18456), .ZN(
        n18453) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18458), .B1(
        n18457), .B2(n18738), .ZN(n18452) );
  OAI211_X1 U21557 ( .C1(n18742), .C2(n18521), .A(n18453), .B(n18452), .ZN(
        P3_U2905) );
  AOI22_X1 U21558 ( .A1(n18457), .A2(n18743), .B1(n18744), .B2(n18456), .ZN(
        n18455) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18458), .B1(
        n18480), .B2(n18745), .ZN(n18454) );
  OAI211_X1 U21560 ( .C1(n18748), .C2(n18521), .A(n18455), .B(n18454), .ZN(
        P3_U2906) );
  AOI22_X1 U21561 ( .A1(n18457), .A2(n18754), .B1(n18750), .B2(n18456), .ZN(
        n18460) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18458), .B1(
        n18480), .B2(n18752), .ZN(n18459) );
  OAI211_X1 U21563 ( .C1(n18758), .C2(n18521), .A(n18460), .B(n18459), .ZN(
        P3_U2907) );
  NOR2_X1 U21564 ( .A1(n18553), .A2(n18485), .ZN(n18479) );
  AOI22_X1 U21565 ( .A1(n18480), .A2(n18672), .B1(n18700), .B2(n18479), .ZN(
        n18465) );
  AOI22_X1 U21566 ( .A1(n18705), .A2(n18462), .B1(n18461), .B2(n18509), .ZN(
        n18481) );
  INV_X1 U21567 ( .A(n18463), .ZN(n18556) );
  NOR2_X2 U21568 ( .A1(n18556), .A2(n18485), .ZN(n18548) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18481), .B1(
        n18706), .B2(n18548), .ZN(n18464) );
  OAI211_X1 U21570 ( .C1(n18679), .C2(n18491), .A(n18465), .B(n18464), .ZN(
        P3_U2908) );
  INV_X1 U21571 ( .A(n18548), .ZN(n18484) );
  AOI22_X1 U21572 ( .A1(n18712), .A2(n18505), .B1(n18711), .B2(n18479), .ZN(
        n18467) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18713), .ZN(n18466) );
  OAI211_X1 U21574 ( .C1(n18716), .C2(n18484), .A(n18467), .B(n18466), .ZN(
        P3_U2909) );
  AOI22_X1 U21575 ( .A1(n18480), .A2(n18719), .B1(n18717), .B2(n18479), .ZN(
        n18469) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18481), .B1(
        n18718), .B2(n18505), .ZN(n18468) );
  OAI211_X1 U21577 ( .C1(n18722), .C2(n18484), .A(n18469), .B(n18468), .ZN(
        P3_U2910) );
  AOI22_X1 U21578 ( .A1(n18480), .A2(n18725), .B1(n18723), .B2(n18479), .ZN(
        n18471) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18481), .B1(
        n18724), .B2(n18505), .ZN(n18470) );
  OAI211_X1 U21580 ( .C1(n18728), .C2(n18484), .A(n18471), .B(n18470), .ZN(
        P3_U2911) );
  AOI22_X1 U21581 ( .A1(n18657), .A2(n18505), .B1(n18729), .B2(n18479), .ZN(
        n18473) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18481), .B1(
        n18731), .B2(n18548), .ZN(n18472) );
  OAI211_X1 U21583 ( .C1(n18474), .C2(n18661), .A(n18473), .B(n18472), .ZN(
        P3_U2912) );
  AOI22_X1 U21584 ( .A1(n18739), .A2(n18505), .B1(n18737), .B2(n18479), .ZN(
        n18476) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18738), .ZN(n18475) );
  OAI211_X1 U21586 ( .C1(n18742), .C2(n18484), .A(n18476), .B(n18475), .ZN(
        P3_U2913) );
  AOI22_X1 U21587 ( .A1(n18745), .A2(n18505), .B1(n18744), .B2(n18479), .ZN(
        n18478) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18743), .ZN(n18477) );
  OAI211_X1 U21589 ( .C1(n18748), .C2(n18484), .A(n18478), .B(n18477), .ZN(
        P3_U2914) );
  AOI22_X1 U21590 ( .A1(n18480), .A2(n18754), .B1(n18750), .B2(n18479), .ZN(
        n18483) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18481), .B1(
        n18752), .B2(n18505), .ZN(n18482) );
  OAI211_X1 U21592 ( .C1(n18758), .C2(n18484), .A(n18483), .B(n18482), .ZN(
        P3_U2915) );
  NOR2_X2 U21593 ( .A1(n18486), .A2(n18485), .ZN(n18573) );
  NOR2_X1 U21594 ( .A1(n18548), .A2(n18573), .ZN(n18531) );
  NOR2_X1 U21595 ( .A1(n18820), .A2(n18531), .ZN(n18504) );
  AOI22_X1 U21596 ( .A1(n18701), .A2(n18527), .B1(n18700), .B2(n18504), .ZN(
        n18490) );
  NOR2_X1 U21597 ( .A1(n18505), .A2(n18527), .ZN(n18487) );
  OAI21_X1 U21598 ( .B1(n18487), .B2(n18579), .A(n18531), .ZN(n18488) );
  OAI211_X1 U21599 ( .C1(n18573), .C2(n18920), .A(n18626), .B(n18488), .ZN(
        n18506) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18506), .B1(
        n18706), .B2(n18573), .ZN(n18489) );
  OAI211_X1 U21601 ( .C1(n18710), .C2(n18491), .A(n18490), .B(n18489), .ZN(
        P3_U2916) );
  INV_X1 U21602 ( .A(n18573), .ZN(n18567) );
  AOI22_X1 U21603 ( .A1(n18712), .A2(n18527), .B1(n18711), .B2(n18504), .ZN(
        n18493) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18506), .B1(
        n18713), .B2(n18505), .ZN(n18492) );
  OAI211_X1 U21605 ( .C1(n18716), .C2(n18567), .A(n18493), .B(n18492), .ZN(
        P3_U2917) );
  AOI22_X1 U21606 ( .A1(n18717), .A2(n18504), .B1(n18719), .B2(n18505), .ZN(
        n18495) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18506), .B1(
        n18718), .B2(n18527), .ZN(n18494) );
  OAI211_X1 U21608 ( .C1(n18722), .C2(n18567), .A(n18495), .B(n18494), .ZN(
        P3_U2918) );
  AOI22_X1 U21609 ( .A1(n18723), .A2(n18504), .B1(n18725), .B2(n18505), .ZN(
        n18497) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18506), .B1(
        n18724), .B2(n18527), .ZN(n18496) );
  OAI211_X1 U21611 ( .C1(n18728), .C2(n18567), .A(n18497), .B(n18496), .ZN(
        P3_U2919) );
  AOI22_X1 U21612 ( .A1(n18730), .A2(n18505), .B1(n18729), .B2(n18504), .ZN(
        n18499) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18506), .B1(
        n18731), .B2(n18573), .ZN(n18498) );
  OAI211_X1 U21614 ( .C1(n18736), .C2(n18521), .A(n18499), .B(n18498), .ZN(
        P3_U2920) );
  AOI22_X1 U21615 ( .A1(n18738), .A2(n18505), .B1(n18737), .B2(n18504), .ZN(
        n18501) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18506), .B1(
        n18739), .B2(n18527), .ZN(n18500) );
  OAI211_X1 U21617 ( .C1(n18742), .C2(n18567), .A(n18501), .B(n18500), .ZN(
        P3_U2921) );
  AOI22_X1 U21618 ( .A1(n18745), .A2(n18527), .B1(n18744), .B2(n18504), .ZN(
        n18503) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18506), .B1(
        n18743), .B2(n18505), .ZN(n18502) );
  OAI211_X1 U21620 ( .C1(n18748), .C2(n18567), .A(n18503), .B(n18502), .ZN(
        P3_U2922) );
  AOI22_X1 U21621 ( .A1(n18754), .A2(n18505), .B1(n18750), .B2(n18504), .ZN(
        n18508) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18506), .B1(
        n18752), .B2(n18527), .ZN(n18507) );
  OAI211_X1 U21623 ( .C1(n18758), .C2(n18567), .A(n18508), .B(n18507), .ZN(
        P3_U2923) );
  AOI22_X1 U21624 ( .A1(n18701), .A2(n18548), .B1(n18700), .B2(n18526), .ZN(
        n18512) );
  NAND2_X1 U21625 ( .A1(n18510), .A2(n18509), .ZN(n18528) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18528), .B1(
        n18706), .B2(n18598), .ZN(n18511) );
  OAI211_X1 U21627 ( .C1(n18710), .C2(n18521), .A(n18512), .B(n18511), .ZN(
        P3_U2924) );
  INV_X1 U21628 ( .A(n18598), .ZN(n18592) );
  AOI22_X1 U21629 ( .A1(n18712), .A2(n18548), .B1(n18711), .B2(n18526), .ZN(
        n18514) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18528), .B1(
        n18713), .B2(n18527), .ZN(n18513) );
  OAI211_X1 U21631 ( .C1(n18716), .C2(n18592), .A(n18514), .B(n18513), .ZN(
        P3_U2925) );
  AOI22_X1 U21632 ( .A1(n18717), .A2(n18526), .B1(n18719), .B2(n18527), .ZN(
        n18516) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18528), .B1(
        n18718), .B2(n18548), .ZN(n18515) );
  OAI211_X1 U21634 ( .C1(n18722), .C2(n18592), .A(n18516), .B(n18515), .ZN(
        P3_U2926) );
  AOI22_X1 U21635 ( .A1(n18723), .A2(n18526), .B1(n18725), .B2(n18527), .ZN(
        n18518) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18528), .B1(
        n18724), .B2(n18548), .ZN(n18517) );
  OAI211_X1 U21637 ( .C1(n18728), .C2(n18592), .A(n18518), .B(n18517), .ZN(
        P3_U2927) );
  AOI22_X1 U21638 ( .A1(n18657), .A2(n18548), .B1(n18729), .B2(n18526), .ZN(
        n18520) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18528), .B1(
        n18731), .B2(n18598), .ZN(n18519) );
  OAI211_X1 U21640 ( .C1(n18661), .C2(n18521), .A(n18520), .B(n18519), .ZN(
        P3_U2928) );
  AOI22_X1 U21641 ( .A1(n18738), .A2(n18527), .B1(n18737), .B2(n18526), .ZN(
        n18523) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18528), .B1(
        n18739), .B2(n18548), .ZN(n18522) );
  OAI211_X1 U21643 ( .C1(n18742), .C2(n18592), .A(n18523), .B(n18522), .ZN(
        P3_U2929) );
  AOI22_X1 U21644 ( .A1(n18744), .A2(n18526), .B1(n18743), .B2(n18527), .ZN(
        n18525) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18528), .B1(
        n18745), .B2(n18548), .ZN(n18524) );
  OAI211_X1 U21646 ( .C1(n18748), .C2(n18592), .A(n18525), .B(n18524), .ZN(
        P3_U2930) );
  AOI22_X1 U21647 ( .A1(n18752), .A2(n18548), .B1(n18750), .B2(n18526), .ZN(
        n18530) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18528), .B1(
        n18754), .B2(n18527), .ZN(n18529) );
  OAI211_X1 U21649 ( .C1(n18758), .C2(n18592), .A(n18530), .B(n18529), .ZN(
        P3_U2931) );
  NOR2_X2 U21650 ( .A1(n18794), .A2(n18602), .ZN(n18619) );
  NOR2_X1 U21651 ( .A1(n18598), .A2(n18619), .ZN(n18580) );
  OAI21_X1 U21652 ( .B1(n18531), .B2(n18579), .A(n18580), .ZN(n18532) );
  OAI211_X1 U21653 ( .C1(n18619), .C2(n18920), .A(n18626), .B(n18532), .ZN(
        n18549) );
  NOR2_X1 U21654 ( .A1(n18820), .A2(n18580), .ZN(n18547) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18549), .B1(
        n18700), .B2(n18547), .ZN(n18534) );
  AOI22_X1 U21656 ( .A1(n18672), .A2(n18548), .B1(n18706), .B2(n18619), .ZN(
        n18533) );
  OAI211_X1 U21657 ( .C1(n18679), .C2(n18567), .A(n18534), .B(n18533), .ZN(
        P3_U2932) );
  INV_X1 U21658 ( .A(n18619), .ZN(n18552) );
  AOI22_X1 U21659 ( .A1(n18712), .A2(n18573), .B1(n18711), .B2(n18547), .ZN(
        n18536) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18549), .B1(
        n18713), .B2(n18548), .ZN(n18535) );
  OAI211_X1 U21661 ( .C1(n18716), .C2(n18552), .A(n18536), .B(n18535), .ZN(
        P3_U2933) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18549), .B1(
        n18717), .B2(n18547), .ZN(n18538) );
  AOI22_X1 U21663 ( .A1(n18718), .A2(n18573), .B1(n18719), .B2(n18548), .ZN(
        n18537) );
  OAI211_X1 U21664 ( .C1(n18722), .C2(n18552), .A(n18538), .B(n18537), .ZN(
        P3_U2934) );
  AOI22_X1 U21665 ( .A1(n18724), .A2(n18573), .B1(n18723), .B2(n18547), .ZN(
        n18540) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18549), .B1(
        n18725), .B2(n18548), .ZN(n18539) );
  OAI211_X1 U21667 ( .C1(n18728), .C2(n18552), .A(n18540), .B(n18539), .ZN(
        P3_U2935) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18549), .B1(
        n18729), .B2(n18547), .ZN(n18542) );
  AOI22_X1 U21669 ( .A1(n18730), .A2(n18548), .B1(n18731), .B2(n18619), .ZN(
        n18541) );
  OAI211_X1 U21670 ( .C1(n18736), .C2(n18567), .A(n18542), .B(n18541), .ZN(
        P3_U2936) );
  AOI22_X1 U21671 ( .A1(n18738), .A2(n18548), .B1(n18737), .B2(n18547), .ZN(
        n18544) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18549), .B1(
        n18739), .B2(n18573), .ZN(n18543) );
  OAI211_X1 U21673 ( .C1(n18742), .C2(n18552), .A(n18544), .B(n18543), .ZN(
        P3_U2937) );
  AOI22_X1 U21674 ( .A1(n18745), .A2(n18573), .B1(n18744), .B2(n18547), .ZN(
        n18546) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18549), .B1(
        n18743), .B2(n18548), .ZN(n18545) );
  OAI211_X1 U21676 ( .C1(n18748), .C2(n18552), .A(n18546), .B(n18545), .ZN(
        P3_U2938) );
  AOI22_X1 U21677 ( .A1(n18752), .A2(n18573), .B1(n18750), .B2(n18547), .ZN(
        n18551) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18549), .B1(
        n18754), .B2(n18548), .ZN(n18550) );
  OAI211_X1 U21679 ( .C1(n18758), .C2(n18552), .A(n18551), .B(n18550), .ZN(
        P3_U2939) );
  NOR2_X1 U21680 ( .A1(n18553), .A2(n18602), .ZN(n18572) );
  AOI22_X1 U21681 ( .A1(n18672), .A2(n18573), .B1(n18700), .B2(n18572), .ZN(
        n18558) );
  NOR2_X1 U21682 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18554), .ZN(
        n18555) );
  NOR2_X1 U21683 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18602), .ZN(
        n18603) );
  AOI22_X1 U21684 ( .A1(n18705), .A2(n18555), .B1(n18702), .B2(n18603), .ZN(
        n18574) );
  NOR2_X2 U21685 ( .A1(n18556), .A2(n18602), .ZN(n18644) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18574), .B1(
        n18706), .B2(n18644), .ZN(n18557) );
  OAI211_X1 U21687 ( .C1(n18679), .C2(n18592), .A(n18558), .B(n18557), .ZN(
        P3_U2940) );
  AOI22_X1 U21688 ( .A1(n18713), .A2(n18573), .B1(n18711), .B2(n18572), .ZN(
        n18560) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18574), .B1(
        n18712), .B2(n18598), .ZN(n18559) );
  OAI211_X1 U21690 ( .C1(n18716), .C2(n18637), .A(n18560), .B(n18559), .ZN(
        P3_U2941) );
  AOI22_X1 U21691 ( .A1(n18718), .A2(n18598), .B1(n18717), .B2(n18572), .ZN(
        n18562) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18574), .B1(
        n18719), .B2(n18573), .ZN(n18561) );
  OAI211_X1 U21693 ( .C1(n18722), .C2(n18637), .A(n18562), .B(n18561), .ZN(
        P3_U2942) );
  AOI22_X1 U21694 ( .A1(n18723), .A2(n18572), .B1(n18725), .B2(n18573), .ZN(
        n18564) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18574), .B1(
        n18724), .B2(n18598), .ZN(n18563) );
  OAI211_X1 U21696 ( .C1(n18728), .C2(n18637), .A(n18564), .B(n18563), .ZN(
        P3_U2943) );
  AOI22_X1 U21697 ( .A1(n18657), .A2(n18598), .B1(n18729), .B2(n18572), .ZN(
        n18566) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18574), .B1(
        n18731), .B2(n18644), .ZN(n18565) );
  OAI211_X1 U21699 ( .C1(n18661), .C2(n18567), .A(n18566), .B(n18565), .ZN(
        P3_U2944) );
  AOI22_X1 U21700 ( .A1(n18738), .A2(n18573), .B1(n18737), .B2(n18572), .ZN(
        n18569) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18574), .B1(
        n18739), .B2(n18598), .ZN(n18568) );
  OAI211_X1 U21702 ( .C1(n18742), .C2(n18637), .A(n18569), .B(n18568), .ZN(
        P3_U2945) );
  AOI22_X1 U21703 ( .A1(n18744), .A2(n18572), .B1(n18743), .B2(n18573), .ZN(
        n18571) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18574), .B1(
        n18745), .B2(n18598), .ZN(n18570) );
  OAI211_X1 U21705 ( .C1(n18748), .C2(n18637), .A(n18571), .B(n18570), .ZN(
        P3_U2946) );
  AOI22_X1 U21706 ( .A1(n18752), .A2(n18598), .B1(n18750), .B2(n18572), .ZN(
        n18576) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18574), .B1(
        n18754), .B2(n18573), .ZN(n18575) );
  OAI211_X1 U21708 ( .C1(n18758), .C2(n18637), .A(n18576), .B(n18575), .ZN(
        P3_U2947) );
  NAND2_X1 U21709 ( .A1(n18578), .A2(n18577), .ZN(n18660) );
  AOI21_X1 U21710 ( .B1(n18637), .B2(n18660), .A(n18820), .ZN(n18597) );
  AOI22_X1 U21711 ( .A1(n18701), .A2(n18619), .B1(n18700), .B2(n18597), .ZN(
        n18583) );
  OAI211_X1 U21712 ( .C1(n18580), .C2(n18579), .A(n18637), .B(n18660), .ZN(
        n18581) );
  OAI211_X1 U21713 ( .C1(n18667), .C2(n18920), .A(n18626), .B(n18581), .ZN(
        n18599) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18599), .B1(
        n18706), .B2(n18667), .ZN(n18582) );
  OAI211_X1 U21715 ( .C1(n18710), .C2(n18592), .A(n18583), .B(n18582), .ZN(
        P3_U2948) );
  AOI22_X1 U21716 ( .A1(n18713), .A2(n18598), .B1(n18711), .B2(n18597), .ZN(
        n18585) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18599), .B1(
        n18712), .B2(n18619), .ZN(n18584) );
  OAI211_X1 U21718 ( .C1(n18716), .C2(n18660), .A(n18585), .B(n18584), .ZN(
        P3_U2949) );
  AOI22_X1 U21719 ( .A1(n18718), .A2(n18619), .B1(n18717), .B2(n18597), .ZN(
        n18587) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18599), .B1(
        n18719), .B2(n18598), .ZN(n18586) );
  OAI211_X1 U21721 ( .C1(n18722), .C2(n18660), .A(n18587), .B(n18586), .ZN(
        P3_U2950) );
  AOI22_X1 U21722 ( .A1(n18723), .A2(n18597), .B1(n18725), .B2(n18598), .ZN(
        n18589) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18599), .B1(
        n18724), .B2(n18619), .ZN(n18588) );
  OAI211_X1 U21724 ( .C1(n18728), .C2(n18660), .A(n18589), .B(n18588), .ZN(
        P3_U2951) );
  AOI22_X1 U21725 ( .A1(n18657), .A2(n18619), .B1(n18729), .B2(n18597), .ZN(
        n18591) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18599), .B1(
        n18731), .B2(n18667), .ZN(n18590) );
  OAI211_X1 U21727 ( .C1(n18661), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U2952) );
  AOI22_X1 U21728 ( .A1(n18738), .A2(n18598), .B1(n18737), .B2(n18597), .ZN(
        n18594) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18599), .B1(
        n18739), .B2(n18619), .ZN(n18593) );
  OAI211_X1 U21730 ( .C1(n18742), .C2(n18660), .A(n18594), .B(n18593), .ZN(
        P3_U2953) );
  AOI22_X1 U21731 ( .A1(n18745), .A2(n18619), .B1(n18744), .B2(n18597), .ZN(
        n18596) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18599), .B1(
        n18743), .B2(n18598), .ZN(n18595) );
  OAI211_X1 U21733 ( .C1(n18748), .C2(n18660), .A(n18596), .B(n18595), .ZN(
        P3_U2954) );
  AOI22_X1 U21734 ( .A1(n18754), .A2(n18598), .B1(n18750), .B2(n18597), .ZN(
        n18601) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18599), .B1(
        n18752), .B2(n18619), .ZN(n18600) );
  OAI211_X1 U21736 ( .C1(n18758), .C2(n18660), .A(n18601), .B(n18600), .ZN(
        P3_U2955) );
  NOR2_X1 U21737 ( .A1(n18793), .A2(n18602), .ZN(n18647) );
  AND2_X1 U21738 ( .A1(n18699), .A2(n18647), .ZN(n18618) );
  AOI22_X1 U21739 ( .A1(n18672), .A2(n18619), .B1(n18700), .B2(n18618), .ZN(
        n18605) );
  AOI22_X1 U21740 ( .A1(n18705), .A2(n18603), .B1(n18702), .B2(n18647), .ZN(
        n18620) );
  NAND2_X1 U21741 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18647), .ZN(
        n18650) );
  INV_X1 U21742 ( .A(n18650), .ZN(n18694) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18620), .B1(
        n18706), .B2(n18694), .ZN(n18604) );
  OAI211_X1 U21744 ( .C1(n18679), .C2(n18637), .A(n18605), .B(n18604), .ZN(
        P3_U2956) );
  AOI22_X1 U21745 ( .A1(n18713), .A2(n18619), .B1(n18711), .B2(n18618), .ZN(
        n18607) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18620), .B1(
        n18712), .B2(n18644), .ZN(n18606) );
  OAI211_X1 U21747 ( .C1(n18716), .C2(n18650), .A(n18607), .B(n18606), .ZN(
        P3_U2957) );
  AOI22_X1 U21748 ( .A1(n18717), .A2(n18618), .B1(n18719), .B2(n18619), .ZN(
        n18609) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18620), .B1(
        n18718), .B2(n18644), .ZN(n18608) );
  OAI211_X1 U21750 ( .C1(n18722), .C2(n18650), .A(n18609), .B(n18608), .ZN(
        P3_U2958) );
  AOI22_X1 U21751 ( .A1(n18723), .A2(n18618), .B1(n18725), .B2(n18619), .ZN(
        n18611) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18620), .B1(
        n18724), .B2(n18644), .ZN(n18610) );
  OAI211_X1 U21753 ( .C1(n18728), .C2(n18650), .A(n18611), .B(n18610), .ZN(
        P3_U2959) );
  AOI22_X1 U21754 ( .A1(n18730), .A2(n18619), .B1(n18729), .B2(n18618), .ZN(
        n18613) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18620), .B1(
        n18731), .B2(n18694), .ZN(n18612) );
  OAI211_X1 U21756 ( .C1(n18736), .C2(n18637), .A(n18613), .B(n18612), .ZN(
        P3_U2960) );
  AOI22_X1 U21757 ( .A1(n18738), .A2(n18619), .B1(n18737), .B2(n18618), .ZN(
        n18615) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18620), .B1(
        n18739), .B2(n18644), .ZN(n18614) );
  OAI211_X1 U21759 ( .C1(n18742), .C2(n18650), .A(n18615), .B(n18614), .ZN(
        P3_U2961) );
  AOI22_X1 U21760 ( .A1(n18744), .A2(n18618), .B1(n18743), .B2(n18619), .ZN(
        n18617) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18620), .B1(
        n18745), .B2(n18644), .ZN(n18616) );
  OAI211_X1 U21762 ( .C1(n18748), .C2(n18650), .A(n18617), .B(n18616), .ZN(
        P3_U2962) );
  AOI22_X1 U21763 ( .A1(n18754), .A2(n18619), .B1(n18750), .B2(n18618), .ZN(
        n18622) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18620), .B1(
        n18752), .B2(n18644), .ZN(n18621) );
  OAI211_X1 U21765 ( .C1(n18758), .C2(n18650), .A(n18622), .B(n18621), .ZN(
        P3_U2963) );
  NAND2_X1 U21766 ( .A1(n18791), .A2(n18704), .ZN(n18709) );
  INV_X1 U21767 ( .A(n18709), .ZN(n18753) );
  NOR2_X1 U21768 ( .A1(n18694), .A2(n18753), .ZN(n18675) );
  NOR2_X1 U21769 ( .A1(n18820), .A2(n18675), .ZN(n18642) );
  AOI22_X1 U21770 ( .A1(n18672), .A2(n18644), .B1(n18700), .B2(n18642), .ZN(
        n18628) );
  OAI21_X1 U21771 ( .B1(n18624), .B2(n18623), .A(n18675), .ZN(n18625) );
  OAI211_X1 U21772 ( .C1(n18753), .C2(n18920), .A(n18626), .B(n18625), .ZN(
        n18643) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18643), .B1(
        n18706), .B2(n18753), .ZN(n18627) );
  OAI211_X1 U21774 ( .C1(n18679), .C2(n18660), .A(n18628), .B(n18627), .ZN(
        P3_U2964) );
  AOI22_X1 U21775 ( .A1(n18712), .A2(n18667), .B1(n18711), .B2(n18642), .ZN(
        n18630) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18643), .B1(
        n18713), .B2(n18644), .ZN(n18629) );
  OAI211_X1 U21777 ( .C1(n18716), .C2(n18709), .A(n18630), .B(n18629), .ZN(
        P3_U2965) );
  AOI22_X1 U21778 ( .A1(n18717), .A2(n18642), .B1(n18719), .B2(n18644), .ZN(
        n18632) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18643), .B1(
        n18718), .B2(n18667), .ZN(n18631) );
  OAI211_X1 U21780 ( .C1(n18722), .C2(n18709), .A(n18632), .B(n18631), .ZN(
        P3_U2966) );
  AOI22_X1 U21781 ( .A1(n18723), .A2(n18642), .B1(n18725), .B2(n18644), .ZN(
        n18634) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18643), .B1(
        n18724), .B2(n18667), .ZN(n18633) );
  OAI211_X1 U21783 ( .C1(n18728), .C2(n18709), .A(n18634), .B(n18633), .ZN(
        P3_U2967) );
  AOI22_X1 U21784 ( .A1(n18657), .A2(n18667), .B1(n18729), .B2(n18642), .ZN(
        n18636) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18643), .B1(
        n18731), .B2(n18753), .ZN(n18635) );
  OAI211_X1 U21786 ( .C1(n18661), .C2(n18637), .A(n18636), .B(n18635), .ZN(
        P3_U2968) );
  AOI22_X1 U21787 ( .A1(n18738), .A2(n18644), .B1(n18737), .B2(n18642), .ZN(
        n18639) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18643), .B1(
        n18739), .B2(n18667), .ZN(n18638) );
  OAI211_X1 U21789 ( .C1(n18742), .C2(n18709), .A(n18639), .B(n18638), .ZN(
        P3_U2969) );
  AOI22_X1 U21790 ( .A1(n18744), .A2(n18642), .B1(n18743), .B2(n18644), .ZN(
        n18641) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18643), .B1(
        n18745), .B2(n18667), .ZN(n18640) );
  OAI211_X1 U21792 ( .C1(n18748), .C2(n18709), .A(n18641), .B(n18640), .ZN(
        P3_U2970) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18643), .B1(
        n18750), .B2(n18642), .ZN(n18646) );
  AOI22_X1 U21794 ( .A1(n18752), .A2(n18667), .B1(n18754), .B2(n18644), .ZN(
        n18645) );
  OAI211_X1 U21795 ( .C1(n18758), .C2(n18709), .A(n18646), .B(n18645), .ZN(
        P3_U2971) );
  AND2_X1 U21796 ( .A1(n18699), .A2(n18704), .ZN(n18666) );
  AOI22_X1 U21797 ( .A1(n18672), .A2(n18667), .B1(n18700), .B2(n18666), .ZN(
        n18649) );
  AOI22_X1 U21798 ( .A1(n18705), .A2(n18647), .B1(n18704), .B2(n18702), .ZN(
        n18668) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18668), .B1(
        n18706), .B2(n18751), .ZN(n18648) );
  OAI211_X1 U21800 ( .C1(n18679), .C2(n18650), .A(n18649), .B(n18648), .ZN(
        P3_U2972) );
  AOI22_X1 U21801 ( .A1(n18712), .A2(n18694), .B1(n18711), .B2(n18666), .ZN(
        n18652) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18668), .B1(
        n18713), .B2(n18667), .ZN(n18651) );
  OAI211_X1 U21803 ( .C1(n18716), .C2(n18735), .A(n18652), .B(n18651), .ZN(
        P3_U2973) );
  AOI22_X1 U21804 ( .A1(n18717), .A2(n18666), .B1(n18719), .B2(n18667), .ZN(
        n18654) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18668), .B1(
        n18718), .B2(n18694), .ZN(n18653) );
  OAI211_X1 U21806 ( .C1(n18722), .C2(n18735), .A(n18654), .B(n18653), .ZN(
        P3_U2974) );
  AOI22_X1 U21807 ( .A1(n18723), .A2(n18666), .B1(n18725), .B2(n18667), .ZN(
        n18656) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18668), .B1(
        n18724), .B2(n18694), .ZN(n18655) );
  OAI211_X1 U21809 ( .C1(n18728), .C2(n18735), .A(n18656), .B(n18655), .ZN(
        P3_U2975) );
  AOI22_X1 U21810 ( .A1(n18657), .A2(n18694), .B1(n18729), .B2(n18666), .ZN(
        n18659) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18668), .B1(
        n18731), .B2(n18751), .ZN(n18658) );
  OAI211_X1 U21812 ( .C1(n18661), .C2(n18660), .A(n18659), .B(n18658), .ZN(
        P3_U2976) );
  AOI22_X1 U21813 ( .A1(n18738), .A2(n18667), .B1(n18737), .B2(n18666), .ZN(
        n18663) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18668), .B1(
        n18739), .B2(n18694), .ZN(n18662) );
  OAI211_X1 U21815 ( .C1(n18742), .C2(n18735), .A(n18663), .B(n18662), .ZN(
        P3_U2977) );
  AOI22_X1 U21816 ( .A1(n18744), .A2(n18666), .B1(n18743), .B2(n18667), .ZN(
        n18665) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18668), .B1(
        n18745), .B2(n18694), .ZN(n18664) );
  OAI211_X1 U21818 ( .C1(n18748), .C2(n18735), .A(n18665), .B(n18664), .ZN(
        P3_U2978) );
  AOI22_X1 U21819 ( .A1(n18754), .A2(n18667), .B1(n18750), .B2(n18666), .ZN(
        n18670) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18668), .B1(
        n18752), .B2(n18694), .ZN(n18669) );
  OAI211_X1 U21821 ( .C1(n18758), .C2(n18735), .A(n18670), .B(n18669), .ZN(
        P3_U2979) );
  INV_X1 U21822 ( .A(n18671), .ZN(n18673) );
  NOR2_X1 U21823 ( .A1(n18820), .A2(n18673), .ZN(n18693) );
  AOI22_X1 U21824 ( .A1(n18672), .A2(n18694), .B1(n18700), .B2(n18693), .ZN(
        n18678) );
  OAI22_X1 U21825 ( .A1(n18675), .A2(n18364), .B1(n18674), .B2(n18673), .ZN(
        n18676) );
  OAI21_X1 U21826 ( .B1(n18686), .B2(n18920), .A(n18676), .ZN(n18695) );
  AOI22_X1 U21827 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18695), .B1(
        n18706), .B2(n18686), .ZN(n18677) );
  OAI211_X1 U21828 ( .C1(n18679), .C2(n18709), .A(n18678), .B(n18677), .ZN(
        P3_U2980) );
  AOI22_X1 U21829 ( .A1(n18712), .A2(n18753), .B1(n18711), .B2(n18693), .ZN(
        n18681) );
  AOI22_X1 U21830 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18695), .B1(
        n18713), .B2(n18694), .ZN(n18680) );
  OAI211_X1 U21831 ( .C1(n18716), .C2(n18698), .A(n18681), .B(n18680), .ZN(
        P3_U2981) );
  AOI22_X1 U21832 ( .A1(n18718), .A2(n18753), .B1(n18717), .B2(n18693), .ZN(
        n18683) );
  AOI22_X1 U21833 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18695), .B1(
        n18719), .B2(n18694), .ZN(n18682) );
  OAI211_X1 U21834 ( .C1(n18722), .C2(n18698), .A(n18683), .B(n18682), .ZN(
        P3_U2982) );
  AOI22_X1 U21835 ( .A1(n18724), .A2(n18753), .B1(n18723), .B2(n18693), .ZN(
        n18685) );
  AOI22_X1 U21836 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18695), .B1(
        n18725), .B2(n18694), .ZN(n18684) );
  OAI211_X1 U21837 ( .C1(n18728), .C2(n18698), .A(n18685), .B(n18684), .ZN(
        P3_U2983) );
  AOI22_X1 U21838 ( .A1(n18730), .A2(n18694), .B1(n18729), .B2(n18693), .ZN(
        n18688) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18695), .B1(
        n18731), .B2(n18686), .ZN(n18687) );
  OAI211_X1 U21840 ( .C1(n18736), .C2(n18709), .A(n18688), .B(n18687), .ZN(
        P3_U2984) );
  AOI22_X1 U21841 ( .A1(n18739), .A2(n18753), .B1(n18737), .B2(n18693), .ZN(
        n18690) );
  AOI22_X1 U21842 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18695), .B1(
        n18738), .B2(n18694), .ZN(n18689) );
  OAI211_X1 U21843 ( .C1(n18742), .C2(n18698), .A(n18690), .B(n18689), .ZN(
        P3_U2985) );
  AOI22_X1 U21844 ( .A1(n18745), .A2(n18753), .B1(n18744), .B2(n18693), .ZN(
        n18692) );
  AOI22_X1 U21845 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18695), .B1(
        n18743), .B2(n18694), .ZN(n18691) );
  OAI211_X1 U21846 ( .C1(n18748), .C2(n18698), .A(n18692), .B(n18691), .ZN(
        P3_U2986) );
  AOI22_X1 U21847 ( .A1(n18752), .A2(n18753), .B1(n18750), .B2(n18693), .ZN(
        n18697) );
  AOI22_X1 U21848 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18695), .B1(
        n18754), .B2(n18694), .ZN(n18696) );
  OAI211_X1 U21849 ( .C1(n18758), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        P3_U2987) );
  AND2_X1 U21850 ( .A1(n18699), .A2(n18703), .ZN(n18749) );
  AOI22_X1 U21851 ( .A1(n18701), .A2(n18751), .B1(n18700), .B2(n18749), .ZN(
        n18708) );
  AOI22_X1 U21852 ( .A1(n18705), .A2(n18704), .B1(n18703), .B2(n18702), .ZN(
        n18755) );
  AOI22_X1 U21853 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18755), .B1(
        n18732), .B2(n18706), .ZN(n18707) );
  OAI211_X1 U21854 ( .C1(n18710), .C2(n18709), .A(n18708), .B(n18707), .ZN(
        P3_U2988) );
  AOI22_X1 U21855 ( .A1(n18712), .A2(n18751), .B1(n18711), .B2(n18749), .ZN(
        n18715) );
  AOI22_X1 U21856 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18755), .B1(
        n18713), .B2(n18753), .ZN(n18714) );
  OAI211_X1 U21857 ( .C1(n18759), .C2(n18716), .A(n18715), .B(n18714), .ZN(
        P3_U2989) );
  AOI22_X1 U21858 ( .A1(n18718), .A2(n18751), .B1(n18717), .B2(n18749), .ZN(
        n18721) );
  AOI22_X1 U21859 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18755), .B1(
        n18719), .B2(n18753), .ZN(n18720) );
  OAI211_X1 U21860 ( .C1(n18759), .C2(n18722), .A(n18721), .B(n18720), .ZN(
        P3_U2990) );
  AOI22_X1 U21861 ( .A1(n18724), .A2(n18751), .B1(n18723), .B2(n18749), .ZN(
        n18727) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18755), .B1(
        n18725), .B2(n18753), .ZN(n18726) );
  OAI211_X1 U21863 ( .C1(n18759), .C2(n18728), .A(n18727), .B(n18726), .ZN(
        P3_U2991) );
  AOI22_X1 U21864 ( .A1(n18730), .A2(n18753), .B1(n18729), .B2(n18749), .ZN(
        n18734) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18755), .B1(
        n18732), .B2(n18731), .ZN(n18733) );
  OAI211_X1 U21866 ( .C1(n18736), .C2(n18735), .A(n18734), .B(n18733), .ZN(
        P3_U2992) );
  AOI22_X1 U21867 ( .A1(n18738), .A2(n18753), .B1(n18737), .B2(n18749), .ZN(
        n18741) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18755), .B1(
        n18739), .B2(n18751), .ZN(n18740) );
  OAI211_X1 U21869 ( .C1(n18759), .C2(n18742), .A(n18741), .B(n18740), .ZN(
        P3_U2993) );
  AOI22_X1 U21870 ( .A1(n18744), .A2(n18749), .B1(n18743), .B2(n18753), .ZN(
        n18747) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18755), .B1(
        n18745), .B2(n18751), .ZN(n18746) );
  OAI211_X1 U21872 ( .C1(n18759), .C2(n18748), .A(n18747), .B(n18746), .ZN(
        P3_U2994) );
  AOI22_X1 U21873 ( .A1(n18752), .A2(n18751), .B1(n18750), .B2(n18749), .ZN(
        n18757) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18755), .B1(
        n18754), .B2(n18753), .ZN(n18756) );
  OAI211_X1 U21875 ( .C1(n18759), .C2(n18758), .A(n18757), .B(n18756), .ZN(
        P3_U2995) );
  NAND2_X1 U21876 ( .A1(n18761), .A2(n18760), .ZN(n18762) );
  AOI22_X1 U21877 ( .A1(n18784), .A2(n18958), .B1(n18763), .B2(n18762), .ZN(
        n18961) );
  AOI221_X1 U21878 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18765), .C1(
        P3_MORE_REG_SCAN_IN), .C2(n18765), .A(n18764), .ZN(n18766) );
  OAI211_X1 U21879 ( .C1(n18767), .C2(n18785), .A(n18961), .B(n18766), .ZN(
        n18807) );
  AOI21_X1 U21880 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18786), .A(
        n18768), .ZN(n18789) );
  OAI22_X1 U21881 ( .A1(n18776), .A2(n18770), .B1(n18769), .B2(n18789), .ZN(
        n18771) );
  INV_X1 U21882 ( .A(n18771), .ZN(n18778) );
  AOI21_X1 U21883 ( .B1(n18774), .B2(n18773), .A(n18772), .ZN(n18779) );
  AOI222_X1 U21884 ( .A1(n18781), .A2(n18779), .B1(n18781), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C1(n18779), .C2(n18788), .ZN(
        n18775) );
  NOR2_X1 U21885 ( .A1(n18776), .A2(n18775), .ZN(n18777) );
  MUX2_X1 U21886 ( .A(n18778), .B(n18777), .S(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n18922) );
  INV_X1 U21887 ( .A(n18785), .ZN(n18796) );
  MUX2_X1 U21888 ( .A(n18922), .B(n18925), .S(n18796), .Z(n18805) );
  NOR3_X1 U21889 ( .A1(n18780), .A2(n18779), .A3(n12415), .ZN(n18783) );
  AOI211_X1 U21890 ( .C1(n12415), .C2(n12414), .A(n18781), .B(n18789), .ZN(
        n18782) );
  AOI211_X1 U21891 ( .C1(n18784), .C2(n18929), .A(n18783), .B(n18782), .ZN(
        n18931) );
  AOI22_X1 U21892 ( .A1(n18796), .A2(n12415), .B1(n18931), .B2(n18785), .ZN(
        n18800) );
  NOR2_X1 U21893 ( .A1(n18787), .A2(n18786), .ZN(n18790) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18788), .B1(
        n18790), .B2(n12413), .ZN(n18942) );
  OAI22_X1 U21895 ( .A1(n18790), .A2(n18934), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18789), .ZN(n18939) );
  OR3_X1 U21896 ( .A1(n18942), .A2(n18793), .A3(n18791), .ZN(n18792) );
  AOI22_X1 U21897 ( .A1(n18942), .A2(n18793), .B1(n18939), .B2(n18792), .ZN(
        n18795) );
  OAI21_X1 U21898 ( .B1(n18796), .B2(n18795), .A(n18794), .ZN(n18799) );
  AND2_X1 U21899 ( .A1(n18800), .A2(n18799), .ZN(n18797) );
  OAI221_X1 U21900 ( .B1(n18800), .B2(n18799), .C1(n18798), .C2(n18797), .A(
        n18802), .ZN(n18804) );
  AOI21_X1 U21901 ( .B1(n18802), .B2(n18801), .A(n18800), .ZN(n18803) );
  AOI222_X1 U21902 ( .A1(n18805), .A2(n18804), .B1(n18805), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18804), .C2(n18803), .ZN(
        n18806) );
  NOR4_X1 U21903 ( .A1(n18959), .A2(n18808), .A3(n18807), .A4(n18806), .ZN(
        n18818) );
  NOR2_X1 U21904 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18975) );
  AOI22_X1 U21905 ( .A1(n18941), .A2(n18975), .B1(n18836), .B2(n17576), .ZN(
        n18809) );
  INV_X1 U21906 ( .A(n18809), .ZN(n18814) );
  OAI211_X1 U21907 ( .C1(n18811), .C2(n18810), .A(n18967), .B(n18818), .ZN(
        n18919) );
  OAI21_X1 U21908 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18973), .A(n18919), 
        .ZN(n18821) );
  NOR2_X1 U21909 ( .A1(n18812), .A2(n18821), .ZN(n18813) );
  MUX2_X1 U21910 ( .A(n18814), .B(n18813), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18816) );
  OAI211_X1 U21911 ( .C1(n18818), .C2(n18817), .A(n18816), .B(n18815), .ZN(
        P3_U2996) );
  NAND2_X1 U21912 ( .A1(n18836), .A2(n17576), .ZN(n18824) );
  NAND4_X1 U21913 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18836), .A4(n18819), .ZN(n18826) );
  OR3_X1 U21914 ( .A1(n18822), .A2(n18821), .A3(n18820), .ZN(n18823) );
  NAND4_X1 U21915 ( .A1(n18825), .A2(n18824), .A3(n18826), .A4(n18823), .ZN(
        P3_U2997) );
  INV_X1 U21916 ( .A(n18826), .ZN(n18828) );
  INV_X1 U21917 ( .A(n18918), .ZN(n18827) );
  NOR4_X1 U21918 ( .A1(n18975), .A2(n18829), .A3(n18828), .A4(n18827), .ZN(
        P3_U2998) );
  AND2_X1 U21919 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18915), .ZN(
        P3_U2999) );
  AND2_X1 U21920 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18915), .ZN(
        P3_U3000) );
  AND2_X1 U21921 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18915), .ZN(
        P3_U3001) );
  AND2_X1 U21922 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18915), .ZN(
        P3_U3002) );
  AND2_X1 U21923 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18915), .ZN(
        P3_U3003) );
  AND2_X1 U21924 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18915), .ZN(
        P3_U3004) );
  AND2_X1 U21925 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18915), .ZN(
        P3_U3005) );
  AND2_X1 U21926 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18915), .ZN(
        P3_U3006) );
  AND2_X1 U21927 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18915), .ZN(
        P3_U3007) );
  AND2_X1 U21928 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18915), .ZN(
        P3_U3008) );
  INV_X1 U21929 ( .A(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21119) );
  NOR2_X1 U21930 ( .A1(n21119), .A2(n18917), .ZN(P3_U3009) );
  AND2_X1 U21931 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18915), .ZN(
        P3_U3010) );
  AND2_X1 U21932 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18915), .ZN(
        P3_U3011) );
  AND2_X1 U21933 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18915), .ZN(
        P3_U3012) );
  AND2_X1 U21934 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18915), .ZN(
        P3_U3013) );
  AND2_X1 U21935 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18915), .ZN(
        P3_U3014) );
  AND2_X1 U21936 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18915), .ZN(
        P3_U3015) );
  AND2_X1 U21937 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18915), .ZN(
        P3_U3016) );
  AND2_X1 U21938 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18915), .ZN(
        P3_U3017) );
  AND2_X1 U21939 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18915), .ZN(
        P3_U3018) );
  INV_X1 U21940 ( .A(P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21251) );
  NOR2_X1 U21941 ( .A1(n21251), .A2(n18917), .ZN(P3_U3019) );
  AND2_X1 U21942 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18915), .ZN(
        P3_U3020) );
  AND2_X1 U21943 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18915), .ZN(P3_U3021) );
  AND2_X1 U21944 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18915), .ZN(P3_U3022) );
  AND2_X1 U21945 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18915), .ZN(P3_U3023) );
  AND2_X1 U21946 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18915), .ZN(P3_U3024) );
  AND2_X1 U21947 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18915), .ZN(P3_U3025) );
  AND2_X1 U21948 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18915), .ZN(P3_U3026) );
  AND2_X1 U21949 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18915), .ZN(P3_U3027) );
  AND2_X1 U21950 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18915), .ZN(P3_U3028) );
  OAI21_X1 U21951 ( .B1(n18830), .B2(n20866), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18831) );
  AOI22_X1 U21952 ( .A1(n18845), .A2(n18847), .B1(n18981), .B2(n18831), .ZN(
        n18832) );
  NAND3_X1 U21953 ( .A1(NA), .A2(n18845), .A3(n18838), .ZN(n18839) );
  OAI211_X1 U21954 ( .C1(n18833), .C2(n18973), .A(n18832), .B(n18839), .ZN(
        P3_U3029) );
  AOI21_X1 U21955 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18834) );
  AOI21_X1 U21956 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18834), .ZN(
        n18835) );
  AOI22_X1 U21957 ( .A1(n18836), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18835), .ZN(n18837) );
  NAND2_X1 U21958 ( .A1(n18837), .A2(n18970), .ZN(P3_U3030) );
  NOR2_X1 U21959 ( .A1(n18973), .A2(n18838), .ZN(n18840) );
  AOI21_X1 U21960 ( .B1(n18845), .B2(n18839), .A(n18840), .ZN(n18846) );
  NOR2_X1 U21961 ( .A1(n18847), .A2(n20866), .ZN(n18843) );
  INV_X1 U21962 ( .A(n18840), .ZN(n18841) );
  OAI22_X1 U21963 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18841), .ZN(n18842) );
  OAI22_X1 U21964 ( .A1(n18843), .A2(n18842), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18844) );
  OAI22_X1 U21965 ( .A1(n18846), .A2(n18847), .B1(n18845), .B2(n18844), .ZN(
        P3_U3031) );
  INV_X1 U21966 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18849) );
  OAI222_X1 U21967 ( .A1(n18849), .A2(n18908), .B1(n18848), .B2(n18957), .C1(
        n18850), .C2(n18905), .ZN(P3_U3032) );
  OAI222_X1 U21968 ( .A1(n18905), .A2(n18852), .B1(n18851), .B2(n18957), .C1(
        n18850), .C2(n18908), .ZN(P3_U3033) );
  OAI222_X1 U21969 ( .A1(n18905), .A2(n18854), .B1(n18853), .B2(n18957), .C1(
        n18852), .C2(n18908), .ZN(P3_U3034) );
  OAI222_X1 U21970 ( .A1(n18905), .A2(n18856), .B1(n18855), .B2(n18957), .C1(
        n18854), .C2(n18908), .ZN(P3_U3035) );
  OAI222_X1 U21971 ( .A1(n18905), .A2(n18858), .B1(n18857), .B2(n18957), .C1(
        n18856), .C2(n18908), .ZN(P3_U3036) );
  OAI222_X1 U21972 ( .A1(n18905), .A2(n18860), .B1(n18859), .B2(n18957), .C1(
        n18858), .C2(n18908), .ZN(P3_U3037) );
  OAI222_X1 U21973 ( .A1(n18905), .A2(n18863), .B1(n18861), .B2(n18957), .C1(
        n18860), .C2(n18908), .ZN(P3_U3038) );
  OAI222_X1 U21974 ( .A1(n18863), .A2(n18908), .B1(n18862), .B2(n18957), .C1(
        n18864), .C2(n18905), .ZN(P3_U3039) );
  OAI222_X1 U21975 ( .A1(n18905), .A2(n18866), .B1(n18865), .B2(n18957), .C1(
        n18864), .C2(n18908), .ZN(P3_U3040) );
  OAI222_X1 U21976 ( .A1(n18905), .A2(n18868), .B1(n18867), .B2(n18957), .C1(
        n18866), .C2(n18908), .ZN(P3_U3041) );
  INV_X1 U21977 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18870) );
  OAI222_X1 U21978 ( .A1(n18905), .A2(n18870), .B1(n18869), .B2(n18957), .C1(
        n18868), .C2(n18908), .ZN(P3_U3042) );
  OAI222_X1 U21979 ( .A1(n18905), .A2(n18872), .B1(n18871), .B2(n18957), .C1(
        n18870), .C2(n18908), .ZN(P3_U3043) );
  OAI222_X1 U21980 ( .A1(n18905), .A2(n18875), .B1(n18873), .B2(n18980), .C1(
        n18872), .C2(n18908), .ZN(P3_U3044) );
  OAI222_X1 U21981 ( .A1(n18875), .A2(n18908), .B1(n18874), .B2(n18980), .C1(
        n18876), .C2(n18905), .ZN(P3_U3045) );
  INV_X1 U21982 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18878) );
  OAI222_X1 U21983 ( .A1(n18905), .A2(n18878), .B1(n18877), .B2(n18980), .C1(
        n18876), .C2(n18908), .ZN(P3_U3046) );
  OAI222_X1 U21984 ( .A1(n18905), .A2(n18881), .B1(n18879), .B2(n18980), .C1(
        n18878), .C2(n18908), .ZN(P3_U3047) );
  OAI222_X1 U21985 ( .A1(n18881), .A2(n18908), .B1(n18880), .B2(n18980), .C1(
        n18882), .C2(n18905), .ZN(P3_U3048) );
  INV_X1 U21986 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18884) );
  OAI222_X1 U21987 ( .A1(n18905), .A2(n18884), .B1(n18883), .B2(n18980), .C1(
        n18882), .C2(n18908), .ZN(P3_U3049) );
  OAI222_X1 U21988 ( .A1(n18905), .A2(n18886), .B1(n18885), .B2(n18980), .C1(
        n18884), .C2(n18908), .ZN(P3_U3050) );
  OAI222_X1 U21989 ( .A1(n18905), .A2(n18889), .B1(n18887), .B2(n18980), .C1(
        n18886), .C2(n18908), .ZN(P3_U3051) );
  OAI222_X1 U21990 ( .A1(n18889), .A2(n18908), .B1(n18888), .B2(n18980), .C1(
        n18890), .C2(n18905), .ZN(P3_U3052) );
  OAI222_X1 U21991 ( .A1(n18905), .A2(n18893), .B1(n18891), .B2(n18980), .C1(
        n18890), .C2(n18908), .ZN(P3_U3053) );
  OAI222_X1 U21992 ( .A1(n18893), .A2(n18908), .B1(n18892), .B2(n18980), .C1(
        n18894), .C2(n18905), .ZN(P3_U3054) );
  OAI222_X1 U21993 ( .A1(n18905), .A2(n18896), .B1(n18895), .B2(n18980), .C1(
        n18894), .C2(n18908), .ZN(P3_U3055) );
  OAI222_X1 U21994 ( .A1(n18905), .A2(n18898), .B1(n18897), .B2(n18957), .C1(
        n18896), .C2(n18908), .ZN(P3_U3056) );
  OAI222_X1 U21995 ( .A1(n18905), .A2(n21163), .B1(n18899), .B2(n18957), .C1(
        n18898), .C2(n18908), .ZN(P3_U3057) );
  OAI222_X1 U21996 ( .A1(n18905), .A2(n18901), .B1(n18900), .B2(n18957), .C1(
        n21163), .C2(n18908), .ZN(P3_U3058) );
  OAI222_X1 U21997 ( .A1(n18905), .A2(n18903), .B1(n18902), .B2(n18957), .C1(
        n18901), .C2(n18908), .ZN(P3_U3059) );
  OAI222_X1 U21998 ( .A1(n18905), .A2(n18907), .B1(n18904), .B2(n18957), .C1(
        n18903), .C2(n18908), .ZN(P3_U3060) );
  OAI222_X1 U21999 ( .A1(n18908), .A2(n18907), .B1(n18906), .B2(n18957), .C1(
        n21196), .C2(n18905), .ZN(P3_U3061) );
  INV_X1 U22000 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18909) );
  INV_X1 U22001 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n21236) );
  AOI22_X1 U22002 ( .A1(n18980), .A2(n18909), .B1(n21236), .B2(n18981), .ZN(
        P3_U3274) );
  INV_X1 U22003 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21084) );
  INV_X1 U22004 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18910) );
  AOI22_X1 U22005 ( .A1(n18980), .A2(n21084), .B1(n18910), .B2(n18981), .ZN(
        P3_U3275) );
  INV_X1 U22006 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18911) );
  AOI22_X1 U22007 ( .A1(n18980), .A2(n18912), .B1(n18911), .B2(n18981), .ZN(
        P3_U3276) );
  INV_X1 U22008 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18952) );
  INV_X1 U22009 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18913) );
  AOI22_X1 U22010 ( .A1(n18980), .A2(n18952), .B1(n18913), .B2(n18981), .ZN(
        P3_U3277) );
  INV_X1 U22011 ( .A(n18916), .ZN(n18914) );
  AOI21_X1 U22012 ( .B1(n18915), .B2(n21254), .A(n18914), .ZN(P3_U3280) );
  OAI21_X1 U22013 ( .B1(n18917), .B2(n21102), .A(n18916), .ZN(P3_U3281) );
  OAI221_X1 U22014 ( .B1(n18920), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18920), 
        .C2(n18919), .A(n18918), .ZN(P3_U3282) );
  OAI22_X1 U22015 ( .A1(n18983), .A2(n18922), .B1(n18930), .B2(n18921), .ZN(
        n18923) );
  INV_X1 U22016 ( .A(n18923), .ZN(n18924) );
  AOI22_X1 U22017 ( .A1(n18947), .A2(n18925), .B1(n18924), .B2(n18945), .ZN(
        P3_U3285) );
  AOI22_X1 U22018 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18927), .B2(n18926), .ZN(
        n18935) );
  NOR2_X1 U22019 ( .A1(n18928), .A2(n18944), .ZN(n18936) );
  OAI22_X1 U22020 ( .A1(n18931), .A2(n18983), .B1(n18930), .B2(n18929), .ZN(
        n18932) );
  AOI21_X1 U22021 ( .B1(n18935), .B2(n18936), .A(n18932), .ZN(n18933) );
  AOI22_X1 U22022 ( .A1(n18947), .A2(n12415), .B1(n18933), .B2(n18945), .ZN(
        P3_U3288) );
  INV_X1 U22023 ( .A(n18934), .ZN(n18938) );
  INV_X1 U22024 ( .A(n18935), .ZN(n18937) );
  AOI222_X1 U22025 ( .A1(n18939), .A2(n18943), .B1(n18941), .B2(n18938), .C1(
        n18937), .C2(n18936), .ZN(n18940) );
  AOI22_X1 U22026 ( .A1(n18947), .A2(n12414), .B1(n18940), .B2(n18945), .ZN(
        P3_U3289) );
  AOI222_X1 U22027 ( .A1(n18944), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18943), 
        .B2(n18942), .C1(n12413), .C2(n18941), .ZN(n18946) );
  AOI22_X1 U22028 ( .A1(n18947), .A2(n12413), .B1(n18946), .B2(n18945), .ZN(
        P3_U3290) );
  NAND2_X1 U22029 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18951) );
  INV_X1 U22030 ( .A(n18955), .ZN(n18948) );
  AOI211_X1 U22031 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18948), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18949) );
  AOI21_X1 U22032 ( .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n18953), .A(n18949), 
        .ZN(n18950) );
  OAI21_X1 U22033 ( .B1(n18951), .B2(n18953), .A(n18950), .ZN(P3_U3292) );
  AOI22_X1 U22034 ( .A1(n18955), .A2(n18954), .B1(n18953), .B2(n18952), .ZN(
        P3_U3293) );
  INV_X1 U22035 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18956) );
  AOI22_X1 U22036 ( .A1(n18957), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18956), 
        .B2(n18981), .ZN(P3_U3294) );
  NAND2_X1 U22037 ( .A1(n18959), .A2(n18958), .ZN(n18960) );
  OAI211_X1 U22038 ( .C1(n18963), .C2(n18962), .A(n18961), .B(n18960), .ZN(
        n18965) );
  MUX2_X1 U22039 ( .A(P3_MORE_REG_SCAN_IN), .B(n18965), .S(n18964), .Z(
        P3_U3295) );
  OAI21_X1 U22040 ( .B1(n18967), .B2(n18966), .A(n18985), .ZN(n18968) );
  AOI21_X1 U22041 ( .B1(n17576), .B2(n18973), .A(n18968), .ZN(n18979) );
  INV_X1 U22042 ( .A(n18969), .ZN(n18984) );
  AOI21_X1 U22043 ( .B1(n18972), .B2(n18971), .A(n18970), .ZN(n18974) );
  OAI211_X1 U22044 ( .C1(n18984), .C2(n18974), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18973), .ZN(n18976) );
  AOI21_X1 U22045 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18976), .A(n18975), 
        .ZN(n18978) );
  NAND2_X1 U22046 ( .A1(n18979), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18977) );
  OAI21_X1 U22047 ( .B1(n18979), .B2(n18978), .A(n18977), .ZN(P3_U3296) );
  OAI22_X1 U22048 ( .A1(n18981), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18980), .ZN(n18982) );
  INV_X1 U22049 ( .A(n18982), .ZN(P3_U3297) );
  OAI21_X1 U22050 ( .B1(n18983), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18985), 
        .ZN(n18988) );
  OAI22_X1 U22051 ( .A1(n18988), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18985), 
        .B2(n18984), .ZN(n18986) );
  INV_X1 U22052 ( .A(n18986), .ZN(P3_U3298) );
  OAI21_X1 U22053 ( .B1(n18988), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18987), 
        .ZN(n18989) );
  INV_X1 U22054 ( .A(n18989), .ZN(P3_U3299) );
  INV_X1 U22055 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18991) );
  NAND2_X1 U22056 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19908), .ZN(n19901) );
  NAND2_X1 U22057 ( .A1(n19897), .A2(n18990), .ZN(n19898) );
  OAI21_X1 U22058 ( .B1(n19897), .B2(n19901), .A(n19898), .ZN(n19959) );
  OAI21_X1 U22059 ( .B1(n19897), .B2(n18991), .A(n19892), .ZN(P2_U2815) );
  INV_X1 U22060 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18993) );
  OAI22_X1 U22061 ( .A1(n20019), .A2(n18993), .B1(n19237), .B2(n18992), .ZN(
        P2_U2816) );
  AOI21_X1 U22062 ( .B1(n19897), .B2(n19908), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18994) );
  AOI22_X1 U22063 ( .A1(n20039), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18994), 
        .B2(n20036), .ZN(P2_U2817) );
  INV_X1 U22064 ( .A(n19902), .ZN(n18995) );
  OAI21_X1 U22065 ( .B1(n18995), .B2(BS16), .A(n19959), .ZN(n19957) );
  OAI21_X1 U22066 ( .B1(n19959), .B2(n15893), .A(n19957), .ZN(P2_U2818) );
  NOR4_X1 U22067 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19005) );
  NOR4_X1 U22068 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19004) );
  NOR4_X1 U22069 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18996) );
  INV_X1 U22070 ( .A(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n21054) );
  INV_X1 U22071 ( .A(P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21173) );
  NAND3_X1 U22072 ( .A1(n18996), .A2(n21054), .A3(n21173), .ZN(n19002) );
  NOR4_X1 U22073 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19000) );
  NOR4_X1 U22074 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n18999) );
  NOR4_X1 U22075 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18998) );
  NOR4_X1 U22076 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_23__SCAN_IN), .A3(P2_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18997) );
  NAND4_X1 U22077 ( .A1(n19000), .A2(n18999), .A3(n18998), .A4(n18997), .ZN(
        n19001) );
  AOI211_X1 U22078 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19002), .B(n19001), .ZN(n19003) );
  NAND3_X1 U22079 ( .A1(n19005), .A2(n19004), .A3(n19003), .ZN(n19012) );
  NOR2_X1 U22080 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19012), .ZN(n19006) );
  INV_X1 U22081 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U22082 ( .A1(n19006), .A2(n19007), .B1(n19012), .B2(n19955), .ZN(
        P2_U2820) );
  OR3_X1 U22083 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19011) );
  INV_X1 U22084 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19954) );
  AOI22_X1 U22085 ( .A1(n19006), .A2(n19011), .B1(n19012), .B2(n19954), .ZN(
        P2_U2821) );
  INV_X1 U22086 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19958) );
  NAND2_X1 U22087 ( .A1(n19006), .A2(n19958), .ZN(n19010) );
  INV_X1 U22088 ( .A(n19012), .ZN(n19013) );
  OAI21_X1 U22089 ( .B1(n11471), .B2(n19007), .A(n19013), .ZN(n19008) );
  OAI21_X1 U22090 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19013), .A(n19008), 
        .ZN(n19009) );
  OAI221_X1 U22091 ( .B1(n19010), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19010), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19009), .ZN(P2_U2822) );
  INV_X1 U22092 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19952) );
  OAI221_X1 U22093 ( .B1(n19013), .B2(n19952), .C1(n19012), .C2(n19011), .A(
        n19010), .ZN(P2_U2823) );
  NAND2_X1 U22094 ( .A1(n11321), .A2(n19014), .ZN(n19015) );
  XOR2_X1 U22095 ( .A(n19016), .B(n19015), .Z(n19027) );
  OAI21_X1 U22096 ( .B1(n19928), .B2(n19110), .A(n19124), .ZN(n19020) );
  OAI22_X1 U22097 ( .A1(n19018), .A2(n19145), .B1(n19017), .B2(n19155), .ZN(
        n19019) );
  AOI211_X1 U22098 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19147), .A(n19020), .B(
        n19019), .ZN(n19026) );
  INV_X1 U22099 ( .A(n19021), .ZN(n19022) );
  OAI22_X1 U22100 ( .A1(n19023), .A2(n19149), .B1(n19022), .B2(n19143), .ZN(
        n19024) );
  INV_X1 U22101 ( .A(n19024), .ZN(n19025) );
  OAI211_X1 U22102 ( .C1(n19888), .C2(n19027), .A(n19026), .B(n19025), .ZN(
        P2_U2836) );
  AOI22_X1 U22103 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19042), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19147), .ZN(n19028) );
  OAI211_X1 U22104 ( .C1(n19036), .C2(n19154), .A(n19028), .B(n19324), .ZN(
        n19029) );
  AOI21_X1 U22105 ( .B1(n19030), .B2(n19135), .A(n19029), .ZN(n19031) );
  OAI21_X1 U22106 ( .B1(n19110), .B2(n19925), .A(n19031), .ZN(n19032) );
  AOI21_X1 U22107 ( .B1(n19033), .B2(n19102), .A(n19032), .ZN(n19039) );
  INV_X1 U22108 ( .A(n19034), .ZN(n19037) );
  OAI211_X1 U22109 ( .C1(n19037), .C2(n19036), .A(n19136), .B(n19035), .ZN(
        n19038) );
  OAI211_X1 U22110 ( .C1(n19143), .C2(n19040), .A(n19039), .B(n19038), .ZN(
        P2_U2838) );
  INV_X1 U22111 ( .A(n19041), .ZN(n19049) );
  AOI22_X1 U22112 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19042), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n19147), .ZN(n19043) );
  OAI211_X1 U22113 ( .C1(n19044), .C2(n19149), .A(n19043), .B(n19324), .ZN(
        n19045) );
  AOI21_X1 U22114 ( .B1(n19046), .B2(n19051), .A(n19045), .ZN(n19047) );
  OAI21_X1 U22115 ( .B1(n19110), .B2(n11956), .A(n19047), .ZN(n19048) );
  AOI21_X1 U22116 ( .B1(n19049), .B2(n19102), .A(n19048), .ZN(n19056) );
  INV_X1 U22117 ( .A(n19050), .ZN(n19054) );
  INV_X1 U22118 ( .A(n19051), .ZN(n19053) );
  OAI21_X1 U22119 ( .B1(n19054), .B2(n19053), .A(n19052), .ZN(n19055) );
  OAI211_X1 U22120 ( .C1(n19143), .C2(n19177), .A(n19056), .B(n19055), .ZN(
        P2_U2840) );
  NAND2_X1 U22121 ( .A1(n11321), .A2(n19057), .ZN(n19059) );
  XOR2_X1 U22122 ( .A(n19059), .B(n19058), .Z(n19067) );
  AOI22_X1 U22123 ( .A1(n19060), .A2(n19102), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n19147), .ZN(n19061) );
  OAI211_X1 U22124 ( .C1(n11903), .C2(n19110), .A(n19061), .B(n19324), .ZN(
        n19065) );
  INV_X1 U22125 ( .A(n19062), .ZN(n19063) );
  OAI22_X1 U22126 ( .A1(n19063), .A2(n19149), .B1(n19143), .B2(n19182), .ZN(
        n19064) );
  AOI211_X1 U22127 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n19115), .A(
        n19065), .B(n19064), .ZN(n19066) );
  OAI21_X1 U22128 ( .B1(n19067), .B2(n19888), .A(n19066), .ZN(P2_U2842) );
  NAND2_X1 U22129 ( .A1(n11321), .A2(n19068), .ZN(n19070) );
  XOR2_X1 U22130 ( .A(n19070), .B(n19069), .Z(n19077) );
  AOI22_X1 U22131 ( .A1(n19071), .A2(n19102), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n19147), .ZN(n19072) );
  OAI211_X1 U22132 ( .C1(n11862), .C2(n19110), .A(n19072), .B(n19324), .ZN(
        n19075) );
  OAI22_X1 U22133 ( .A1(n19187), .A2(n19143), .B1(n19149), .B2(n19073), .ZN(
        n19074) );
  AOI211_X1 U22134 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19115), .A(
        n19075), .B(n19074), .ZN(n19076) );
  OAI21_X1 U22135 ( .B1(n19077), .B2(n19888), .A(n19076), .ZN(P2_U2844) );
  OAI21_X1 U22136 ( .B1(n11845), .B2(n19110), .A(n19124), .ZN(n19081) );
  OAI22_X1 U22137 ( .A1(n19079), .A2(n19145), .B1(n19126), .B2(n19078), .ZN(
        n19080) );
  AOI211_X1 U22138 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19115), .A(
        n19081), .B(n19080), .ZN(n19088) );
  NOR2_X1 U22139 ( .A1(n19117), .A2(n19082), .ZN(n19084) );
  XNOR2_X1 U22140 ( .A(n19084), .B(n19083), .ZN(n19086) );
  AOI22_X1 U22141 ( .A1(n19086), .A2(n19136), .B1(n19135), .B2(n19085), .ZN(
        n19087) );
  OAI211_X1 U22142 ( .C1(n19190), .C2(n19143), .A(n19088), .B(n19087), .ZN(
        P2_U2845) );
  NAND2_X1 U22143 ( .A1(n11321), .A2(n19089), .ZN(n19091) );
  XOR2_X1 U22144 ( .A(n19091), .B(n19090), .Z(n19098) );
  AOI22_X1 U22145 ( .A1(n19092), .A2(n19102), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19147), .ZN(n19093) );
  OAI211_X1 U22146 ( .C1(n15608), .C2(n19110), .A(n19093), .B(n19324), .ZN(
        n19096) );
  OAI22_X1 U22147 ( .A1(n19192), .A2(n19143), .B1(n19149), .B2(n19094), .ZN(
        n19095) );
  AOI211_X1 U22148 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19115), .A(
        n19096), .B(n19095), .ZN(n19097) );
  OAI21_X1 U22149 ( .B1(n19098), .B2(n19888), .A(n19097), .ZN(P2_U2846) );
  NAND2_X1 U22150 ( .A1(n11321), .A2(n19099), .ZN(n19101) );
  XOR2_X1 U22151 ( .A(n19101), .B(n19100), .Z(n19109) );
  AOI22_X1 U22152 ( .A1(n19103), .A2(n19102), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19147), .ZN(n19104) );
  OAI211_X1 U22153 ( .C1(n11535), .C2(n19110), .A(n19104), .B(n19324), .ZN(
        n19107) );
  OAI22_X1 U22154 ( .A1(n19143), .A2(n19196), .B1(n19105), .B2(n19149), .ZN(
        n19106) );
  AOI211_X1 U22155 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19115), .A(
        n19107), .B(n19106), .ZN(n19108) );
  OAI21_X1 U22156 ( .B1(n19109), .B2(n19888), .A(n19108), .ZN(P2_U2848) );
  OAI21_X1 U22157 ( .B1(n11529), .B2(n19110), .A(n19124), .ZN(n19114) );
  OAI22_X1 U22158 ( .A1(n19112), .A2(n19145), .B1(n19126), .B2(n19111), .ZN(
        n19113) );
  AOI211_X1 U22159 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19115), .A(
        n19114), .B(n19113), .ZN(n19123) );
  NOR2_X1 U22160 ( .A1(n19117), .A2(n19116), .ZN(n19119) );
  XNOR2_X1 U22161 ( .A(n19119), .B(n19118), .ZN(n19121) );
  AOI22_X1 U22162 ( .A1(n19121), .A2(n19136), .B1(n19135), .B2(n19120), .ZN(
        n19122) );
  OAI211_X1 U22163 ( .C1(n19143), .C2(n19199), .A(n19123), .B(n19122), .ZN(
        P2_U2849) );
  OAI21_X1 U22164 ( .B1(n19126), .B2(n19125), .A(n19124), .ZN(n19130) );
  OAI22_X1 U22165 ( .A1(n19145), .A2(n19128), .B1(n19127), .B2(n19155), .ZN(
        n19129) );
  AOI211_X1 U22166 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n9962), .A(n19130), .B(
        n19129), .ZN(n19139) );
  NAND2_X1 U22167 ( .A1(n11321), .A2(n19131), .ZN(n19132) );
  XNOR2_X1 U22168 ( .A(n19133), .B(n19132), .ZN(n19137) );
  AOI22_X1 U22169 ( .A1(n19137), .A2(n19136), .B1(n19135), .B2(n19134), .ZN(
        n19138) );
  OAI211_X1 U22170 ( .C1(n19143), .C2(n19206), .A(n19139), .B(n19138), .ZN(
        P2_U2850) );
  INV_X1 U22171 ( .A(n19140), .ZN(n19162) );
  INV_X1 U22172 ( .A(n19141), .ZN(n19142) );
  OAI22_X1 U22173 ( .A1(n19145), .A2(n19144), .B1(n19143), .B2(n19142), .ZN(
        n19146) );
  AOI21_X1 U22174 ( .B1(n19147), .B2(P2_EBX_REG_0__SCAN_IN), .A(n19146), .ZN(
        n19148) );
  OAI21_X1 U22175 ( .B1(n19150), .B2(n19149), .A(n19148), .ZN(n19151) );
  AOI21_X1 U22176 ( .B1(n9962), .B2(P2_REIP_REG_0__SCAN_IN), .A(n19151), .ZN(
        n19160) );
  AOI21_X1 U22177 ( .B1(n19155), .B2(n19154), .A(n19153), .ZN(n19156) );
  AOI21_X1 U22178 ( .B1(n19158), .B2(n19157), .A(n19156), .ZN(n19159) );
  OAI211_X1 U22179 ( .C1(n19162), .C2(n19161), .A(n19160), .B(n19159), .ZN(
        P2_U2855) );
  AOI22_X1 U22180 ( .A1(n19223), .A2(n19163), .B1(n19169), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19165) );
  AOI22_X1 U22181 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19222), .B1(n19168), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19164) );
  NAND2_X1 U22182 ( .A1(n19165), .A2(n19164), .ZN(P2_U2888) );
  AOI22_X1 U22183 ( .A1(n19167), .A2(n19166), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19222), .ZN(n19175) );
  AOI22_X1 U22184 ( .A1(n19169), .A2(BUF1_REG_16__SCAN_IN), .B1(n19168), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19174) );
  INV_X1 U22185 ( .A(n19170), .ZN(n19171) );
  AOI22_X1 U22186 ( .A1(n19172), .A2(n19210), .B1(n19223), .B2(n19171), .ZN(
        n19173) );
  NAND3_X1 U22187 ( .A1(n19175), .A2(n19174), .A3(n19173), .ZN(P2_U2903) );
  OAI222_X1 U22188 ( .A1(n19177), .A2(n19207), .B1(n13081), .B2(n19198), .C1(
        n19176), .C2(n19231), .ZN(P2_U2904) );
  INV_X1 U22189 ( .A(n19178), .ZN(n19180) );
  AOI22_X1 U22190 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19222), .B1(n19302), 
        .B2(n19200), .ZN(n19179) );
  OAI21_X1 U22191 ( .B1(n19207), .B2(n19180), .A(n19179), .ZN(P2_U2905) );
  INV_X1 U22192 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19274) );
  OAI222_X1 U22193 ( .A1(n19182), .A2(n19207), .B1(n19274), .B2(n19198), .C1(
        n19231), .C2(n19181), .ZN(P2_U2906) );
  AOI22_X1 U22194 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19222), .B1(n19183), 
        .B2(n19200), .ZN(n19184) );
  OAI21_X1 U22195 ( .B1(n19207), .B2(n19185), .A(n19184), .ZN(P2_U2907) );
  INV_X1 U22196 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19278) );
  OAI222_X1 U22197 ( .A1(n19187), .A2(n19207), .B1(n19278), .B2(n19198), .C1(
        n19231), .C2(n19186), .ZN(P2_U2908) );
  AOI22_X1 U22198 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19222), .B1(n19188), 
        .B2(n19200), .ZN(n19189) );
  OAI21_X1 U22199 ( .B1(n19207), .B2(n19190), .A(n19189), .ZN(P2_U2909) );
  INV_X1 U22200 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19282) );
  OAI222_X1 U22201 ( .A1(n19192), .A2(n19207), .B1(n19282), .B2(n19198), .C1(
        n19231), .C2(n19191), .ZN(P2_U2910) );
  AOI22_X1 U22202 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19222), .B1(n19193), .B2(
        n19200), .ZN(n19194) );
  OAI21_X1 U22203 ( .B1(n19207), .B2(n19195), .A(n19194), .ZN(P2_U2911) );
  INV_X1 U22204 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n21269) );
  OAI222_X1 U22205 ( .A1(n19196), .A2(n19207), .B1(n21269), .B2(n19198), .C1(
        n19231), .C2(n19357), .ZN(P2_U2912) );
  INV_X1 U22206 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19287) );
  INV_X1 U22207 ( .A(n19197), .ZN(n19348) );
  OAI222_X1 U22208 ( .A1(n19199), .A2(n19207), .B1(n19287), .B2(n19198), .C1(
        n19231), .C2(n19348), .ZN(P2_U2913) );
  AOI22_X1 U22209 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19222), .B1(n19201), .B2(
        n19200), .ZN(n19205) );
  AOI21_X1 U22210 ( .B1(n19983), .B2(n19981), .A(n19202), .ZN(n19217) );
  XNOR2_X1 U22211 ( .A(n19972), .B(n19214), .ZN(n19216) );
  NOR2_X1 U22212 ( .A1(n19217), .A2(n19216), .ZN(n19215) );
  AOI21_X1 U22213 ( .B1(n19214), .B2(n19972), .A(n19215), .ZN(n19203) );
  NOR2_X1 U22214 ( .A1(n19203), .A2(n19309), .ZN(n19208) );
  OR3_X1 U22215 ( .A1(n19208), .A2(n19209), .A3(n19227), .ZN(n19204) );
  OAI211_X1 U22216 ( .C1(n19207), .C2(n19206), .A(n19205), .B(n19204), .ZN(
        P2_U2914) );
  AOI22_X1 U22217 ( .A1(n19223), .A2(n19309), .B1(n19222), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19213) );
  XOR2_X1 U22218 ( .A(n19209), .B(n19208), .Z(n19211) );
  NAND2_X1 U22219 ( .A1(n19211), .A2(n19210), .ZN(n19212) );
  OAI211_X1 U22220 ( .C1(n19338), .C2(n19231), .A(n19213), .B(n19212), .ZN(
        P2_U2915) );
  INV_X1 U22221 ( .A(n19214), .ZN(n19978) );
  AOI22_X1 U22222 ( .A1(n19223), .A2(n19978), .B1(n19222), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19220) );
  AOI21_X1 U22223 ( .B1(n19217), .B2(n19216), .A(n19215), .ZN(n19218) );
  OR2_X1 U22224 ( .A1(n19218), .A2(n19227), .ZN(n19219) );
  OAI211_X1 U22225 ( .C1(n19221), .C2(n19231), .A(n19220), .B(n19219), .ZN(
        P2_U2916) );
  AOI22_X1 U22226 ( .A1(n19223), .A2(n19994), .B1(n19222), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19230) );
  AOI21_X1 U22227 ( .B1(n19226), .B2(n19225), .A(n19224), .ZN(n19228) );
  OR2_X1 U22228 ( .A1(n19228), .A2(n19227), .ZN(n19229) );
  OAI211_X1 U22229 ( .C1(n19232), .C2(n19231), .A(n19230), .B(n19229), .ZN(
        P2_U2918) );
  NAND2_X1 U22230 ( .A1(n19238), .A2(n19237), .ZN(n20022) );
  NOR2_X1 U22231 ( .A1(n19256), .A2(n21176), .ZN(P2_U2920) );
  INV_X1 U22232 ( .A(n19268), .ZN(n19254) );
  AOI22_X1 U22233 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19254), .B1(n19299), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19240) );
  OAI21_X1 U22234 ( .B1(n21222), .B2(n19256), .A(n19240), .ZN(P2_U2921) );
  AOI22_X1 U22235 ( .A1(n19299), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19241) );
  OAI21_X1 U22236 ( .B1(n19242), .B2(n19268), .A(n19241), .ZN(P2_U2922) );
  AOI22_X1 U22237 ( .A1(n19299), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19243) );
  OAI21_X1 U22238 ( .B1(n19244), .B2(n19268), .A(n19243), .ZN(P2_U2923) );
  AOI22_X1 U22239 ( .A1(n19299), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19245) );
  OAI21_X1 U22240 ( .B1(n21193), .B2(n19268), .A(n19245), .ZN(P2_U2924) );
  AOI22_X1 U22241 ( .A1(n19299), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19246) );
  OAI21_X1 U22242 ( .B1(n19247), .B2(n19268), .A(n19246), .ZN(P2_U2925) );
  AOI22_X1 U22243 ( .A1(n19299), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19248) );
  OAI21_X1 U22244 ( .B1(n19249), .B2(n19268), .A(n19248), .ZN(P2_U2926) );
  AOI22_X1 U22245 ( .A1(n19299), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19250) );
  OAI21_X1 U22246 ( .B1(n19251), .B2(n19268), .A(n19250), .ZN(P2_U2927) );
  AOI22_X1 U22247 ( .A1(n19299), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19252) );
  OAI21_X1 U22248 ( .B1(n19253), .B2(n19268), .A(n19252), .ZN(P2_U2928) );
  AOI22_X1 U22249 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n19254), .B1(n19299), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n19255) );
  OAI21_X1 U22250 ( .B1(n19256), .B2(n21180), .A(n19255), .ZN(P2_U2929) );
  AOI22_X1 U22251 ( .A1(n19299), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19257) );
  OAI21_X1 U22252 ( .B1(n19258), .B2(n19268), .A(n19257), .ZN(P2_U2930) );
  INV_X1 U22253 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19260) );
  AOI22_X1 U22254 ( .A1(n19299), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19259) );
  OAI21_X1 U22255 ( .B1(n19260), .B2(n19268), .A(n19259), .ZN(P2_U2931) );
  AOI22_X1 U22256 ( .A1(n19299), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19261) );
  OAI21_X1 U22257 ( .B1(n19262), .B2(n19268), .A(n19261), .ZN(P2_U2932) );
  INV_X1 U22258 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19264) );
  AOI22_X1 U22259 ( .A1(n19299), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19263) );
  OAI21_X1 U22260 ( .B1(n19264), .B2(n19268), .A(n19263), .ZN(P2_U2933) );
  AOI22_X1 U22261 ( .A1(n19299), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19265) );
  OAI21_X1 U22262 ( .B1(n19266), .B2(n19268), .A(n19265), .ZN(P2_U2934) );
  AOI22_X1 U22263 ( .A1(n19299), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19267) );
  OAI21_X1 U22264 ( .B1(n19269), .B2(n19268), .A(n19267), .ZN(P2_U2935) );
  AOI22_X1 U22265 ( .A1(n19299), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19270) );
  OAI21_X1 U22266 ( .B1(n13081), .B2(n19301), .A(n19270), .ZN(P2_U2936) );
  INV_X1 U22267 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19272) );
  AOI22_X1 U22268 ( .A1(n19299), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19271) );
  OAI21_X1 U22269 ( .B1(n19272), .B2(n19301), .A(n19271), .ZN(P2_U2937) );
  AOI22_X1 U22270 ( .A1(n19299), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19273) );
  OAI21_X1 U22271 ( .B1(n19274), .B2(n19301), .A(n19273), .ZN(P2_U2938) );
  AOI22_X1 U22272 ( .A1(n19299), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19275) );
  OAI21_X1 U22273 ( .B1(n19276), .B2(n19301), .A(n19275), .ZN(P2_U2939) );
  AOI22_X1 U22274 ( .A1(n19299), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19277) );
  OAI21_X1 U22275 ( .B1(n19278), .B2(n19301), .A(n19277), .ZN(P2_U2940) );
  AOI22_X1 U22276 ( .A1(n19299), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19279) );
  OAI21_X1 U22277 ( .B1(n19280), .B2(n19301), .A(n19279), .ZN(P2_U2941) );
  AOI22_X1 U22278 ( .A1(n19299), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19281) );
  OAI21_X1 U22279 ( .B1(n19282), .B2(n19301), .A(n19281), .ZN(P2_U2942) );
  AOI22_X1 U22280 ( .A1(n19299), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19283) );
  OAI21_X1 U22281 ( .B1(n19284), .B2(n19301), .A(n19283), .ZN(P2_U2943) );
  AOI22_X1 U22282 ( .A1(n19299), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19285) );
  OAI21_X1 U22283 ( .B1(n21269), .B2(n19301), .A(n19285), .ZN(P2_U2944) );
  AOI22_X1 U22284 ( .A1(n19299), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19286) );
  OAI21_X1 U22285 ( .B1(n19287), .B2(n19301), .A(n19286), .ZN(P2_U2945) );
  INV_X1 U22286 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19290) );
  AOI22_X1 U22287 ( .A1(n19299), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19289) );
  OAI21_X1 U22288 ( .B1(n19290), .B2(n19301), .A(n19289), .ZN(P2_U2946) );
  INV_X1 U22289 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19292) );
  AOI22_X1 U22290 ( .A1(n19299), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19291) );
  OAI21_X1 U22291 ( .B1(n19292), .B2(n19301), .A(n19291), .ZN(P2_U2947) );
  INV_X1 U22292 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19294) );
  AOI22_X1 U22293 ( .A1(n19299), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19293) );
  OAI21_X1 U22294 ( .B1(n19294), .B2(n19301), .A(n19293), .ZN(P2_U2948) );
  INV_X1 U22295 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19296) );
  AOI22_X1 U22296 ( .A1(n19299), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19295) );
  OAI21_X1 U22297 ( .B1(n19296), .B2(n19301), .A(n19295), .ZN(P2_U2949) );
  INV_X1 U22298 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19298) );
  AOI22_X1 U22299 ( .A1(n19299), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19297) );
  OAI21_X1 U22300 ( .B1(n19298), .B2(n19301), .A(n19297), .ZN(P2_U2950) );
  AOI22_X1 U22301 ( .A1(n19299), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19288), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19300) );
  OAI21_X1 U22302 ( .B1(n13083), .B2(n19301), .A(n19300), .ZN(P2_U2951) );
  AOI22_X1 U22303 ( .A1(n19306), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19305), .ZN(n19304) );
  NAND2_X1 U22304 ( .A1(n19303), .A2(n19302), .ZN(n19307) );
  NAND2_X1 U22305 ( .A1(n19304), .A2(n19307), .ZN(P2_U2966) );
  AOI22_X1 U22306 ( .A1(n19306), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19305), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19308) );
  NAND2_X1 U22307 ( .A1(n19308), .A2(n19307), .ZN(P2_U2981) );
  AOI22_X1 U22308 ( .A1(n19311), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19310), .B2(n19309), .ZN(n19323) );
  OAI22_X1 U22309 ( .A1(n19314), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19313), .B2(n19312), .ZN(n19321) );
  INV_X1 U22310 ( .A(n19315), .ZN(n19319) );
  OAI22_X1 U22311 ( .A1(n19319), .A2(n19318), .B1(n19317), .B2(n19316), .ZN(
        n19320) );
  NOR2_X1 U22312 ( .A1(n19321), .A2(n19320), .ZN(n19322) );
  OAI211_X1 U22313 ( .C1(n11650), .C2(n19324), .A(n19323), .B(n19322), .ZN(
        P2_U3042) );
  INV_X1 U22314 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19330) );
  AOI22_X2 U22315 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19352), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19353), .ZN(n19838) );
  INV_X1 U22316 ( .A(n19838), .ZN(n19664) );
  AOI22_X1 U22317 ( .A1(n19664), .A2(n19879), .B1(n19356), .B2(n19827), .ZN(
        n19329) );
  AOI22_X1 U22318 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19352), .ZN(n19327) );
  AOI22_X1 U22319 ( .A1(n19326), .A2(n19360), .B1(n19400), .B2(n19835), .ZN(
        n19328) );
  OAI211_X1 U22320 ( .C1(n19364), .C2(n19330), .A(n19329), .B(n19328), .ZN(
        P2_U3048) );
  AOI22_X1 U22321 ( .A1(n19700), .A2(n19879), .B1(n19839), .B2(n19356), .ZN(
        n19332) );
  AOI22_X1 U22322 ( .A1(n15917), .A2(n19360), .B1(n19400), .B2(n19840), .ZN(
        n19331) );
  OAI211_X1 U22323 ( .C1(n19364), .C2(n19333), .A(n19332), .B(n19331), .ZN(
        P2_U3049) );
  INV_X1 U22324 ( .A(n19855), .ZN(n19800) );
  AOI22_X1 U22325 ( .A1(n19800), .A2(n19879), .B1(n19356), .B2(n19850), .ZN(
        n19335) );
  AOI22_X1 U22326 ( .A1(n19851), .A2(n19360), .B1(n19400), .B2(n19852), .ZN(
        n19334) );
  OAI211_X1 U22327 ( .C1(n19364), .C2(n19336), .A(n19335), .B(n19334), .ZN(
        P2_U3051) );
  OAI22_X2 U22328 ( .A1(n20314), .A2(n19359), .B1(n21189), .B2(n19358), .ZN(
        n19804) );
  NOR2_X2 U22329 ( .A1(n19337), .A2(n19342), .ZN(n19856) );
  AOI22_X1 U22330 ( .A1(n19804), .A2(n19879), .B1(n19356), .B2(n19856), .ZN(
        n19340) );
  NOR2_X2 U22331 ( .A1(n19338), .A2(n19576), .ZN(n19857) );
  AOI22_X1 U22332 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19352), .ZN(n19807) );
  INV_X1 U22333 ( .A(n19807), .ZN(n19858) );
  AOI22_X1 U22334 ( .A1(n19857), .A2(n19360), .B1(n19400), .B2(n19858), .ZN(
        n19339) );
  OAI211_X1 U22335 ( .C1(n19364), .C2(n19341), .A(n19340), .B(n19339), .ZN(
        P2_U3052) );
  AOI22_X1 U22336 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19352), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19353), .ZN(n19867) );
  INV_X1 U22337 ( .A(n19867), .ZN(n19676) );
  NOR2_X2 U22338 ( .A1(n12883), .A2(n19342), .ZN(n19862) );
  AOI22_X1 U22339 ( .A1(n19676), .A2(n19879), .B1(n19356), .B2(n19862), .ZN(
        n19345) );
  NOR2_X2 U22340 ( .A1(n19343), .A2(n19576), .ZN(n19863) );
  OAI22_X2 U22341 ( .A1(n15457), .A2(n19359), .B1(n15455), .B2(n19358), .ZN(
        n19864) );
  AOI22_X1 U22342 ( .A1(n19863), .A2(n19360), .B1(n19400), .B2(n19864), .ZN(
        n19344) );
  OAI211_X1 U22343 ( .C1(n19364), .C2(n13423), .A(n19345), .B(n19344), .ZN(
        P2_U3053) );
  OAI22_X2 U22344 ( .A1(n20330), .A2(n19359), .B1(n19346), .B2(n19358), .ZN(
        n19812) );
  AOI22_X1 U22345 ( .A1(n19812), .A2(n19879), .B1(n19356), .B2(n19868), .ZN(
        n19350) );
  NOR2_X2 U22346 ( .A1(n19348), .A2(n19576), .ZN(n19869) );
  AOI22_X1 U22347 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19352), .ZN(n19815) );
  INV_X1 U22348 ( .A(n19815), .ZN(n19870) );
  AOI22_X1 U22349 ( .A1(n19869), .A2(n19360), .B1(n19400), .B2(n19870), .ZN(
        n19349) );
  OAI211_X1 U22350 ( .C1(n19364), .C2(n19351), .A(n19350), .B(n19349), .ZN(
        P2_U3054) );
  AOI22_X1 U22351 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19353), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19352), .ZN(n19884) );
  INV_X1 U22352 ( .A(n19884), .ZN(n19818) );
  AOI22_X1 U22353 ( .A1(n19818), .A2(n19879), .B1(n19356), .B2(n19875), .ZN(
        n19362) );
  NOR2_X2 U22354 ( .A1(n19357), .A2(n19576), .ZN(n19876) );
  AOI22_X1 U22355 ( .A1(n19876), .A2(n19360), .B1(n19400), .B2(n19878), .ZN(
        n19361) );
  OAI211_X1 U22356 ( .C1(n19364), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        P2_U3055) );
  INV_X1 U22357 ( .A(n19400), .ZN(n19387) );
  NAND2_X1 U22358 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19996), .ZN(
        n19634) );
  INV_X1 U22359 ( .A(n19438), .ZN(n19437) );
  NOR2_X1 U22360 ( .A1(n19634), .A2(n19437), .ZN(n19375) );
  OR2_X1 U22361 ( .A1(n19375), .A2(n20017), .ZN(n19365) );
  NOR2_X1 U22362 ( .A1(n19366), .A2(n19365), .ZN(n19371) );
  INV_X1 U22363 ( .A(n19372), .ZN(n19367) );
  NOR2_X1 U22364 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19367), .ZN(n19369) );
  INV_X1 U22365 ( .A(n19368), .ZN(n19574) );
  INV_X1 U22366 ( .A(n19326), .ZN(n19476) );
  INV_X1 U22367 ( .A(n19827), .ZN(n19475) );
  INV_X1 U22368 ( .A(n19375), .ZN(n19397) );
  OAI22_X1 U22369 ( .A1(n19398), .A2(n19476), .B1(n19475), .B2(n19397), .ZN(
        n19370) );
  INV_X1 U22370 ( .A(n19370), .ZN(n19377) );
  NAND2_X1 U22371 ( .A1(n19575), .A2(n19635), .ZN(n19373) );
  AOI21_X1 U22372 ( .B1(n19373), .B2(n19372), .A(n19371), .ZN(n19374) );
  OAI211_X1 U22373 ( .C1(n19375), .C2(n19825), .A(n19374), .B(n19833), .ZN(
        n19401) );
  INV_X1 U22374 ( .A(n19435), .ZN(n19427) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19401), .B1(
        n19427), .B2(n19835), .ZN(n19376) );
  OAI211_X1 U22376 ( .C1(n19838), .C2(n19387), .A(n19377), .B(n19376), .ZN(
        P2_U3056) );
  INV_X1 U22377 ( .A(n15917), .ZN(n19485) );
  OAI22_X1 U22378 ( .A1(n19398), .A2(n19485), .B1(n19484), .B2(n19397), .ZN(
        n19378) );
  INV_X1 U22379 ( .A(n19378), .ZN(n19380) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19700), .ZN(n19379) );
  OAI211_X1 U22381 ( .C1(n19703), .C2(n19435), .A(n19380), .B(n19379), .ZN(
        P2_U3057) );
  INV_X1 U22382 ( .A(n19845), .ZN(n19490) );
  INV_X1 U22383 ( .A(n19844), .ZN(n19489) );
  OAI22_X1 U22384 ( .A1(n19398), .A2(n19490), .B1(n19489), .B2(n19397), .ZN(
        n19381) );
  INV_X1 U22385 ( .A(n19381), .ZN(n19383) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19401), .B1(
        n19427), .B2(n19846), .ZN(n19382) );
  OAI211_X1 U22387 ( .C1(n19849), .C2(n19387), .A(n19383), .B(n19382), .ZN(
        P2_U3058) );
  INV_X1 U22388 ( .A(n19851), .ZN(n19495) );
  INV_X1 U22389 ( .A(n19850), .ZN(n19494) );
  OAI22_X1 U22390 ( .A1(n19398), .A2(n19495), .B1(n19494), .B2(n19397), .ZN(
        n19384) );
  INV_X1 U22391 ( .A(n19384), .ZN(n19386) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19401), .B1(
        n19427), .B2(n19852), .ZN(n19385) );
  OAI211_X1 U22393 ( .C1(n19855), .C2(n19387), .A(n19386), .B(n19385), .ZN(
        P2_U3059) );
  INV_X1 U22394 ( .A(n19857), .ZN(n19500) );
  INV_X1 U22395 ( .A(n19856), .ZN(n19499) );
  OAI22_X1 U22396 ( .A1(n19398), .A2(n19500), .B1(n19499), .B2(n19397), .ZN(
        n19388) );
  INV_X1 U22397 ( .A(n19388), .ZN(n19390) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19804), .ZN(n19389) );
  OAI211_X1 U22399 ( .C1(n19807), .C2(n19435), .A(n19390), .B(n19389), .ZN(
        P2_U3060) );
  INV_X1 U22400 ( .A(n19864), .ZN(n19564) );
  INV_X1 U22401 ( .A(n19863), .ZN(n19505) );
  INV_X1 U22402 ( .A(n19862), .ZN(n19504) );
  OAI22_X1 U22403 ( .A1(n19398), .A2(n19505), .B1(n19504), .B2(n19397), .ZN(
        n19391) );
  INV_X1 U22404 ( .A(n19391), .ZN(n19393) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19676), .ZN(n19392) );
  OAI211_X1 U22406 ( .C1(n19564), .C2(n19435), .A(n19393), .B(n19392), .ZN(
        P2_U3061) );
  INV_X1 U22407 ( .A(n19869), .ZN(n19510) );
  INV_X1 U22408 ( .A(n19868), .ZN(n19509) );
  OAI22_X1 U22409 ( .A1(n19398), .A2(n19510), .B1(n19509), .B2(n19397), .ZN(
        n19394) );
  INV_X1 U22410 ( .A(n19394), .ZN(n19396) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19812), .ZN(n19395) );
  OAI211_X1 U22412 ( .C1(n19815), .C2(n19435), .A(n19396), .B(n19395), .ZN(
        P2_U3062) );
  INV_X1 U22413 ( .A(n19876), .ZN(n19517) );
  INV_X1 U22414 ( .A(n19875), .ZN(n19516) );
  OAI22_X1 U22415 ( .A1(n19398), .A2(n19517), .B1(n19516), .B2(n19397), .ZN(
        n19399) );
  INV_X1 U22416 ( .A(n19399), .ZN(n19403) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19818), .ZN(n19402) );
  OAI211_X1 U22418 ( .C1(n19823), .C2(n19435), .A(n19403), .B(n19402), .ZN(
        P2_U3063) );
  NAND2_X1 U22419 ( .A1(n19404), .A2(n19438), .ZN(n19408) );
  AOI21_X1 U22420 ( .B1(n19405), .B2(n19408), .A(n20017), .ZN(n19407) );
  NOR2_X1 U22421 ( .A1(n19406), .A2(n19437), .ZN(n19409) );
  OR2_X1 U22422 ( .A1(n19407), .A2(n19409), .ZN(n19431) );
  INV_X1 U22423 ( .A(n19408), .ZN(n19430) );
  AOI22_X1 U22424 ( .A1(n19431), .A2(n19326), .B1(n19827), .B2(n19430), .ZN(
        n19416) );
  NAND2_X1 U22425 ( .A1(n19461), .A2(n19435), .ZN(n19410) );
  AOI21_X1 U22426 ( .B1(n19410), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19409), 
        .ZN(n19413) );
  AOI21_X1 U22427 ( .B1(n19411), .B2(n19825), .A(n19430), .ZN(n19412) );
  MUX2_X1 U22428 ( .A(n19413), .B(n19412), .S(n19974), .Z(n19414) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19432), .B1(
        n19463), .B2(n19835), .ZN(n19415) );
  OAI211_X1 U22430 ( .C1(n19838), .C2(n19435), .A(n19416), .B(n19415), .ZN(
        P2_U3064) );
  AOI22_X1 U22431 ( .A1(n19431), .A2(n15917), .B1(n19839), .B2(n19430), .ZN(
        n19418) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19432), .B1(
        n19463), .B2(n19840), .ZN(n19417) );
  OAI211_X1 U22433 ( .C1(n19843), .C2(n19435), .A(n19418), .B(n19417), .ZN(
        P2_U3065) );
  AOI22_X1 U22434 ( .A1(n19431), .A2(n19845), .B1(n19844), .B2(n19430), .ZN(
        n19420) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19432), .B1(
        n19463), .B2(n19846), .ZN(n19419) );
  OAI211_X1 U22436 ( .C1(n19849), .C2(n19435), .A(n19420), .B(n19419), .ZN(
        P2_U3066) );
  AOI22_X1 U22437 ( .A1(n19431), .A2(n19851), .B1(n19850), .B2(n19430), .ZN(
        n19422) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19432), .B1(
        n19463), .B2(n19852), .ZN(n19421) );
  OAI211_X1 U22439 ( .C1(n19855), .C2(n19435), .A(n19422), .B(n19421), .ZN(
        P2_U3067) );
  AOI22_X1 U22440 ( .A1(n19431), .A2(n19857), .B1(n19856), .B2(n19430), .ZN(
        n19424) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19432), .B1(
        n19427), .B2(n19804), .ZN(n19423) );
  OAI211_X1 U22442 ( .C1(n19807), .C2(n19461), .A(n19424), .B(n19423), .ZN(
        P2_U3068) );
  AOI22_X1 U22443 ( .A1(n19431), .A2(n19863), .B1(n19862), .B2(n19430), .ZN(
        n19426) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19432), .B1(
        n19463), .B2(n19864), .ZN(n19425) );
  OAI211_X1 U22445 ( .C1(n19867), .C2(n19435), .A(n19426), .B(n19425), .ZN(
        P2_U3069) );
  AOI22_X1 U22446 ( .A1(n19431), .A2(n19869), .B1(n19868), .B2(n19430), .ZN(
        n19429) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19432), .B1(
        n19427), .B2(n19812), .ZN(n19428) );
  OAI211_X1 U22448 ( .C1(n19815), .C2(n19461), .A(n19429), .B(n19428), .ZN(
        P2_U3070) );
  AOI22_X1 U22449 ( .A1(n19431), .A2(n19876), .B1(n19875), .B2(n19430), .ZN(
        n19434) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19432), .B1(
        n19463), .B2(n19878), .ZN(n19433) );
  OAI211_X1 U22451 ( .C1(n19884), .C2(n19435), .A(n19434), .B(n19433), .ZN(
        P2_U3071) );
  NOR2_X1 U22452 ( .A1(n19688), .A2(n19437), .ZN(n19462) );
  AOI22_X1 U22453 ( .A1(n19835), .A2(n19512), .B1(n19462), .B2(n19827), .ZN(
        n19448) );
  INV_X1 U22454 ( .A(n19575), .ZN(n19975) );
  OAI21_X1 U22455 ( .B1(n19975), .B2(n19694), .A(n19971), .ZN(n19446) );
  NAND2_X1 U22456 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19438), .ZN(
        n19445) );
  INV_X1 U22457 ( .A(n19445), .ZN(n19441) );
  INV_X1 U22458 ( .A(n19462), .ZN(n19439) );
  OAI211_X1 U22459 ( .C1(n19442), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19974), 
        .B(n19439), .ZN(n19440) );
  OAI211_X1 U22460 ( .C1(n19446), .C2(n19441), .A(n19833), .B(n19440), .ZN(
        n19465) );
  INV_X1 U22461 ( .A(n19442), .ZN(n19443) );
  OAI21_X1 U22462 ( .B1(n19443), .B2(n19462), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19444) );
  OAI21_X1 U22463 ( .B1(n19446), .B2(n19445), .A(n19444), .ZN(n19464) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19465), .B1(
        n19326), .B2(n19464), .ZN(n19447) );
  OAI211_X1 U22465 ( .C1(n19838), .C2(n19461), .A(n19448), .B(n19447), .ZN(
        P2_U3072) );
  AOI22_X1 U22466 ( .A1(n19700), .A2(n19463), .B1(n19839), .B2(n19462), .ZN(
        n19450) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19465), .B1(
        n15917), .B2(n19464), .ZN(n19449) );
  OAI211_X1 U22468 ( .C1(n19703), .C2(n19523), .A(n19450), .B(n19449), .ZN(
        P2_U3073) );
  AOI22_X1 U22469 ( .A1(n19846), .A2(n19512), .B1(n19844), .B2(n19462), .ZN(
        n19452) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19465), .B1(
        n19845), .B2(n19464), .ZN(n19451) );
  OAI211_X1 U22471 ( .C1(n19849), .C2(n19461), .A(n19452), .B(n19451), .ZN(
        P2_U3074) );
  INV_X1 U22472 ( .A(n19852), .ZN(n19803) );
  AOI22_X1 U22473 ( .A1(n19800), .A2(n19463), .B1(n19850), .B2(n19462), .ZN(
        n19454) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19465), .B1(
        n19851), .B2(n19464), .ZN(n19453) );
  OAI211_X1 U22475 ( .C1(n19803), .C2(n19523), .A(n19454), .B(n19453), .ZN(
        P2_U3075) );
  AOI22_X1 U22476 ( .A1(n19804), .A2(n19463), .B1(n19462), .B2(n19856), .ZN(
        n19456) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19465), .B1(
        n19857), .B2(n19464), .ZN(n19455) );
  OAI211_X1 U22478 ( .C1(n19807), .C2(n19523), .A(n19456), .B(n19455), .ZN(
        P2_U3076) );
  AOI22_X1 U22479 ( .A1(n19676), .A2(n19463), .B1(n19462), .B2(n19862), .ZN(
        n19458) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19465), .B1(
        n19863), .B2(n19464), .ZN(n19457) );
  OAI211_X1 U22481 ( .C1(n19564), .C2(n19523), .A(n19458), .B(n19457), .ZN(
        P2_U3077) );
  INV_X1 U22482 ( .A(n19812), .ZN(n19873) );
  AOI22_X1 U22483 ( .A1(n19870), .A2(n19512), .B1(n19462), .B2(n19868), .ZN(
        n19460) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19465), .B1(
        n19869), .B2(n19464), .ZN(n19459) );
  OAI211_X1 U22485 ( .C1(n19873), .C2(n19461), .A(n19460), .B(n19459), .ZN(
        P2_U3078) );
  AOI22_X1 U22486 ( .A1(n19818), .A2(n19463), .B1(n19462), .B2(n19875), .ZN(
        n19467) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19465), .B1(
        n19876), .B2(n19464), .ZN(n19466) );
  OAI211_X1 U22488 ( .C1(n19823), .C2(n19523), .A(n19467), .B(n19466), .ZN(
        P2_U3079) );
  INV_X1 U22489 ( .A(n19468), .ZN(n19470) );
  NOR2_X1 U22490 ( .A1(n19470), .A2(n19469), .ZN(n19726) );
  AND2_X1 U22491 ( .A1(n19726), .A2(n19980), .ZN(n19480) );
  NAND2_X1 U22492 ( .A1(n19825), .A2(n19480), .ZN(n19473) );
  NOR2_X1 U22493 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19471), .ZN(
        n19474) );
  NOR2_X1 U22494 ( .A1(n12632), .A2(n19474), .ZN(n19472) );
  MUX2_X1 U22495 ( .A(n19473), .B(n19472), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19518) );
  INV_X1 U22496 ( .A(n19474), .ZN(n19515) );
  OAI22_X1 U22497 ( .A1(n19518), .A2(n19476), .B1(n19475), .B2(n19515), .ZN(
        n19477) );
  INV_X1 U22498 ( .A(n19477), .ZN(n19483) );
  AOI21_X1 U22499 ( .B1(n19523), .B2(n19534), .A(n15893), .ZN(n19481) );
  OAI21_X1 U22500 ( .B1(n12632), .B2(n20017), .A(n19825), .ZN(n19478) );
  NAND2_X1 U22501 ( .A1(n19478), .A2(n19515), .ZN(n19479) );
  OAI211_X1 U22502 ( .C1(n19481), .C2(n19480), .A(n19479), .B(n19833), .ZN(
        n19520) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19835), .ZN(n19482) );
  OAI211_X1 U22504 ( .C1(n19838), .C2(n19523), .A(n19483), .B(n19482), .ZN(
        P2_U3080) );
  OAI22_X1 U22505 ( .A1(n19518), .A2(n19485), .B1(n19484), .B2(n19515), .ZN(
        n19486) );
  INV_X1 U22506 ( .A(n19486), .ZN(n19488) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19520), .B1(
        n19512), .B2(n19700), .ZN(n19487) );
  OAI211_X1 U22508 ( .C1(n19703), .C2(n19534), .A(n19488), .B(n19487), .ZN(
        P2_U3081) );
  OAI22_X1 U22509 ( .A1(n19518), .A2(n19490), .B1(n19489), .B2(n19515), .ZN(
        n19491) );
  INV_X1 U22510 ( .A(n19491), .ZN(n19493) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19846), .ZN(n19492) );
  OAI211_X1 U22512 ( .C1(n19849), .C2(n19523), .A(n19493), .B(n19492), .ZN(
        P2_U3082) );
  OAI22_X1 U22513 ( .A1(n19518), .A2(n19495), .B1(n19494), .B2(n19515), .ZN(
        n19496) );
  INV_X1 U22514 ( .A(n19496), .ZN(n19498) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19520), .B1(
        n19512), .B2(n19800), .ZN(n19497) );
  OAI211_X1 U22516 ( .C1(n19803), .C2(n19534), .A(n19498), .B(n19497), .ZN(
        P2_U3083) );
  OAI22_X1 U22517 ( .A1(n19518), .A2(n19500), .B1(n19499), .B2(n19515), .ZN(
        n19501) );
  INV_X1 U22518 ( .A(n19501), .ZN(n19503) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19520), .B1(
        n19512), .B2(n19804), .ZN(n19502) );
  OAI211_X1 U22520 ( .C1(n19807), .C2(n19534), .A(n19503), .B(n19502), .ZN(
        P2_U3084) );
  OAI22_X1 U22521 ( .A1(n19518), .A2(n19505), .B1(n19504), .B2(n19515), .ZN(
        n19506) );
  INV_X1 U22522 ( .A(n19506), .ZN(n19508) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19520), .B1(
        n19512), .B2(n19676), .ZN(n19507) );
  OAI211_X1 U22524 ( .C1(n19564), .C2(n19534), .A(n19508), .B(n19507), .ZN(
        P2_U3085) );
  OAI22_X1 U22525 ( .A1(n19518), .A2(n19510), .B1(n19509), .B2(n19515), .ZN(
        n19511) );
  INV_X1 U22526 ( .A(n19511), .ZN(n19514) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19520), .B1(
        n19512), .B2(n19812), .ZN(n19513) );
  OAI211_X1 U22528 ( .C1(n19815), .C2(n19534), .A(n19514), .B(n19513), .ZN(
        P2_U3086) );
  OAI22_X1 U22529 ( .A1(n19518), .A2(n19517), .B1(n19516), .B2(n19515), .ZN(
        n19519) );
  INV_X1 U22530 ( .A(n19519), .ZN(n19522) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19878), .ZN(n19521) );
  OAI211_X1 U22532 ( .C1(n19884), .C2(n19523), .A(n19522), .B(n19521), .ZN(
        P2_U3087) );
  AOI22_X1 U22533 ( .A1(n19569), .A2(n19835), .B1(n19544), .B2(n19827), .ZN(
        n19525) );
  AOI22_X1 U22534 ( .A1(n19326), .A2(n19540), .B1(n19539), .B2(n19664), .ZN(
        n19524) );
  OAI211_X1 U22535 ( .C1(n19527), .C2(n19526), .A(n19525), .B(n19524), .ZN(
        P2_U3088) );
  AOI22_X1 U22536 ( .A1(n19840), .A2(n19569), .B1(n19839), .B2(n19544), .ZN(
        n19529) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19541), .B1(
        n15917), .B2(n19540), .ZN(n19528) );
  OAI211_X1 U22538 ( .C1(n19843), .C2(n19534), .A(n19529), .B(n19528), .ZN(
        P2_U3089) );
  AOI22_X1 U22539 ( .A1(n19846), .A2(n19569), .B1(n19844), .B2(n19544), .ZN(
        n19531) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19541), .B1(
        n19845), .B2(n19540), .ZN(n19530) );
  OAI211_X1 U22541 ( .C1(n19849), .C2(n19534), .A(n19531), .B(n19530), .ZN(
        P2_U3090) );
  AOI22_X1 U22542 ( .A1(n19858), .A2(n19569), .B1(n19544), .B2(n19856), .ZN(
        n19533) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19541), .B1(
        n19857), .B2(n19540), .ZN(n19532) );
  OAI211_X1 U22544 ( .C1(n19861), .C2(n19534), .A(n19533), .B(n19532), .ZN(
        P2_U3092) );
  AOI22_X1 U22545 ( .A1(n19676), .A2(n19539), .B1(n19544), .B2(n19862), .ZN(
        n19536) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19541), .B1(
        n19863), .B2(n19540), .ZN(n19535) );
  OAI211_X1 U22547 ( .C1(n19564), .C2(n19559), .A(n19536), .B(n19535), .ZN(
        P2_U3093) );
  AOI22_X1 U22548 ( .A1(n19812), .A2(n19539), .B1(n19544), .B2(n19868), .ZN(
        n19538) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19541), .B1(
        n19869), .B2(n19540), .ZN(n19537) );
  OAI211_X1 U22550 ( .C1(n19815), .C2(n19559), .A(n19538), .B(n19537), .ZN(
        P2_U3094) );
  AOI22_X1 U22551 ( .A1(n19818), .A2(n19539), .B1(n19544), .B2(n19875), .ZN(
        n19543) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19541), .B1(
        n19876), .B2(n19540), .ZN(n19542) );
  OAI211_X1 U22553 ( .C1(n19823), .C2(n19559), .A(n19543), .B(n19542), .ZN(
        P2_U3095) );
  NOR2_X1 U22554 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19578), .ZN(
        n19567) );
  NOR2_X1 U22555 ( .A1(n19544), .A2(n19567), .ZN(n19548) );
  OAI21_X1 U22556 ( .B1(n12625), .B2(n19567), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19545) );
  OAI21_X1 U22557 ( .B1(n19548), .B2(n19974), .A(n19545), .ZN(n19568) );
  AOI22_X1 U22558 ( .A1(n19568), .A2(n19326), .B1(n19827), .B2(n19567), .ZN(
        n19552) );
  OAI21_X1 U22559 ( .B1(n19569), .B2(n19594), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19549) );
  AOI211_X1 U22560 ( .C1(n12625), .C2(n19825), .A(n19971), .B(n19567), .ZN(
        n19547) );
  AOI211_X1 U22561 ( .C1(n19549), .C2(n19548), .A(n19547), .B(n19576), .ZN(
        n19550) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19570), .B1(
        n19594), .B2(n19835), .ZN(n19551) );
  OAI211_X1 U22563 ( .C1(n19838), .C2(n19559), .A(n19552), .B(n19551), .ZN(
        P2_U3096) );
  AOI22_X1 U22564 ( .A1(n19568), .A2(n15917), .B1(n19839), .B2(n19567), .ZN(
        n19554) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19700), .ZN(n19553) );
  OAI211_X1 U22566 ( .C1(n19703), .C2(n19601), .A(n19554), .B(n19553), .ZN(
        P2_U3097) );
  AOI22_X1 U22567 ( .A1(n19568), .A2(n19845), .B1(n19844), .B2(n19567), .ZN(
        n19556) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19796), .ZN(n19555) );
  OAI211_X1 U22569 ( .C1(n19799), .C2(n19601), .A(n19556), .B(n19555), .ZN(
        P2_U3098) );
  AOI22_X1 U22570 ( .A1(n19568), .A2(n19851), .B1(n19850), .B2(n19567), .ZN(
        n19558) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19570), .B1(
        n19594), .B2(n19852), .ZN(n19557) );
  OAI211_X1 U22572 ( .C1(n19855), .C2(n19559), .A(n19558), .B(n19557), .ZN(
        P2_U3099) );
  AOI22_X1 U22573 ( .A1(n19568), .A2(n19857), .B1(n19856), .B2(n19567), .ZN(
        n19561) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19804), .ZN(n19560) );
  OAI211_X1 U22575 ( .C1(n19807), .C2(n19601), .A(n19561), .B(n19560), .ZN(
        P2_U3100) );
  AOI22_X1 U22576 ( .A1(n19568), .A2(n19863), .B1(n19862), .B2(n19567), .ZN(
        n19563) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19676), .ZN(n19562) );
  OAI211_X1 U22578 ( .C1(n19564), .C2(n19601), .A(n19563), .B(n19562), .ZN(
        P2_U3101) );
  AOI22_X1 U22579 ( .A1(n19568), .A2(n19869), .B1(n19868), .B2(n19567), .ZN(
        n19566) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19812), .ZN(n19565) );
  OAI211_X1 U22581 ( .C1(n19815), .C2(n19601), .A(n19566), .B(n19565), .ZN(
        P2_U3102) );
  AOI22_X1 U22582 ( .A1(n19568), .A2(n19876), .B1(n19875), .B2(n19567), .ZN(
        n19572) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19818), .ZN(n19571) );
  OAI211_X1 U22584 ( .C1(n19823), .C2(n19601), .A(n19572), .B(n19571), .ZN(
        P2_U3103) );
  NOR3_X1 U22585 ( .A1(n19573), .A2(n19609), .A3(n20017), .ZN(n19577) );
  AOI211_X2 U22586 ( .C1(n19578), .C2(n20017), .A(n19574), .B(n19577), .ZN(
        n19597) );
  AOI22_X1 U22587 ( .A1(n19597), .A2(n19326), .B1(n19609), .B2(n19827), .ZN(
        n19583) );
  INV_X1 U22588 ( .A(n19973), .ZN(n19828) );
  NAND2_X1 U22589 ( .A1(n19575), .A2(n19828), .ZN(n19579) );
  AOI211_X1 U22590 ( .C1(n19579), .C2(n19578), .A(n19577), .B(n19576), .ZN(
        n19580) );
  OAI21_X1 U22591 ( .B1(n19609), .B2(n19825), .A(n19580), .ZN(n19598) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19598), .B1(
        n19624), .B2(n19835), .ZN(n19582) );
  OAI211_X1 U22593 ( .C1(n19838), .C2(n19601), .A(n19583), .B(n19582), .ZN(
        P2_U3104) );
  AOI22_X1 U22594 ( .A1(n19597), .A2(n15917), .B1(n19609), .B2(n19839), .ZN(
        n19585) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19598), .B1(
        n19594), .B2(n19700), .ZN(n19584) );
  OAI211_X1 U22596 ( .C1(n19703), .C2(n19632), .A(n19585), .B(n19584), .ZN(
        P2_U3105) );
  AOI22_X1 U22597 ( .A1(n19597), .A2(n19845), .B1(n19609), .B2(n19844), .ZN(
        n19587) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19598), .B1(
        n19594), .B2(n19796), .ZN(n19586) );
  OAI211_X1 U22599 ( .C1(n19799), .C2(n19632), .A(n19587), .B(n19586), .ZN(
        P2_U3106) );
  AOI22_X1 U22600 ( .A1(n19597), .A2(n19851), .B1(n19609), .B2(n19850), .ZN(
        n19589) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19598), .B1(
        n19624), .B2(n19852), .ZN(n19588) );
  OAI211_X1 U22602 ( .C1(n19855), .C2(n19601), .A(n19589), .B(n19588), .ZN(
        P2_U3107) );
  AOI22_X1 U22603 ( .A1(n19597), .A2(n19857), .B1(n19609), .B2(n19856), .ZN(
        n19591) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19598), .B1(
        n19624), .B2(n19858), .ZN(n19590) );
  OAI211_X1 U22605 ( .C1(n19861), .C2(n19601), .A(n19591), .B(n19590), .ZN(
        P2_U3108) );
  AOI22_X1 U22606 ( .A1(n19597), .A2(n19863), .B1(n19609), .B2(n19862), .ZN(
        n19593) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19598), .B1(
        n19624), .B2(n19864), .ZN(n19592) );
  OAI211_X1 U22608 ( .C1(n19867), .C2(n19601), .A(n19593), .B(n19592), .ZN(
        P2_U3109) );
  AOI22_X1 U22609 ( .A1(n19597), .A2(n19869), .B1(n19609), .B2(n19868), .ZN(
        n19596) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19598), .B1(
        n19594), .B2(n19812), .ZN(n19595) );
  OAI211_X1 U22611 ( .C1(n19815), .C2(n19632), .A(n19596), .B(n19595), .ZN(
        P2_U3110) );
  AOI22_X1 U22612 ( .A1(n19597), .A2(n19876), .B1(n19609), .B2(n19875), .ZN(
        n19600) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19598), .B1(
        n19624), .B2(n19878), .ZN(n19599) );
  OAI211_X1 U22614 ( .C1(n19884), .C2(n19601), .A(n19600), .B(n19599), .ZN(
        P2_U3111) );
  NAND2_X1 U22615 ( .A1(n19690), .A2(n19996), .ZN(n19640) );
  NOR2_X1 U22616 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19640), .ZN(
        n19627) );
  AOI22_X1 U22617 ( .A1(n19658), .A2(n19835), .B1(n19627), .B2(n19827), .ZN(
        n19613) );
  NAND2_X1 U22618 ( .A1(n19632), .A2(n19971), .ZN(n19604) );
  INV_X1 U22619 ( .A(n19970), .ZN(n19603) );
  OAI21_X1 U22620 ( .B1(n19604), .B2(n19658), .A(n19603), .ZN(n19608) );
  OAI21_X1 U22621 ( .B1(n12631), .B2(n20017), .A(n19825), .ZN(n19605) );
  AOI21_X1 U22622 ( .B1(n19608), .B2(n19606), .A(n19605), .ZN(n19607) );
  OAI21_X1 U22623 ( .B1(n19627), .B2(n19607), .A(n19833), .ZN(n19629) );
  OAI21_X1 U22624 ( .B1(n19609), .B2(n19627), .A(n19608), .ZN(n19611) );
  OAI21_X1 U22625 ( .B1(n12631), .B2(n19627), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19610) );
  NAND2_X1 U22626 ( .A1(n19611), .A2(n19610), .ZN(n19628) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19629), .B1(
        n19326), .B2(n19628), .ZN(n19612) );
  OAI211_X1 U22628 ( .C1(n19838), .C2(n19632), .A(n19613), .B(n19612), .ZN(
        P2_U3112) );
  AOI22_X1 U22629 ( .A1(n19840), .A2(n19658), .B1(n19839), .B2(n19627), .ZN(
        n19615) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n15917), .ZN(n19614) );
  OAI211_X1 U22631 ( .C1(n19843), .C2(n19632), .A(n19615), .B(n19614), .ZN(
        P2_U3113) );
  AOI22_X1 U22632 ( .A1(n19846), .A2(n19658), .B1(n19844), .B2(n19627), .ZN(
        n19617) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19845), .ZN(n19616) );
  OAI211_X1 U22634 ( .C1(n19849), .C2(n19632), .A(n19617), .B(n19616), .ZN(
        P2_U3114) );
  AOI22_X1 U22635 ( .A1(n19852), .A2(n19658), .B1(n19850), .B2(n19627), .ZN(
        n19619) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19851), .ZN(n19618) );
  OAI211_X1 U22637 ( .C1(n19855), .C2(n19632), .A(n19619), .B(n19618), .ZN(
        P2_U3115) );
  AOI22_X1 U22638 ( .A1(n19804), .A2(n19624), .B1(n19856), .B2(n19627), .ZN(
        n19621) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19857), .ZN(n19620) );
  OAI211_X1 U22640 ( .C1(n19807), .C2(n19654), .A(n19621), .B(n19620), .ZN(
        P2_U3116) );
  AOI22_X1 U22641 ( .A1(n19864), .A2(n19658), .B1(n19627), .B2(n19862), .ZN(
        n19623) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19863), .ZN(n19622) );
  OAI211_X1 U22643 ( .C1(n19867), .C2(n19632), .A(n19623), .B(n19622), .ZN(
        P2_U3117) );
  AOI22_X1 U22644 ( .A1(n19812), .A2(n19624), .B1(n19627), .B2(n19868), .ZN(
        n19626) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19869), .ZN(n19625) );
  OAI211_X1 U22646 ( .C1(n19815), .C2(n19654), .A(n19626), .B(n19625), .ZN(
        P2_U3118) );
  AOI22_X1 U22647 ( .A1(n19878), .A2(n19658), .B1(n19627), .B2(n19875), .ZN(
        n19631) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19876), .ZN(n19630) );
  OAI211_X1 U22649 ( .C1(n19884), .C2(n19632), .A(n19631), .B(n19630), .ZN(
        P2_U3119) );
  INV_X1 U22650 ( .A(n19690), .ZN(n19633) );
  NOR2_X1 U22651 ( .A1(n19634), .A2(n19633), .ZN(n19657) );
  AOI22_X1 U22652 ( .A1(n19682), .A2(n19835), .B1(n19827), .B2(n19657), .ZN(
        n19643) );
  NOR2_X1 U22653 ( .A1(n19972), .A2(n15893), .ZN(n19829) );
  AOI21_X1 U22654 ( .B1(n19829), .B2(n19635), .A(n19974), .ZN(n19638) );
  NOR2_X1 U22655 ( .A1(n19636), .A2(n19657), .ZN(n19639) );
  AOI22_X1 U22656 ( .A1(n19638), .A2(n19640), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19639), .ZN(n19637) );
  OAI211_X1 U22657 ( .C1(n19657), .C2(n19825), .A(n19637), .B(n19833), .ZN(
        n19660) );
  INV_X1 U22658 ( .A(n19638), .ZN(n19641) );
  OAI22_X1 U22659 ( .A1(n19641), .A2(n19640), .B1(n19639), .B2(n20017), .ZN(
        n19659) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19660), .B1(
        n19326), .B2(n19659), .ZN(n19642) );
  OAI211_X1 U22661 ( .C1(n19838), .C2(n19654), .A(n19643), .B(n19642), .ZN(
        P2_U3120) );
  INV_X1 U22662 ( .A(n19682), .ZN(n19663) );
  AOI22_X1 U22663 ( .A1(n19700), .A2(n19658), .B1(n19839), .B2(n19657), .ZN(
        n19645) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19660), .B1(
        n15917), .B2(n19659), .ZN(n19644) );
  OAI211_X1 U22665 ( .C1(n19703), .C2(n19663), .A(n19645), .B(n19644), .ZN(
        P2_U3121) );
  AOI22_X1 U22666 ( .A1(n19796), .A2(n19658), .B1(n19844), .B2(n19657), .ZN(
        n19647) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19660), .B1(
        n19845), .B2(n19659), .ZN(n19646) );
  OAI211_X1 U22668 ( .C1(n19799), .C2(n19663), .A(n19647), .B(n19646), .ZN(
        P2_U3122) );
  AOI22_X1 U22669 ( .A1(n19852), .A2(n19682), .B1(n19850), .B2(n19657), .ZN(
        n19649) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19660), .B1(
        n19851), .B2(n19659), .ZN(n19648) );
  OAI211_X1 U22671 ( .C1(n19855), .C2(n19654), .A(n19649), .B(n19648), .ZN(
        P2_U3123) );
  AOI22_X1 U22672 ( .A1(n19804), .A2(n19658), .B1(n19856), .B2(n19657), .ZN(
        n19651) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19660), .B1(
        n19857), .B2(n19659), .ZN(n19650) );
  OAI211_X1 U22674 ( .C1(n19807), .C2(n19663), .A(n19651), .B(n19650), .ZN(
        P2_U3124) );
  AOI22_X1 U22675 ( .A1(n19864), .A2(n19682), .B1(n19862), .B2(n19657), .ZN(
        n19653) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19660), .B1(
        n19863), .B2(n19659), .ZN(n19652) );
  OAI211_X1 U22677 ( .C1(n19867), .C2(n19654), .A(n19653), .B(n19652), .ZN(
        P2_U3125) );
  AOI22_X1 U22678 ( .A1(n19812), .A2(n19658), .B1(n19868), .B2(n19657), .ZN(
        n19656) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19660), .B1(
        n19869), .B2(n19659), .ZN(n19655) );
  OAI211_X1 U22680 ( .C1(n19815), .C2(n19663), .A(n19656), .B(n19655), .ZN(
        P2_U3126) );
  AOI22_X1 U22681 ( .A1(n19818), .A2(n19658), .B1(n19875), .B2(n19657), .ZN(
        n19662) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19660), .B1(
        n19876), .B2(n19659), .ZN(n19661) );
  OAI211_X1 U22683 ( .C1(n19823), .C2(n19663), .A(n19662), .B(n19661), .ZN(
        P2_U3127) );
  INV_X1 U22684 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19667) );
  AOI22_X1 U22685 ( .A1(n19664), .A2(n19682), .B1(n19681), .B2(n19827), .ZN(
        n19666) );
  AOI22_X1 U22686 ( .A1(n19326), .A2(n19683), .B1(n19717), .B2(n19835), .ZN(
        n19665) );
  OAI211_X1 U22687 ( .C1(n19687), .C2(n19667), .A(n19666), .B(n19665), .ZN(
        P2_U3128) );
  INV_X1 U22688 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n19670) );
  AOI22_X1 U22689 ( .A1(n19796), .A2(n19682), .B1(n19681), .B2(n19844), .ZN(
        n19669) );
  AOI22_X1 U22690 ( .A1(n19845), .A2(n19683), .B1(n19717), .B2(n19846), .ZN(
        n19668) );
  OAI211_X1 U22691 ( .C1(n19687), .C2(n19670), .A(n19669), .B(n19668), .ZN(
        P2_U3130) );
  AOI22_X1 U22692 ( .A1(n19852), .A2(n19717), .B1(n19681), .B2(n19850), .ZN(
        n19672) );
  AOI22_X1 U22693 ( .A1(n19851), .A2(n19683), .B1(n19682), .B2(n19800), .ZN(
        n19671) );
  OAI211_X1 U22694 ( .C1(n19687), .C2(n12587), .A(n19672), .B(n19671), .ZN(
        P2_U3131) );
  INV_X1 U22695 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n19675) );
  AOI22_X1 U22696 ( .A1(n19804), .A2(n19682), .B1(n19681), .B2(n19856), .ZN(
        n19674) );
  AOI22_X1 U22697 ( .A1(n19857), .A2(n19683), .B1(n19717), .B2(n19858), .ZN(
        n19673) );
  OAI211_X1 U22698 ( .C1(n19687), .C2(n19675), .A(n19674), .B(n19673), .ZN(
        P2_U3132) );
  AOI22_X1 U22699 ( .A1(n19864), .A2(n19717), .B1(n19681), .B2(n19862), .ZN(
        n19678) );
  AOI22_X1 U22700 ( .A1(n19863), .A2(n19683), .B1(n19682), .B2(n19676), .ZN(
        n19677) );
  OAI211_X1 U22701 ( .C1(n19687), .C2(n12628), .A(n19678), .B(n19677), .ZN(
        P2_U3133) );
  AOI22_X1 U22702 ( .A1(n19870), .A2(n19717), .B1(n19681), .B2(n19868), .ZN(
        n19680) );
  AOI22_X1 U22703 ( .A1(n19869), .A2(n19683), .B1(n19682), .B2(n19812), .ZN(
        n19679) );
  OAI211_X1 U22704 ( .C1(n19687), .C2(n15100), .A(n19680), .B(n19679), .ZN(
        P2_U3134) );
  INV_X1 U22705 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19686) );
  AOI22_X1 U22706 ( .A1(n19818), .A2(n19682), .B1(n19681), .B2(n19875), .ZN(
        n19685) );
  AOI22_X1 U22707 ( .A1(n19876), .A2(n19683), .B1(n19717), .B2(n19878), .ZN(
        n19684) );
  OAI211_X1 U22708 ( .C1(n19687), .C2(n19686), .A(n19685), .B(n19684), .ZN(
        P2_U3135) );
  INV_X1 U22709 ( .A(n19688), .ZN(n19689) );
  NAND2_X1 U22710 ( .A1(n19689), .A2(n19690), .ZN(n19692) );
  NAND3_X1 U22711 ( .A1(n12619), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19692), 
        .ZN(n19695) );
  NAND2_X1 U22712 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19690), .ZN(
        n19693) );
  OAI21_X1 U22713 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19693), .A(n20017), 
        .ZN(n19691) );
  INV_X1 U22714 ( .A(n19692), .ZN(n19715) );
  AOI22_X1 U22715 ( .A1(n19716), .A2(n19326), .B1(n19827), .B2(n19715), .ZN(
        n19699) );
  NAND2_X1 U22716 ( .A1(n19829), .A2(n19825), .ZN(n19754) );
  NOR2_X1 U22717 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19825), .ZN(
        n20003) );
  OAI22_X1 U22718 ( .A1(n19694), .A2(n19754), .B1(n20003), .B2(n19693), .ZN(
        n19696) );
  NAND3_X1 U22719 ( .A1(n19696), .A2(n19833), .A3(n19695), .ZN(n19718) );
  INV_X1 U22720 ( .A(n19750), .ZN(n19725) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19718), .B1(
        n19725), .B2(n19835), .ZN(n19698) );
  OAI211_X1 U22722 ( .C1(n19838), .C2(n19714), .A(n19699), .B(n19698), .ZN(
        P2_U3136) );
  AOI22_X1 U22723 ( .A1(n19716), .A2(n15917), .B1(n19839), .B2(n19715), .ZN(
        n19702) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19700), .ZN(n19701) );
  OAI211_X1 U22725 ( .C1(n19703), .C2(n19750), .A(n19702), .B(n19701), .ZN(
        P2_U3137) );
  AOI22_X1 U22726 ( .A1(n19716), .A2(n19845), .B1(n19844), .B2(n19715), .ZN(
        n19705) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19796), .ZN(n19704) );
  OAI211_X1 U22728 ( .C1(n19799), .C2(n19750), .A(n19705), .B(n19704), .ZN(
        P2_U3138) );
  AOI22_X1 U22729 ( .A1(n19716), .A2(n19851), .B1(n19850), .B2(n19715), .ZN(
        n19707) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19800), .ZN(n19706) );
  OAI211_X1 U22731 ( .C1(n19803), .C2(n19750), .A(n19707), .B(n19706), .ZN(
        P2_U3139) );
  AOI22_X1 U22732 ( .A1(n19716), .A2(n19857), .B1(n19856), .B2(n19715), .ZN(
        n19709) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19718), .B1(
        n19725), .B2(n19858), .ZN(n19708) );
  OAI211_X1 U22734 ( .C1(n19861), .C2(n19714), .A(n19709), .B(n19708), .ZN(
        P2_U3140) );
  AOI22_X1 U22735 ( .A1(n19716), .A2(n19863), .B1(n19862), .B2(n19715), .ZN(
        n19711) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19718), .B1(
        n19725), .B2(n19864), .ZN(n19710) );
  OAI211_X1 U22737 ( .C1(n19867), .C2(n19714), .A(n19711), .B(n19710), .ZN(
        P2_U3141) );
  AOI22_X1 U22738 ( .A1(n19716), .A2(n19869), .B1(n19868), .B2(n19715), .ZN(
        n19713) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19718), .B1(
        n19725), .B2(n19870), .ZN(n19712) );
  OAI211_X1 U22740 ( .C1(n19873), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P2_U3142) );
  AOI22_X1 U22741 ( .A1(n19716), .A2(n19876), .B1(n19875), .B2(n19715), .ZN(
        n19720) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19718), .B1(
        n19717), .B2(n19818), .ZN(n19719) );
  OAI211_X1 U22743 ( .C1(n19823), .C2(n19750), .A(n19720), .B(n19719), .ZN(
        P2_U3143) );
  NAND3_X1 U22744 ( .A1(n19996), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19753) );
  NOR2_X1 U22745 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19753), .ZN(
        n19745) );
  NOR2_X1 U22746 ( .A1(n19721), .A2(n19745), .ZN(n19727) );
  INV_X1 U22747 ( .A(n19722), .ZN(n19724) );
  INV_X1 U22748 ( .A(n19726), .ZN(n19723) );
  OAI22_X1 U22749 ( .A1(n19727), .A2(n20017), .B1(n19724), .B2(n19723), .ZN(
        n19746) );
  AOI22_X1 U22750 ( .A1(n19746), .A2(n19326), .B1(n19827), .B2(n19745), .ZN(
        n19732) );
  NOR2_X2 U22751 ( .A1(n19780), .A2(n19755), .ZN(n19772) );
  OAI21_X1 U22752 ( .B1(n19772), .B2(n19725), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19729) );
  NAND2_X1 U22753 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19726), .ZN(
        n19728) );
  AOI22_X1 U22754 ( .A1(n19729), .A2(n19728), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19727), .ZN(n19730) );
  OAI211_X1 U22755 ( .C1(n19745), .C2(n19825), .A(n19730), .B(n19833), .ZN(
        n19747) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19835), .ZN(n19731) );
  OAI211_X1 U22757 ( .C1(n19838), .C2(n19750), .A(n19732), .B(n19731), .ZN(
        P2_U3144) );
  AOI22_X1 U22758 ( .A1(n19746), .A2(n15917), .B1(n19839), .B2(n19745), .ZN(
        n19734) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19840), .ZN(n19733) );
  OAI211_X1 U22760 ( .C1(n19843), .C2(n19750), .A(n19734), .B(n19733), .ZN(
        P2_U3145) );
  AOI22_X1 U22761 ( .A1(n19746), .A2(n19845), .B1(n19844), .B2(n19745), .ZN(
        n19736) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19846), .ZN(n19735) );
  OAI211_X1 U22763 ( .C1(n19849), .C2(n19750), .A(n19736), .B(n19735), .ZN(
        P2_U3146) );
  AOI22_X1 U22764 ( .A1(n19746), .A2(n19851), .B1(n19850), .B2(n19745), .ZN(
        n19738) );
  AOI22_X1 U22765 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19852), .ZN(n19737) );
  OAI211_X1 U22766 ( .C1(n19855), .C2(n19750), .A(n19738), .B(n19737), .ZN(
        P2_U3147) );
  AOI22_X1 U22767 ( .A1(n19746), .A2(n19857), .B1(n19856), .B2(n19745), .ZN(
        n19740) );
  AOI22_X1 U22768 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19858), .ZN(n19739) );
  OAI211_X1 U22769 ( .C1(n19861), .C2(n19750), .A(n19740), .B(n19739), .ZN(
        P2_U3148) );
  AOI22_X1 U22770 ( .A1(n19746), .A2(n19863), .B1(n19862), .B2(n19745), .ZN(
        n19742) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19864), .ZN(n19741) );
  OAI211_X1 U22772 ( .C1(n19867), .C2(n19750), .A(n19742), .B(n19741), .ZN(
        P2_U3149) );
  AOI22_X1 U22773 ( .A1(n19746), .A2(n19869), .B1(n19868), .B2(n19745), .ZN(
        n19744) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19870), .ZN(n19743) );
  OAI211_X1 U22775 ( .C1(n19873), .C2(n19750), .A(n19744), .B(n19743), .ZN(
        P2_U3150) );
  AOI22_X1 U22776 ( .A1(n19746), .A2(n19876), .B1(n19875), .B2(n19745), .ZN(
        n19749) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19747), .B1(
        n19772), .B2(n19878), .ZN(n19748) );
  OAI211_X1 U22778 ( .C1(n19884), .C2(n19750), .A(n19749), .B(n19748), .ZN(
        P2_U3151) );
  NOR2_X1 U22779 ( .A1(n20006), .A2(n19753), .ZN(n19783) );
  INV_X1 U22780 ( .A(n19783), .ZN(n19751) );
  NAND3_X1 U22781 ( .A1(n12620), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19751), 
        .ZN(n19756) );
  OAI21_X1 U22782 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19753), .A(n20017), 
        .ZN(n19752) );
  AOI22_X1 U22783 ( .A1(n19775), .A2(n19326), .B1(n19827), .B2(n19783), .ZN(
        n19761) );
  OAI22_X1 U22784 ( .A1(n19755), .A2(n19754), .B1(n20003), .B2(n19753), .ZN(
        n19757) );
  NAND3_X1 U22785 ( .A1(n19757), .A2(n19833), .A3(n19756), .ZN(n19776) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19776), .B1(
        n19817), .B2(n19835), .ZN(n19760) );
  OAI211_X1 U22787 ( .C1(n19838), .C2(n19779), .A(n19761), .B(n19760), .ZN(
        P2_U3152) );
  AOI22_X1 U22788 ( .A1(n19775), .A2(n15917), .B1(n19839), .B2(n19783), .ZN(
        n19763) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19776), .B1(
        n19817), .B2(n19840), .ZN(n19762) );
  OAI211_X1 U22790 ( .C1(n19843), .C2(n19779), .A(n19763), .B(n19762), .ZN(
        P2_U3153) );
  AOI22_X1 U22791 ( .A1(n19775), .A2(n19845), .B1(n19844), .B2(n19783), .ZN(
        n19765) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19776), .B1(
        n19772), .B2(n19796), .ZN(n19764) );
  OAI211_X1 U22793 ( .C1(n19799), .C2(n19811), .A(n19765), .B(n19764), .ZN(
        P2_U3154) );
  AOI22_X1 U22794 ( .A1(n19775), .A2(n19851), .B1(n19850), .B2(n19783), .ZN(
        n19767) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19776), .B1(
        n19772), .B2(n19800), .ZN(n19766) );
  OAI211_X1 U22796 ( .C1(n19803), .C2(n19811), .A(n19767), .B(n19766), .ZN(
        P2_U3155) );
  AOI22_X1 U22797 ( .A1(n19775), .A2(n19857), .B1(n19856), .B2(n19783), .ZN(
        n19769) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19776), .B1(
        n19817), .B2(n19858), .ZN(n19768) );
  OAI211_X1 U22799 ( .C1(n19861), .C2(n19779), .A(n19769), .B(n19768), .ZN(
        P2_U3156) );
  AOI22_X1 U22800 ( .A1(n19775), .A2(n19863), .B1(n19862), .B2(n19783), .ZN(
        n19771) );
  AOI22_X1 U22801 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19776), .B1(
        n19817), .B2(n19864), .ZN(n19770) );
  OAI211_X1 U22802 ( .C1(n19867), .C2(n19779), .A(n19771), .B(n19770), .ZN(
        P2_U3157) );
  AOI22_X1 U22803 ( .A1(n19775), .A2(n19869), .B1(n19868), .B2(n19783), .ZN(
        n19774) );
  AOI22_X1 U22804 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19776), .B1(
        n19772), .B2(n19812), .ZN(n19773) );
  OAI211_X1 U22805 ( .C1(n19815), .C2(n19811), .A(n19774), .B(n19773), .ZN(
        P2_U3158) );
  AOI22_X1 U22806 ( .A1(n19775), .A2(n19876), .B1(n19875), .B2(n19783), .ZN(
        n19778) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19776), .B1(
        n19817), .B2(n19878), .ZN(n19777) );
  OAI211_X1 U22808 ( .C1(n19884), .C2(n19779), .A(n19778), .B(n19777), .ZN(
        P2_U3159) );
  NAND2_X1 U22809 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19781), .ZN(
        n19831) );
  NOR2_X1 U22810 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19831), .ZN(
        n19816) );
  AOI22_X1 U22811 ( .A1(n19808), .A2(n19835), .B1(n19827), .B2(n19816), .ZN(
        n19793) );
  NOR3_X1 U22812 ( .A1(n19817), .A2(n19808), .A3(n19974), .ZN(n19782) );
  NOR2_X1 U22813 ( .A1(n19782), .A2(n19970), .ZN(n19791) );
  NOR2_X1 U22814 ( .A1(n19816), .A2(n19783), .ZN(n19790) );
  INV_X1 U22815 ( .A(n19790), .ZN(n19787) );
  INV_X1 U22816 ( .A(n19816), .ZN(n19784) );
  OAI211_X1 U22817 ( .C1(n19785), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19974), 
        .B(n19784), .ZN(n19786) );
  OAI211_X1 U22818 ( .C1(n19791), .C2(n19787), .A(n19833), .B(n19786), .ZN(
        n19820) );
  OAI21_X1 U22819 ( .B1(n19788), .B2(n19816), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19789) );
  AOI22_X1 U22820 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19820), .B1(
        n19326), .B2(n19819), .ZN(n19792) );
  OAI211_X1 U22821 ( .C1(n19838), .C2(n19811), .A(n19793), .B(n19792), .ZN(
        P2_U3160) );
  AOI22_X1 U22822 ( .A1(n19840), .A2(n19808), .B1(n19839), .B2(n19816), .ZN(
        n19795) );
  AOI22_X1 U22823 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19820), .B1(
        n15917), .B2(n19819), .ZN(n19794) );
  OAI211_X1 U22824 ( .C1(n19843), .C2(n19811), .A(n19795), .B(n19794), .ZN(
        P2_U3161) );
  AOI22_X1 U22825 ( .A1(n19796), .A2(n19817), .B1(n19844), .B2(n19816), .ZN(
        n19798) );
  AOI22_X1 U22826 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19820), .B1(
        n19845), .B2(n19819), .ZN(n19797) );
  OAI211_X1 U22827 ( .C1(n19799), .C2(n19883), .A(n19798), .B(n19797), .ZN(
        P2_U3162) );
  AOI22_X1 U22828 ( .A1(n19800), .A2(n19817), .B1(n19850), .B2(n19816), .ZN(
        n19802) );
  AOI22_X1 U22829 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19820), .B1(
        n19851), .B2(n19819), .ZN(n19801) );
  OAI211_X1 U22830 ( .C1(n19803), .C2(n19883), .A(n19802), .B(n19801), .ZN(
        P2_U3163) );
  AOI22_X1 U22831 ( .A1(n19804), .A2(n19817), .B1(n19856), .B2(n19816), .ZN(
        n19806) );
  AOI22_X1 U22832 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19820), .B1(
        n19857), .B2(n19819), .ZN(n19805) );
  OAI211_X1 U22833 ( .C1(n19807), .C2(n19883), .A(n19806), .B(n19805), .ZN(
        P2_U3164) );
  AOI22_X1 U22834 ( .A1(n19864), .A2(n19808), .B1(n19862), .B2(n19816), .ZN(
        n19810) );
  AOI22_X1 U22835 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19820), .B1(
        n19863), .B2(n19819), .ZN(n19809) );
  OAI211_X1 U22836 ( .C1(n19867), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P2_U3165) );
  AOI22_X1 U22837 ( .A1(n19812), .A2(n19817), .B1(n19868), .B2(n19816), .ZN(
        n19814) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19820), .B1(
        n19869), .B2(n19819), .ZN(n19813) );
  OAI211_X1 U22839 ( .C1(n19815), .C2(n19883), .A(n19814), .B(n19813), .ZN(
        P2_U3166) );
  AOI22_X1 U22840 ( .A1(n19818), .A2(n19817), .B1(n19875), .B2(n19816), .ZN(
        n19822) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19820), .B1(
        n19876), .B2(n19819), .ZN(n19821) );
  OAI211_X1 U22842 ( .C1(n19823), .C2(n19883), .A(n19822), .B(n19821), .ZN(
        P2_U3167) );
  NOR3_X1 U22843 ( .A1(n12634), .A2(n19874), .A3(n20017), .ZN(n19830) );
  INV_X1 U22844 ( .A(n19831), .ZN(n19824) );
  AOI21_X1 U22845 ( .B1(n19825), .B2(n19824), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19826) );
  NOR2_X1 U22846 ( .A1(n19830), .A2(n19826), .ZN(n19877) );
  AOI22_X1 U22847 ( .A1(n19877), .A2(n19326), .B1(n19827), .B2(n19874), .ZN(
        n19837) );
  NAND2_X1 U22848 ( .A1(n19829), .A2(n19828), .ZN(n19832) );
  AOI21_X1 U22849 ( .B1(n19832), .B2(n19831), .A(n19830), .ZN(n19834) );
  OAI211_X1 U22850 ( .C1(n19874), .C2(n19825), .A(n19834), .B(n19833), .ZN(
        n19880) );
  AOI22_X1 U22851 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19835), .ZN(n19836) );
  OAI211_X1 U22852 ( .C1(n19838), .C2(n19883), .A(n19837), .B(n19836), .ZN(
        P2_U3168) );
  AOI22_X1 U22853 ( .A1(n19877), .A2(n15917), .B1(n19839), .B2(n19874), .ZN(
        n19842) );
  AOI22_X1 U22854 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19840), .ZN(n19841) );
  OAI211_X1 U22855 ( .C1(n19843), .C2(n19883), .A(n19842), .B(n19841), .ZN(
        P2_U3169) );
  AOI22_X1 U22856 ( .A1(n19877), .A2(n19845), .B1(n19844), .B2(n19874), .ZN(
        n19848) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19846), .ZN(n19847) );
  OAI211_X1 U22858 ( .C1(n19849), .C2(n19883), .A(n19848), .B(n19847), .ZN(
        P2_U3170) );
  AOI22_X1 U22859 ( .A1(n19877), .A2(n19851), .B1(n19850), .B2(n19874), .ZN(
        n19854) );
  AOI22_X1 U22860 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19852), .ZN(n19853) );
  OAI211_X1 U22861 ( .C1(n19855), .C2(n19883), .A(n19854), .B(n19853), .ZN(
        P2_U3171) );
  AOI22_X1 U22862 ( .A1(n19877), .A2(n19857), .B1(n19856), .B2(n19874), .ZN(
        n19860) );
  AOI22_X1 U22863 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19858), .ZN(n19859) );
  OAI211_X1 U22864 ( .C1(n19861), .C2(n19883), .A(n19860), .B(n19859), .ZN(
        P2_U3172) );
  AOI22_X1 U22865 ( .A1(n19877), .A2(n19863), .B1(n19862), .B2(n19874), .ZN(
        n19866) );
  AOI22_X1 U22866 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19864), .ZN(n19865) );
  OAI211_X1 U22867 ( .C1(n19867), .C2(n19883), .A(n19866), .B(n19865), .ZN(
        P2_U3173) );
  AOI22_X1 U22868 ( .A1(n19877), .A2(n19869), .B1(n19868), .B2(n19874), .ZN(
        n19872) );
  AOI22_X1 U22869 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19870), .ZN(n19871) );
  OAI211_X1 U22870 ( .C1(n19873), .C2(n19883), .A(n19872), .B(n19871), .ZN(
        P2_U3174) );
  AOI22_X1 U22871 ( .A1(n19877), .A2(n19876), .B1(n19875), .B2(n19874), .ZN(
        n19882) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19878), .ZN(n19881) );
  OAI211_X1 U22873 ( .C1(n19884), .C2(n19883), .A(n19882), .B(n19881), .ZN(
        P2_U3175) );
  OAI221_X1 U22874 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19825), .C1(
        P2_STATE2_REG_2__SCAN_IN), .C2(n20026), .A(n19885), .ZN(n19890) );
  OAI21_X1 U22875 ( .B1(n19887), .B2(n19886), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19889) );
  OAI211_X1 U22876 ( .C1(n19891), .C2(n19890), .A(n19889), .B(n19888), .ZN(
        P2_U3177) );
  AND2_X1 U22877 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19892), .ZN(
        P2_U3179) );
  AND2_X1 U22878 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19892), .ZN(
        P2_U3180) );
  NOR2_X1 U22879 ( .A1(n21054), .A2(n19959), .ZN(P2_U3181) );
  AND2_X1 U22880 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19892), .ZN(
        P2_U3182) );
  AND2_X1 U22881 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19892), .ZN(
        P2_U3183) );
  AND2_X1 U22882 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19892), .ZN(
        P2_U3184) );
  NOR2_X1 U22883 ( .A1(n21173), .A2(n19959), .ZN(P2_U3185) );
  AND2_X1 U22884 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19892), .ZN(
        P2_U3186) );
  AND2_X1 U22885 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19892), .ZN(
        P2_U3187) );
  AND2_X1 U22886 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19892), .ZN(
        P2_U3188) );
  AND2_X1 U22887 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19892), .ZN(
        P2_U3189) );
  AND2_X1 U22888 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19892), .ZN(
        P2_U3190) );
  AND2_X1 U22889 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19892), .ZN(
        P2_U3191) );
  AND2_X1 U22890 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19892), .ZN(
        P2_U3192) );
  AND2_X1 U22891 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19892), .ZN(
        P2_U3193) );
  AND2_X1 U22892 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19892), .ZN(
        P2_U3194) );
  AND2_X1 U22893 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19892), .ZN(
        P2_U3195) );
  AND2_X1 U22894 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19892), .ZN(
        P2_U3196) );
  AND2_X1 U22895 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19892), .ZN(
        P2_U3197) );
  AND2_X1 U22896 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19892), .ZN(
        P2_U3198) );
  AND2_X1 U22897 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19892), .ZN(
        P2_U3199) );
  AND2_X1 U22898 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19892), .ZN(
        P2_U3200) );
  AND2_X1 U22899 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19892), .ZN(P2_U3201) );
  AND2_X1 U22900 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19892), .ZN(P2_U3202) );
  AND2_X1 U22901 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19892), .ZN(P2_U3203) );
  AND2_X1 U22902 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19892), .ZN(P2_U3204) );
  AND2_X1 U22903 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19892), .ZN(P2_U3205) );
  AND2_X1 U22904 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19892), .ZN(P2_U3206) );
  AND2_X1 U22905 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19892), .ZN(P2_U3207) );
  AND2_X1 U22906 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19892), .ZN(P2_U3208) );
  INV_X1 U22907 ( .A(NA), .ZN(n20871) );
  OAI21_X1 U22908 ( .B1(n20871), .B2(n19898), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19907) );
  INV_X1 U22909 ( .A(n19907), .ZN(n19895) );
  NAND2_X1 U22910 ( .A1(n20023), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19905) );
  INV_X1 U22911 ( .A(n19905), .ZN(n19896) );
  INV_X1 U22912 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20034) );
  NOR3_X1 U22913 ( .A1(n19896), .A2(n20034), .A3(n19897), .ZN(n19894) );
  OAI211_X1 U22914 ( .C1(HOLD), .C2(n20034), .A(n20036), .B(n19902), .ZN(
        n19893) );
  OAI21_X1 U22915 ( .B1(n19895), .B2(n19894), .A(n19893), .ZN(P2_U3209) );
  NOR2_X1 U22916 ( .A1(n20027), .A2(n19896), .ZN(n19900) );
  NOR2_X1 U22917 ( .A1(HOLD), .A2(n19897), .ZN(n19906) );
  OAI211_X1 U22918 ( .C1(n19906), .C2(n19908), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19898), .ZN(n19899) );
  OAI211_X1 U22919 ( .C1(n19901), .C2(n20866), .A(n19900), .B(n19899), .ZN(
        P2_U3210) );
  OAI22_X1 U22920 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19902), .B1(NA), 
        .B2(n19905), .ZN(n19903) );
  OAI211_X1 U22921 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19903), .ZN(n19904) );
  OAI221_X1 U22922 ( .B1(n19907), .B2(n19906), .C1(n19907), .C2(n19905), .A(
        n19904), .ZN(P2_U3211) );
  NAND2_X1 U22923 ( .A1(n20039), .A2(n19908), .ZN(n19950) );
  OAI222_X1 U22924 ( .A1(n19947), .A2(n11500), .B1(n19909), .B2(n20039), .C1(
        n11471), .C2(n19948), .ZN(P2_U3212) );
  OAI222_X1 U22925 ( .A1(n19950), .A2(n11513), .B1(n19910), .B2(n20039), .C1(
        n11500), .C2(n19948), .ZN(P2_U3213) );
  OAI222_X1 U22926 ( .A1(n19950), .A2(n11650), .B1(n19911), .B2(n20039), .C1(
        n11513), .C2(n19948), .ZN(P2_U3214) );
  OAI222_X1 U22927 ( .A1(n19950), .A2(n11753), .B1(n19912), .B2(n20039), .C1(
        n11650), .C2(n19948), .ZN(P2_U3215) );
  OAI222_X1 U22928 ( .A1(n19950), .A2(n11529), .B1(n19913), .B2(n20039), .C1(
        n11753), .C2(n19948), .ZN(P2_U3216) );
  OAI222_X1 U22929 ( .A1(n19950), .A2(n11535), .B1(n19914), .B2(n20039), .C1(
        n11529), .C2(n19948), .ZN(P2_U3217) );
  OAI222_X1 U22930 ( .A1(n19947), .A2(n13838), .B1(n19915), .B2(n20039), .C1(
        n11535), .C2(n19948), .ZN(P2_U3218) );
  OAI222_X1 U22931 ( .A1(n19947), .A2(n15608), .B1(n19916), .B2(n20039), .C1(
        n13838), .C2(n19948), .ZN(P2_U3219) );
  OAI222_X1 U22932 ( .A1(n19947), .A2(n11845), .B1(n19917), .B2(n20039), .C1(
        n15608), .C2(n19948), .ZN(P2_U3220) );
  OAI222_X1 U22933 ( .A1(n19947), .A2(n11862), .B1(n19918), .B2(n20039), .C1(
        n11845), .C2(n19948), .ZN(P2_U3221) );
  OAI222_X1 U22934 ( .A1(n19947), .A2(n11883), .B1(n19919), .B2(n20039), .C1(
        n11862), .C2(n19948), .ZN(P2_U3222) );
  OAI222_X1 U22935 ( .A1(n19947), .A2(n11903), .B1(n19920), .B2(n20039), .C1(
        n11883), .C2(n19948), .ZN(P2_U3223) );
  OAI222_X1 U22936 ( .A1(n19950), .A2(n11930), .B1(n19921), .B2(n20039), .C1(
        n11903), .C2(n19948), .ZN(P2_U3224) );
  OAI222_X1 U22937 ( .A1(n19950), .A2(n11956), .B1(n19922), .B2(n20039), .C1(
        n11930), .C2(n19948), .ZN(P2_U3225) );
  OAI222_X1 U22938 ( .A1(n19950), .A2(n15769), .B1(n19923), .B2(n20039), .C1(
        n11956), .C2(n19948), .ZN(P2_U3226) );
  OAI222_X1 U22939 ( .A1(n19950), .A2(n19925), .B1(n19924), .B2(n20039), .C1(
        n15769), .C2(n19948), .ZN(P2_U3227) );
  OAI222_X1 U22940 ( .A1(n19950), .A2(n15576), .B1(n19926), .B2(n20039), .C1(
        n19925), .C2(n19948), .ZN(P2_U3228) );
  OAI222_X1 U22941 ( .A1(n19950), .A2(n19928), .B1(n19927), .B2(n20039), .C1(
        n15576), .C2(n19948), .ZN(P2_U3229) );
  OAI222_X1 U22942 ( .A1(n19947), .A2(n19930), .B1(n19929), .B2(n20039), .C1(
        n19928), .C2(n19948), .ZN(P2_U3230) );
  OAI222_X1 U22943 ( .A1(n19947), .A2(n19932), .B1(n19931), .B2(n20039), .C1(
        n19930), .C2(n19948), .ZN(P2_U3231) );
  OAI222_X1 U22944 ( .A1(n19947), .A2(n11966), .B1(n19933), .B2(n20039), .C1(
        n19932), .C2(n19948), .ZN(P2_U3232) );
  OAI222_X1 U22945 ( .A1(n19947), .A2(n19935), .B1(n19934), .B2(n20039), .C1(
        n11966), .C2(n19948), .ZN(P2_U3233) );
  OAI222_X1 U22946 ( .A1(n19947), .A2(n19937), .B1(n19936), .B2(n20039), .C1(
        n19935), .C2(n19948), .ZN(P2_U3234) );
  OAI222_X1 U22947 ( .A1(n19947), .A2(n19939), .B1(n19938), .B2(n20039), .C1(
        n19937), .C2(n19948), .ZN(P2_U3235) );
  OAI222_X1 U22948 ( .A1(n19947), .A2(n19941), .B1(n19940), .B2(n20039), .C1(
        n19939), .C2(n19948), .ZN(P2_U3236) );
  INV_X1 U22949 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19943) );
  OAI222_X1 U22950 ( .A1(n19947), .A2(n19943), .B1(n21231), .B2(n20039), .C1(
        n19941), .C2(n19948), .ZN(P2_U3237) );
  OAI222_X1 U22951 ( .A1(n19948), .A2(n19943), .B1(n19942), .B2(n20039), .C1(
        n11588), .C2(n19947), .ZN(P2_U3238) );
  OAI222_X1 U22952 ( .A1(n19947), .A2(n19945), .B1(n19944), .B2(n20039), .C1(
        n11588), .C2(n19948), .ZN(P2_U3239) );
  OAI222_X1 U22953 ( .A1(n19947), .A2(n14356), .B1(n19946), .B2(n20039), .C1(
        n19945), .C2(n19948), .ZN(P2_U3240) );
  OAI222_X1 U22954 ( .A1(n19950), .A2(n14370), .B1(n19949), .B2(n20039), .C1(
        n14356), .C2(n19948), .ZN(P2_U3241) );
  INV_X1 U22955 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U22956 ( .A1(n20039), .A2(n19952), .B1(n19951), .B2(n20036), .ZN(
        P2_U3585) );
  MUX2_X1 U22957 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20039), .Z(P2_U3586) );
  INV_X1 U22958 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U22959 ( .A1(n20039), .A2(n19954), .B1(n19953), .B2(n20036), .ZN(
        P2_U3587) );
  INV_X1 U22960 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U22961 ( .A1(n20039), .A2(n19955), .B1(n21195), .B2(n20036), .ZN(
        P2_U3588) );
  OAI21_X1 U22962 ( .B1(n19959), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19957), 
        .ZN(n19956) );
  INV_X1 U22963 ( .A(n19956), .ZN(P2_U3591) );
  OAI21_X1 U22964 ( .B1(n19959), .B2(n19958), .A(n19957), .ZN(P2_U3592) );
  INV_X1 U22965 ( .A(n19960), .ZN(n19961) );
  OAI222_X1 U22966 ( .A1(n19981), .A2(n19965), .B1(n19964), .B2(n19963), .C1(
        n19962), .C2(n19961), .ZN(n19967) );
  MUX2_X1 U22967 ( .A(n19967), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19966), .Z(P2_U3599) );
  INV_X1 U22968 ( .A(n20007), .ZN(n19997) );
  AND2_X1 U22969 ( .A1(n19971), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19991) );
  NAND2_X1 U22970 ( .A1(n19968), .A2(n19991), .ZN(n19988) );
  OR2_X1 U22971 ( .A1(n19970), .A2(n19969), .ZN(n19992) );
  AOI21_X1 U22972 ( .B1(n19990), .B2(n19971), .A(n19992), .ZN(n19982) );
  AOI21_X1 U22973 ( .B1(n19988), .B2(n19982), .A(n19972), .ZN(n19977) );
  NOR3_X1 U22974 ( .A1(n19975), .A2(n19974), .A3(n19973), .ZN(n19976) );
  AOI211_X1 U22975 ( .C1(n19978), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19977), 
        .B(n19976), .ZN(n19979) );
  AOI22_X1 U22976 ( .A1(n19997), .A2(n19980), .B1(n19979), .B2(n20007), .ZN(
        P2_U3602) );
  INV_X1 U22977 ( .A(n19981), .ZN(n19986) );
  INV_X1 U22978 ( .A(n19982), .ZN(n19985) );
  NOR2_X1 U22979 ( .A1(n19983), .A2(n19825), .ZN(n19984) );
  AOI21_X1 U22980 ( .B1(n19986), .B2(n19985), .A(n19984), .ZN(n19987) );
  AND2_X1 U22981 ( .A1(n19988), .A2(n19987), .ZN(n19989) );
  AOI22_X1 U22982 ( .A1(n19997), .A2(n16505), .B1(n19989), .B2(n20007), .ZN(
        P2_U3603) );
  MUX2_X1 U22983 ( .A(n19992), .B(n19991), .S(n19990), .Z(n19993) );
  AOI21_X1 U22984 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19994), .A(n19993), 
        .ZN(n19995) );
  AOI22_X1 U22985 ( .A1(n19997), .A2(n19996), .B1(n19995), .B2(n20007), .ZN(
        P2_U3604) );
  INV_X1 U22986 ( .A(n19998), .ZN(n20001) );
  OAI22_X1 U22987 ( .A1(n20002), .A2(n20001), .B1(n20000), .B2(n19999), .ZN(
        n20004) );
  OAI21_X1 U22988 ( .B1(n20004), .B2(n20003), .A(n20007), .ZN(n20005) );
  OAI21_X1 U22989 ( .B1(n20007), .B2(n20006), .A(n20005), .ZN(P2_U3605) );
  INV_X1 U22990 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20008) );
  AOI22_X1 U22991 ( .A1(n20039), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20008), 
        .B2(n20036), .ZN(P2_U3608) );
  AOI22_X1 U22992 ( .A1(n20012), .A2(n20011), .B1(n20010), .B2(n20009), .ZN(
        n20013) );
  NAND2_X1 U22993 ( .A1(n20014), .A2(n20013), .ZN(n20016) );
  MUX2_X1 U22994 ( .A(P2_MORE_REG_SCAN_IN), .B(n20016), .S(n20015), .Z(
        P2_U3609) );
  OAI21_X1 U22995 ( .B1(n20018), .B2(n20017), .A(n19825), .ZN(n20021) );
  INV_X1 U22996 ( .A(n20019), .ZN(n20020) );
  OAI211_X1 U22997 ( .C1(n20023), .C2(n20022), .A(n20021), .B(n20020), .ZN(
        n20035) );
  INV_X1 U22998 ( .A(n20024), .ZN(n20025) );
  AOI21_X1 U22999 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20026), .A(n20025), 
        .ZN(n20032) );
  OAI21_X1 U23000 ( .B1(n20028), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20027), 
        .ZN(n20029) );
  AND3_X1 U23001 ( .A1(n20030), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20029), 
        .ZN(n20031) );
  OAI21_X1 U23002 ( .B1(n20032), .B2(n20031), .A(n20035), .ZN(n20033) );
  OAI21_X1 U23003 ( .B1(n20035), .B2(n20034), .A(n20033), .ZN(P2_U3610) );
  INV_X1 U23004 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20037) );
  AOI22_X1 U23005 ( .A1(n20039), .A2(n20038), .B1(n20037), .B2(n20036), .ZN(
        P2_U3611) );
  AOI21_X1 U23006 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20874), .A(n20865), 
        .ZN(n20867) );
  INV_X1 U23007 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20040) );
  AOI21_X1 U23008 ( .B1(n20867), .B2(n20040), .A(n20976), .ZN(P1_U2802) );
  INV_X1 U23009 ( .A(n20041), .ZN(n20043) );
  OAI21_X1 U23010 ( .B1(n20043), .B2(n20042), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20044) );
  OAI21_X1 U23011 ( .B1(n20045), .B2(n20968), .A(n20044), .ZN(P1_U2803) );
  NOR2_X1 U23012 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20047) );
  OAI21_X1 U23013 ( .B1(n20047), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20961), .ZN(
        n20046) );
  OAI21_X1 U23014 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20961), .A(n20046), 
        .ZN(P1_U2804) );
  OAI21_X1 U23015 ( .B1(BS16), .B2(n20047), .A(n20933), .ZN(n20931) );
  OAI21_X1 U23016 ( .B1(n20933), .B2(n20965), .A(n20931), .ZN(P1_U2805) );
  OAI21_X1 U23017 ( .B1(n20050), .B2(n20049), .A(n20048), .ZN(P1_U2806) );
  NOR4_X1 U23018 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20054) );
  NOR4_X1 U23019 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20053) );
  NOR4_X1 U23020 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20052) );
  NOR4_X1 U23021 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20051) );
  NAND4_X1 U23022 ( .A1(n20054), .A2(n20053), .A3(n20052), .A4(n20051), .ZN(
        n20060) );
  NOR4_X1 U23023 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20058) );
  AOI211_X1 U23024 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_11__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20057) );
  NOR4_X1 U23025 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20056) );
  NOR4_X1 U23026 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20055) );
  NAND4_X1 U23027 ( .A1(n20058), .A2(n20057), .A3(n20056), .A4(n20055), .ZN(
        n20059) );
  NOR2_X1 U23028 ( .A1(n20060), .A2(n20059), .ZN(n20958) );
  INV_X1 U23029 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20926) );
  NOR3_X1 U23030 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20062) );
  OAI21_X1 U23031 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20062), .A(n20958), .ZN(
        n20061) );
  OAI21_X1 U23032 ( .B1(n20958), .B2(n20926), .A(n20061), .ZN(P1_U2807) );
  INV_X1 U23033 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20932) );
  AOI21_X1 U23034 ( .B1(n20954), .B2(n20932), .A(n20062), .ZN(n20063) );
  INV_X1 U23035 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20923) );
  INV_X1 U23036 ( .A(n20958), .ZN(n20960) );
  AOI22_X1 U23037 ( .A1(n20958), .A2(n20063), .B1(n20923), .B2(n20960), .ZN(
        P1_U2808) );
  OAI22_X1 U23038 ( .A1(n20100), .A2(n20065), .B1(n20144), .B2(n20064), .ZN(
        n20066) );
  AOI211_X1 U23039 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20067), .A(n20110), .B(
        n20066), .ZN(n20073) );
  AOI22_X1 U23040 ( .A1(n20142), .A2(n20089), .B1(n20136), .B2(n20068), .ZN(
        n20072) );
  INV_X1 U23041 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20886) );
  NAND3_X1 U23042 ( .A1(n20069), .A2(n20094), .A3(n20886), .ZN(n20071) );
  NAND2_X1 U23043 ( .A1(n20097), .A2(n20141), .ZN(n20070) );
  NAND4_X1 U23044 ( .A1(n20073), .A2(n20072), .A3(n20071), .A4(n20070), .ZN(
        P1_U2831) );
  NAND2_X1 U23045 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20079) );
  NOR2_X1 U23046 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20079), .ZN(n20078) );
  AOI22_X1 U23047 ( .A1(n20074), .A2(n20097), .B1(n20125), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20075) );
  OAI211_X1 U23048 ( .C1(n20100), .C2(n20076), .A(n20075), .B(n20098), .ZN(
        n20077) );
  AOI21_X1 U23049 ( .B1(n20078), .B2(n20094), .A(n20077), .ZN(n20082) );
  INV_X1 U23050 ( .A(n20079), .ZN(n20080) );
  AOI21_X1 U23051 ( .B1(n20080), .B2(n20095), .A(n20096), .ZN(n20088) );
  AOI22_X1 U23052 ( .A1(n20148), .A2(n20089), .B1(n20088), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n20081) );
  OAI211_X1 U23053 ( .C1(n20083), .C2(n20114), .A(n20082), .B(n20081), .ZN(
        P1_U2833) );
  NAND2_X1 U23054 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20094), .ZN(n20086) );
  AOI22_X1 U23055 ( .A1(n20084), .A2(n20097), .B1(n20125), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20085) );
  OAI21_X1 U23056 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20086), .A(n20085), .ZN(
        n20087) );
  AOI211_X1 U23057 ( .C1(n20126), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20110), .B(n20087), .ZN(n20092) );
  AOI22_X1 U23058 ( .A1(n20090), .A2(n20089), .B1(n20088), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n20091) );
  OAI211_X1 U23059 ( .C1(n20093), .C2(n20114), .A(n20092), .B(n20091), .ZN(
        P1_U2834) );
  INV_X1 U23060 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20880) );
  AOI22_X1 U23061 ( .A1(n20094), .A2(n20880), .B1(n20125), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20104) );
  NOR2_X1 U23062 ( .A1(n20096), .A2(n20095), .ZN(n20109) );
  AOI22_X1 U23063 ( .A1(n20097), .A2(n20151), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20109), .ZN(n20099) );
  OAI211_X1 U23064 ( .C1(n20101), .C2(n20100), .A(n20099), .B(n20098), .ZN(
        n20102) );
  AOI21_X1 U23065 ( .B1(n20117), .B2(n20154), .A(n20102), .ZN(n20103) );
  OAI211_X1 U23066 ( .C1(n20105), .C2(n20114), .A(n20104), .B(n20103), .ZN(
        P1_U2835) );
  NAND3_X1 U23067 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20106) );
  NOR3_X1 U23068 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20107), .A3(n20106), .ZN(
        n20108) );
  AOI21_X1 U23069 ( .B1(n20109), .B2(P1_REIP_REG_4__SCAN_IN), .A(n20108), .ZN(
        n20119) );
  AOI21_X1 U23070 ( .B1(n20125), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20110), .ZN(
        n20112) );
  NAND2_X1 U23071 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20111) );
  OAI211_X1 U23072 ( .C1(n20113), .C2(n20130), .A(n20112), .B(n20111), .ZN(
        n20116) );
  NOR2_X1 U23073 ( .A1(n20114), .A2(n20229), .ZN(n20115) );
  AOI211_X1 U23074 ( .C1(n20224), .C2(n20117), .A(n20116), .B(n20115), .ZN(
        n20118) );
  OAI211_X1 U23075 ( .C1(n20140), .C2(n20120), .A(n20119), .B(n20118), .ZN(
        P1_U2836) );
  AOI21_X1 U23076 ( .B1(n20123), .B2(n20122), .A(n20121), .ZN(n20124) );
  AOI21_X1 U23077 ( .B1(n20125), .B2(P1_EBX_REG_2__SCAN_IN), .A(n20124), .ZN(
        n20139) );
  NAND2_X1 U23078 ( .A1(n20126), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n20129) );
  NAND3_X1 U23079 ( .A1(n20127), .A2(n20121), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n20128) );
  OAI211_X1 U23080 ( .C1(n20684), .C2(n20130), .A(n20129), .B(n20128), .ZN(
        n20131) );
  INV_X1 U23081 ( .A(n20131), .ZN(n20132) );
  OAI21_X1 U23082 ( .B1(n20134), .B2(n20133), .A(n20132), .ZN(n20135) );
  AOI21_X1 U23083 ( .B1(n20137), .B2(n20136), .A(n20135), .ZN(n20138) );
  OAI211_X1 U23084 ( .C1(n20140), .C2(n20253), .A(n20139), .B(n20138), .ZN(
        P1_U2838) );
  AOI22_X1 U23085 ( .A1(n20142), .A2(n20153), .B1(n20152), .B2(n20141), .ZN(
        n20143) );
  OAI21_X1 U23086 ( .B1(n20157), .B2(n20144), .A(n20143), .ZN(P1_U2863) );
  NOR2_X1 U23087 ( .A1(n20146), .A2(n20145), .ZN(n20147) );
  AOI21_X1 U23088 ( .B1(n20148), .B2(n20153), .A(n20147), .ZN(n20149) );
  OAI21_X1 U23089 ( .B1(n20157), .B2(n20150), .A(n20149), .ZN(P1_U2865) );
  AOI22_X1 U23090 ( .A1(n20154), .A2(n20153), .B1(n20152), .B2(n20151), .ZN(
        n20155) );
  OAI21_X1 U23091 ( .B1(n20157), .B2(n20156), .A(n20155), .ZN(P1_U2867) );
  AOI22_X1 U23092 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20170), .B1(n20175), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20158) );
  OAI21_X1 U23093 ( .B1(n20159), .B2(n20172), .A(n20158), .ZN(P1_U2921) );
  INV_X1 U23094 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U23095 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20160) );
  OAI21_X1 U23096 ( .B1(n20161), .B2(n20188), .A(n20160), .ZN(P1_U2922) );
  INV_X1 U23097 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20163) );
  AOI22_X1 U23098 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20162) );
  OAI21_X1 U23099 ( .B1(n20163), .B2(n20188), .A(n20162), .ZN(P1_U2923) );
  AOI22_X1 U23100 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20164) );
  OAI21_X1 U23101 ( .B1(n14080), .B2(n20188), .A(n20164), .ZN(P1_U2924) );
  AOI22_X1 U23102 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20165) );
  OAI21_X1 U23103 ( .B1(n14066), .B2(n20188), .A(n20165), .ZN(P1_U2925) );
  INV_X1 U23104 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20167) );
  AOI22_X1 U23105 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20166) );
  OAI21_X1 U23106 ( .B1(n20167), .B2(n20188), .A(n20166), .ZN(P1_U2926) );
  INV_X1 U23107 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20169) );
  AOI22_X1 U23108 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20973), .B1(n20175), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20168) );
  OAI21_X1 U23109 ( .B1(n20169), .B2(n20188), .A(n20168), .ZN(P1_U2927) );
  INV_X1 U23110 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n21275) );
  AOI22_X1 U23111 ( .A1(P1_EAX_REG_8__SCAN_IN), .A2(n20170), .B1(n20175), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n20171) );
  OAI21_X1 U23112 ( .B1(n21275), .B2(n20172), .A(n20171), .ZN(P1_U2928) );
  AOI22_X1 U23113 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20173) );
  OAI21_X1 U23114 ( .B1(n20174), .B2(n20188), .A(n20173), .ZN(P1_U2929) );
  AOI22_X1 U23115 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20176) );
  OAI21_X1 U23116 ( .B1(n10675), .B2(n20188), .A(n20176), .ZN(P1_U2930) );
  AOI22_X1 U23117 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20177) );
  OAI21_X1 U23118 ( .B1(n10657), .B2(n20188), .A(n20177), .ZN(P1_U2931) );
  INV_X1 U23119 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20179) );
  AOI22_X1 U23120 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20178) );
  OAI21_X1 U23121 ( .B1(n20179), .B2(n20188), .A(n20178), .ZN(P1_U2932) );
  AOI22_X1 U23122 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20180) );
  OAI21_X1 U23123 ( .B1(n20181), .B2(n20188), .A(n20180), .ZN(P1_U2933) );
  AOI22_X1 U23124 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20182) );
  OAI21_X1 U23125 ( .B1(n20183), .B2(n20188), .A(n20182), .ZN(P1_U2934) );
  AOI22_X1 U23126 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20184) );
  OAI21_X1 U23127 ( .B1(n20185), .B2(n20188), .A(n20184), .ZN(P1_U2935) );
  AOI22_X1 U23128 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20186), .B1(n20175), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20187) );
  OAI21_X1 U23129 ( .B1(n20189), .B2(n20188), .A(n20187), .ZN(P1_U2936) );
  AOI22_X1 U23130 ( .A1(n20192), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20195), .ZN(n20191) );
  NAND2_X1 U23131 ( .A1(n20203), .A2(n20190), .ZN(n20205) );
  NAND2_X1 U23132 ( .A1(n20191), .A2(n20205), .ZN(P1_U2945) );
  AOI22_X1 U23133 ( .A1(n20192), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20195), .ZN(n20194) );
  NAND2_X1 U23134 ( .A1(n20203), .A2(n20193), .ZN(n20209) );
  NAND2_X1 U23135 ( .A1(n20194), .A2(n20209), .ZN(P1_U2947) );
  AOI22_X1 U23136 ( .A1(n20218), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20195), .ZN(n20197) );
  NAND2_X1 U23137 ( .A1(n20203), .A2(n20196), .ZN(n20211) );
  NAND2_X1 U23138 ( .A1(n20197), .A2(n20211), .ZN(P1_U2948) );
  AOI22_X1 U23139 ( .A1(n20218), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20215), .ZN(n20199) );
  NAND2_X1 U23140 ( .A1(n20203), .A2(n20198), .ZN(n20213) );
  NAND2_X1 U23141 ( .A1(n20199), .A2(n20213), .ZN(P1_U2949) );
  AOI22_X1 U23142 ( .A1(n20218), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20215), .ZN(n20201) );
  NAND2_X1 U23143 ( .A1(n20203), .A2(n20200), .ZN(n20216) );
  NAND2_X1 U23144 ( .A1(n20201), .A2(n20216), .ZN(P1_U2950) );
  AOI22_X1 U23145 ( .A1(n20218), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20215), .ZN(n20204) );
  NAND2_X1 U23146 ( .A1(n20203), .A2(n20202), .ZN(n20219) );
  NAND2_X1 U23147 ( .A1(n20204), .A2(n20219), .ZN(P1_U2951) );
  AOI22_X1 U23148 ( .A1(n20218), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20215), .ZN(n20206) );
  NAND2_X1 U23149 ( .A1(n20206), .A2(n20205), .ZN(P1_U2960) );
  AOI22_X1 U23150 ( .A1(n20218), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20215), .ZN(n20208) );
  NAND2_X1 U23151 ( .A1(n20208), .A2(n20207), .ZN(P1_U2961) );
  AOI22_X1 U23152 ( .A1(n20218), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20215), .ZN(n20210) );
  NAND2_X1 U23153 ( .A1(n20210), .A2(n20209), .ZN(P1_U2962) );
  AOI22_X1 U23154 ( .A1(n20218), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20215), .ZN(n20212) );
  NAND2_X1 U23155 ( .A1(n20212), .A2(n20211), .ZN(P1_U2963) );
  AOI22_X1 U23156 ( .A1(n20218), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20215), .ZN(n20214) );
  NAND2_X1 U23157 ( .A1(n20214), .A2(n20213), .ZN(P1_U2964) );
  AOI22_X1 U23158 ( .A1(n20218), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20215), .ZN(n20217) );
  NAND2_X1 U23159 ( .A1(n20217), .A2(n20216), .ZN(P1_U2965) );
  AOI22_X1 U23160 ( .A1(n20218), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20215), .ZN(n20220) );
  NAND2_X1 U23161 ( .A1(n20220), .A2(n20219), .ZN(P1_U2966) );
  AOI22_X1 U23162 ( .A1(n20222), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20221), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20228) );
  INV_X1 U23163 ( .A(n20223), .ZN(n20226) );
  AOI22_X1 U23164 ( .A1(n20226), .A2(n20225), .B1(n16192), .B2(n20224), .ZN(
        n20227) );
  OAI211_X1 U23165 ( .C1(n20230), .C2(n20229), .A(n20228), .B(n20227), .ZN(
        P1_U2995) );
  INV_X1 U23166 ( .A(n20231), .ZN(n20233) );
  AOI21_X1 U23167 ( .B1(n20234), .B2(n20233), .A(n20232), .ZN(n20240) );
  INV_X1 U23168 ( .A(n20235), .ZN(n20238) );
  AOI22_X1 U23169 ( .A1(n20238), .A2(n20237), .B1(n20241), .B2(n20236), .ZN(
        n20239) );
  OAI211_X1 U23170 ( .C1(n20242), .C2(n20241), .A(n20240), .B(n20239), .ZN(
        P1_U3028) );
  NAND2_X1 U23171 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20243), .ZN(
        n20262) );
  NOR3_X1 U23172 ( .A1(n20245), .A2(n20249), .A3(n20244), .ZN(n20247) );
  AOI211_X1 U23173 ( .C1(n20249), .C2(n20248), .A(n20247), .B(n20246), .ZN(
        n20260) );
  NOR2_X1 U23174 ( .A1(n20251), .A2(n20250), .ZN(n20258) );
  OAI22_X1 U23175 ( .A1(n20254), .A2(n20253), .B1(n20121), .B2(n20252), .ZN(
        n20255) );
  AOI211_X1 U23176 ( .C1(n20258), .C2(n20257), .A(n20256), .B(n20255), .ZN(
        n20259) );
  OAI221_X1 U23177 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20262), .C1(
        n20261), .C2(n20260), .A(n20259), .ZN(P1_U3029) );
  NOR2_X1 U23178 ( .A1(n20263), .A2(n20953), .ZN(P1_U3032) );
  NAND2_X1 U23179 ( .A1(n20560), .A2(n20620), .ZN(n20450) );
  NAND2_X1 U23180 ( .A1(n20277), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20759) );
  NAND2_X1 U23181 ( .A1(n20346), .A2(n20759), .ZN(n20563) );
  OAI21_X1 U23182 ( .B1(n20374), .B2(n20851), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20266) );
  NAND2_X1 U23183 ( .A1(n20266), .A2(n20680), .ZN(n20279) );
  INV_X1 U23184 ( .A(n20684), .ZN(n20267) );
  OR2_X1 U23185 ( .A1(n20558), .A2(n20267), .ZN(n20414) );
  OR2_X1 U23186 ( .A1(n20414), .A2(n10546), .ZN(n20278) );
  INV_X1 U23187 ( .A(n20278), .ZN(n20268) );
  NAND3_X1 U23188 ( .A1(n20945), .A2(n15974), .A3(n20687), .ZN(n20354) );
  NOR2_X1 U23189 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20354), .ZN(
        n20344) );
  OAI22_X1 U23190 ( .A1(n20279), .A2(n20268), .B1(n20344), .B2(n20694), .ZN(
        n20269) );
  AOI211_X1 U23191 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20450), .A(n20563), 
        .B(n20269), .ZN(n20290) );
  INV_X1 U23192 ( .A(DATAI_24_), .ZN(n21230) );
  OAI22_X2 U23193 ( .A1(n20272), .A2(n20338), .B1(n21230), .B2(n20340), .ZN(
        n20804) );
  INV_X1 U23194 ( .A(n20804), .ZN(n20595) );
  NOR2_X2 U23195 ( .A1(n20343), .A2(n20274), .ZN(n20798) );
  INV_X1 U23196 ( .A(n20798), .ZN(n20379) );
  INV_X1 U23197 ( .A(n20344), .ZN(n20331) );
  OAI22_X1 U23198 ( .A1(n20838), .A2(n20595), .B1(n20379), .B2(n20331), .ZN(
        n20275) );
  INV_X1 U23199 ( .A(n20275), .ZN(n20283) );
  NAND2_X1 U23200 ( .A1(n20346), .A2(n20276), .ZN(n20698) );
  INV_X1 U23201 ( .A(n20698), .ZN(n20797) );
  NOR2_X1 U23202 ( .A1(n20277), .A2(n20964), .ZN(n20622) );
  INV_X1 U23203 ( .A(n20622), .ZN(n20562) );
  INV_X1 U23204 ( .A(DATAI_16_), .ZN(n20280) );
  OAI22_X1 U23205 ( .A1(n20281), .A2(n20338), .B1(n20280), .B2(n20340), .ZN(
        n20688) );
  AOI22_X1 U23206 ( .A1(n20797), .A2(n20347), .B1(n20374), .B2(n20688), .ZN(
        n20282) );
  OAI211_X1 U23207 ( .C1(n20290), .C2(n21187), .A(n20283), .B(n20282), .ZN(
        P1_U3033) );
  INV_X1 U23208 ( .A(DATAI_17_), .ZN(n20284) );
  OAI22_X1 U23209 ( .A1(n20284), .A2(n20340), .B1(n13792), .B2(n20338), .ZN(
        n20699) );
  INV_X1 U23210 ( .A(n20699), .ZN(n20813) );
  INV_X1 U23211 ( .A(DATAI_25_), .ZN(n20285) );
  OAI22_X2 U23212 ( .A1(n20286), .A2(n20338), .B1(n20285), .B2(n20340), .ZN(
        n20810) );
  INV_X1 U23213 ( .A(n20810), .ZN(n20598) );
  INV_X1 U23214 ( .A(n20809), .ZN(n20288) );
  OAI22_X1 U23215 ( .A1(n20838), .A2(n20598), .B1(n20288), .B2(n20331), .ZN(
        n20289) );
  INV_X1 U23216 ( .A(n20289), .ZN(n20293) );
  INV_X1 U23217 ( .A(n20290), .ZN(n20348) );
  NAND2_X1 U23218 ( .A1(n20346), .A2(n20291), .ZN(n20702) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20348), .B1(
        n20808), .B2(n20347), .ZN(n20292) );
  OAI211_X1 U23220 ( .C1(n20813), .C2(n20351), .A(n20293), .B(n20292), .ZN(
        P1_U3034) );
  INV_X1 U23221 ( .A(DATAI_18_), .ZN(n20295) );
  OAI22_X1 U23222 ( .A1(n20295), .A2(n20340), .B1(n20294), .B2(n20338), .ZN(
        n20703) );
  INV_X1 U23223 ( .A(n20703), .ZN(n20819) );
  INV_X1 U23224 ( .A(DATAI_26_), .ZN(n20296) );
  OAI22_X2 U23225 ( .A1(n20297), .A2(n20338), .B1(n20296), .B2(n20340), .ZN(
        n20816) );
  INV_X1 U23226 ( .A(n20816), .ZN(n20601) );
  NOR2_X2 U23227 ( .A1(n20343), .A2(n20298), .ZN(n20815) );
  INV_X1 U23228 ( .A(n20815), .ZN(n20389) );
  OAI22_X1 U23229 ( .A1(n20838), .A2(n20601), .B1(n20389), .B2(n20331), .ZN(
        n20299) );
  INV_X1 U23230 ( .A(n20299), .ZN(n20302) );
  NAND2_X1 U23231 ( .A1(n20346), .A2(n20300), .ZN(n20706) );
  INV_X1 U23232 ( .A(n20706), .ZN(n20814) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20348), .B1(
        n20814), .B2(n20347), .ZN(n20301) );
  OAI211_X1 U23234 ( .C1(n20819), .C2(n20351), .A(n20302), .B(n20301), .ZN(
        P1_U3035) );
  INV_X1 U23235 ( .A(DATAI_19_), .ZN(n20303) );
  OAI22_X1 U23236 ( .A1(n20304), .A2(n20338), .B1(n20303), .B2(n20340), .ZN(
        n20707) );
  INV_X1 U23237 ( .A(DATAI_27_), .ZN(n20305) );
  OAI22_X2 U23238 ( .A1(n20306), .A2(n20338), .B1(n20305), .B2(n20340), .ZN(
        n20822) );
  INV_X1 U23239 ( .A(n20822), .ZN(n20604) );
  NOR2_X2 U23240 ( .A1(n20343), .A2(n20307), .ZN(n20821) );
  INV_X1 U23241 ( .A(n20821), .ZN(n20393) );
  OAI22_X1 U23242 ( .A1(n20838), .A2(n20604), .B1(n20393), .B2(n20331), .ZN(
        n20308) );
  INV_X1 U23243 ( .A(n20308), .ZN(n20311) );
  NAND2_X1 U23244 ( .A1(n20346), .A2(n20309), .ZN(n20710) );
  INV_X1 U23245 ( .A(n20710), .ZN(n20820) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20348), .B1(
        n20820), .B2(n20347), .ZN(n20310) );
  OAI211_X1 U23247 ( .C1(n20825), .C2(n20351), .A(n20311), .B(n20310), .ZN(
        P1_U3036) );
  INV_X1 U23248 ( .A(DATAI_20_), .ZN(n20312) );
  OAI22_X1 U23249 ( .A1(n20312), .A2(n20340), .B1(n14594), .B2(n20338), .ZN(
        n20828) );
  INV_X1 U23250 ( .A(n20828), .ZN(n20778) );
  INV_X1 U23251 ( .A(DATAI_28_), .ZN(n20313) );
  OAI22_X2 U23252 ( .A1(n20314), .A2(n20338), .B1(n20313), .B2(n20340), .ZN(
        n20775) );
  INV_X1 U23253 ( .A(n20775), .ZN(n20831) );
  NOR2_X2 U23254 ( .A1(n20343), .A2(n10412), .ZN(n20827) );
  INV_X1 U23255 ( .A(n20827), .ZN(n20315) );
  OAI22_X1 U23256 ( .A1(n20838), .A2(n20831), .B1(n20315), .B2(n20331), .ZN(
        n20316) );
  INV_X1 U23257 ( .A(n20316), .ZN(n20319) );
  NAND2_X1 U23258 ( .A1(n20346), .A2(n20317), .ZN(n20713) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20348), .B1(
        n20826), .B2(n20347), .ZN(n20318) );
  OAI211_X1 U23260 ( .C1(n20778), .C2(n20351), .A(n20319), .B(n20318), .ZN(
        P1_U3037) );
  INV_X1 U23261 ( .A(DATAI_21_), .ZN(n20320) );
  OAI22_X1 U23262 ( .A1(n20320), .A2(n20340), .B1(n15457), .B2(n20338), .ZN(
        n20714) );
  INV_X1 U23263 ( .A(n20714), .ZN(n20839) );
  INV_X1 U23264 ( .A(DATAI_29_), .ZN(n20321) );
  OAI22_X2 U23265 ( .A1(n20322), .A2(n20338), .B1(n20321), .B2(n20340), .ZN(
        n20834) );
  NOR2_X2 U23266 ( .A1(n20343), .A2(n20323), .ZN(n20833) );
  AOI22_X1 U23267 ( .A1(n20851), .A2(n20834), .B1(n20833), .B2(n20344), .ZN(
        n20326) );
  NAND2_X1 U23268 ( .A1(n20346), .A2(n20324), .ZN(n20717) );
  INV_X1 U23269 ( .A(n20717), .ZN(n20832) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20348), .B1(
        n20832), .B2(n20347), .ZN(n20325) );
  OAI211_X1 U23271 ( .C1(n20839), .C2(n20351), .A(n20326), .B(n20325), .ZN(
        P1_U3038) );
  INV_X1 U23272 ( .A(DATAI_22_), .ZN(n20328) );
  OAI22_X1 U23273 ( .A1(n20328), .A2(n20340), .B1(n20327), .B2(n20338), .ZN(
        n20842) );
  INV_X1 U23274 ( .A(DATAI_30_), .ZN(n20329) );
  OAI22_X2 U23275 ( .A1(n20330), .A2(n20338), .B1(n20329), .B2(n20340), .ZN(
        n20781) );
  INV_X1 U23276 ( .A(n20781), .ZN(n20845) );
  NOR2_X2 U23277 ( .A1(n20343), .A2(n10446), .ZN(n20841) );
  INV_X1 U23278 ( .A(n20841), .ZN(n20401) );
  OAI22_X1 U23279 ( .A1(n20838), .A2(n20845), .B1(n20401), .B2(n20331), .ZN(
        n20332) );
  INV_X1 U23280 ( .A(n20332), .ZN(n20335) );
  NAND2_X1 U23281 ( .A1(n20346), .A2(n20333), .ZN(n20720) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20348), .B1(
        n20840), .B2(n20347), .ZN(n20334) );
  OAI211_X1 U23283 ( .C1(n20784), .C2(n20351), .A(n20335), .B(n20334), .ZN(
        P1_U3039) );
  INV_X1 U23284 ( .A(DATAI_23_), .ZN(n20337) );
  OAI22_X1 U23285 ( .A1(n20337), .A2(n20340), .B1(n20336), .B2(n20338), .ZN(
        n20850) );
  INV_X1 U23286 ( .A(n20850), .ZN(n20792) );
  INV_X1 U23287 ( .A(DATAI_31_), .ZN(n20341) );
  OAI22_X2 U23288 ( .A1(n20341), .A2(n20340), .B1(n20339), .B2(n20338), .ZN(
        n20787) );
  NOR2_X2 U23289 ( .A1(n20343), .A2(n20342), .ZN(n20849) );
  AOI22_X1 U23290 ( .A1(n20851), .A2(n20787), .B1(n20849), .B2(n20344), .ZN(
        n20350) );
  NAND2_X1 U23291 ( .A1(n20346), .A2(n20345), .ZN(n20726) );
  INV_X1 U23292 ( .A(n20726), .ZN(n20846) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20348), .B1(
        n20846), .B2(n20347), .ZN(n20349) );
  OAI211_X1 U23294 ( .C1(n20792), .C2(n20351), .A(n20350), .B(n20349), .ZN(
        P1_U3040) );
  INV_X1 U23295 ( .A(n20688), .ZN(n20807) );
  INV_X1 U23296 ( .A(n20414), .ZN(n20353) );
  INV_X1 U23297 ( .A(n20352), .ZN(n20730) );
  NOR2_X1 U23298 ( .A1(n20952), .A2(n20354), .ZN(n20372) );
  AOI21_X1 U23299 ( .B1(n20353), .B2(n20730), .A(n20372), .ZN(n20355) );
  OAI22_X1 U23300 ( .A1(n20355), .A2(n20948), .B1(n20354), .B2(n20964), .ZN(
        n20373) );
  AOI22_X1 U23301 ( .A1(n20373), .A2(n20797), .B1(n20798), .B2(n20372), .ZN(
        n20359) );
  INV_X1 U23302 ( .A(n20354), .ZN(n20357) );
  OAI21_X1 U23303 ( .B1(n20426), .B2(n20965), .A(n20355), .ZN(n20356) );
  OAI221_X1 U23304 ( .B1(n20680), .B2(n20357), .C1(n20948), .C2(n20356), .A(
        n20801), .ZN(n20375) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20804), .ZN(n20358) );
  OAI211_X1 U23306 ( .C1(n20807), .C2(n20403), .A(n20359), .B(n20358), .ZN(
        P1_U3041) );
  AOI22_X1 U23307 ( .A1(n20373), .A2(n20808), .B1(n20809), .B2(n20372), .ZN(
        n20361) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20810), .ZN(n20360) );
  OAI211_X1 U23309 ( .C1(n20813), .C2(n20403), .A(n20361), .B(n20360), .ZN(
        P1_U3042) );
  AOI22_X1 U23310 ( .A1(n20373), .A2(n20814), .B1(n20815), .B2(n20372), .ZN(
        n20363) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20816), .ZN(n20362) );
  OAI211_X1 U23312 ( .C1(n20819), .C2(n20403), .A(n20363), .B(n20362), .ZN(
        P1_U3043) );
  AOI22_X1 U23313 ( .A1(n20373), .A2(n20820), .B1(n20821), .B2(n20372), .ZN(
        n20365) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20822), .ZN(n20364) );
  OAI211_X1 U23315 ( .C1(n20825), .C2(n20403), .A(n20365), .B(n20364), .ZN(
        P1_U3044) );
  AOI22_X1 U23316 ( .A1(n20373), .A2(n20826), .B1(n20827), .B2(n20372), .ZN(
        n20367) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20775), .ZN(n20366) );
  OAI211_X1 U23318 ( .C1(n20778), .C2(n20403), .A(n20367), .B(n20366), .ZN(
        P1_U3045) );
  AOI22_X1 U23319 ( .A1(n20373), .A2(n20832), .B1(n20833), .B2(n20372), .ZN(
        n20369) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20834), .ZN(n20368) );
  OAI211_X1 U23321 ( .C1(n20839), .C2(n20403), .A(n20369), .B(n20368), .ZN(
        P1_U3046) );
  AOI22_X1 U23322 ( .A1(n20373), .A2(n20840), .B1(n20841), .B2(n20372), .ZN(
        n20371) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20781), .ZN(n20370) );
  OAI211_X1 U23324 ( .C1(n20784), .C2(n20403), .A(n20371), .B(n20370), .ZN(
        P1_U3047) );
  AOI22_X1 U23325 ( .A1(n20373), .A2(n20846), .B1(n20849), .B2(n20372), .ZN(
        n20377) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20787), .ZN(n20376) );
  OAI211_X1 U23327 ( .C1(n20792), .C2(n20403), .A(n20377), .B(n20376), .ZN(
        P1_U3048) );
  NAND2_X1 U23328 ( .A1(n20403), .A2(n20680), .ZN(n20378) );
  OAI21_X1 U23329 ( .B1(n20442), .B2(n20378), .A(n20936), .ZN(n20381) );
  NOR2_X1 U23330 ( .A1(n20414), .A2(n20559), .ZN(n20383) );
  NOR3_X1 U23331 ( .A1(n20687), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20421) );
  NAND2_X1 U23332 ( .A1(n20952), .A2(n20421), .ZN(n20402) );
  OAI22_X1 U23333 ( .A1(n20403), .A2(n20595), .B1(n20379), .B2(n20402), .ZN(
        n20380) );
  INV_X1 U23334 ( .A(n20380), .ZN(n20386) );
  INV_X1 U23335 ( .A(n20381), .ZN(n20384) );
  NOR2_X1 U23336 ( .A1(n10294), .A2(n20964), .ZN(n20503) );
  AOI211_X1 U23337 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20402), .A(n20503), 
        .B(n20563), .ZN(n20382) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20409), .B1(
        n20442), .B2(n20688), .ZN(n20385) );
  OAI211_X1 U23339 ( .C1(n20412), .C2(n20698), .A(n20386), .B(n20385), .ZN(
        P1_U3049) );
  INV_X1 U23340 ( .A(n20402), .ZN(n20407) );
  AOI22_X1 U23341 ( .A1(n20442), .A2(n20699), .B1(n20809), .B2(n20407), .ZN(
        n20388) );
  INV_X1 U23342 ( .A(n20403), .ZN(n20408) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20409), .B1(
        n20408), .B2(n20810), .ZN(n20387) );
  OAI211_X1 U23344 ( .C1(n20412), .C2(n20702), .A(n20388), .B(n20387), .ZN(
        P1_U3050) );
  OAI22_X1 U23345 ( .A1(n20403), .A2(n20601), .B1(n20402), .B2(n20389), .ZN(
        n20390) );
  INV_X1 U23346 ( .A(n20390), .ZN(n20392) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20409), .B1(
        n20442), .B2(n20703), .ZN(n20391) );
  OAI211_X1 U23348 ( .C1(n20412), .C2(n20706), .A(n20392), .B(n20391), .ZN(
        P1_U3051) );
  OAI22_X1 U23349 ( .A1(n20403), .A2(n20604), .B1(n20393), .B2(n20402), .ZN(
        n20394) );
  INV_X1 U23350 ( .A(n20394), .ZN(n20396) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20409), .B1(
        n20442), .B2(n20707), .ZN(n20395) );
  OAI211_X1 U23352 ( .C1(n20412), .C2(n20710), .A(n20396), .B(n20395), .ZN(
        P1_U3052) );
  AOI22_X1 U23353 ( .A1(n20442), .A2(n20828), .B1(n20827), .B2(n20407), .ZN(
        n20398) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20409), .B1(
        n20408), .B2(n20775), .ZN(n20397) );
  OAI211_X1 U23355 ( .C1(n20412), .C2(n20713), .A(n20398), .B(n20397), .ZN(
        P1_U3053) );
  AOI22_X1 U23356 ( .A1(n20442), .A2(n20714), .B1(n20833), .B2(n20407), .ZN(
        n20400) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20409), .B1(
        n20408), .B2(n20834), .ZN(n20399) );
  OAI211_X1 U23358 ( .C1(n20412), .C2(n20717), .A(n20400), .B(n20399), .ZN(
        P1_U3054) );
  OAI22_X1 U23359 ( .A1(n20403), .A2(n20845), .B1(n20402), .B2(n20401), .ZN(
        n20404) );
  INV_X1 U23360 ( .A(n20404), .ZN(n20406) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20409), .B1(
        n20442), .B2(n20842), .ZN(n20405) );
  OAI211_X1 U23362 ( .C1(n20412), .C2(n20720), .A(n20406), .B(n20405), .ZN(
        P1_U3055) );
  AOI22_X1 U23363 ( .A1(n20408), .A2(n20787), .B1(n20849), .B2(n20407), .ZN(
        n20411) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20409), .B1(
        n20442), .B2(n20850), .ZN(n20410) );
  OAI211_X1 U23365 ( .C1(n20412), .C2(n20726), .A(n20411), .B(n20410), .ZN(
        P1_U3056) );
  NAND2_X1 U23366 ( .A1(n10573), .A2(n20413), .ZN(n20529) );
  OR2_X1 U23367 ( .A1(n20414), .A2(n20529), .ZN(n20416) );
  NOR2_X1 U23368 ( .A1(n20651), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20441) );
  INV_X1 U23369 ( .A(n20441), .ZN(n20415) );
  AND2_X1 U23370 ( .A1(n20416), .A2(n20415), .ZN(n20423) );
  INV_X1 U23371 ( .A(n20423), .ZN(n20420) );
  INV_X1 U23372 ( .A(n20426), .ZN(n20419) );
  INV_X1 U23373 ( .A(n20417), .ZN(n20418) );
  AOI21_X1 U23374 ( .B1(n20419), .B2(n20418), .A(n20948), .ZN(n20424) );
  AOI22_X1 U23375 ( .A1(n20442), .A2(n20804), .B1(n20441), .B2(n20798), .ZN(
        n20428) );
  OAI21_X1 U23376 ( .B1(n20680), .B2(n20421), .A(n20801), .ZN(n20422) );
  AOI21_X1 U23377 ( .B1(n20424), .B2(n20423), .A(n20422), .ZN(n20425) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20443), .B1(
        n20472), .B2(n20688), .ZN(n20427) );
  OAI211_X1 U23379 ( .C1(n20446), .C2(n20698), .A(n20428), .B(n20427), .ZN(
        P1_U3057) );
  AOI22_X1 U23380 ( .A1(n20472), .A2(n20699), .B1(n20809), .B2(n20441), .ZN(
        n20430) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20810), .ZN(n20429) );
  OAI211_X1 U23382 ( .C1(n20446), .C2(n20702), .A(n20430), .B(n20429), .ZN(
        P1_U3058) );
  AOI22_X1 U23383 ( .A1(n20442), .A2(n20816), .B1(n20441), .B2(n20815), .ZN(
        n20432) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20443), .B1(
        n20472), .B2(n20703), .ZN(n20431) );
  OAI211_X1 U23385 ( .C1(n20446), .C2(n20706), .A(n20432), .B(n20431), .ZN(
        P1_U3059) );
  AOI22_X1 U23386 ( .A1(n20472), .A2(n20707), .B1(n20441), .B2(n20821), .ZN(
        n20434) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20822), .ZN(n20433) );
  OAI211_X1 U23388 ( .C1(n20446), .C2(n20710), .A(n20434), .B(n20433), .ZN(
        P1_U3060) );
  AOI22_X1 U23389 ( .A1(n20472), .A2(n20828), .B1(n20441), .B2(n20827), .ZN(
        n20436) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20775), .ZN(n20435) );
  OAI211_X1 U23391 ( .C1(n20446), .C2(n20713), .A(n20436), .B(n20435), .ZN(
        P1_U3061) );
  AOI22_X1 U23392 ( .A1(n20472), .A2(n20714), .B1(n20441), .B2(n20833), .ZN(
        n20438) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20834), .ZN(n20437) );
  OAI211_X1 U23394 ( .C1(n20446), .C2(n20717), .A(n20438), .B(n20437), .ZN(
        P1_U3062) );
  AOI22_X1 U23395 ( .A1(n20442), .A2(n20781), .B1(n20441), .B2(n20841), .ZN(
        n20440) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20443), .B1(
        n20472), .B2(n20842), .ZN(n20439) );
  OAI211_X1 U23397 ( .C1(n20446), .C2(n20720), .A(n20440), .B(n20439), .ZN(
        P1_U3063) );
  AOI22_X1 U23398 ( .A1(n20472), .A2(n20850), .B1(n20441), .B2(n20849), .ZN(
        n20445) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20787), .ZN(n20444) );
  OAI211_X1 U23400 ( .C1(n20446), .C2(n20726), .A(n20445), .B(n20444), .ZN(
        P1_U3064) );
  NAND3_X1 U23401 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20945), .A3(
        n20687), .ZN(n20476) );
  NOR2_X1 U23402 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20476), .ZN(
        n20471) );
  NOR2_X1 U23403 ( .A1(n20684), .A2(n20448), .ZN(n20530) );
  NAND3_X1 U23404 ( .A1(n20530), .A2(n20680), .A3(n20559), .ZN(n20449) );
  OAI21_X1 U23405 ( .B1(n20759), .B2(n20450), .A(n20449), .ZN(n20470) );
  AOI22_X1 U23406 ( .A1(n20798), .A2(n20471), .B1(n20797), .B2(n20470), .ZN(
        n20457) );
  INV_X1 U23407 ( .A(n20472), .ZN(n20451) );
  AOI21_X1 U23408 ( .B1(n20451), .B2(n20499), .A(n20965), .ZN(n20452) );
  AOI21_X1 U23409 ( .B1(n20530), .B2(n20559), .A(n20452), .ZN(n20453) );
  NOR2_X1 U23410 ( .A1(n20453), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20455) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20804), .ZN(n20456) );
  OAI211_X1 U23412 ( .C1(n20807), .C2(n20499), .A(n20457), .B(n20456), .ZN(
        P1_U3065) );
  AOI22_X1 U23413 ( .A1(n20809), .A2(n20471), .B1(n20808), .B2(n20470), .ZN(
        n20459) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20810), .ZN(n20458) );
  OAI211_X1 U23415 ( .C1(n20813), .C2(n20499), .A(n20459), .B(n20458), .ZN(
        P1_U3066) );
  AOI22_X1 U23416 ( .A1(n20815), .A2(n20471), .B1(n20814), .B2(n20470), .ZN(
        n20461) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20816), .ZN(n20460) );
  OAI211_X1 U23418 ( .C1(n20819), .C2(n20499), .A(n20461), .B(n20460), .ZN(
        P1_U3067) );
  AOI22_X1 U23419 ( .A1(n20821), .A2(n20471), .B1(n20820), .B2(n20470), .ZN(
        n20463) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20822), .ZN(n20462) );
  OAI211_X1 U23421 ( .C1(n20825), .C2(n20499), .A(n20463), .B(n20462), .ZN(
        P1_U3068) );
  AOI22_X1 U23422 ( .A1(n20827), .A2(n20471), .B1(n20826), .B2(n20470), .ZN(
        n20465) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20775), .ZN(n20464) );
  OAI211_X1 U23424 ( .C1(n20778), .C2(n20499), .A(n20465), .B(n20464), .ZN(
        P1_U3069) );
  AOI22_X1 U23425 ( .A1(n20833), .A2(n20471), .B1(n20832), .B2(n20470), .ZN(
        n20467) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20834), .ZN(n20466) );
  OAI211_X1 U23427 ( .C1(n20839), .C2(n20499), .A(n20467), .B(n20466), .ZN(
        P1_U3070) );
  AOI22_X1 U23428 ( .A1(n20841), .A2(n20471), .B1(n20840), .B2(n20470), .ZN(
        n20469) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20781), .ZN(n20468) );
  OAI211_X1 U23430 ( .C1(n20784), .C2(n20499), .A(n20469), .B(n20468), .ZN(
        P1_U3071) );
  AOI22_X1 U23431 ( .A1(n20849), .A2(n20471), .B1(n20846), .B2(n20470), .ZN(
        n20475) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20787), .ZN(n20474) );
  OAI211_X1 U23433 ( .C1(n20792), .C2(n20499), .A(n20475), .B(n20474), .ZN(
        P1_U3072) );
  NOR2_X1 U23434 ( .A1(n20952), .A2(n20476), .ZN(n20494) );
  AOI21_X1 U23435 ( .B1(n20530), .B2(n20730), .A(n20494), .ZN(n20477) );
  OAI22_X1 U23436 ( .A1(n20477), .A2(n20948), .B1(n20476), .B2(n20964), .ZN(
        n20495) );
  AOI22_X1 U23437 ( .A1(n20495), .A2(n20797), .B1(n20798), .B2(n20494), .ZN(
        n20481) );
  INV_X1 U23438 ( .A(n20476), .ZN(n20479) );
  OAI21_X1 U23439 ( .B1(n20534), .B2(n20965), .A(n20477), .ZN(n20478) );
  OAI221_X1 U23440 ( .B1(n20680), .B2(n20479), .C1(n20948), .C2(n20478), .A(
        n20801), .ZN(n20496) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20688), .ZN(n20480) );
  OAI211_X1 U23442 ( .C1(n20595), .C2(n20499), .A(n20481), .B(n20480), .ZN(
        P1_U3073) );
  AOI22_X1 U23443 ( .A1(n20495), .A2(n20808), .B1(n20809), .B2(n20494), .ZN(
        n20483) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20699), .ZN(n20482) );
  OAI211_X1 U23445 ( .C1(n20598), .C2(n20499), .A(n20483), .B(n20482), .ZN(
        P1_U3074) );
  AOI22_X1 U23446 ( .A1(n20495), .A2(n20814), .B1(n20815), .B2(n20494), .ZN(
        n20485) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20703), .ZN(n20484) );
  OAI211_X1 U23448 ( .C1(n20601), .C2(n20499), .A(n20485), .B(n20484), .ZN(
        P1_U3075) );
  AOI22_X1 U23449 ( .A1(n20495), .A2(n20820), .B1(n20821), .B2(n20494), .ZN(
        n20487) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20707), .ZN(n20486) );
  OAI211_X1 U23451 ( .C1(n20604), .C2(n20499), .A(n20487), .B(n20486), .ZN(
        P1_U3076) );
  AOI22_X1 U23452 ( .A1(n20495), .A2(n20826), .B1(n20827), .B2(n20494), .ZN(
        n20489) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20828), .ZN(n20488) );
  OAI211_X1 U23454 ( .C1(n20831), .C2(n20499), .A(n20489), .B(n20488), .ZN(
        P1_U3077) );
  INV_X1 U23455 ( .A(n20834), .ZN(n20609) );
  AOI22_X1 U23456 ( .A1(n20495), .A2(n20832), .B1(n20833), .B2(n20494), .ZN(
        n20491) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20714), .ZN(n20490) );
  OAI211_X1 U23458 ( .C1(n20609), .C2(n20499), .A(n20491), .B(n20490), .ZN(
        P1_U3078) );
  AOI22_X1 U23459 ( .A1(n20495), .A2(n20840), .B1(n20841), .B2(n20494), .ZN(
        n20493) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20842), .ZN(n20492) );
  OAI211_X1 U23461 ( .C1(n20845), .C2(n20499), .A(n20493), .B(n20492), .ZN(
        P1_U3079) );
  INV_X1 U23462 ( .A(n20787), .ZN(n20856) );
  AOI22_X1 U23463 ( .A1(n20495), .A2(n20846), .B1(n20849), .B2(n20494), .ZN(
        n20498) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20496), .B1(
        n20522), .B2(n20850), .ZN(n20497) );
  OAI211_X1 U23465 ( .C1(n20856), .C2(n20499), .A(n20498), .B(n20497), .ZN(
        P1_U3080) );
  INV_X1 U23466 ( .A(n20522), .ZN(n20500) );
  NAND2_X1 U23467 ( .A1(n20500), .A2(n20680), .ZN(n20501) );
  OAI21_X1 U23468 ( .B1(n20501), .B2(n20552), .A(n20936), .ZN(n20505) );
  AND2_X1 U23469 ( .A1(n20530), .A2(n10546), .ZN(n20502) );
  INV_X1 U23470 ( .A(n20759), .ZN(n20686) );
  INV_X1 U23471 ( .A(n20535), .ZN(n20531) );
  NOR2_X1 U23472 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20531), .ZN(
        n20521) );
  AOI22_X1 U23473 ( .A1(n20552), .A2(n20688), .B1(n20798), .B2(n20521), .ZN(
        n20508) );
  INV_X1 U23474 ( .A(n20502), .ZN(n20504) );
  AOI21_X1 U23475 ( .B1(n20505), .B2(n20504), .A(n20503), .ZN(n20506) );
  OAI211_X1 U23476 ( .C1(n20521), .C2(n20694), .A(n20765), .B(n20506), .ZN(
        n20523) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(n20804), .ZN(n20507) );
  OAI211_X1 U23478 ( .C1(n20526), .C2(n20698), .A(n20508), .B(n20507), .ZN(
        P1_U3081) );
  AOI22_X1 U23479 ( .A1(n20552), .A2(n20699), .B1(n20809), .B2(n20521), .ZN(
        n20510) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(n20810), .ZN(n20509) );
  OAI211_X1 U23481 ( .C1(n20526), .C2(n20702), .A(n20510), .B(n20509), .ZN(
        P1_U3082) );
  AOI22_X1 U23482 ( .A1(n20522), .A2(n20816), .B1(n20815), .B2(n20521), .ZN(
        n20512) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20523), .B1(
        n20552), .B2(n20703), .ZN(n20511) );
  OAI211_X1 U23484 ( .C1(n20526), .C2(n20706), .A(n20512), .B(n20511), .ZN(
        P1_U3083) );
  AOI22_X1 U23485 ( .A1(n20522), .A2(n20822), .B1(n20821), .B2(n20521), .ZN(
        n20514) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20523), .B1(
        n20552), .B2(n20707), .ZN(n20513) );
  OAI211_X1 U23487 ( .C1(n20526), .C2(n20710), .A(n20514), .B(n20513), .ZN(
        P1_U3084) );
  AOI22_X1 U23488 ( .A1(n20522), .A2(n20775), .B1(n20827), .B2(n20521), .ZN(
        n20516) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20523), .B1(
        n20552), .B2(n20828), .ZN(n20515) );
  OAI211_X1 U23490 ( .C1(n20526), .C2(n20713), .A(n20516), .B(n20515), .ZN(
        P1_U3085) );
  AOI22_X1 U23491 ( .A1(n20522), .A2(n20834), .B1(n20833), .B2(n20521), .ZN(
        n20518) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20523), .B1(
        n20552), .B2(n20714), .ZN(n20517) );
  OAI211_X1 U23493 ( .C1(n20526), .C2(n20717), .A(n20518), .B(n20517), .ZN(
        P1_U3086) );
  AOI22_X1 U23494 ( .A1(n20522), .A2(n20781), .B1(n20841), .B2(n20521), .ZN(
        n20520) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20523), .B1(
        n20552), .B2(n20842), .ZN(n20519) );
  OAI211_X1 U23496 ( .C1(n20526), .C2(n20720), .A(n20520), .B(n20519), .ZN(
        P1_U3087) );
  AOI22_X1 U23497 ( .A1(n20552), .A2(n20850), .B1(n20849), .B2(n20521), .ZN(
        n20525) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(n20787), .ZN(n20524) );
  OAI211_X1 U23499 ( .C1(n20526), .C2(n20726), .A(n20525), .B(n20524), .ZN(
        P1_U3088) );
  OR2_X1 U23500 ( .A1(n20529), .A2(n20948), .ZN(n20793) );
  INV_X1 U23501 ( .A(n20530), .ZN(n20532) );
  OAI222_X1 U23502 ( .A1(n20793), .A2(n20532), .B1(n20964), .B2(n20531), .C1(
        n20533), .C2(n20948), .ZN(n20551) );
  INV_X1 U23503 ( .A(n20533), .ZN(n20550) );
  AOI22_X1 U23504 ( .A1(n20551), .A2(n20797), .B1(n20798), .B2(n20550), .ZN(
        n20537) );
  NOR2_X1 U23505 ( .A1(n20534), .A2(n20799), .ZN(n20937) );
  OAI21_X1 U23506 ( .B1(n20535), .B2(n20937), .A(n20801), .ZN(n20553) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20804), .ZN(n20536) );
  OAI211_X1 U23508 ( .C1(n20807), .C2(n20564), .A(n20537), .B(n20536), .ZN(
        P1_U3089) );
  AOI22_X1 U23509 ( .A1(n20551), .A2(n20808), .B1(n20809), .B2(n20550), .ZN(
        n20539) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20810), .ZN(n20538) );
  OAI211_X1 U23511 ( .C1(n20813), .C2(n20564), .A(n20539), .B(n20538), .ZN(
        P1_U3090) );
  AOI22_X1 U23512 ( .A1(n20551), .A2(n20814), .B1(n20815), .B2(n20550), .ZN(
        n20541) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20816), .ZN(n20540) );
  OAI211_X1 U23514 ( .C1(n20819), .C2(n20564), .A(n20541), .B(n20540), .ZN(
        P1_U3091) );
  AOI22_X1 U23515 ( .A1(n20551), .A2(n20820), .B1(n20821), .B2(n20550), .ZN(
        n20543) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20822), .ZN(n20542) );
  OAI211_X1 U23517 ( .C1(n20825), .C2(n20564), .A(n20543), .B(n20542), .ZN(
        P1_U3092) );
  AOI22_X1 U23518 ( .A1(n20551), .A2(n20826), .B1(n20827), .B2(n20550), .ZN(
        n20545) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20775), .ZN(n20544) );
  OAI211_X1 U23520 ( .C1(n20778), .C2(n20564), .A(n20545), .B(n20544), .ZN(
        P1_U3093) );
  AOI22_X1 U23521 ( .A1(n20551), .A2(n20832), .B1(n20833), .B2(n20550), .ZN(
        n20547) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20834), .ZN(n20546) );
  OAI211_X1 U23523 ( .C1(n20839), .C2(n20564), .A(n20547), .B(n20546), .ZN(
        P1_U3094) );
  AOI22_X1 U23524 ( .A1(n20551), .A2(n20840), .B1(n20841), .B2(n20550), .ZN(
        n20549) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20781), .ZN(n20548) );
  OAI211_X1 U23526 ( .C1(n20784), .C2(n20564), .A(n20549), .B(n20548), .ZN(
        P1_U3095) );
  AOI22_X1 U23527 ( .A1(n20551), .A2(n20846), .B1(n20849), .B2(n20550), .ZN(
        n20555) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20787), .ZN(n20554) );
  OAI211_X1 U23529 ( .C1(n20792), .C2(n20564), .A(n20555), .B(n20554), .ZN(
        P1_U3096) );
  INV_X1 U23530 ( .A(n11190), .ZN(n20556) );
  INV_X1 U23531 ( .A(n20655), .ZN(n20939) );
  AND2_X1 U23532 ( .A1(n20558), .A2(n20684), .ZN(n20650) );
  NAND3_X1 U23533 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15974), .A3(
        n20687), .ZN(n20589) );
  NOR2_X1 U23534 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20589), .ZN(
        n20583) );
  AOI21_X1 U23535 ( .B1(n20650), .B2(n20559), .A(n20583), .ZN(n20566) );
  INV_X1 U23536 ( .A(n20560), .ZN(n20561) );
  AND2_X1 U23537 ( .A1(n20561), .A2(n20620), .ZN(n20685) );
  INV_X1 U23538 ( .A(n20685), .ZN(n20690) );
  OAI22_X1 U23539 ( .A1(n20566), .A2(n20948), .B1(n20562), .B2(n20690), .ZN(
        n20584) );
  AOI22_X1 U23540 ( .A1(n20584), .A2(n20797), .B1(n20798), .B2(n20583), .ZN(
        n20570) );
  INV_X1 U23541 ( .A(n20563), .ZN(n20624) );
  INV_X1 U23542 ( .A(n20617), .ZN(n20565) );
  OAI21_X1 U23543 ( .B1(n20565), .B2(n20585), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20567) );
  NAND2_X1 U23544 ( .A1(n20567), .A2(n20566), .ZN(n20568) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20804), .ZN(n20569) );
  OAI211_X1 U23546 ( .C1(n20807), .C2(n20617), .A(n20570), .B(n20569), .ZN(
        P1_U3097) );
  AOI22_X1 U23547 ( .A1(n20584), .A2(n20808), .B1(n20809), .B2(n20583), .ZN(
        n20572) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20810), .ZN(n20571) );
  OAI211_X1 U23549 ( .C1(n20813), .C2(n20617), .A(n20572), .B(n20571), .ZN(
        P1_U3098) );
  AOI22_X1 U23550 ( .A1(n20584), .A2(n20814), .B1(n20815), .B2(n20583), .ZN(
        n20574) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20816), .ZN(n20573) );
  OAI211_X1 U23552 ( .C1(n20819), .C2(n20617), .A(n20574), .B(n20573), .ZN(
        P1_U3099) );
  AOI22_X1 U23553 ( .A1(n20584), .A2(n20820), .B1(n20821), .B2(n20583), .ZN(
        n20576) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20822), .ZN(n20575) );
  OAI211_X1 U23555 ( .C1(n20825), .C2(n20617), .A(n20576), .B(n20575), .ZN(
        P1_U3100) );
  AOI22_X1 U23556 ( .A1(n20584), .A2(n20826), .B1(n20827), .B2(n20583), .ZN(
        n20578) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20775), .ZN(n20577) );
  OAI211_X1 U23558 ( .C1(n20778), .C2(n20617), .A(n20578), .B(n20577), .ZN(
        P1_U3101) );
  AOI22_X1 U23559 ( .A1(n20584), .A2(n20832), .B1(n20833), .B2(n20583), .ZN(
        n20580) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20834), .ZN(n20579) );
  OAI211_X1 U23561 ( .C1(n20839), .C2(n20617), .A(n20580), .B(n20579), .ZN(
        P1_U3102) );
  AOI22_X1 U23562 ( .A1(n20584), .A2(n20840), .B1(n20841), .B2(n20583), .ZN(
        n20582) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20781), .ZN(n20581) );
  OAI211_X1 U23564 ( .C1(n20784), .C2(n20617), .A(n20582), .B(n20581), .ZN(
        P1_U3103) );
  AOI22_X1 U23565 ( .A1(n20584), .A2(n20846), .B1(n20849), .B2(n20583), .ZN(
        n20588) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20586), .B1(
        n20585), .B2(n20787), .ZN(n20587) );
  OAI211_X1 U23567 ( .C1(n20792), .C2(n20617), .A(n20588), .B(n20587), .ZN(
        P1_U3104) );
  NOR2_X1 U23568 ( .A1(n20952), .A2(n20589), .ZN(n20612) );
  AOI21_X1 U23569 ( .B1(n20650), .B2(n20730), .A(n20612), .ZN(n20590) );
  OAI22_X1 U23570 ( .A1(n20590), .A2(n20948), .B1(n20589), .B2(n20964), .ZN(
        n20613) );
  AOI22_X1 U23571 ( .A1(n20613), .A2(n20797), .B1(n20798), .B2(n20612), .ZN(
        n20594) );
  INV_X1 U23572 ( .A(n20589), .ZN(n20592) );
  OAI21_X1 U23573 ( .B1(n20655), .B2(n20965), .A(n20590), .ZN(n20591) );
  OAI221_X1 U23574 ( .B1(n20680), .B2(n20592), .C1(n20948), .C2(n20591), .A(
        n20801), .ZN(n20614) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20688), .ZN(n20593) );
  OAI211_X1 U23576 ( .C1(n20595), .C2(n20617), .A(n20594), .B(n20593), .ZN(
        P1_U3105) );
  AOI22_X1 U23577 ( .A1(n20613), .A2(n20808), .B1(n20809), .B2(n20612), .ZN(
        n20597) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20699), .ZN(n20596) );
  OAI211_X1 U23579 ( .C1(n20598), .C2(n20617), .A(n20597), .B(n20596), .ZN(
        P1_U3106) );
  AOI22_X1 U23580 ( .A1(n20613), .A2(n20814), .B1(n20815), .B2(n20612), .ZN(
        n20600) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20703), .ZN(n20599) );
  OAI211_X1 U23582 ( .C1(n20601), .C2(n20617), .A(n20600), .B(n20599), .ZN(
        P1_U3107) );
  AOI22_X1 U23583 ( .A1(n20613), .A2(n20820), .B1(n20821), .B2(n20612), .ZN(
        n20603) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20707), .ZN(n20602) );
  OAI211_X1 U23585 ( .C1(n20604), .C2(n20617), .A(n20603), .B(n20602), .ZN(
        P1_U3108) );
  AOI22_X1 U23586 ( .A1(n20613), .A2(n20826), .B1(n20827), .B2(n20612), .ZN(
        n20606) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20828), .ZN(n20605) );
  OAI211_X1 U23588 ( .C1(n20831), .C2(n20617), .A(n20606), .B(n20605), .ZN(
        P1_U3109) );
  AOI22_X1 U23589 ( .A1(n20613), .A2(n20832), .B1(n20833), .B2(n20612), .ZN(
        n20608) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20714), .ZN(n20607) );
  OAI211_X1 U23591 ( .C1(n20609), .C2(n20617), .A(n20608), .B(n20607), .ZN(
        P1_U3110) );
  AOI22_X1 U23592 ( .A1(n20613), .A2(n20840), .B1(n20841), .B2(n20612), .ZN(
        n20611) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20842), .ZN(n20610) );
  OAI211_X1 U23594 ( .C1(n20845), .C2(n20617), .A(n20611), .B(n20610), .ZN(
        P1_U3111) );
  AOI22_X1 U23595 ( .A1(n20613), .A2(n20846), .B1(n20849), .B2(n20612), .ZN(
        n20616) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20614), .B1(
        n20644), .B2(n20850), .ZN(n20615) );
  OAI211_X1 U23597 ( .C1(n20856), .C2(n20617), .A(n20616), .B(n20615), .ZN(
        P1_U3112) );
  INV_X1 U23598 ( .A(n20644), .ZN(n20618) );
  NAND2_X1 U23599 ( .A1(n20618), .A2(n20680), .ZN(n20619) );
  OAI21_X1 U23600 ( .B1(n20619), .B2(n20675), .A(n20936), .ZN(n20627) );
  AND2_X1 U23601 ( .A1(n20650), .A2(n10546), .ZN(n20623) );
  OR2_X1 U23602 ( .A1(n20620), .A2(n20945), .ZN(n20760) );
  INV_X1 U23603 ( .A(n20760), .ZN(n20621) );
  NAND3_X1 U23604 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n15974), .ZN(n20656) );
  NOR2_X1 U23605 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20656), .ZN(
        n20643) );
  AOI22_X1 U23606 ( .A1(n20644), .A2(n20804), .B1(n20798), .B2(n20643), .ZN(
        n20630) );
  INV_X1 U23607 ( .A(n20623), .ZN(n20626) );
  NAND2_X1 U23608 ( .A1(n20760), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20764) );
  OAI211_X1 U23609 ( .C1(n20694), .C2(n20643), .A(n20764), .B(n20624), .ZN(
        n20625) );
  AOI21_X1 U23610 ( .B1(n20627), .B2(n20626), .A(n20625), .ZN(n20628) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20645), .B1(
        n20675), .B2(n20688), .ZN(n20629) );
  OAI211_X1 U23612 ( .C1(n20648), .C2(n20698), .A(n20630), .B(n20629), .ZN(
        P1_U3113) );
  AOI22_X1 U23613 ( .A1(n20675), .A2(n20699), .B1(n20809), .B2(n20643), .ZN(
        n20632) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20810), .ZN(n20631) );
  OAI211_X1 U23615 ( .C1(n20648), .C2(n20702), .A(n20632), .B(n20631), .ZN(
        P1_U3114) );
  AOI22_X1 U23616 ( .A1(n20644), .A2(n20816), .B1(n20815), .B2(n20643), .ZN(
        n20634) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20645), .B1(
        n20675), .B2(n20703), .ZN(n20633) );
  OAI211_X1 U23618 ( .C1(n20648), .C2(n20706), .A(n20634), .B(n20633), .ZN(
        P1_U3115) );
  AOI22_X1 U23619 ( .A1(n20644), .A2(n20822), .B1(n20821), .B2(n20643), .ZN(
        n20636) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20645), .B1(
        n20675), .B2(n20707), .ZN(n20635) );
  OAI211_X1 U23621 ( .C1(n20648), .C2(n20710), .A(n20636), .B(n20635), .ZN(
        P1_U3116) );
  AOI22_X1 U23622 ( .A1(n20644), .A2(n20775), .B1(n20827), .B2(n20643), .ZN(
        n20638) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20645), .B1(
        n20675), .B2(n20828), .ZN(n20637) );
  OAI211_X1 U23624 ( .C1(n20648), .C2(n20713), .A(n20638), .B(n20637), .ZN(
        P1_U3117) );
  AOI22_X1 U23625 ( .A1(n20675), .A2(n20714), .B1(n20833), .B2(n20643), .ZN(
        n20640) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20834), .ZN(n20639) );
  OAI211_X1 U23627 ( .C1(n20648), .C2(n20717), .A(n20640), .B(n20639), .ZN(
        P1_U3118) );
  AOI22_X1 U23628 ( .A1(n20644), .A2(n20781), .B1(n20841), .B2(n20643), .ZN(
        n20642) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20645), .B1(
        n20675), .B2(n20842), .ZN(n20641) );
  OAI211_X1 U23630 ( .C1(n20648), .C2(n20720), .A(n20642), .B(n20641), .ZN(
        P1_U3119) );
  AOI22_X1 U23631 ( .A1(n20675), .A2(n20850), .B1(n20849), .B2(n20643), .ZN(
        n20647) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20787), .ZN(n20646) );
  OAI211_X1 U23633 ( .C1(n20648), .C2(n20726), .A(n20647), .B(n20646), .ZN(
        P1_U3120) );
  INV_X1 U23634 ( .A(n20650), .ZN(n20653) );
  INV_X1 U23635 ( .A(n20651), .ZN(n20652) );
  NAND2_X1 U23636 ( .A1(n20652), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20654) );
  OAI222_X1 U23637 ( .A1(n20793), .A2(n20653), .B1(n20964), .B2(n20656), .C1(
        n20948), .C2(n20654), .ZN(n20674) );
  INV_X1 U23638 ( .A(n20654), .ZN(n20673) );
  AOI22_X1 U23639 ( .A1(n20674), .A2(n20797), .B1(n20798), .B2(n20673), .ZN(
        n20660) );
  NOR2_X1 U23640 ( .A1(n20655), .A2(n20799), .ZN(n20658) );
  INV_X1 U23641 ( .A(n20656), .ZN(n20657) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20804), .ZN(n20659) );
  OAI211_X1 U23643 ( .C1(n20807), .C2(n20695), .A(n20660), .B(n20659), .ZN(
        P1_U3121) );
  AOI22_X1 U23644 ( .A1(n20674), .A2(n20808), .B1(n20809), .B2(n20673), .ZN(
        n20662) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20810), .ZN(n20661) );
  OAI211_X1 U23646 ( .C1(n20813), .C2(n20695), .A(n20662), .B(n20661), .ZN(
        P1_U3122) );
  AOI22_X1 U23647 ( .A1(n20674), .A2(n20814), .B1(n20815), .B2(n20673), .ZN(
        n20664) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20816), .ZN(n20663) );
  OAI211_X1 U23649 ( .C1(n20819), .C2(n20695), .A(n20664), .B(n20663), .ZN(
        P1_U3123) );
  AOI22_X1 U23650 ( .A1(n20674), .A2(n20820), .B1(n20821), .B2(n20673), .ZN(
        n20666) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20822), .ZN(n20665) );
  OAI211_X1 U23652 ( .C1(n20825), .C2(n20695), .A(n20666), .B(n20665), .ZN(
        P1_U3124) );
  AOI22_X1 U23653 ( .A1(n20674), .A2(n20826), .B1(n20827), .B2(n20673), .ZN(
        n20668) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20775), .ZN(n20667) );
  OAI211_X1 U23655 ( .C1(n20778), .C2(n20695), .A(n20668), .B(n20667), .ZN(
        P1_U3125) );
  AOI22_X1 U23656 ( .A1(n20674), .A2(n20832), .B1(n20833), .B2(n20673), .ZN(
        n20670) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20834), .ZN(n20669) );
  OAI211_X1 U23658 ( .C1(n20839), .C2(n20695), .A(n20670), .B(n20669), .ZN(
        P1_U3126) );
  AOI22_X1 U23659 ( .A1(n20674), .A2(n20840), .B1(n20841), .B2(n20673), .ZN(
        n20672) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20781), .ZN(n20671) );
  OAI211_X1 U23661 ( .C1(n20784), .C2(n20695), .A(n20672), .B(n20671), .ZN(
        P1_U3127) );
  AOI22_X1 U23662 ( .A1(n20674), .A2(n20846), .B1(n20849), .B2(n20673), .ZN(
        n20678) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20676), .B1(
        n20675), .B2(n20787), .ZN(n20677) );
  OAI211_X1 U23664 ( .C1(n20792), .C2(n20695), .A(n20678), .B(n20677), .ZN(
        P1_U3128) );
  INV_X1 U23665 ( .A(n20751), .ZN(n20681) );
  NAND3_X1 U23666 ( .A1(n20681), .A2(n20680), .A3(n20695), .ZN(n20682) );
  NAND2_X1 U23667 ( .A1(n20682), .A2(n20936), .ZN(n20692) );
  OR2_X1 U23668 ( .A1(n20684), .A2(n20683), .ZN(n20794) );
  NOR2_X1 U23669 ( .A1(n20794), .A2(n10546), .ZN(n20689) );
  NAND3_X1 U23670 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20687), .ZN(n20732) );
  NOR2_X1 U23671 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20732), .ZN(
        n20721) );
  AOI22_X1 U23672 ( .A1(n20751), .A2(n20688), .B1(n20798), .B2(n20721), .ZN(
        n20697) );
  INV_X1 U23673 ( .A(n20689), .ZN(n20691) );
  AOI22_X1 U23674 ( .A1(n20692), .A2(n20691), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20690), .ZN(n20693) );
  OAI211_X1 U23675 ( .C1(n20721), .C2(n20694), .A(n20765), .B(n20693), .ZN(
        n20723) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20804), .ZN(n20696) );
  OAI211_X1 U23677 ( .C1(n20727), .C2(n20698), .A(n20697), .B(n20696), .ZN(
        P1_U3129) );
  AOI22_X1 U23678 ( .A1(n20751), .A2(n20699), .B1(n20809), .B2(n20721), .ZN(
        n20701) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20810), .ZN(n20700) );
  OAI211_X1 U23680 ( .C1(n20727), .C2(n20702), .A(n20701), .B(n20700), .ZN(
        P1_U3130) );
  AOI22_X1 U23681 ( .A1(n20751), .A2(n20703), .B1(n20815), .B2(n20721), .ZN(
        n20705) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20816), .ZN(n20704) );
  OAI211_X1 U23683 ( .C1(n20727), .C2(n20706), .A(n20705), .B(n20704), .ZN(
        P1_U3131) );
  AOI22_X1 U23684 ( .A1(n20751), .A2(n20707), .B1(n20821), .B2(n20721), .ZN(
        n20709) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20822), .ZN(n20708) );
  OAI211_X1 U23686 ( .C1(n20727), .C2(n20710), .A(n20709), .B(n20708), .ZN(
        P1_U3132) );
  AOI22_X1 U23687 ( .A1(n20751), .A2(n20828), .B1(n20827), .B2(n20721), .ZN(
        n20712) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20775), .ZN(n20711) );
  OAI211_X1 U23689 ( .C1(n20727), .C2(n20713), .A(n20712), .B(n20711), .ZN(
        P1_U3133) );
  AOI22_X1 U23690 ( .A1(n20751), .A2(n20714), .B1(n20833), .B2(n20721), .ZN(
        n20716) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20834), .ZN(n20715) );
  OAI211_X1 U23692 ( .C1(n20727), .C2(n20717), .A(n20716), .B(n20715), .ZN(
        P1_U3134) );
  AOI22_X1 U23693 ( .A1(n20751), .A2(n20842), .B1(n20841), .B2(n20721), .ZN(
        n20719) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20781), .ZN(n20718) );
  OAI211_X1 U23695 ( .C1(n20727), .C2(n20720), .A(n20719), .B(n20718), .ZN(
        P1_U3135) );
  AOI22_X1 U23696 ( .A1(n20751), .A2(n20850), .B1(n20849), .B2(n20721), .ZN(
        n20725) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20723), .B1(
        n20722), .B2(n20787), .ZN(n20724) );
  OAI211_X1 U23698 ( .C1(n20727), .C2(n20726), .A(n20725), .B(n20724), .ZN(
        P1_U3136) );
  INV_X1 U23699 ( .A(n20728), .ZN(n20729) );
  INV_X1 U23700 ( .A(n20794), .ZN(n20758) );
  NOR2_X1 U23701 ( .A1(n20952), .A2(n20732), .ZN(n20749) );
  AOI21_X1 U23702 ( .B1(n20758), .B2(n20730), .A(n20749), .ZN(n20731) );
  OAI22_X1 U23703 ( .A1(n20731), .A2(n20948), .B1(n20732), .B2(n20964), .ZN(
        n20750) );
  AOI22_X1 U23704 ( .A1(n20750), .A2(n20797), .B1(n20798), .B2(n20749), .ZN(
        n20736) );
  INV_X1 U23705 ( .A(n20732), .ZN(n20734) );
  AND2_X1 U23706 ( .A1(n20757), .A2(n20733), .ZN(n20941) );
  OAI21_X1 U23707 ( .B1(n20734), .B2(n20941), .A(n20801), .ZN(n20752) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20804), .ZN(n20735) );
  OAI211_X1 U23709 ( .C1(n20807), .C2(n20761), .A(n20736), .B(n20735), .ZN(
        P1_U3137) );
  AOI22_X1 U23710 ( .A1(n20750), .A2(n20808), .B1(n20809), .B2(n20749), .ZN(
        n20738) );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20810), .ZN(n20737) );
  OAI211_X1 U23712 ( .C1(n20813), .C2(n20761), .A(n20738), .B(n20737), .ZN(
        P1_U3138) );
  AOI22_X1 U23713 ( .A1(n20750), .A2(n20814), .B1(n20815), .B2(n20749), .ZN(
        n20740) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20816), .ZN(n20739) );
  OAI211_X1 U23715 ( .C1(n20819), .C2(n20761), .A(n20740), .B(n20739), .ZN(
        P1_U3139) );
  AOI22_X1 U23716 ( .A1(n20750), .A2(n20820), .B1(n20821), .B2(n20749), .ZN(
        n20742) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20822), .ZN(n20741) );
  OAI211_X1 U23718 ( .C1(n20825), .C2(n20761), .A(n20742), .B(n20741), .ZN(
        P1_U3140) );
  AOI22_X1 U23719 ( .A1(n20750), .A2(n20826), .B1(n20827), .B2(n20749), .ZN(
        n20744) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20775), .ZN(n20743) );
  OAI211_X1 U23721 ( .C1(n20778), .C2(n20761), .A(n20744), .B(n20743), .ZN(
        P1_U3141) );
  AOI22_X1 U23722 ( .A1(n20750), .A2(n20832), .B1(n20833), .B2(n20749), .ZN(
        n20746) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20834), .ZN(n20745) );
  OAI211_X1 U23724 ( .C1(n20839), .C2(n20761), .A(n20746), .B(n20745), .ZN(
        P1_U3142) );
  AOI22_X1 U23725 ( .A1(n20750), .A2(n20840), .B1(n20841), .B2(n20749), .ZN(
        n20748) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20781), .ZN(n20747) );
  OAI211_X1 U23727 ( .C1(n20784), .C2(n20761), .A(n20748), .B(n20747), .ZN(
        P1_U3143) );
  AOI22_X1 U23728 ( .A1(n20750), .A2(n20846), .B1(n20849), .B2(n20749), .ZN(
        n20754) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20787), .ZN(n20753) );
  OAI211_X1 U23730 ( .C1(n20792), .C2(n20761), .A(n20754), .B(n20753), .ZN(
        P1_U3144) );
  INV_X1 U23731 ( .A(n20755), .ZN(n20756) );
  NAND2_X1 U23732 ( .A1(n20758), .A2(n10546), .ZN(n20762) );
  OAI22_X1 U23733 ( .A1(n20762), .A2(n20948), .B1(n20760), .B2(n20759), .ZN(
        n20786) );
  NOR2_X1 U23734 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20795), .ZN(
        n20785) );
  AOI22_X1 U23735 ( .A1(n20797), .A2(n20786), .B1(n20798), .B2(n20785), .ZN(
        n20768) );
  OAI21_X1 U23736 ( .B1(n20835), .B2(n20788), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20763) );
  AOI21_X1 U23737 ( .B1(n20763), .B2(n20762), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20766) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20804), .ZN(n20767) );
  OAI211_X1 U23739 ( .C1(n20807), .C2(n20855), .A(n20768), .B(n20767), .ZN(
        P1_U3145) );
  AOI22_X1 U23740 ( .A1(n20808), .A2(n20786), .B1(n20809), .B2(n20785), .ZN(
        n20770) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20810), .ZN(n20769) );
  OAI211_X1 U23742 ( .C1(n20813), .C2(n20855), .A(n20770), .B(n20769), .ZN(
        P1_U3146) );
  AOI22_X1 U23743 ( .A1(n20814), .A2(n20786), .B1(n20815), .B2(n20785), .ZN(
        n20772) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20816), .ZN(n20771) );
  OAI211_X1 U23745 ( .C1(n20819), .C2(n20855), .A(n20772), .B(n20771), .ZN(
        P1_U3147) );
  AOI22_X1 U23746 ( .A1(n20820), .A2(n20786), .B1(n20821), .B2(n20785), .ZN(
        n20774) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20822), .ZN(n20773) );
  OAI211_X1 U23748 ( .C1(n20825), .C2(n20855), .A(n20774), .B(n20773), .ZN(
        P1_U3148) );
  AOI22_X1 U23749 ( .A1(n20826), .A2(n20786), .B1(n20827), .B2(n20785), .ZN(
        n20777) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20775), .ZN(n20776) );
  OAI211_X1 U23751 ( .C1(n20778), .C2(n20855), .A(n20777), .B(n20776), .ZN(
        P1_U3149) );
  AOI22_X1 U23752 ( .A1(n20832), .A2(n20786), .B1(n20833), .B2(n20785), .ZN(
        n20780) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20834), .ZN(n20779) );
  OAI211_X1 U23754 ( .C1(n20839), .C2(n20855), .A(n20780), .B(n20779), .ZN(
        P1_U3150) );
  AOI22_X1 U23755 ( .A1(n20840), .A2(n20786), .B1(n20841), .B2(n20785), .ZN(
        n20783) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20781), .ZN(n20782) );
  OAI211_X1 U23757 ( .C1(n20784), .C2(n20855), .A(n20783), .B(n20782), .ZN(
        P1_U3151) );
  AOI22_X1 U23758 ( .A1(n20846), .A2(n20786), .B1(n20849), .B2(n20785), .ZN(
        n20791) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20789), .B1(
        n20788), .B2(n20787), .ZN(n20790) );
  OAI211_X1 U23760 ( .C1(n20792), .C2(n20855), .A(n20791), .B(n20790), .ZN(
        P1_U3152) );
  INV_X1 U23761 ( .A(n20796), .ZN(n20848) );
  OAI222_X1 U23762 ( .A1(n20948), .A2(n20796), .B1(n20964), .B2(n20795), .C1(
        n20794), .C2(n20793), .ZN(n20847) );
  AOI22_X1 U23763 ( .A1(n20798), .A2(n20848), .B1(n20847), .B2(n20797), .ZN(
        n20806) );
  NOR2_X1 U23764 ( .A1(n20800), .A2(n20799), .ZN(n20803) );
  OAI21_X1 U23765 ( .B1(n20803), .B2(n20802), .A(n20801), .ZN(n20852) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20852), .B1(
        n20835), .B2(n20804), .ZN(n20805) );
  OAI211_X1 U23767 ( .C1(n20807), .C2(n20838), .A(n20806), .B(n20805), .ZN(
        P1_U3153) );
  AOI22_X1 U23768 ( .A1(n20809), .A2(n20848), .B1(n20847), .B2(n20808), .ZN(
        n20812) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20852), .B1(
        n20835), .B2(n20810), .ZN(n20811) );
  OAI211_X1 U23770 ( .C1(n20813), .C2(n20838), .A(n20812), .B(n20811), .ZN(
        P1_U3154) );
  AOI22_X1 U23771 ( .A1(n20815), .A2(n20848), .B1(n20847), .B2(n20814), .ZN(
        n20818) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20852), .B1(
        n20835), .B2(n20816), .ZN(n20817) );
  OAI211_X1 U23773 ( .C1(n20819), .C2(n20838), .A(n20818), .B(n20817), .ZN(
        P1_U3155) );
  AOI22_X1 U23774 ( .A1(n20821), .A2(n20848), .B1(n20847), .B2(n20820), .ZN(
        n20824) );
  AOI22_X1 U23775 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20852), .B1(
        n20835), .B2(n20822), .ZN(n20823) );
  OAI211_X1 U23776 ( .C1(n20825), .C2(n20838), .A(n20824), .B(n20823), .ZN(
        P1_U3156) );
  AOI22_X1 U23777 ( .A1(n20827), .A2(n20848), .B1(n20847), .B2(n20826), .ZN(
        n20830) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20852), .B1(
        n20851), .B2(n20828), .ZN(n20829) );
  OAI211_X1 U23779 ( .C1(n20831), .C2(n20855), .A(n20830), .B(n20829), .ZN(
        P1_U3157) );
  AOI22_X1 U23780 ( .A1(n20833), .A2(n20848), .B1(n20847), .B2(n20832), .ZN(
        n20837) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20852), .B1(
        n20835), .B2(n20834), .ZN(n20836) );
  OAI211_X1 U23782 ( .C1(n20839), .C2(n20838), .A(n20837), .B(n20836), .ZN(
        P1_U3158) );
  AOI22_X1 U23783 ( .A1(n20841), .A2(n20848), .B1(n20847), .B2(n20840), .ZN(
        n20844) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20852), .B1(
        n20851), .B2(n20842), .ZN(n20843) );
  OAI211_X1 U23785 ( .C1(n20845), .C2(n20855), .A(n20844), .B(n20843), .ZN(
        P1_U3159) );
  AOI22_X1 U23786 ( .A1(n20849), .A2(n20848), .B1(n20847), .B2(n20846), .ZN(
        n20854) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20852), .B1(
        n20851), .B2(n20850), .ZN(n20853) );
  OAI211_X1 U23788 ( .C1(n20856), .C2(n20855), .A(n20854), .B(n20853), .ZN(
        P1_U3160) );
  NOR2_X1 U23789 ( .A1(n20968), .A2(n20857), .ZN(n20859) );
  OAI21_X1 U23790 ( .B1(n20859), .B2(n20964), .A(n20858), .ZN(P1_U3163) );
  INV_X1 U23791 ( .A(n20933), .ZN(n20929) );
  AND2_X1 U23792 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20929), .ZN(
        P1_U3164) );
  AND2_X1 U23793 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20929), .ZN(
        P1_U3165) );
  AND2_X1 U23794 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20929), .ZN(
        P1_U3166) );
  AND2_X1 U23795 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20929), .ZN(
        P1_U3167) );
  AND2_X1 U23796 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20929), .ZN(
        P1_U3168) );
  AND2_X1 U23797 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20929), .ZN(
        P1_U3169) );
  AND2_X1 U23798 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20929), .ZN(
        P1_U3170) );
  AND2_X1 U23799 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20929), .ZN(
        P1_U3171) );
  AND2_X1 U23800 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20929), .ZN(
        P1_U3172) );
  AND2_X1 U23801 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20929), .ZN(
        P1_U3173) );
  AND2_X1 U23802 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20929), .ZN(
        P1_U3174) );
  AND2_X1 U23803 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20929), .ZN(
        P1_U3175) );
  AND2_X1 U23804 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20929), .ZN(
        P1_U3176) );
  AND2_X1 U23805 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20929), .ZN(
        P1_U3177) );
  AND2_X1 U23806 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20929), .ZN(
        P1_U3178) );
  AND2_X1 U23807 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20929), .ZN(
        P1_U3179) );
  AND2_X1 U23808 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20929), .ZN(
        P1_U3180) );
  AND2_X1 U23809 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20929), .ZN(
        P1_U3181) );
  INV_X1 U23810 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21181) );
  NOR2_X1 U23811 ( .A1(n20933), .A2(n21181), .ZN(P1_U3182) );
  AND2_X1 U23812 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20929), .ZN(
        P1_U3183) );
  AND2_X1 U23813 ( .A1(n20929), .A2(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P1_U3184) );
  AND2_X1 U23814 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20929), .ZN(
        P1_U3185) );
  AND2_X1 U23815 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20929), .ZN(P1_U3186) );
  AND2_X1 U23816 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20929), .ZN(P1_U3187) );
  AND2_X1 U23817 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20929), .ZN(P1_U3188) );
  AND2_X1 U23818 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20929), .ZN(P1_U3189) );
  AND2_X1 U23819 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20929), .ZN(P1_U3190) );
  AND2_X1 U23820 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20929), .ZN(P1_U3191) );
  INV_X1 U23821 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21112) );
  NOR2_X1 U23822 ( .A1(n20933), .A2(n21112), .ZN(P1_U3192) );
  AND2_X1 U23823 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20929), .ZN(P1_U3193) );
  NAND2_X1 U23824 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20864), .ZN(n20870) );
  INV_X1 U23825 ( .A(n20870), .ZN(n20863) );
  OAI21_X1 U23826 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20871), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20860) );
  AOI211_X1 U23827 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20861), .B(
        n20860), .ZN(n20862) );
  OAI22_X1 U23828 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20863), .B1(n20976), 
        .B2(n20862), .ZN(P1_U3194) );
  NOR3_X1 U23829 ( .A1(NA), .A2(n20865), .A3(n20864), .ZN(n20869) );
  AOI21_X1 U23830 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20874), .A(n20866), .ZN(n20868) );
  AOI222_X1 U23831 ( .A1(n20869), .A2(n20868), .B1(n20869), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(n20868), .C2(n20867), .ZN(n20873)
         );
  OAI211_X1 U23832 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20871), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20870), .ZN(n20872) );
  NAND2_X1 U23833 ( .A1(n20873), .A2(n20872), .ZN(P1_U3196) );
  NAND2_X1 U23834 ( .A1(n20976), .A2(n20874), .ZN(n20917) );
  INV_X1 U23835 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20875) );
  NAND2_X1 U23836 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20976), .ZN(n20921) );
  OAI222_X1 U23837 ( .A1(n20917), .A2(n20121), .B1(n20875), .B2(n20976), .C1(
        n20954), .C2(n20921), .ZN(P1_U3197) );
  INV_X1 U23838 ( .A(n20921), .ZN(n20903) );
  AOI222_X1 U23839 ( .A1(n20903), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20961), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20902), .ZN(n20876) );
  INV_X1 U23840 ( .A(n20876), .ZN(P1_U3198) );
  AOI222_X1 U23841 ( .A1(n20903), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20961), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20902), .ZN(n20877) );
  INV_X1 U23842 ( .A(n20877), .ZN(P1_U3199) );
  AOI222_X1 U23843 ( .A1(n20902), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20961), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20903), .ZN(n20878) );
  INV_X1 U23844 ( .A(n20878), .ZN(P1_U3200) );
  AOI22_X1 U23845 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20902), .ZN(n20879) );
  OAI21_X1 U23846 ( .B1(n20880), .B2(n20921), .A(n20879), .ZN(P1_U3201) );
  INV_X1 U23847 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U23848 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20902), .ZN(n20881) );
  OAI21_X1 U23849 ( .B1(n20882), .B2(n20921), .A(n20881), .ZN(P1_U3202) );
  AOI22_X1 U23850 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20903), .ZN(n20883) );
  OAI21_X1 U23851 ( .B1(n21118), .B2(n20917), .A(n20883), .ZN(P1_U3203) );
  INV_X1 U23852 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20884) );
  OAI222_X1 U23853 ( .A1(n20921), .A2(n21118), .B1(n20884), .B2(n20976), .C1(
        n20886), .C2(n20917), .ZN(P1_U3204) );
  INV_X1 U23854 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20885) );
  OAI222_X1 U23855 ( .A1(n20921), .A2(n20886), .B1(n20885), .B2(n20976), .C1(
        n20887), .C2(n20917), .ZN(P1_U3205) );
  INV_X1 U23856 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20888) );
  OAI222_X1 U23857 ( .A1(n20917), .A2(n20890), .B1(n20888), .B2(n20976), .C1(
        n20887), .C2(n20921), .ZN(P1_U3206) );
  AOI22_X1 U23858 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20902), .ZN(n20889) );
  OAI21_X1 U23859 ( .B1(n20890), .B2(n20921), .A(n20889), .ZN(P1_U3207) );
  AOI22_X1 U23860 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20903), .ZN(n20891) );
  OAI21_X1 U23861 ( .B1(n20893), .B2(n20917), .A(n20891), .ZN(P1_U3208) );
  AOI22_X1 U23862 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20902), .ZN(n20892) );
  OAI21_X1 U23863 ( .B1(n20893), .B2(n20921), .A(n20892), .ZN(P1_U3209) );
  AOI22_X1 U23864 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20903), .ZN(n20894) );
  OAI21_X1 U23865 ( .B1(n20895), .B2(n20917), .A(n20894), .ZN(P1_U3210) );
  INV_X1 U23866 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21078) );
  OAI222_X1 U23867 ( .A1(n20921), .A2(n20895), .B1(n21078), .B2(n20976), .C1(
        n14708), .C2(n20917), .ZN(P1_U3211) );
  AOI22_X1 U23868 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20902), .ZN(n20896) );
  OAI21_X1 U23869 ( .B1(n14708), .B2(n20921), .A(n20896), .ZN(P1_U3212) );
  AOI22_X1 U23870 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20961), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20903), .ZN(n20897) );
  OAI21_X1 U23871 ( .B1(n20900), .B2(n20917), .A(n20897), .ZN(P1_U3213) );
  INV_X1 U23872 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20899) );
  OAI222_X1 U23873 ( .A1(n20921), .A2(n20900), .B1(n20899), .B2(n20976), .C1(
        n20898), .C2(n20917), .ZN(P1_U3214) );
  AOI222_X1 U23874 ( .A1(n20902), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20961), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20903), .ZN(n20901) );
  INV_X1 U23875 ( .A(n20901), .ZN(P1_U3215) );
  AOI222_X1 U23876 ( .A1(n20903), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20961), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20902), .ZN(n20904) );
  INV_X1 U23877 ( .A(n20904), .ZN(P1_U3216) );
  INV_X1 U23878 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20905) );
  OAI222_X1 U23879 ( .A1(n20921), .A2(n14680), .B1(n20905), .B2(n20976), .C1(
        n21166), .C2(n20917), .ZN(P1_U3217) );
  INV_X1 U23880 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20906) );
  OAI222_X1 U23881 ( .A1(n20921), .A2(n21166), .B1(n20906), .B2(n20976), .C1(
        n14664), .C2(n20917), .ZN(P1_U3218) );
  INV_X1 U23882 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20907) );
  OAI222_X1 U23883 ( .A1(n20921), .A2(n14664), .B1(n20907), .B2(n20976), .C1(
        n21260), .C2(n20917), .ZN(P1_U3219) );
  INV_X1 U23884 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20908) );
  OAI222_X1 U23885 ( .A1(n20921), .A2(n21260), .B1(n20908), .B2(n20976), .C1(
        n20909), .C2(n20917), .ZN(P1_U3220) );
  INV_X1 U23886 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21157) );
  OAI222_X1 U23887 ( .A1(n20921), .A2(n20909), .B1(n21157), .B2(n20976), .C1(
        n20911), .C2(n20917), .ZN(P1_U3221) );
  INV_X1 U23888 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20910) );
  OAI222_X1 U23889 ( .A1(n20921), .A2(n20911), .B1(n20910), .B2(n20976), .C1(
        n21202), .C2(n20917), .ZN(P1_U3222) );
  INV_X1 U23890 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20912) );
  OAI222_X1 U23891 ( .A1(n20921), .A2(n21202), .B1(n20912), .B2(n20976), .C1(
        n20914), .C2(n20917), .ZN(P1_U3223) );
  INV_X1 U23892 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20913) );
  OAI222_X1 U23893 ( .A1(n20921), .A2(n20914), .B1(n20913), .B2(n20919), .C1(
        n20916), .C2(n20917), .ZN(P1_U3224) );
  INV_X1 U23894 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20915) );
  OAI222_X1 U23895 ( .A1(n20921), .A2(n20916), .B1(n20915), .B2(n20919), .C1(
        n12147), .C2(n20917), .ZN(P1_U3225) );
  INV_X1 U23896 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20920) );
  OAI222_X1 U23897 ( .A1(n20921), .A2(n12147), .B1(n20920), .B2(n20919), .C1(
        n20918), .C2(n20917), .ZN(P1_U3226) );
  INV_X1 U23898 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20922) );
  AOI22_X1 U23899 ( .A1(n20976), .A2(n20923), .B1(n20922), .B2(n20961), .ZN(
        P1_U3458) );
  INV_X1 U23900 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20956) );
  INV_X1 U23901 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U23902 ( .A1(n20976), .A2(n20956), .B1(n20924), .B2(n20961), .ZN(
        P1_U3459) );
  INV_X1 U23903 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20925) );
  AOI22_X1 U23904 ( .A1(n20976), .A2(n20926), .B1(n20925), .B2(n20961), .ZN(
        P1_U3460) );
  INV_X1 U23905 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21165) );
  INV_X1 U23906 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U23907 ( .A1(n20976), .A2(n21165), .B1(n20927), .B2(n20961), .ZN(
        P1_U3461) );
  INV_X1 U23908 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20930) );
  INV_X1 U23909 ( .A(n20931), .ZN(n20928) );
  AOI21_X1 U23910 ( .B1(n20930), .B2(n20929), .A(n20928), .ZN(P1_U3464) );
  OAI21_X1 U23911 ( .B1(n20933), .B2(n20932), .A(n20931), .ZN(P1_U3465) );
  INV_X1 U23912 ( .A(n20953), .ZN(n20944) );
  INV_X1 U23913 ( .A(n20934), .ZN(n20940) );
  OAI22_X1 U23914 ( .A1(n11190), .A2(n20936), .B1(n20935), .B2(n20947), .ZN(
        n20938) );
  AOI211_X1 U23915 ( .C1(n20940), .C2(n20939), .A(n20938), .B(n20937), .ZN(
        n20943) );
  NOR2_X1 U23916 ( .A1(n20944), .A2(n20941), .ZN(n20942) );
  AOI22_X1 U23917 ( .A1(n20945), .A2(n20944), .B1(n20943), .B2(n20942), .ZN(
        P1_U3475) );
  OAI22_X1 U23918 ( .A1(n11174), .A2(n20948), .B1(n20947), .B2(n20946), .ZN(
        n20949) );
  OAI21_X1 U23919 ( .B1(n20950), .B2(n20949), .A(n20953), .ZN(n20951) );
  OAI21_X1 U23920 ( .B1(n20953), .B2(n20952), .A(n20951), .ZN(P1_U3478) );
  AOI21_X1 U23921 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20955) );
  AOI22_X1 U23922 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20955), .B2(n20954), .ZN(n20957) );
  AOI22_X1 U23923 ( .A1(n20958), .A2(n20957), .B1(n20956), .B2(n20960), .ZN(
        P1_U3481) );
  NOR2_X1 U23924 ( .A1(n20960), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20959) );
  AOI22_X1 U23925 ( .A1(n21165), .A2(n20960), .B1(n13336), .B2(n20959), .ZN(
        P1_U3482) );
  AOI22_X1 U23926 ( .A1(n20976), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20962), 
        .B2(n20961), .ZN(P1_U3483) );
  AOI211_X1 U23927 ( .C1(n20966), .C2(n20965), .A(n20964), .B(n20963), .ZN(
        n20969) );
  OAI21_X1 U23928 ( .B1(n20969), .B2(n20968), .A(n20967), .ZN(n20975) );
  AOI211_X1 U23929 ( .C1(n20973), .C2(n20972), .A(n20971), .B(n20970), .ZN(
        n20974) );
  MUX2_X1 U23930 ( .A(n20975), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20974), 
        .Z(P1_U3485) );
  MUX2_X1 U23931 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20976), .Z(P1_U3486) );
  AOI222_X1 U23932 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20978), .B1(n17576), 
        .B2(P3_UWORD_REG_2__SCAN_IN), .C1(n20977), .C2(
        P3_DATAO_REG_18__SCAN_IN), .ZN(n21363) );
  AOI22_X1 U23933 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(keyinput164), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(keyinput182), .ZN(n20979) );
  OAI221_X1 U23934 ( .B1(P3_BE_N_REG_3__SCAN_IN), .B2(keyinput164), .C1(
        P2_EAX_REG_7__SCAN_IN), .C2(keyinput182), .A(n20979), .ZN(n20986) );
  AOI22_X1 U23935 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput167), .B1(
        P1_INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput152), .ZN(n20980) );
  OAI221_X1 U23936 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput167), .C1(
        P1_INSTQUEUE_REG_3__2__SCAN_IN), .C2(keyinput152), .A(n20980), .ZN(
        n20985) );
  AOI22_X1 U23937 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(keyinput186), .B1(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput184), .ZN(n20981) );
  OAI221_X1 U23938 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(keyinput186), .C1(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput184), .A(n20981), .ZN(
        n20984) );
  AOI22_X1 U23939 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput128), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(keyinput176), .ZN(n20982) );
  OAI221_X1 U23940 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput128), 
        .C1(P2_EAX_REG_4__SCAN_IN), .C2(keyinput176), .A(n20982), .ZN(n20983)
         );
  NOR4_X1 U23941 ( .A1(n20986), .A2(n20985), .A3(n20984), .A4(n20983), .ZN(
        n21014) );
  AOI22_X1 U23942 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput207), .B1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput170), .ZN(n20987) );
  OAI221_X1 U23943 ( .B1(P1_DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput207), .C1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(keyinput170), .A(n20987), .ZN(
        n20994) );
  AOI22_X1 U23944 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput229), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput135), .ZN(n20988) );
  OAI221_X1 U23945 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput229), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput135), .A(n20988), .ZN(n20993) );
  AOI22_X1 U23946 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(keyinput203), .B1(
        P3_EAX_REG_10__SCAN_IN), .B2(keyinput139), .ZN(n20989) );
  OAI221_X1 U23947 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(keyinput203), .C1(
        P3_EAX_REG_10__SCAN_IN), .C2(keyinput139), .A(n20989), .ZN(n20992) );
  AOI22_X1 U23948 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(keyinput159), 
        .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput242), .ZN(n20990) );
  OAI221_X1 U23949 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput159), 
        .C1(P1_REIP_REG_23__SCAN_IN), .C2(keyinput242), .A(n20990), .ZN(n20991) );
  NOR4_X1 U23950 ( .A1(n20994), .A2(n20993), .A3(n20992), .A4(n20991), .ZN(
        n21013) );
  AOI22_X1 U23951 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput189), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput173), .ZN(n20995) );
  OAI221_X1 U23952 ( .B1(P3_DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput189), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput173), .A(n20995), .ZN(
        n21002) );
  AOI22_X1 U23953 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(keyinput147), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput154), .ZN(n20996) );
  OAI221_X1 U23954 ( .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput147), .C1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(keyinput154), .A(n20996), 
        .ZN(n21001) );
  AOI22_X1 U23955 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(keyinput192), .B1(
        P3_FLUSH_REG_SCAN_IN), .B2(keyinput195), .ZN(n20997) );
  OAI221_X1 U23956 ( .B1(P2_D_C_N_REG_SCAN_IN), .B2(keyinput192), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(keyinput195), .A(n20997), .ZN(n21000) );
  AOI22_X1 U23957 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput185), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput171), .ZN(n20998) );
  OAI221_X1 U23958 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput185), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput171), .A(n20998), .ZN(n20999)
         );
  NOR4_X1 U23959 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21012) );
  AOI22_X1 U23960 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(keyinput198), .B1(
        BUF2_REG_5__SCAN_IN), .B2(keyinput129), .ZN(n21003) );
  OAI221_X1 U23961 ( .B1(P1_DATAO_REG_24__SCAN_IN), .B2(keyinput198), .C1(
        BUF2_REG_5__SCAN_IN), .C2(keyinput129), .A(n21003), .ZN(n21010) );
  AOI22_X1 U23962 ( .A1(DATAI_24_), .A2(keyinput161), .B1(
        P2_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput236), .ZN(n21004) );
  OAI221_X1 U23963 ( .B1(DATAI_24_), .B2(keyinput161), .C1(
        P2_INSTQUEUE_REG_9__2__SCAN_IN), .C2(keyinput236), .A(n21004), .ZN(
        n21009) );
  AOI22_X1 U23964 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(keyinput168), 
        .B1(P2_REIP_REG_5__SCAN_IN), .B2(keyinput174), .ZN(n21005) );
  OAI221_X1 U23965 ( .B1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B2(keyinput168), 
        .C1(P2_REIP_REG_5__SCAN_IN), .C2(keyinput174), .A(n21005), .ZN(n21008)
         );
  AOI22_X1 U23966 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(keyinput132), .B1(
        BUF2_REG_21__SCAN_IN), .B2(keyinput249), .ZN(n21006) );
  OAI221_X1 U23967 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(keyinput132), .C1(
        BUF2_REG_21__SCAN_IN), .C2(keyinput249), .A(n21006), .ZN(n21007) );
  NOR4_X1 U23968 ( .A1(n21010), .A2(n21009), .A3(n21008), .A4(n21007), .ZN(
        n21011) );
  NAND4_X1 U23969 ( .A1(n21014), .A2(n21013), .A3(n21012), .A4(n21011), .ZN(
        n21154) );
  AOI22_X1 U23970 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(keyinput245), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput232), .ZN(n21015) );
  OAI221_X1 U23971 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(keyinput245), .C1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput232), .A(n21015), 
        .ZN(n21022) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(keyinput241), 
        .B1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput208), .ZN(n21016) );
  OAI221_X1 U23973 ( .B1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B2(keyinput241), 
        .C1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .C2(keyinput208), .A(n21016), 
        .ZN(n21021) );
  AOI22_X1 U23974 ( .A1(P3_LWORD_REG_11__SCAN_IN), .A2(keyinput230), .B1(
        DATAI_19_), .B2(keyinput177), .ZN(n21017) );
  OAI221_X1 U23975 ( .B1(P3_LWORD_REG_11__SCAN_IN), .B2(keyinput230), .C1(
        DATAI_19_), .C2(keyinput177), .A(n21017), .ZN(n21020) );
  AOI22_X1 U23976 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput201), .B1(
        P3_DATAO_REG_18__SCAN_IN), .B2(keyinput158), .ZN(n21018) );
  OAI221_X1 U23977 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput201), .C1(
        P3_DATAO_REG_18__SCAN_IN), .C2(keyinput158), .A(n21018), .ZN(n21019)
         );
  NOR4_X1 U23978 ( .A1(n21022), .A2(n21021), .A3(n21020), .A4(n21019), .ZN(
        n21050) );
  AOI22_X1 U23979 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(keyinput193), 
        .B1(P2_EAX_REG_2__SCAN_IN), .B2(keyinput227), .ZN(n21023) );
  OAI221_X1 U23980 ( .B1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput193), 
        .C1(P2_EAX_REG_2__SCAN_IN), .C2(keyinput227), .A(n21023), .ZN(n21030)
         );
  AOI22_X1 U23981 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(keyinput224), .B1(
        P3_EAX_REG_28__SCAN_IN), .B2(keyinput228), .ZN(n21024) );
  OAI221_X1 U23982 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(keyinput224), .C1(
        P3_EAX_REG_28__SCAN_IN), .C2(keyinput228), .A(n21024), .ZN(n21029) );
  AOI22_X1 U23983 ( .A1(BUF2_REG_28__SCAN_IN), .A2(keyinput191), .B1(
        BUF2_REG_29__SCAN_IN), .B2(keyinput155), .ZN(n21025) );
  OAI221_X1 U23984 ( .B1(BUF2_REG_28__SCAN_IN), .B2(keyinput191), .C1(
        BUF2_REG_29__SCAN_IN), .C2(keyinput155), .A(n21025), .ZN(n21028) );
  AOI22_X1 U23985 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(keyinput178), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(keyinput130), .ZN(n21026) );
  OAI221_X1 U23986 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(keyinput178), .C1(
        P1_ADDRESS_REG_24__SCAN_IN), .C2(keyinput130), .A(n21026), .ZN(n21027)
         );
  NOR4_X1 U23987 ( .A1(n21030), .A2(n21029), .A3(n21028), .A4(n21027), .ZN(
        n21049) );
  AOI22_X1 U23988 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(keyinput140), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(keyinput199), .ZN(n21031) );
  OAI221_X1 U23989 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(keyinput140), .C1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .C2(keyinput199), .A(n21031), .ZN(
        n21038) );
  AOI22_X1 U23990 ( .A1(BUF1_REG_10__SCAN_IN), .A2(keyinput226), .B1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput145), .ZN(n21032) );
  OAI221_X1 U23991 ( .B1(BUF1_REG_10__SCAN_IN), .B2(keyinput226), .C1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .C2(keyinput145), .A(n21032), .ZN(
        n21037) );
  AOI22_X1 U23992 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput169), .B1(
        P1_EBX_REG_23__SCAN_IN), .B2(keyinput244), .ZN(n21033) );
  OAI221_X1 U23993 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput169), .C1(
        P1_EBX_REG_23__SCAN_IN), .C2(keyinput244), .A(n21033), .ZN(n21036) );
  AOI22_X1 U23994 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(keyinput157), .B1(
        P2_ADDRESS_REG_23__SCAN_IN), .B2(keyinput211), .ZN(n21034) );
  OAI221_X1 U23995 ( .B1(P2_ADDRESS_REG_19__SCAN_IN), .B2(keyinput157), .C1(
        P2_ADDRESS_REG_23__SCAN_IN), .C2(keyinput211), .A(n21034), .ZN(n21035)
         );
  NOR4_X1 U23996 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21048) );
  AOI22_X1 U23997 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(keyinput190), .B1(
        P3_INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput213), .ZN(n21039) );
  OAI221_X1 U23998 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(keyinput190), .C1(
        P3_INSTQUEUE_REG_5__4__SCAN_IN), .C2(keyinput213), .A(n21039), .ZN(
        n21046) );
  AOI22_X1 U23999 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput150), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput134), .ZN(n21040) );
  OAI221_X1 U24000 ( .B1(P1_DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput150), .C1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput134), .A(n21040), .ZN(
        n21045) );
  AOI22_X1 U24001 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput235), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(keyinput181), .ZN(n21041) );
  OAI221_X1 U24002 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput235), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput181), .A(n21041), .ZN(n21044)
         );
  AOI22_X1 U24003 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput146), .B1(
        P1_INSTQUEUE_REG_11__7__SCAN_IN), .B2(keyinput243), .ZN(n21042) );
  OAI221_X1 U24004 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput146), .C1(
        P1_INSTQUEUE_REG_11__7__SCAN_IN), .C2(keyinput243), .A(n21042), .ZN(
        n21043) );
  NOR4_X1 U24005 ( .A1(n21046), .A2(n21045), .A3(n21044), .A4(n21043), .ZN(
        n21047) );
  NAND4_X1 U24006 ( .A1(n21050), .A2(n21049), .A3(n21048), .A4(n21047), .ZN(
        n21153) );
  AOI22_X1 U24007 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput197), .B1(
        P1_INSTQUEUE_REG_1__4__SCAN_IN), .B2(keyinput247), .ZN(n21051) );
  OAI221_X1 U24008 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput197), .C1(
        P1_INSTQUEUE_REG_1__4__SCAN_IN), .C2(keyinput247), .A(n21051), .ZN(
        n21060) );
  AOI22_X1 U24009 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput142), .B1(
        P2_UWORD_REG_5__SCAN_IN), .B2(keyinput160), .ZN(n21052) );
  OAI221_X1 U24010 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput142), .C1(
        P2_UWORD_REG_5__SCAN_IN), .C2(keyinput160), .A(n21052), .ZN(n21059) );
  AOI22_X1 U24011 ( .A1(n21254), .A2(keyinput234), .B1(keyinput196), .B2(
        n21054), .ZN(n21053) );
  OAI221_X1 U24012 ( .B1(n21254), .B2(keyinput234), .C1(n21054), .C2(
        keyinput196), .A(n21053), .ZN(n21058) );
  AOI22_X1 U24013 ( .A1(n21056), .A2(keyinput149), .B1(n21178), .B2(
        keyinput246), .ZN(n21055) );
  OAI221_X1 U24014 ( .B1(n21056), .B2(keyinput149), .C1(n21178), .C2(
        keyinput246), .A(n21055), .ZN(n21057) );
  NOR4_X1 U24015 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21098) );
  AOI22_X1 U24016 ( .A1(n13792), .A2(keyinput210), .B1(keyinput248), .B2(
        n21062), .ZN(n21061) );
  OAI221_X1 U24017 ( .B1(n13792), .B2(keyinput210), .C1(n21062), .C2(
        keyinput248), .A(n21061), .ZN(n21065) );
  XNOR2_X1 U24018 ( .A(n10315), .B(keyinput220), .ZN(n21064) );
  INV_X1 U24019 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n21160) );
  XNOR2_X1 U24020 ( .A(n21160), .B(keyinput172), .ZN(n21063) );
  OR3_X1 U24021 ( .A1(n21065), .A2(n21064), .A3(n21063), .ZN(n21071) );
  INV_X1 U24022 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21067) );
  AOI22_X1 U24023 ( .A1(n21067), .A2(keyinput252), .B1(keyinput148), .B2(
        n21162), .ZN(n21066) );
  OAI221_X1 U24024 ( .B1(n21067), .B2(keyinput252), .C1(n21162), .C2(
        keyinput148), .A(n21066), .ZN(n21070) );
  AOI22_X1 U24025 ( .A1(n21237), .A2(keyinput187), .B1(keyinput206), .B2(
        n10657), .ZN(n21068) );
  OAI221_X1 U24026 ( .B1(n21237), .B2(keyinput187), .C1(n10657), .C2(
        keyinput206), .A(n21068), .ZN(n21069) );
  NOR3_X1 U24027 ( .A1(n21071), .A2(n21070), .A3(n21069), .ZN(n21097) );
  AOI22_X1 U24028 ( .A1(n12680), .A2(keyinput254), .B1(keyinput251), .B2(
        n21212), .ZN(n21072) );
  OAI221_X1 U24029 ( .B1(n12680), .B2(keyinput254), .C1(n21212), .C2(
        keyinput251), .A(n21072), .ZN(n21075) );
  XOR2_X1 U24030 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B(keyinput231), .Z(
        n21074) );
  XNOR2_X1 U24031 ( .A(n21195), .B(keyinput250), .ZN(n21073) );
  OR3_X1 U24032 ( .A1(n21075), .A2(n21074), .A3(n21073), .ZN(n21081) );
  AOI22_X1 U24033 ( .A1(n14593), .A2(keyinput151), .B1(n14356), .B2(
        keyinput202), .ZN(n21076) );
  OAI221_X1 U24034 ( .B1(n14593), .B2(keyinput151), .C1(n14356), .C2(
        keyinput202), .A(n21076), .ZN(n21080) );
  AOI22_X1 U24035 ( .A1(n21268), .A2(keyinput163), .B1(n21078), .B2(
        keyinput239), .ZN(n21077) );
  OAI221_X1 U24036 ( .B1(n21268), .B2(keyinput163), .C1(n21078), .C2(
        keyinput239), .A(n21077), .ZN(n21079) );
  NOR3_X1 U24037 ( .A1(n21081), .A2(n21080), .A3(n21079), .ZN(n21096) );
  AOI22_X1 U24038 ( .A1(n21084), .A2(keyinput143), .B1(n21083), .B2(
        keyinput233), .ZN(n21082) );
  OAI221_X1 U24039 ( .B1(n21084), .B2(keyinput143), .C1(n21083), .C2(
        keyinput233), .A(n21082), .ZN(n21094) );
  AOI22_X1 U24040 ( .A1(n21209), .A2(keyinput183), .B1(keyinput144), .B2(
        n21086), .ZN(n21085) );
  OAI221_X1 U24041 ( .B1(n21209), .B2(keyinput183), .C1(n21086), .C2(
        keyinput144), .A(n21085), .ZN(n21093) );
  AOI22_X1 U24042 ( .A1(n21227), .A2(keyinput209), .B1(keyinput219), .B2(
        n21088), .ZN(n21087) );
  OAI221_X1 U24043 ( .B1(n21227), .B2(keyinput209), .C1(n21088), .C2(
        keyinput219), .A(n21087), .ZN(n21092) );
  INV_X1 U24044 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n21090) );
  AOI22_X1 U24045 ( .A1(n21090), .A2(keyinput165), .B1(keyinput175), .B2(
        n21193), .ZN(n21089) );
  OAI221_X1 U24046 ( .B1(n21090), .B2(keyinput165), .C1(n21193), .C2(
        keyinput175), .A(n21089), .ZN(n21091) );
  NOR4_X1 U24047 ( .A1(n21094), .A2(n21093), .A3(n21092), .A4(n21091), .ZN(
        n21095) );
  NAND4_X1 U24048 ( .A1(n21098), .A2(n21097), .A3(n21096), .A4(n21095), .ZN(
        n21152) );
  AOI22_X1 U24049 ( .A1(n21100), .A2(keyinput131), .B1(keyinput188), .B2(
        n21274), .ZN(n21099) );
  OAI221_X1 U24050 ( .B1(n21100), .B2(keyinput131), .C1(n21274), .C2(
        keyinput188), .A(n21099), .ZN(n21110) );
  INV_X1 U24051 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n21224) );
  AOI22_X1 U24052 ( .A1(n21102), .A2(keyinput212), .B1(n21224), .B2(
        keyinput153), .ZN(n21101) );
  OAI221_X1 U24053 ( .B1(n21102), .B2(keyinput212), .C1(n21224), .C2(
        keyinput153), .A(n21101), .ZN(n21109) );
  INV_X1 U24054 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21104) );
  AOI22_X1 U24055 ( .A1(n21173), .A2(keyinput222), .B1(n21104), .B2(
        keyinput162), .ZN(n21103) );
  OAI221_X1 U24056 ( .B1(n21173), .B2(keyinput222), .C1(n21104), .C2(
        keyinput162), .A(n21103), .ZN(n21108) );
  XNOR2_X1 U24057 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput221), .ZN(
        n21106) );
  XNOR2_X1 U24058 ( .A(keyinput255), .B(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n21105) );
  NAND2_X1 U24059 ( .A1(n21106), .A2(n21105), .ZN(n21107) );
  NOR4_X1 U24060 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21150) );
  AOI22_X1 U24061 ( .A1(n21196), .A2(keyinput215), .B1(n21260), .B2(
        keyinput214), .ZN(n21111) );
  OAI221_X1 U24062 ( .B1(n21196), .B2(keyinput215), .C1(n21260), .C2(
        keyinput214), .A(n21111), .ZN(n21115) );
  XNOR2_X1 U24063 ( .A(n21112), .B(keyinput179), .ZN(n21114) );
  XOR2_X1 U24064 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B(keyinput253), .Z(
        n21113) );
  OR3_X1 U24065 ( .A1(n21115), .A2(n21114), .A3(n21113), .ZN(n21122) );
  AOI22_X1 U24066 ( .A1(n21231), .A2(keyinput216), .B1(keyinput180), .B2(
        n21271), .ZN(n21116) );
  OAI221_X1 U24067 ( .B1(n21231), .B2(keyinput216), .C1(n21271), .C2(
        keyinput180), .A(n21116), .ZN(n21121) );
  AOI22_X1 U24068 ( .A1(n21119), .A2(keyinput200), .B1(n21118), .B2(
        keyinput166), .ZN(n21117) );
  OAI221_X1 U24069 ( .B1(n21119), .B2(keyinput200), .C1(n21118), .C2(
        keyinput166), .A(n21117), .ZN(n21120) );
  NOR3_X1 U24070 ( .A1(n21122), .A2(n21121), .A3(n21120), .ZN(n21149) );
  INV_X1 U24071 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21124) );
  AOI22_X1 U24072 ( .A1(n21124), .A2(keyinput137), .B1(n12754), .B2(
        keyinput136), .ZN(n21123) );
  OAI221_X1 U24073 ( .B1(n21124), .B2(keyinput137), .C1(n12754), .C2(
        keyinput136), .A(n21123), .ZN(n21133) );
  INV_X1 U24074 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21257) );
  AOI22_X1 U24075 ( .A1(n21257), .A2(keyinput133), .B1(keyinput223), .B2(
        n21222), .ZN(n21125) );
  OAI221_X1 U24076 ( .B1(n21257), .B2(keyinput133), .C1(n21222), .C2(
        keyinput223), .A(n21125), .ZN(n21132) );
  AOI22_X1 U24077 ( .A1(n21127), .A2(keyinput238), .B1(n21204), .B2(
        keyinput240), .ZN(n21126) );
  OAI221_X1 U24078 ( .B1(n21127), .B2(keyinput238), .C1(n21204), .C2(
        keyinput240), .A(n21126), .ZN(n21131) );
  AOI22_X1 U24079 ( .A1(n21129), .A2(keyinput204), .B1(n11903), .B2(
        keyinput225), .ZN(n21128) );
  OAI221_X1 U24080 ( .B1(n21129), .B2(keyinput204), .C1(n11903), .C2(
        keyinput225), .A(n21128), .ZN(n21130) );
  NOR4_X1 U24081 ( .A1(n21133), .A2(n21132), .A3(n21131), .A4(n21130), .ZN(
        n21148) );
  INV_X1 U24082 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n21135) );
  AOI22_X1 U24083 ( .A1(n21135), .A2(keyinput237), .B1(keyinput138), .B2(
        n21192), .ZN(n21134) );
  OAI221_X1 U24084 ( .B1(n21135), .B2(keyinput237), .C1(n21192), .C2(
        keyinput138), .A(n21134), .ZN(n21146) );
  AOI22_X1 U24085 ( .A1(n21138), .A2(keyinput218), .B1(keyinput194), .B2(
        n21137), .ZN(n21136) );
  OAI221_X1 U24086 ( .B1(n21138), .B2(keyinput218), .C1(n21137), .C2(
        keyinput194), .A(n21136), .ZN(n21145) );
  AOI22_X1 U24087 ( .A1(n14246), .A2(keyinput156), .B1(keyinput205), .B2(
        n21140), .ZN(n21139) );
  OAI221_X1 U24088 ( .B1(n14246), .B2(keyinput156), .C1(n21140), .C2(
        keyinput205), .A(n21139), .ZN(n21144) );
  AOI22_X1 U24089 ( .A1(n21142), .A2(keyinput141), .B1(n11500), .B2(
        keyinput217), .ZN(n21141) );
  OAI221_X1 U24090 ( .B1(n21142), .B2(keyinput141), .C1(n11500), .C2(
        keyinput217), .A(n21141), .ZN(n21143) );
  NOR4_X1 U24091 ( .A1(n21146), .A2(n21145), .A3(n21144), .A4(n21143), .ZN(
        n21147) );
  NAND4_X1 U24092 ( .A1(n21150), .A2(n21149), .A3(n21148), .A4(n21147), .ZN(
        n21151) );
  NOR4_X1 U24093 ( .A1(n21154), .A2(n21153), .A3(n21152), .A4(n21151), .ZN(
        n21361) );
  AOI22_X1 U24094 ( .A1(n21157), .A2(keyinput2), .B1(keyinput19), .B2(n21156), 
        .ZN(n21155) );
  OAI221_X1 U24095 ( .B1(n21157), .B2(keyinput2), .C1(n21156), .C2(keyinput19), 
        .A(n21155), .ZN(n21170) );
  AOI22_X1 U24096 ( .A1(n21160), .A2(keyinput44), .B1(n21159), .B2(keyinput42), 
        .ZN(n21158) );
  OAI221_X1 U24097 ( .B1(n21160), .B2(keyinput44), .C1(n21159), .C2(keyinput42), .A(n21158), .ZN(n21169) );
  AOI22_X1 U24098 ( .A1(n21163), .A2(keyinput62), .B1(n21162), .B2(keyinput20), 
        .ZN(n21161) );
  OAI221_X1 U24099 ( .B1(n21163), .B2(keyinput62), .C1(n21162), .C2(keyinput20), .A(n21161), .ZN(n21168) );
  AOI22_X1 U24100 ( .A1(n21166), .A2(keyinput69), .B1(keyinput45), .B2(n21165), 
        .ZN(n21164) );
  OAI221_X1 U24101 ( .B1(n21166), .B2(keyinput69), .C1(n21165), .C2(keyinput45), .A(n21164), .ZN(n21167) );
  NOR4_X1 U24102 ( .A1(n21170), .A2(n21169), .A3(n21168), .A4(n21167), .ZN(
        n21220) );
  INV_X1 U24103 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n21172) );
  AOI22_X1 U24104 ( .A1(n21173), .A2(keyinput94), .B1(n21172), .B2(keyinput30), 
        .ZN(n21171) );
  OAI221_X1 U24105 ( .B1(n21173), .B2(keyinput94), .C1(n21172), .C2(keyinput30), .A(n21171), .ZN(n21185) );
  AOI22_X1 U24106 ( .A1(n21176), .A2(keyinput53), .B1(n21175), .B2(keyinput113), .ZN(n21174) );
  OAI221_X1 U24107 ( .B1(n21176), .B2(keyinput53), .C1(n21175), .C2(
        keyinput113), .A(n21174), .ZN(n21184) );
  AOI22_X1 U24108 ( .A1(n14593), .A2(keyinput23), .B1(keyinput118), .B2(n21178), .ZN(n21177) );
  OAI221_X1 U24109 ( .B1(n14593), .B2(keyinput23), .C1(n21178), .C2(
        keyinput118), .A(n21177), .ZN(n21183) );
  AOI22_X1 U24110 ( .A1(n21181), .A2(keyinput22), .B1(n21180), .B2(keyinput43), 
        .ZN(n21179) );
  OAI221_X1 U24111 ( .B1(n21181), .B2(keyinput22), .C1(n21180), .C2(keyinput43), .A(n21179), .ZN(n21182) );
  NOR4_X1 U24112 ( .A1(n21185), .A2(n21184), .A3(n21183), .A4(n21182), .ZN(
        n21219) );
  AOI22_X1 U24113 ( .A1(n21187), .A2(keyinput17), .B1(keyinput82), .B2(n13792), 
        .ZN(n21186) );
  OAI221_X1 U24114 ( .B1(n21187), .B2(keyinput17), .C1(n13792), .C2(keyinput82), .A(n21186), .ZN(n21200) );
  AOI22_X1 U24115 ( .A1(n21190), .A2(keyinput85), .B1(n21189), .B2(keyinput63), 
        .ZN(n21188) );
  OAI221_X1 U24116 ( .B1(n21190), .B2(keyinput85), .C1(n21189), .C2(keyinput63), .A(n21188), .ZN(n21199) );
  AOI22_X1 U24117 ( .A1(n21193), .A2(keyinput47), .B1(keyinput10), .B2(n21192), 
        .ZN(n21191) );
  OAI221_X1 U24118 ( .B1(n21193), .B2(keyinput47), .C1(n21192), .C2(keyinput10), .A(n21191), .ZN(n21198) );
  AOI22_X1 U24119 ( .A1(n21196), .A2(keyinput87), .B1(keyinput122), .B2(n21195), .ZN(n21194) );
  OAI221_X1 U24120 ( .B1(n21196), .B2(keyinput87), .C1(n21195), .C2(
        keyinput122), .A(n21194), .ZN(n21197) );
  NOR4_X1 U24121 ( .A1(n21200), .A2(n21199), .A3(n21198), .A4(n21197), .ZN(
        n21218) );
  AOI22_X1 U24122 ( .A1(n21203), .A2(keyinput100), .B1(n21202), .B2(keyinput41), .ZN(n21201) );
  OAI221_X1 U24123 ( .B1(n21203), .B2(keyinput100), .C1(n21202), .C2(
        keyinput41), .A(n21201), .ZN(n21207) );
  XNOR2_X1 U24124 ( .A(n21204), .B(keyinput112), .ZN(n21206) );
  XOR2_X1 U24125 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput93), .Z(
        n21205) );
  OR3_X1 U24126 ( .A1(n21207), .A2(n21206), .A3(n21205), .ZN(n21216) );
  AOI22_X1 U24127 ( .A1(n21210), .A2(keyinput67), .B1(n21209), .B2(keyinput55), 
        .ZN(n21208) );
  OAI221_X1 U24128 ( .B1(n21210), .B2(keyinput67), .C1(n21209), .C2(keyinput55), .A(n21208), .ZN(n21215) );
  AOI22_X1 U24129 ( .A1(n21213), .A2(keyinput127), .B1(keyinput123), .B2(
        n21212), .ZN(n21211) );
  OAI221_X1 U24130 ( .B1(n21213), .B2(keyinput127), .C1(n21212), .C2(
        keyinput123), .A(n21211), .ZN(n21214) );
  NOR3_X1 U24131 ( .A1(n21216), .A2(n21215), .A3(n21214), .ZN(n21217) );
  NAND4_X1 U24132 ( .A1(n21220), .A2(n21219), .A3(n21218), .A4(n21217), .ZN(
        n21360) );
  AOI22_X1 U24133 ( .A1(n21222), .A2(keyinput95), .B1(n12147), .B2(keyinput7), 
        .ZN(n21221) );
  OAI221_X1 U24134 ( .B1(n21222), .B2(keyinput95), .C1(n12147), .C2(keyinput7), 
        .A(n21221), .ZN(n21235) );
  INV_X1 U24135 ( .A(P3_LWORD_REG_11__SCAN_IN), .ZN(n21225) );
  AOI22_X1 U24136 ( .A1(n21225), .A2(keyinput102), .B1(n21224), .B2(keyinput25), .ZN(n21223) );
  OAI221_X1 U24137 ( .B1(n21225), .B2(keyinput102), .C1(n21224), .C2(
        keyinput25), .A(n21223), .ZN(n21234) );
  AOI22_X1 U24138 ( .A1(n21228), .A2(keyinput31), .B1(keyinput81), .B2(n21227), 
        .ZN(n21226) );
  OAI221_X1 U24139 ( .B1(n21228), .B2(keyinput31), .C1(n21227), .C2(keyinput81), .A(n21226), .ZN(n21233) );
  AOI22_X1 U24140 ( .A1(n21231), .A2(keyinput88), .B1(keyinput33), .B2(n21230), 
        .ZN(n21229) );
  OAI221_X1 U24141 ( .B1(n21231), .B2(keyinput88), .C1(n21230), .C2(keyinput33), .A(n21229), .ZN(n21232) );
  NOR4_X1 U24142 ( .A1(n21235), .A2(n21234), .A3(n21233), .A4(n21232), .ZN(
        n21358) );
  XNOR2_X1 U24143 ( .A(n21236), .B(keyinput36), .ZN(n21241) );
  XOR2_X1 U24144 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput24), .Z(
        n21240) );
  XOR2_X1 U24145 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B(keyinput80), .Z(
        n21239) );
  XNOR2_X1 U24146 ( .A(n21237), .B(keyinput59), .ZN(n21238) );
  NOR4_X1 U24147 ( .A1(n21241), .A2(n21240), .A3(n21239), .A4(n21238), .ZN(
        n21249) );
  OAI22_X1 U24148 ( .A1(n14664), .A2(keyinput114), .B1(n21243), .B2(keyinput65), .ZN(n21242) );
  AOI221_X1 U24149 ( .B1(n14664), .B2(keyinput114), .C1(keyinput65), .C2(
        n21243), .A(n21242), .ZN(n21248) );
  INV_X1 U24150 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n21245) );
  OAI22_X1 U24151 ( .A1(n21246), .A2(keyinput1), .B1(n21245), .B2(keyinput75), 
        .ZN(n21244) );
  AOI221_X1 U24152 ( .B1(n21246), .B2(keyinput1), .C1(keyinput75), .C2(n21245), 
        .A(n21244), .ZN(n21247) );
  NAND3_X1 U24153 ( .A1(n21249), .A2(n21248), .A3(n21247), .ZN(n21282) );
  OAI22_X1 U24154 ( .A1(n21252), .A2(keyinput11), .B1(n21251), .B2(keyinput61), 
        .ZN(n21250) );
  AOI221_X1 U24155 ( .B1(n21252), .B2(keyinput11), .C1(keyinput61), .C2(n21251), .A(n21250), .ZN(n21264) );
  INV_X1 U24156 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n21255) );
  OAI22_X1 U24157 ( .A1(n21255), .A2(keyinput117), .B1(n21254), .B2(
        keyinput106), .ZN(n21253) );
  AOI221_X1 U24158 ( .B1(n21255), .B2(keyinput117), .C1(keyinput106), .C2(
        n21254), .A(n21253), .ZN(n21263) );
  OAI22_X1 U24159 ( .A1(n10657), .A2(keyinput78), .B1(n21257), .B2(keyinput5), 
        .ZN(n21256) );
  AOI221_X1 U24160 ( .B1(n10657), .B2(keyinput78), .C1(keyinput5), .C2(n21257), 
        .A(n21256), .ZN(n21262) );
  OAI22_X1 U24161 ( .A1(n21260), .A2(keyinput86), .B1(n21259), .B2(keyinput14), 
        .ZN(n21258) );
  AOI221_X1 U24162 ( .B1(n21260), .B2(keyinput86), .C1(keyinput14), .C2(n21259), .A(n21258), .ZN(n21261) );
  NAND4_X1 U24163 ( .A1(n21264), .A2(n21263), .A3(n21262), .A4(n21261), .ZN(
        n21281) );
  INV_X1 U24164 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n21266) );
  AOI22_X1 U24165 ( .A1(n21266), .A2(keyinput12), .B1(n11500), .B2(keyinput89), 
        .ZN(n21265) );
  OAI221_X1 U24166 ( .B1(n21266), .B2(keyinput12), .C1(n11500), .C2(keyinput89), .A(n21265), .ZN(n21280) );
  OAI22_X1 U24167 ( .A1(n21269), .A2(keyinput54), .B1(n21268), .B2(keyinput35), 
        .ZN(n21267) );
  AOI221_X1 U24168 ( .B1(n21269), .B2(keyinput54), .C1(keyinput35), .C2(n21268), .A(n21267), .ZN(n21278) );
  OAI22_X1 U24169 ( .A1(n21272), .A2(keyinput6), .B1(n21271), .B2(keyinput52), 
        .ZN(n21270) );
  AOI221_X1 U24170 ( .B1(n21272), .B2(keyinput6), .C1(keyinput52), .C2(n21271), 
        .A(n21270), .ZN(n21277) );
  OAI22_X1 U24171 ( .A1(n21275), .A2(keyinput50), .B1(n21274), .B2(keyinput60), 
        .ZN(n21273) );
  AOI221_X1 U24172 ( .B1(n21275), .B2(keyinput50), .C1(keyinput60), .C2(n21274), .A(n21273), .ZN(n21276) );
  NAND3_X1 U24173 ( .A1(n21278), .A2(n21277), .A3(n21276), .ZN(n21279) );
  NOR4_X1 U24174 ( .A1(n21282), .A2(n21281), .A3(n21280), .A4(n21279), .ZN(
        n21357) );
  OAI22_X1 U24175 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(keyinput48), .B1(
        keyinput18), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n21283) );
  AOI221_X1 U24176 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(keyinput48), .C1(
        P1_REIP_REG_16__SCAN_IN), .C2(keyinput18), .A(n21283), .ZN(n21290) );
  OAI22_X1 U24177 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(keyinput8), .B1(
        P3_INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput77), .ZN(n21284) );
  AOI221_X1 U24178 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(keyinput8), .C1(
        keyinput77), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(n21284), .ZN(
        n21289) );
  OAI22_X1 U24179 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(keyinput97), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(keyinput34), .ZN(n21285) );
  AOI221_X1 U24180 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(keyinput97), .C1(
        keyinput34), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21285), .ZN(n21288) );
  OAI22_X1 U24181 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(keyinput119), 
        .B1(keyinput72), .B2(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21286) );
  AOI221_X1 U24182 ( .B1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B2(keyinput119), 
        .C1(P3_DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput72), .A(n21286), .ZN(
        n21287) );
  NAND4_X1 U24183 ( .A1(n21290), .A2(n21289), .A3(n21288), .A4(n21287), .ZN(
        n21318) );
  OAI22_X1 U24184 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(keyinput83), .B1(
        keyinput15), .B2(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21291) );
  AOI221_X1 U24185 ( .B1(P2_ADDRESS_REG_23__SCAN_IN), .B2(keyinput83), .C1(
        P3_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput15), .A(n21291), .ZN(n21298) );
  OAI22_X1 U24186 ( .A1(BUF1_REG_10__SCAN_IN), .A2(keyinput98), .B1(keyinput40), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21292) );
  AOI221_X1 U24187 ( .B1(BUF1_REG_10__SCAN_IN), .B2(keyinput98), .C1(
        P3_INSTQUEUE_REG_14__2__SCAN_IN), .C2(keyinput40), .A(n21292), .ZN(
        n21297) );
  OAI22_X1 U24188 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(keyinput37), .B1(
        keyinput70), .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n21293) );
  AOI221_X1 U24189 ( .B1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput37), 
        .C1(P1_DATAO_REG_24__SCAN_IN), .C2(keyinput70), .A(n21293), .ZN(n21296) );
  OAI22_X1 U24190 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(keyinput99), .B1(
        keyinput68), .B2(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n21294) );
  AOI221_X1 U24191 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(keyinput99), .C1(
        P2_DATAWIDTH_REG_29__SCAN_IN), .C2(keyinput68), .A(n21294), .ZN(n21295) );
  NAND4_X1 U24192 ( .A1(n21298), .A2(n21297), .A3(n21296), .A4(n21295), .ZN(
        n21317) );
  OAI22_X1 U24193 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(keyinput108), 
        .B1(keyinput120), .B2(P3_LWORD_REG_15__SCAN_IN), .ZN(n21299) );
  AOI221_X1 U24194 ( .B1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput108), 
        .C1(P3_LWORD_REG_15__SCAN_IN), .C2(keyinput120), .A(n21299), .ZN(
        n21306) );
  OAI22_X1 U24195 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput38), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(keyinput105), .ZN(n21300) );
  AOI221_X1 U24196 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput38), .C1(
        keyinput105), .C2(P3_EAX_REG_20__SCAN_IN), .A(n21300), .ZN(n21305) );
  OAI22_X1 U24197 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(keyinput29), .B1(
        keyinput9), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21301) );
  AOI221_X1 U24198 ( .B1(P2_ADDRESS_REG_19__SCAN_IN), .B2(keyinput29), .C1(
        P1_INSTQUEUE_REG_14__1__SCAN_IN), .C2(keyinput9), .A(n21301), .ZN(
        n21304) );
  OAI22_X1 U24199 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(keyinput58), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput66), .ZN(n21302) );
  AOI221_X1 U24200 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(keyinput58), .C1(
        keyinput66), .C2(P2_DATAO_REG_15__SCAN_IN), .A(n21302), .ZN(n21303) );
  NAND4_X1 U24201 ( .A1(n21306), .A2(n21305), .A3(n21304), .A4(n21303), .ZN(
        n21316) );
  OAI22_X1 U24202 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput107), .B1(
        P1_DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput79), .ZN(n21307) );
  AOI221_X1 U24203 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput107), .C1(
        keyinput79), .C2(P1_DATAWIDTH_REG_11__SCAN_IN), .A(n21307), .ZN(n21314) );
  OAI22_X1 U24204 ( .A1(BUF2_REG_2__SCAN_IN), .A2(keyinput13), .B1(keyinput91), 
        .B2(P3_UWORD_REG_6__SCAN_IN), .ZN(n21308) );
  AOI221_X1 U24205 ( .B1(BUF2_REG_2__SCAN_IN), .B2(keyinput13), .C1(
        P3_UWORD_REG_6__SCAN_IN), .C2(keyinput91), .A(n21308), .ZN(n21313) );
  OAI22_X1 U24206 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(keyinput92), 
        .B1(keyinput73), .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n21309) );
  AOI221_X1 U24207 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput92), 
        .C1(P3_DATAO_REG_9__SCAN_IN), .C2(keyinput73), .A(n21309), .ZN(n21312)
         );
  OAI22_X1 U24208 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(keyinput124), 
        .B1(keyinput57), .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n21310) );
  AOI221_X1 U24209 ( .B1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput124), 
        .C1(P1_DATAO_REG_19__SCAN_IN), .C2(keyinput57), .A(n21310), .ZN(n21311) );
  NAND4_X1 U24210 ( .A1(n21314), .A2(n21313), .A3(n21312), .A4(n21311), .ZN(
        n21315) );
  NOR4_X1 U24211 ( .A1(n21318), .A2(n21317), .A3(n21316), .A4(n21315), .ZN(
        n21356) );
  OAI22_X1 U24212 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(keyinput125), 
        .B1(keyinput71), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n21319) );
  AOI221_X1 U24213 ( .B1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput125), 
        .C1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .C2(keyinput71), .A(n21319), .ZN(
        n21326) );
  OAI22_X1 U24214 ( .A1(BUF2_REG_29__SCAN_IN), .A2(keyinput27), .B1(
        keyinput101), .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n21320) );
  AOI221_X1 U24215 ( .B1(BUF2_REG_29__SCAN_IN), .B2(keyinput27), .C1(
        P1_DATAO_REG_29__SCAN_IN), .C2(keyinput101), .A(n21320), .ZN(n21325)
         );
  OAI22_X1 U24216 ( .A1(DATAI_19_), .A2(keyinput49), .B1(
        P2_UWORD_REG_5__SCAN_IN), .B2(keyinput32), .ZN(n21321) );
  AOI221_X1 U24217 ( .B1(DATAI_19_), .B2(keyinput49), .C1(keyinput32), .C2(
        P2_UWORD_REG_5__SCAN_IN), .A(n21321), .ZN(n21324) );
  OAI22_X1 U24218 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput104), 
        .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput3), .ZN(n21322) );
  AOI221_X1 U24219 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput104), 
        .C1(keyinput3), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(n21322), 
        .ZN(n21323) );
  NAND4_X1 U24220 ( .A1(n21326), .A2(n21325), .A3(n21324), .A4(n21323), .ZN(
        n21354) );
  OAI22_X1 U24221 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(keyinput26), 
        .B1(keyinput115), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n21327) );
  AOI221_X1 U24222 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput26), 
        .C1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .C2(keyinput115), .A(n21327), 
        .ZN(n21334) );
  OAI22_X1 U24223 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput116), .B1(
        keyinput39), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21328) );
  AOI221_X1 U24224 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput116), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput39), .A(n21328), .ZN(n21333) );
  OAI22_X1 U24225 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(keyinput74), .B1(
        keyinput84), .B2(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21329) );
  AOI221_X1 U24226 ( .B1(P2_REIP_REG_30__SCAN_IN), .B2(keyinput74), .C1(
        P3_DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput84), .A(n21329), .ZN(n21332)
         );
  OAI22_X1 U24227 ( .A1(BUF1_REG_4__SCAN_IN), .A2(keyinput16), .B1(keyinput0), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21330) );
  AOI221_X1 U24228 ( .B1(BUF1_REG_4__SCAN_IN), .B2(keyinput16), .C1(
        P3_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput0), .A(n21330), .ZN(n21331) );
  NAND4_X1 U24229 ( .A1(n21334), .A2(n21333), .A3(n21332), .A4(n21331), .ZN(
        n21353) );
  OAI22_X1 U24230 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput28), 
        .B1(keyinput64), .B2(P2_D_C_N_REG_SCAN_IN), .ZN(n21335) );
  AOI221_X1 U24231 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput28), 
        .C1(P2_D_C_N_REG_SCAN_IN), .C2(keyinput64), .A(n21335), .ZN(n21342) );
  OAI22_X1 U24232 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput56), .B1(
        keyinput51), .B2(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21336) );
  AOI221_X1 U24233 ( .B1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput56), 
        .C1(P1_DATAWIDTH_REG_3__SCAN_IN), .C2(keyinput51), .A(n21336), .ZN(
        n21341) );
  OAI22_X1 U24234 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput90), 
        .B1(BUF2_REG_21__SCAN_IN), .B2(keyinput121), .ZN(n21337) );
  AOI221_X1 U24235 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput90), 
        .C1(keyinput121), .C2(BUF2_REG_21__SCAN_IN), .A(n21337), .ZN(n21340)
         );
  OAI22_X1 U24236 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(keyinput103), 
        .B1(P3_EBX_REG_16__SCAN_IN), .B2(keyinput4), .ZN(n21338) );
  AOI221_X1 U24237 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(keyinput103), 
        .C1(keyinput4), .C2(P3_EBX_REG_16__SCAN_IN), .A(n21338), .ZN(n21339)
         );
  NAND4_X1 U24238 ( .A1(n21342), .A2(n21341), .A3(n21340), .A4(n21339), .ZN(
        n21352) );
  OAI22_X1 U24239 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(keyinput109), 
        .B1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput76), .ZN(n21343) );
  AOI221_X1 U24240 ( .B1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(keyinput109), 
        .C1(keyinput76), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(n21343), 
        .ZN(n21350) );
  OAI22_X1 U24241 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(keyinput126), 
        .B1(keyinput110), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n21344) );
  AOI221_X1 U24242 ( .B1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(keyinput126), 
        .C1(P3_EBX_REG_17__SCAN_IN), .C2(keyinput110), .A(n21344), .ZN(n21349)
         );
  OAI22_X1 U24243 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(keyinput46), .B1(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput21), .ZN(n21345) );
  AOI221_X1 U24244 ( .B1(P2_REIP_REG_5__SCAN_IN), .B2(keyinput46), .C1(
        keyinput21), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n21345), .ZN(
        n21348) );
  OAI22_X1 U24245 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(keyinput111), .B1(
        keyinput96), .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n21346) );
  AOI221_X1 U24246 ( .B1(P1_ADDRESS_REG_14__SCAN_IN), .B2(keyinput111), .C1(
        P1_UWORD_REG_11__SCAN_IN), .C2(keyinput96), .A(n21346), .ZN(n21347) );
  NAND4_X1 U24247 ( .A1(n21350), .A2(n21349), .A3(n21348), .A4(n21347), .ZN(
        n21351) );
  NOR4_X1 U24248 ( .A1(n21354), .A2(n21353), .A3(n21352), .A4(n21351), .ZN(
        n21355) );
  NAND4_X1 U24249 ( .A1(n21358), .A2(n21357), .A3(n21356), .A4(n21355), .ZN(
        n21359) );
  NOR3_X1 U24250 ( .A1(n21361), .A2(n21360), .A3(n21359), .ZN(n21362) );
  XNOR2_X1 U24251 ( .A(n21363), .B(n21362), .ZN(P3_U2749) );
  NAND2_X1 U14456 ( .A1(n20028), .A2(n11988), .ZN(n12904) );
  INV_X1 U12646 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19237) );
  NAND2_X1 U12790 ( .A1(n14670), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11263) );
  CLKBUF_X1 U11262 ( .A(n11687), .Z(n15144) );
  CLKBUF_X1 U11286 ( .A(n13369), .Z(n13379) );
  INV_X1 U11287 ( .A(n17326), .ZN(n17300) );
  AND2_X1 U11311 ( .A1(n11425), .A2(n11458), .ZN(n12945) );
  CLKBUF_X1 U11315 ( .A(n12246), .Z(n9827) );
  INV_X1 U11323 ( .A(n17300), .ZN(n17245) );
  CLKBUF_X1 U11332 ( .A(n10448), .Z(n12513) );
  CLKBUF_X1 U11369 ( .A(n13515), .Z(n9846) );
  CLKBUF_X1 U11376 ( .A(n11510), .Z(n14281) );
  CLKBUF_X1 U11392 ( .A(n14457), .Z(n14516) );
  CLKBUF_X1 U11587 ( .A(n14534), .Z(n14535) );
  NAND2_X2 U11595 ( .A1(n14669), .A2(n11263), .ZN(n11275) );
  CLKBUF_X1 U11819 ( .A(n11446), .Z(n19355) );
  NAND2_X2 U11971 ( .A1(n9871), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18189) );
  CLKBUF_X1 U12167 ( .A(n20919), .Z(n20976) );
  CLKBUF_X1 U12333 ( .A(n16670), .Z(n16684) );
endmodule

