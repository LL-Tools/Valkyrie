

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2949, n2950, n2952, n2953, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771;

  AND2_X1 U3397 ( .A1(n5345), .A2(n2991), .ZN(n5185) );
  OR2_X1 U3398 ( .A1(n5446), .A2(n4099), .ZN(n6095) );
  XOR2_X2 U3399 ( .A(n5686), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .Z(n5680) );
  OR2_X1 U3400 ( .A1(n4181), .A2(n6744), .ZN(n3111) );
  BUF_X1 U3401 ( .A(n3996), .Z(n4087) );
  INV_X1 U3402 ( .A(n4000), .ZN(n4567) );
  CLKBUF_X2 U3403 ( .A(n3989), .Z(n4088) );
  AOI21_X1 U3404 ( .B1(n3393), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3286), 
        .ZN(n3390) );
  CLKBUF_X2 U3405 ( .A(n3293), .Z(n3900) );
  CLKBUF_X2 U3406 ( .A(n3326), .Z(n4585) );
  CLKBUF_X2 U3407 ( .A(n3349), .Z(n3405) );
  CLKBUF_X2 U3408 ( .A(n3891), .Z(n3776) );
  BUF_X2 U3409 ( .A(n3342), .Z(n3890) );
  BUF_X2 U3410 ( .A(n3292), .Z(n3892) );
  CLKBUF_X2 U3411 ( .A(n3287), .Z(n3815) );
  CLKBUF_X2 U3412 ( .A(n3341), .Z(n3846) );
  CLKBUF_X2 U3413 ( .A(n3847), .Z(n3897) );
  CLKBUF_X2 U3414 ( .A(n3294), .Z(n3816) );
  AND3_X1 U3415 ( .A1(n6771), .A2(n3233), .A3(n5445), .ZN(n3234) );
  CLKBUF_X2 U3416 ( .A(n3899), .Z(n3817) );
  AND2_X1 U3417 ( .A1(n3990), .A2(n4735), .ZN(n4251) );
  NOR2_X2 U3418 ( .A1(n4735), .A2(n3232), .ZN(n4499) );
  INV_X1 U3419 ( .A(n3237), .ZN(n3226) );
  AND4_X1 U3420 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3134)
         );
  AND4_X1 U3421 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3135)
         );
  AOI22_X1 U3422 ( .A1(n3292), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3142) );
  AND2_X1 U3423 ( .A1(n4579), .A2(n4510), .ZN(n2950) );
  AND2_X2 U3424 ( .A1(n4507), .A2(n4587), .ZN(n3292) );
  AND2_X2 U3425 ( .A1(n4587), .A2(n4509), .ZN(n3294) );
  AND2_X2 U3426 ( .A1(n4522), .A2(n4582), .ZN(n3847) );
  AND2_X2 U3427 ( .A1(n3044), .A2(n2982), .ZN(n5609) );
  NAND2_X1 U3428 ( .A1(n5664), .A2(n5663), .ZN(n2949) );
  NAND2_X1 U3429 ( .A1(n5664), .A2(n5663), .ZN(n5662) );
  XNOR2_X1 U3430 ( .A(n2995), .B(n5779), .ZN(n5635) );
  AND2_X1 U3431 ( .A1(n4579), .A2(n4510), .ZN(n3400) );
  AND2_X2 U3433 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4579) );
  NOR2_X1 U3434 ( .A1(n4000), .A2(n3991), .ZN(n3996) );
  NAND2_X1 U3436 ( .A1(n3109), .A2(n2964), .ZN(n3232) );
  NAND2_X2 U3437 ( .A1(n3116), .A2(n2966), .ZN(n4141) );
  AND2_X1 U3438 ( .A1(n4158), .A2(n4157), .ZN(n4755) );
  OAI21_X1 U3439 ( .B1(n4145), .B2(n4196), .A(n4144), .ZN(n4545) );
  OR2_X1 U3440 ( .A1(n4500), .A2(n3977), .ZN(n4464) );
  INV_X1 U3442 ( .A(n6073), .ZN(n6108) );
  AND2_X2 U3443 ( .A1(n4509), .A2(n4579), .ZN(n3899) );
  BUF_X2 U3444 ( .A(n3343), .Z(n3344) );
  INV_X4 U34450 ( .A(n3989), .ZN(n3991) );
  OAI21_X4 U34460 ( .B1(n4359), .B2(n4358), .A(n4357), .ZN(n5393) );
  AND2_X4 U34470 ( .A1(n3068), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4582) );
  AOI21_X2 U34480 ( .B1(n5609), .B2(n5171), .A(n4389), .ZN(n4390) );
  NAND2_X2 U3449 ( .A1(n3302), .A2(n3301), .ZN(n3306) );
  AOI22_X1 U3450 ( .A1(n5144), .A2(n5578), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6710), .ZN(n5145) );
  OR2_X1 U34510 ( .A1(n4340), .A2(n5882), .ZN(n4301) );
  NAND2_X1 U34520 ( .A1(n2997), .A2(n2996), .ZN(n5643) );
  NAND2_X1 U34530 ( .A1(n4303), .A2(n4302), .ZN(n5577) );
  AND2_X1 U3454 ( .A1(n4386), .A2(n4388), .ZN(n4389) );
  XNOR2_X1 U34550 ( .A(n4310), .B(n4309), .ZN(n5126) );
  OR2_X1 U34560 ( .A1(n5299), .A2(n5288), .ZN(n5286) );
  OR2_X1 U3457 ( .A1(n5174), .A2(n5301), .ZN(n5299) );
  AND2_X1 U3458 ( .A1(n4420), .A2(n4419), .ZN(n4421) );
  OR2_X1 U34590 ( .A1(n5707), .A2(n3075), .ZN(n3074) );
  NOR2_X1 U34600 ( .A1(n3018), .A2(n3020), .ZN(n3017) );
  CLKBUF_X1 U34610 ( .A(n5226), .Z(n5234) );
  AND2_X1 U34620 ( .A1(n4356), .A2(n4355), .ZN(n6073) );
  OAI211_X1 U34630 ( .C1(n3437), .C2(n3080), .A(n3118), .B(n3078), .ZN(n4180)
         );
  OR2_X1 U34640 ( .A1(n3112), .A2(n5301), .ZN(n3748) );
  OAI21_X1 U34650 ( .B1(n3377), .B2(n3378), .A(n3379), .ZN(n3365) );
  NAND2_X1 U3466 ( .A1(n3371), .A2(n3363), .ZN(n3379) );
  NAND2_X1 U3467 ( .A1(n4030), .A2(n4029), .ZN(n5404) );
  NOR2_X1 U34680 ( .A1(n6129), .A2(n4735), .ZN(n4660) );
  XNOR2_X1 U34690 ( .A(n3392), .B(n3390), .ZN(n4525) );
  OAI21_X1 U34700 ( .B1(n3372), .B2(STATE2_REG_0__SCAN_IN), .A(n3367), .ZN(
        n3362) );
  NAND2_X2 U34710 ( .A1(n3975), .A2(n3974), .ZN(n4680) );
  NAND3_X1 U34720 ( .A1(n3253), .A2(n3278), .A3(n3281), .ZN(n3307) );
  NAND2_X1 U34730 ( .A1(n4005), .A2(n4004), .ZN(n4705) );
  NAND2_X1 U34740 ( .A1(n3263), .A2(n3262), .ZN(n3336) );
  OR2_X1 U3475 ( .A1(n3261), .A2(n3260), .ZN(n3262) );
  NAND2_X1 U3476 ( .A1(n3399), .A2(n3398), .ZN(n3969) );
  AND2_X1 U3477 ( .A1(n3225), .A2(n4416), .ZN(n4265) );
  AND2_X1 U3478 ( .A1(n3026), .A2(n4251), .ZN(n3024) );
  AND2_X1 U3479 ( .A1(n3224), .A2(n4416), .ZN(n3250) );
  NAND2_X1 U3480 ( .A1(n4735), .A2(n4235), .ZN(n5445) );
  INV_X1 U3481 ( .A(n3232), .ZN(n3990) );
  BUF_X2 U3482 ( .A(n3237), .Z(n4247) );
  OR2_X2 U3483 ( .A1(n3172), .A2(n3171), .ZN(n4416) );
  AND4_X1 U3484 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3190)
         );
  AND4_X1 U3485 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3192)
         );
  AND4_X1 U3486 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3189)
         );
  AND4_X1 U3487 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3162)
         );
  AND4_X1 U3488 ( .A1(n3204), .A2(n3203), .A3(n3202), .A4(n3201), .ZN(n3220)
         );
  AND4_X1 U3489 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3219)
         );
  AND4_X1 U3490 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3218)
         );
  AND4_X1 U3491 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3217)
         );
  BUF_X2 U3492 ( .A(n3438), .Z(n3871) );
  BUF_X2 U3493 ( .A(n3889), .Z(n3696) );
  NAND2_X1 U3494 ( .A1(n6733), .A2(n5034), .ZN(n6593) );
  NAND2_X1 U3495 ( .A1(n3365), .A2(n3364), .ZN(n3416) );
  NAND2_X2 U3496 ( .A1(n4149), .A2(n4148), .ZN(n6213) );
  AND2_X1 U3497 ( .A1(n4579), .A2(n4507), .ZN(n2952) );
  AND2_X1 U3498 ( .A1(n4579), .A2(n4507), .ZN(n3343) );
  BUF_X1 U3499 ( .A(n3283), .Z(n3393) );
  AND2_X4 U3500 ( .A1(n4582), .A2(n4510), .ZN(n3891) );
  OAI22_X2 U3501 ( .A1(n4197), .A2(n4196), .B1(n4195), .B2(n6600), .ZN(n4198)
         );
  NAND3_X2 U3502 ( .A1(n3070), .A2(n5723), .A3(n3069), .ZN(n5722) );
  NAND2_X2 U3503 ( .A1(n5722), .A2(n4199), .ZN(n5716) );
  OR2_X1 U3504 ( .A1(n3236), .A2(n4247), .ZN(n3230) );
  NAND2_X1 U3505 ( .A1(n3282), .A2(n3308), .ZN(n3392) );
  BUF_X2 U3506 ( .A(n4124), .Z(n2953) );
  AND2_X4 U3507 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4510) );
  NOR2_X2 U3508 ( .A1(n4320), .A2(n5671), .ZN(n5664) );
  INV_X2 U3509 ( .A(n3926), .ZN(n3231) );
  AND2_X1 U3510 ( .A1(n4587), .A2(n4510), .ZN(n2956) );
  OR2_X1 U3511 ( .A1(n3463), .A2(n3087), .ZN(n3086) );
  OR2_X1 U3512 ( .A1(n4247), .A2(n6513), .ZN(n3398) );
  INV_X1 U3513 ( .A(n4403), .ZN(n3100) );
  AND2_X1 U3514 ( .A1(n3047), .A2(n2981), .ZN(n3046) );
  OR2_X1 U3515 ( .A1(n2965), .A2(n5625), .ZN(n3047) );
  NAND2_X1 U3516 ( .A1(n4680), .A2(n6517), .ZN(n4500) );
  INV_X1 U3517 ( .A(n3462), .ZN(n3087) );
  NAND2_X1 U3519 ( .A1(n3436), .A2(n3435), .ZN(n3463) );
  NOR2_X1 U3520 ( .A1(n4121), .A2(n3106), .ZN(n3105) );
  INV_X1 U3521 ( .A(n5314), .ZN(n3102) );
  NOR3_X1 U3522 ( .A1(n4702), .A2(n4639), .A3(n2977), .ZN(n3004) );
  AND2_X1 U3523 ( .A1(n3104), .A2(n5401), .ZN(n3103) );
  INV_X1 U3524 ( .A(n3986), .ZN(n3828) );
  NOR2_X1 U3525 ( .A1(n4345), .A2(n4086), .ZN(n4350) );
  AND2_X1 U3526 ( .A1(n4567), .A2(n4084), .ZN(n4085) );
  OR2_X2 U3527 ( .A1(n4141), .A2(n4735), .ZN(n4080) );
  INV_X1 U3528 ( .A(n3398), .ZN(n4127) );
  OR2_X1 U3529 ( .A1(n3332), .A2(n3331), .ZN(n4202) );
  NAND2_X1 U3530 ( .A1(n3397), .A2(n3396), .ZN(n4937) );
  AND3_X1 U3531 ( .A1(n4725), .A2(n3231), .A3(n4721), .ZN(n4412) );
  OR2_X1 U3532 ( .A1(n4242), .A2(n5428), .ZN(n4527) );
  AND2_X1 U3533 ( .A1(n5034), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3915) );
  NAND2_X1 U3534 ( .A1(n3508), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3525)
         );
  OR2_X1 U3535 ( .A1(n4350), .A2(n3991), .ZN(n4344) );
  NAND2_X1 U3536 ( .A1(n5686), .A2(n5142), .ZN(n4302) );
  NOR2_X1 U3537 ( .A1(n4054), .A2(n3059), .ZN(n3058) );
  INV_X1 U3538 ( .A(n5316), .ZN(n3059) );
  AOI21_X1 U3539 ( .B1(n3046), .B2(n5625), .A(n2980), .ZN(n3045) );
  NAND2_X1 U3540 ( .A1(n3094), .A2(n3046), .ZN(n3044) );
  NAND2_X1 U3541 ( .A1(n2958), .A2(n2989), .ZN(n3063) );
  NAND2_X2 U3542 ( .A1(n4088), .A2(n4080), .ZN(n4551) );
  OR2_X1 U3543 ( .A1(n4241), .A2(n4772), .ZN(n4276) );
  INV_X1 U3544 ( .A(n2955), .ZN(n4941) );
  NAND2_X1 U3545 ( .A1(n3973), .A2(n3979), .ZN(n3974) );
  AOI21_X1 U3546 ( .B1(n6073), .B2(n6187), .A(n3013), .ZN(n4432) );
  AND2_X1 U3547 ( .A1(n6087), .A2(n6189), .ZN(n3013) );
  INV_X1 U3548 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6648) );
  INV_X1 U3549 ( .A(n5882), .ZN(n6294) );
  AND2_X1 U3550 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  INV_X1 U3551 ( .A(n4430), .ZN(n3104) );
  CLKBUF_X1 U3552 ( .A(n3314), .Z(n3558) );
  XNOR2_X1 U3553 ( .A(n4200), .B(n3503), .ZN(n4192) );
  OR2_X1 U3554 ( .A1(n3475), .A2(n3474), .ZN(n4193) );
  NOR2_X1 U3555 ( .A1(n3082), .A2(n4196), .ZN(n3079) );
  NOR2_X1 U3556 ( .A1(n3083), .A2(n3085), .ZN(n3082) );
  NAND2_X1 U3557 ( .A1(n3086), .A2(n3087), .ZN(n3084) );
  NAND2_X1 U3558 ( .A1(n4141), .A2(n3232), .ZN(n3989) );
  NAND2_X1 U3559 ( .A1(n3236), .A2(n4141), .ZN(n3271) );
  AOI22_X1 U3560 ( .A1(n3438), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3899), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U3561 ( .A1(n3847), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U3562 ( .A1(n3349), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U3563 ( .A1(n3342), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3133) );
  AND2_X1 U3564 ( .A1(n4256), .A2(n4255), .ZN(n4271) );
  NOR2_X1 U3565 ( .A1(n3676), .A2(n5332), .ZN(n3012) );
  INV_X1 U3566 ( .A(n3692), .ZN(n3743) );
  AND2_X1 U3567 ( .A1(n5227), .A2(n3062), .ZN(n3061) );
  INV_X1 U3568 ( .A(n5147), .ZN(n3062) );
  NOR2_X2 U3569 ( .A1(n5246), .A2(n5235), .ZN(n5226) );
  NAND2_X1 U3570 ( .A1(n3091), .A2(n4217), .ZN(n3090) );
  NAND2_X1 U3571 ( .A1(n2965), .A2(n4219), .ZN(n3091) );
  INV_X1 U3572 ( .A(n5289), .ZN(n3057) );
  NOR2_X1 U3573 ( .A1(n3040), .A2(n3041), .ZN(n3039) );
  NOR2_X1 U3574 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3041)
         );
  INV_X1 U3575 ( .A(n4322), .ZN(n3040) );
  INV_X1 U3576 ( .A(n4208), .ZN(n3075) );
  AND2_X1 U3577 ( .A1(n3051), .A2(n4974), .ZN(n3054) );
  INV_X1 U3578 ( .A(n3055), .ZN(n3051) );
  OR2_X1 U3579 ( .A1(n4276), .A2(n4269), .ZN(n4554) );
  OAI21_X1 U3580 ( .B1(n5070), .B2(n3020), .A(n3019), .ZN(n3021) );
  INV_X1 U3581 ( .A(n4175), .ZN(n3018) );
  NAND2_X1 U3582 ( .A1(n3053), .A2(n3054), .ZN(n4980) );
  INV_X1 U3583 ( .A(n4705), .ZN(n3053) );
  INV_X1 U3584 ( .A(n4068), .ZN(n4079) );
  AND2_X1 U3585 ( .A1(n4567), .A2(n3991), .ZN(n4068) );
  OAI211_X1 U3586 ( .C1(n4202), .C2(n3398), .A(n3335), .B(n3334), .ZN(n3378)
         );
  OR2_X1 U3587 ( .A1(n3300), .A2(n3299), .ZN(n4159) );
  NAND2_X1 U3588 ( .A1(n3227), .A2(n3026), .ZN(n3025) );
  AND2_X1 U3589 ( .A1(n6347), .A2(n6446), .ZN(n4847) );
  XNOR2_X1 U3590 ( .A(n3920), .B(n4114), .ZN(n4356) );
  NAND2_X1 U3591 ( .A1(n3919), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3920)
         );
  NOR2_X1 U3592 ( .A1(n3642), .A2(n3591), .ZN(n3609) );
  NAND2_X1 U3593 ( .A1(n5191), .A2(n6513), .ZN(n4312) );
  NAND2_X1 U3594 ( .A1(n4564), .A2(n2972), .ZN(n3387) );
  INV_X1 U3595 ( .A(n5611), .ZN(n3043) );
  AND2_X1 U3596 ( .A1(n4051), .A2(n4323), .ZN(n5303) );
  INV_X1 U3597 ( .A(n3096), .ZN(n4320) );
  NAND2_X1 U3598 ( .A1(n3073), .A2(n2976), .ZN(n3072) );
  NAND2_X1 U3599 ( .A1(n3077), .A2(n4208), .ZN(n3076) );
  INV_X1 U3600 ( .A(n4426), .ZN(n4029) );
  INV_X1 U3601 ( .A(n5819), .ZN(n5872) );
  NAND2_X1 U3602 ( .A1(n5069), .A2(n3111), .ZN(n6197) );
  NAND2_X1 U3603 ( .A1(n6197), .A2(n6196), .ZN(n6195) );
  NAND2_X1 U3604 ( .A1(n4136), .A2(n4201), .ZN(n3015) );
  NAND2_X1 U3605 ( .A1(n3978), .A2(n4467), .ZN(n4662) );
  INV_X1 U3606 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6733) );
  CLKBUF_X1 U3607 ( .A(n4580), .Z(n6347) );
  OR2_X1 U3608 ( .A1(n4936), .A2(n5884), .ZN(n4942) );
  AND3_X1 U3609 ( .A1(n6312), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U3610 ( .A1(n4617), .A2(n6513), .ZN(n5033) );
  NAND2_X1 U3611 ( .A1(n5899), .A2(n4616), .ZN(n4617) );
  AND2_X1 U3612 ( .A1(n4526), .A2(n4846), .ZN(n5039) );
  NOR2_X1 U3613 ( .A1(n4996), .A2(n5034), .ZN(n6396) );
  INV_X2 U3614 ( .A(n3221), .ZN(n4721) );
  AND3_X1 U3615 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n5032) );
  AOI21_X1 U3616 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6390), .A(n5033), .ZN(
        n4944) );
  CLKBUF_X1 U3617 ( .A(n4153), .Z(n4899) );
  INV_X1 U3618 ( .A(n3412), .ZN(n3413) );
  NAND2_X1 U3619 ( .A1(n5884), .A2(n4941), .ZN(n6304) );
  NOR2_X2 U3620 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3986) );
  NOR2_X2 U3621 ( .A1(n4359), .A2(n4097), .ZN(n6082) );
  INV_X1 U3622 ( .A(n6098), .ZN(n6068) );
  INV_X1 U3623 ( .A(n6082), .ZN(n6101) );
  NOR2_X1 U3624 ( .A1(n4356), .A2(n4354), .ZN(n6087) );
  AND2_X1 U3625 ( .A1(n5441), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6098) );
  OAI211_X1 U3626 ( .C1(n4500), .C2(n4527), .A(n4131), .B(n6611), .ZN(n5560)
         );
  XNOR2_X1 U3627 ( .A(n3107), .B(n3917), .ZN(n5166) );
  INV_X1 U3628 ( .A(n3916), .ZN(n3917) );
  INV_X1 U3629 ( .A(n3919), .ZN(n3918) );
  NAND2_X1 U3630 ( .A1(n3002), .A2(n4120), .ZN(n5213) );
  NAND2_X1 U3631 ( .A1(n3003), .A2(n3106), .ZN(n3002) );
  OR2_X1 U3632 ( .A1(n4401), .A2(n4404), .ZN(n5537) );
  NAND2_X1 U3633 ( .A1(n3540), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3541)
         );
  OR2_X1 U3634 ( .A1(n4500), .A2(n4689), .ZN(n6192) );
  INV_X1 U3635 ( .A(n5727), .ZN(n6212) );
  INV_X1 U3636 ( .A(n6192), .ZN(n6219) );
  XNOR2_X1 U3637 ( .A(n4096), .B(n4095), .ZN(n5204) );
  AND2_X1 U3638 ( .A1(n4344), .A2(n4093), .ZN(n4096) );
  AND2_X1 U3639 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5139)
         );
  NAND2_X1 U3640 ( .A1(n4465), .A2(n6513), .ZN(n6211) );
  AND4_X1 U3641 ( .A1(n4679), .A2(n2953), .A3(n4245), .A4(n4244), .ZN(n4246)
         );
  OR2_X1 U3642 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  INV_X1 U3643 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6390) );
  CLKBUF_X1 U3644 ( .A(n4136), .Z(n5884) );
  INV_X1 U3645 ( .A(n6593), .ZN(n6442) );
  CLKBUF_X1 U3646 ( .A(n4525), .Z(n4526) );
  NAND2_X1 U3647 ( .A1(n4900), .A2(n5887), .ZN(n6444) );
  INV_X1 U3648 ( .A(n6347), .ZN(n6384) );
  INV_X1 U3649 ( .A(n5902), .ZN(n5200) );
  AND2_X1 U3650 ( .A1(n3087), .A2(n3463), .ZN(n3085) );
  AND2_X1 U3651 ( .A1(n6390), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3935)
         );
  INV_X1 U3652 ( .A(n3111), .ZN(n3020) );
  INV_X1 U3653 ( .A(n3499), .ZN(n3500) );
  OR2_X1 U3654 ( .A1(n3254), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3257)
         );
  AND2_X1 U3655 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3257), .ZN(n3255) );
  OR2_X1 U3656 ( .A1(n3320), .A2(n3319), .ZN(n4137) );
  NAND2_X1 U3657 ( .A1(n3248), .A2(n3247), .ZN(n4252) );
  INV_X1 U3658 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U3659 ( .A1(n3326), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3660 ( .A1(n3303), .A2(n4201), .ZN(n3963) );
  INV_X1 U3661 ( .A(n3980), .ZN(n3964) );
  OR3_X1 U3662 ( .A1(n3966), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6303), 
        .ZN(n3980) );
  NOR2_X1 U3663 ( .A1(n3863), .A2(n5582), .ZN(n3864) );
  AND2_X1 U3664 ( .A1(n3802), .A2(n3801), .ZN(n3825) );
  NOR2_X1 U3665 ( .A1(n3711), .A2(n3710), .ZN(n3010) );
  NAND2_X1 U3666 ( .A1(n4519), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3910) );
  INV_X1 U3667 ( .A(n3910), .ZN(n3884) );
  OR2_X1 U3668 ( .A1(n3577), .A2(n3576), .ZN(n3590) );
  NOR2_X1 U3669 ( .A1(n6648), .A2(n3007), .ZN(n3006) );
  INV_X1 U3670 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6730) );
  CLKBUF_X1 U3671 ( .A(n3249), .Z(n4264) );
  INV_X1 U3672 ( .A(n5626), .ZN(n3093) );
  INV_X1 U3673 ( .A(n5715), .ZN(n3077) );
  AND2_X1 U3674 ( .A1(n3067), .A2(n5507), .ZN(n3066) );
  INV_X1 U3675 ( .A(n5403), .ZN(n3067) );
  INV_X1 U3676 ( .A(n5404), .ZN(n3065) );
  INV_X1 U3677 ( .A(n4752), .ZN(n3056) );
  NAND2_X1 U3678 ( .A1(n3084), .A2(n4201), .ZN(n3080) );
  INV_X1 U3679 ( .A(n4642), .ZN(n4005) );
  AND2_X1 U3680 ( .A1(n5840), .A2(n4554), .ZN(n5813) );
  AND2_X1 U3681 ( .A1(n3992), .A2(n3049), .ZN(n3048) );
  NAND2_X1 U3682 ( .A1(n3996), .A2(n3993), .ZN(n3050) );
  NAND2_X1 U3683 ( .A1(n3991), .A2(EBX_REG_1__SCAN_IN), .ZN(n3049) );
  OR2_X1 U3684 ( .A1(n3356), .A2(n3355), .ZN(n4142) );
  NOR2_X1 U3685 ( .A1(n3264), .A2(n3275), .ZN(n3276) );
  AND2_X1 U3686 ( .A1(n3241), .A2(n3240), .ZN(n3278) );
  AND2_X1 U3687 ( .A1(n3245), .A2(n4230), .ZN(n3023) );
  OR2_X1 U3688 ( .A1(n3236), .A2(n3592), .ZN(n4663) );
  INV_X1 U3689 ( .A(n3373), .ZN(n6446) );
  NAND4_X1 U3690 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3237)
         );
  AOI22_X1 U3691 ( .A1(n3292), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3132) );
  OR2_X1 U3692 ( .A1(n3411), .A2(n3410), .ZN(n4169) );
  AND2_X1 U3693 ( .A1(n4608), .A2(n4607), .ZN(n4612) );
  INV_X1 U3694 ( .A(n3963), .ZN(n3973) );
  AND2_X1 U3695 ( .A1(n3968), .A2(n3967), .ZN(n3979) );
  OR2_X1 U3696 ( .A1(n3966), .A2(n3965), .ZN(n3968) );
  AND2_X1 U3697 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6303), .ZN(n3965)
         );
  OR2_X1 U3698 ( .A1(n4684), .A2(n4678), .ZN(n4460) );
  INV_X1 U3699 ( .A(n4499), .ZN(n6600) );
  OR2_X1 U3700 ( .A1(n5446), .A2(n4112), .ZN(n4359) );
  INV_X1 U3701 ( .A(n4492), .ZN(n4686) );
  NAND2_X1 U3702 ( .A1(n5441), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5446) );
  INV_X1 U3703 ( .A(n4619), .ZN(n4614) );
  INV_X1 U3704 ( .A(n4464), .ZN(n4498) );
  NOR2_X1 U3705 ( .A1(n4416), .A2(n5034), .ZN(n3573) );
  NOR2_X1 U3706 ( .A1(n3912), .A2(n5573), .ZN(n3919) );
  NAND2_X1 U3707 ( .A1(n3864), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3912)
         );
  OR2_X1 U3708 ( .A1(n2970), .A2(n5595), .ZN(n3809) );
  OR2_X1 U3709 ( .A1(n3809), .A2(n3808), .ZN(n3863) );
  INV_X1 U3710 ( .A(n5258), .ZN(n3099) );
  NAND2_X1 U3711 ( .A1(n3010), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3806)
         );
  NAND2_X1 U3712 ( .A1(n3011), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3711)
         );
  INV_X1 U3713 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3710) );
  INV_X1 U3714 ( .A(n3010), .ZN(n3773) );
  NAND2_X1 U3715 ( .A1(n3012), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3730)
         );
  INV_X1 U3716 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U3717 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3676)
         );
  INV_X1 U3718 ( .A(n3012), .ZN(n3709) );
  NAND2_X1 U3719 ( .A1(n3571), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3642)
         );
  AND2_X1 U3720 ( .A1(n3652), .A2(n3589), .ZN(n5510) );
  AND3_X1 U3721 ( .A1(n3554), .A2(n3553), .A3(n3552), .ZN(n3555) );
  NOR2_X1 U3722 ( .A1(n3525), .A2(n5415), .ZN(n3540) );
  AND2_X1 U3723 ( .A1(n3477), .A2(n2985), .ZN(n3508) );
  NAND2_X1 U3724 ( .A1(n3477), .A2(n2959), .ZN(n3504) );
  NOR2_X1 U3725 ( .A1(n4882), .A2(n4883), .ZN(n4892) );
  NOR2_X1 U3726 ( .A1(n3419), .A2(n6730), .ZN(n3454) );
  NAND2_X1 U3727 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3419) );
  INV_X1 U3728 ( .A(n4344), .ZN(n4352) );
  AND2_X1 U3729 ( .A1(n5226), .A2(n2993), .ZN(n5205) );
  INV_X1 U3730 ( .A(n5206), .ZN(n3060) );
  NAND2_X1 U3731 ( .A1(n3042), .A2(n3088), .ZN(n5141) );
  AND2_X1 U3732 ( .A1(n3090), .A2(n3089), .ZN(n3088) );
  NAND2_X1 U3733 ( .A1(n3092), .A2(n5672), .ZN(n3089) );
  AND2_X1 U3734 ( .A1(n4071), .A2(n4070), .ZN(n5249) );
  NAND2_X1 U3735 ( .A1(n4378), .A2(n4072), .ZN(n5246) );
  INV_X1 U3736 ( .A(n5249), .ZN(n4072) );
  AND2_X1 U3737 ( .A1(n5653), .A2(n5803), .ZN(n2996) );
  INV_X1 U3738 ( .A(n5662), .ZN(n2997) );
  NAND2_X1 U3739 ( .A1(n2949), .A2(n2960), .ZN(n5645) );
  NAND2_X1 U3740 ( .A1(n3065), .A2(n2958), .ZN(n5389) );
  INV_X1 U3741 ( .A(n3074), .ZN(n3036) );
  INV_X1 U3742 ( .A(n4211), .ZN(n3034) );
  NAND2_X1 U3743 ( .A1(n3065), .A2(n3066), .ZN(n5387) );
  AND2_X1 U3744 ( .A1(n4283), .A2(n4282), .ZN(n5843) );
  AND2_X1 U3745 ( .A1(n4028), .A2(n4027), .ZN(n4426) );
  OR2_X1 U3746 ( .A1(n5716), .A2(n3074), .ZN(n3038) );
  AND2_X1 U3747 ( .A1(n4277), .A2(n4572), .ZN(n5866) );
  NAND2_X1 U3748 ( .A1(n6206), .A2(n4175), .ZN(n5071) );
  AOI21_X1 U3749 ( .B1(n4566), .B2(n4567), .A(n3995), .ZN(n4644) );
  OR2_X1 U3750 ( .A1(n4276), .A2(n4681), .ZN(n5867) );
  NOR2_X1 U3751 ( .A1(n6593), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4465) );
  XNOR2_X1 U3752 ( .A(n3379), .B(n3378), .ZN(n3016) );
  AOI22_X1 U3753 ( .A1(n3304), .A2(n4159), .B1(n3303), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3305) );
  INV_X1 U3754 ( .A(n4663), .ZN(n4519) );
  AND2_X1 U3755 ( .A1(n4482), .A2(n4481), .ZN(n4666) );
  NOR2_X1 U3756 ( .A1(n6307), .A2(n5884), .ZN(n4904) );
  OR2_X1 U3757 ( .A1(n5981), .A2(n6347), .ZN(n5087) );
  AND2_X1 U3758 ( .A1(n4904), .A2(n4941), .ZN(n5084) );
  OR2_X1 U3759 ( .A1(n4900), .A2(n4899), .ZN(n6307) );
  OAI21_X1 U3760 ( .B1(n4942), .B2(n6028), .A(n6442), .ZN(n6354) );
  OR2_X1 U3761 ( .A1(n4526), .A2(n4846), .ZN(n5941) );
  NOR2_X1 U3762 ( .A1(n6444), .A2(n5884), .ZN(n4849) );
  AND2_X1 U3763 ( .A1(n5982), .A2(n6347), .ZN(n6447) );
  OR2_X1 U3764 ( .A1(n5033), .A2(n6733), .ZN(n4743) );
  INV_X1 U3765 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6312) );
  AND2_X1 U3766 ( .A1(n5194), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3976) );
  NAND2_X1 U3767 ( .A1(n6513), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4311) );
  AND2_X1 U3768 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4619) );
  OR2_X1 U3769 ( .A1(n4130), .A2(n6600), .ZN(n4698) );
  NOR2_X1 U3770 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6601) );
  INV_X1 U3771 ( .A(n6087), .ZN(n6059) );
  OR2_X1 U3772 ( .A1(n4417), .A2(n5519), .ZN(n4420) );
  INV_X1 U3773 ( .A(n5519), .ZN(n5514) );
  INV_X1 U3774 ( .A(n5517), .ZN(n5504) );
  NAND2_X1 U3775 ( .A1(n4415), .A2(n4414), .ZN(n5517) );
  OR3_X1 U3776 ( .A1(n4680), .A2(n4772), .A3(n4681), .ZN(n4415) );
  NAND2_X1 U3777 ( .A1(n5517), .A2(n5164), .ZN(n5519) );
  AND2_X1 U3778 ( .A1(n5560), .A2(n3250), .ZN(n5554) );
  AND2_X1 U3779 ( .A1(n5560), .A2(n4133), .ZN(n5555) );
  INV_X2 U3780 ( .A(n5560), .ZN(n5564) );
  NAND2_X2 U3781 ( .A1(n5560), .A2(n4132), .ZN(n5567) );
  CLKBUF_X2 U3782 ( .A(n4636), .Z(n6592) );
  INV_X2 U3783 ( .A(n4560), .ZN(n6127) );
  OR3_X2 U3784 ( .A1(n4500), .A2(READY_N), .A3(n4245), .ZN(n6611) );
  INV_X1 U3785 ( .A(n6130), .ZN(n6608) );
  INV_X1 U3786 ( .A(n4308), .ZN(n4309) );
  INV_X1 U3787 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5582) );
  INV_X1 U3788 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5595) );
  INV_X1 U3789 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5604) );
  OAI21_X1 U3790 ( .B1(n5342), .B2(n5330), .A(n3101), .ZN(n5641) );
  NAND2_X1 U3791 ( .A1(n6192), .A2(n4314), .ZN(n5727) );
  INV_X1 U3792 ( .A(n6223), .ZN(n6188) );
  AND2_X1 U3793 ( .A1(n4882), .A2(n4750), .ZN(n6207) );
  INV_X1 U3794 ( .A(n6211), .ZN(n6194) );
  NOR2_X1 U3795 ( .A1(n4376), .A2(n4375), .ZN(n5608) );
  AND2_X1 U3796 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U3797 ( .A(n5173), .B(n3110), .ZN(n5190) );
  AND2_X1 U3798 ( .A1(n5686), .A2(n5169), .ZN(n5170) );
  OR2_X1 U3799 ( .A1(n5799), .A2(n4288), .ZN(n5773) );
  NAND2_X1 U3800 ( .A1(n5345), .A2(n3058), .ZN(n5290) );
  NAND2_X1 U3801 ( .A1(n3044), .A2(n3045), .ZN(n5610) );
  NAND2_X1 U3802 ( .A1(n5345), .A2(n5316), .ZN(n5302) );
  NAND2_X1 U3803 ( .A1(n5645), .A2(n5643), .ZN(n2995) );
  INV_X1 U3804 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U3805 ( .A1(n2949), .A2(n4322), .ZN(n5655) );
  INV_X1 U3806 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U3807 ( .A1(n5843), .A2(n4285), .ZN(n6231) );
  OR2_X1 U3808 ( .A1(n5840), .A2(n4284), .ZN(n4285) );
  NAND2_X1 U3809 ( .A1(n6195), .A2(n4191), .ZN(n5724) );
  INV_X1 U3810 ( .A(n5867), .ZN(n6290) );
  CLKBUF_X1 U3811 ( .A(n3372), .Z(n3373) );
  OR2_X1 U3812 ( .A1(n6593), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5896) );
  INV_X1 U3813 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6303) );
  INV_X1 U3814 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U3815 ( .A1(n4680), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5899) );
  NOR2_X1 U3816 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5191) );
  OR2_X1 U3817 ( .A1(n4489), .A2(n4486), .ZN(n5902) );
  INV_X1 U3818 ( .A(n5939), .ZN(n4931) );
  OAI211_X1 U3819 ( .C1(n6401), .C2(n6400), .A(n6399), .B(n6398), .ZN(n6435)
         );
  INV_X1 U3820 ( .A(n5975), .ZN(n4803) );
  INV_X1 U3821 ( .A(n6438), .ZN(n6393) );
  INV_X1 U3822 ( .A(n5940), .ZN(n5978) );
  NAND2_X1 U3823 ( .A1(n4849), .A2(n4941), .ZN(n5984) );
  INV_X1 U3824 ( .A(n6440), .ZN(n6403) );
  INV_X1 U3825 ( .A(n6480), .ZN(n6419) );
  INV_X1 U3826 ( .A(n5984), .ZN(n6020) );
  INV_X1 U3827 ( .A(n6511), .ZN(n6434) );
  AOI22_X1 U3828 ( .A1(n5986), .A2(n6447), .B1(n6396), .B2(n5983), .ZN(n6025)
         );
  NAND2_X1 U3829 ( .A1(n6217), .A2(DATAI_16_), .ZN(n6457) );
  NOR2_X1 U3830 ( .A1(n5033), .A2(n6154), .ZN(n6454) );
  NAND2_X1 U3831 ( .A1(n6217), .A2(DATAI_17_), .ZN(n6459) );
  NOR2_X1 U3832 ( .A1(n5033), .A2(n6156), .ZN(n6461) );
  NAND2_X1 U3833 ( .A1(n6217), .A2(DATAI_18_), .ZN(n6466) );
  NOR2_X1 U3834 ( .A1(n5033), .A2(n6160), .ZN(n6475) );
  NAND2_X1 U3835 ( .A1(n6217), .A2(DATAI_20_), .ZN(n6485) );
  NOR2_X1 U3836 ( .A1(n5033), .A2(n6162), .ZN(n6482) );
  NOR2_X1 U3837 ( .A1(n5033), .A2(n6164), .ZN(n6489) );
  NAND2_X1 U3838 ( .A1(n6217), .A2(DATAI_22_), .ZN(n6499) );
  NOR2_X1 U3839 ( .A1(n5033), .A2(n6166), .ZN(n6496) );
  OR2_X1 U3840 ( .A1(n6444), .A2(n5979), .ZN(n6510) );
  NAND2_X1 U3841 ( .A1(n6217), .A2(DATAI_23_), .ZN(n6502) );
  OAI211_X1 U3842 ( .C1(n4994), .C2(n4993), .A(n5945), .B(n4992), .ZN(n5020)
         );
  INV_X1 U3843 ( .A(n4816), .ZN(n4841) );
  OAI21_X1 U3844 ( .B1(n5037), .B2(n5036), .A(n5035), .ZN(n5061) );
  INV_X1 U3845 ( .A(n6454), .ZN(n5993) );
  INV_X1 U3846 ( .A(n6468), .ZN(n6001) );
  OR2_X1 U3847 ( .A1(n4743), .A2(n4721), .ZN(n6465) );
  INV_X1 U3848 ( .A(n6475), .ZN(n6005) );
  OR2_X1 U3849 ( .A1(n4743), .A2(n3226), .ZN(n6479) );
  INV_X1 U3850 ( .A(n6482), .ZN(n6009) );
  OR2_X1 U3851 ( .A1(n4743), .A2(n3231), .ZN(n6486) );
  INV_X1 U3852 ( .A(n6489), .ZN(n6013) );
  OR2_X1 U3853 ( .A1(n4743), .A2(n3242), .ZN(n6493) );
  OR2_X1 U3854 ( .A1(n4711), .A2(n4941), .ZN(n5038) );
  NAND2_X1 U3855 ( .A1(n5032), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4744) );
  INV_X1 U3856 ( .A(n6506), .ZN(n6024) );
  OR2_X1 U3857 ( .A1(n4743), .A2(n5164), .ZN(n6501) );
  OAI211_X1 U3858 ( .C1(n5032), .C2(n6442), .A(n4714), .B(n4944), .ZN(n4742)
         );
  AND2_X1 U3859 ( .A1(n4715), .A2(n4899), .ZN(n5936) );
  INV_X1 U3860 ( .A(n6517), .ZN(n4772) );
  INV_X2 U3861 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6513) );
  AND2_X1 U3862 ( .A1(n4458), .A2(n6606), .ZN(n6576) );
  OAI21_X1 U3863 ( .B1(n5204), .B2(n6101), .A(n2973), .ZN(U2796) );
  OR4_X1 U3864 ( .A1(n6097), .A2(n4435), .A3(n4434), .A4(n4433), .ZN(U2816) );
  OAI21_X1 U3865 ( .B1(n5213), .B2(n5732), .A(n3001), .ZN(n3000) );
  INV_X1 U3866 ( .A(n5161), .ZN(n3001) );
  OAI21_X1 U3867 ( .B1(n5537), .B2(n5732), .A(n4407), .ZN(n4408) );
  OAI21_X1 U3868 ( .B1(n5204), .B2(n5873), .A(n4298), .ZN(n4299) );
  AND2_X1 U3869 ( .A1(n4397), .A2(n4396), .ZN(n4398) );
  AND4_X1 U3870 ( .A1(n4881), .A2(n4749), .A3(n4891), .A4(n5029), .ZN(n2957)
         );
  NOR2_X1 U3871 ( .A1(n4429), .A2(n4430), .ZN(n4428) );
  NOR2_X1 U3872 ( .A1(n3101), .A2(n2967), .ZN(n4402) );
  NOR2_X1 U3873 ( .A1(n5329), .A2(n2978), .ZN(n5232) );
  AND2_X1 U3874 ( .A1(n3066), .A2(n3064), .ZN(n2958) );
  NAND2_X1 U3875 ( .A1(n3539), .A2(n3120), .ZN(n4429) );
  AND2_X1 U3876 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n2959) );
  AND2_X1 U3877 ( .A1(n3039), .A2(n2988), .ZN(n2960) );
  OR2_X1 U3878 ( .A1(n2967), .A2(n3100), .ZN(n2961) );
  AND2_X1 U3879 ( .A1(n3006), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n2962)
         );
  INV_X1 U3880 ( .A(n3388), .ZN(n2999) );
  AND2_X2 U3881 ( .A1(n3358), .A2(n3238), .ZN(n3303) );
  NOR2_X1 U3882 ( .A1(n3101), .A2(n2961), .ZN(n4401) );
  AND2_X1 U3883 ( .A1(n3038), .A2(n3072), .ZN(n2963) );
  AND2_X2 U3884 ( .A1(n3129), .A2(n4522), .ZN(n3314) );
  NAND2_X1 U3885 ( .A1(n5232), .A2(n5233), .ZN(n5222) );
  NAND2_X1 U3886 ( .A1(n5509), .A2(n3590), .ZN(n5340) );
  INV_X1 U3887 ( .A(n3250), .ZN(n4225) );
  AND4_X1 U3888 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n2964)
         );
  AND2_X1 U3889 ( .A1(n3115), .A2(n3093), .ZN(n2965) );
  AND4_X1 U3890 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n2966)
         );
  OR2_X1 U3891 ( .A1(n3748), .A2(n3102), .ZN(n2967) );
  OR2_X1 U3892 ( .A1(n2961), .A2(n3099), .ZN(n2968) );
  OAI211_X1 U3893 ( .C1(n4551), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n3050), 
        .B(n3048), .ZN(n3995) );
  INV_X1 U3894 ( .A(n5313), .ZN(n3101) );
  NAND2_X1 U3895 ( .A1(n3094), .A2(n3115), .ZN(n5627) );
  NOR2_X1 U3896 ( .A1(n4386), .A2(n5625), .ZN(n5618) );
  NAND2_X1 U3897 ( .A1(n5714), .A2(n4208), .ZN(n5704) );
  NOR2_X1 U3898 ( .A1(n3025), .A2(n4252), .ZN(n3978) );
  OR2_X1 U3899 ( .A1(n2968), .A2(n3679), .ZN(n2969) );
  OR2_X1 U3900 ( .A1(n3806), .A2(n5604), .ZN(n2970) );
  OR2_X1 U3901 ( .A1(n5680), .A2(n3034), .ZN(n2971) );
  INV_X1 U3902 ( .A(n3242), .ZN(n3026) );
  AND2_X1 U3903 ( .A1(n3094), .A2(n2965), .ZN(n4386) );
  NAND2_X1 U3904 ( .A1(n3244), .A2(n4230), .ZN(n3977) );
  NAND2_X1 U3905 ( .A1(n5716), .A2(n5715), .ZN(n5714) );
  AND2_X1 U3906 ( .A1(n3590), .A2(n3578), .ZN(n5508) );
  NOR2_X1 U3907 ( .A1(n4702), .A2(n4639), .ZN(n4703) );
  AND3_X1 U3908 ( .A1(n3005), .A2(n2957), .A3(n4703), .ZN(n3539) );
  AND2_X1 U3909 ( .A1(n4565), .A2(n3388), .ZN(n2972) );
  AND2_X1 U3910 ( .A1(n4119), .A2(n4118), .ZN(n2973) );
  AND2_X1 U3911 ( .A1(n3464), .A2(n3500), .ZN(n2974) );
  INV_X1 U3912 ( .A(n4215), .ZN(n3095) );
  AND2_X1 U3913 ( .A1(n4023), .A2(n4981), .ZN(n2975) );
  NAND2_X1 U3914 ( .A1(n5705), .A2(n3076), .ZN(n2976) );
  NAND2_X1 U3915 ( .A1(n3103), .A2(n3120), .ZN(n2977) );
  INV_X1 U3916 ( .A(n4217), .ZN(n4218) );
  NAND2_X1 U3917 ( .A1(n5689), .A2(n4216), .ZN(n4217) );
  INV_X1 U3918 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5726) );
  OR2_X1 U3919 ( .A1(n2969), .A2(n5244), .ZN(n2978) );
  NOR2_X1 U3920 ( .A1(n4210), .A2(n5688), .ZN(n2979) );
  NOR2_X1 U3921 ( .A1(n5686), .A2(n5786), .ZN(n2980) );
  INV_X1 U3922 ( .A(n3011), .ZN(n3732) );
  NOR2_X1 U3923 ( .A1(n3730), .A2(n3729), .ZN(n3011) );
  NAND2_X1 U3924 ( .A1(n5226), .A2(n5227), .ZN(n5146) );
  INV_X1 U3925 ( .A(n6189), .ZN(n3014) );
  OR2_X1 U3926 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n2981)
         );
  AND2_X1 U3927 ( .A1(n3045), .A2(n3043), .ZN(n2982) );
  AND2_X1 U3928 ( .A1(n5662), .A2(n3039), .ZN(n2983) );
  NAND2_X1 U3929 ( .A1(n4721), .A2(n4141), .ZN(n4254) );
  INV_X1 U3930 ( .A(n4254), .ZN(n3098) );
  AND2_X1 U3931 ( .A1(n4308), .A2(n3105), .ZN(n2984) );
  NOR2_X1 U3932 ( .A1(n4218), .A2(n4215), .ZN(n3092) );
  AND2_X1 U3933 ( .A1(n2959), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n2985)
         );
  OR2_X1 U3934 ( .A1(n4205), .A2(n4204), .ZN(n2986) );
  INV_X1 U3935 ( .A(n4191), .ZN(n3071) );
  OR2_X1 U3936 ( .A1(n4190), .A2(n6268), .ZN(n4191) );
  OR2_X1 U3937 ( .A1(n4207), .A2(n6252), .ZN(n4208) );
  AND2_X1 U3938 ( .A1(n3540), .A2(n3006), .ZN(n2987) );
  NOR2_X1 U3939 ( .A1(n5404), .A2(n5403), .ZN(n5402) );
  NOR2_X1 U3940 ( .A1(n3052), .A2(n4705), .ZN(n4985) );
  INV_X2 U3941 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5034) );
  NOR2_X1 U3942 ( .A1(n4705), .A2(n3055), .ZN(n4884) );
  AND2_X1 U3943 ( .A1(n3926), .A2(n4235), .ZN(n4201) );
  INV_X1 U3944 ( .A(n5158), .ZN(n3106) );
  AND2_X1 U3945 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n2988)
         );
  NAND2_X1 U3946 ( .A1(n5071), .A2(n5070), .ZN(n5069) );
  AND2_X1 U3947 ( .A1(n5359), .A2(n5375), .ZN(n2989) );
  OR3_X1 U3948 ( .A1(n5689), .A2(n4291), .A3(n4292), .ZN(n2990) );
  INV_X1 U3949 ( .A(n4378), .ZN(n5248) );
  NOR2_X1 U3950 ( .A1(n4377), .A2(n4379), .ZN(n4378) );
  INV_X1 U3951 ( .A(n3008), .ZN(n3571) );
  NAND2_X1 U3952 ( .A1(n3540), .A2(n2962), .ZN(n3008) );
  AND2_X1 U3953 ( .A1(n5185), .A2(n5184), .ZN(n4391) );
  AND2_X1 U3954 ( .A1(n3058), .A2(n3057), .ZN(n2991) );
  INV_X1 U3955 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3007) );
  NOR2_X1 U3956 ( .A1(n4705), .A2(n4752), .ZN(n4751) );
  XNOR2_X1 U3957 ( .A(n3995), .B(n4552), .ZN(n4566) );
  INV_X1 U3958 ( .A(n5388), .ZN(n3064) );
  NAND2_X1 U3959 ( .A1(n3477), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n2992)
         );
  AND2_X1 U3960 ( .A1(n3061), .A2(n3060), .ZN(n2993) );
  OAI33_X1 U3961 ( .A1(n6347), .A2(n6346), .A3(n6593), .B1(n6345), .B2(n6387), 
        .B3(n6344), .ZN(n2994) );
  XNOR2_X1 U3962 ( .A(n6390), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6345)
         );
  AND2_X1 U3963 ( .A1(n3394), .A2(n4744), .ZN(n6344) );
  INV_X4 U3964 ( .A(n2998), .ZN(n5689) );
  NAND2_X1 U3965 ( .A1(n2998), .A2(n2986), .ZN(n4206) );
  NAND2_X2 U3966 ( .A1(n4200), .A2(n4203), .ZN(n2998) );
  OR2_X2 U3967 ( .A1(n5670), .A2(n5672), .ZN(n3096) );
  NAND2_X2 U3968 ( .A1(n3027), .A2(n3028), .ZN(n5670) );
  NAND2_X1 U3969 ( .A1(n4564), .A2(n4565), .ZN(n4563) );
  INV_X1 U3970 ( .A(n3000), .ZN(n5162) );
  INV_X1 U3971 ( .A(n5157), .ZN(n3003) );
  NAND3_X1 U3972 ( .A1(n3005), .A2(n2957), .A3(n3004), .ZN(n3577) );
  INV_X1 U3973 ( .A(n3539), .ZN(n4894) );
  AND2_X1 U3974 ( .A1(n4978), .A2(n3524), .ZN(n3005) );
  OR2_X1 U3975 ( .A1(n5329), .A2(n2969), .ZN(n5243) );
  NOR2_X1 U3976 ( .A1(n5329), .A2(n3679), .ZN(n5313) );
  INV_X1 U3977 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U3978 ( .A1(n3015), .A2(n4140), .ZN(n4570) );
  XNOR2_X1 U3979 ( .A(n3016), .B(n3377), .ZN(n4136) );
  NAND2_X1 U3980 ( .A1(n6206), .A2(n3017), .ZN(n3019) );
  NAND2_X2 U3981 ( .A1(n6204), .A2(n6203), .ZN(n6206) );
  NAND2_X1 U3982 ( .A1(n3021), .A2(n4191), .ZN(n3070) );
  NAND3_X1 U3983 ( .A1(n4248), .A2(n2953), .A3(n3022), .ZN(n3252) );
  NAND2_X1 U3984 ( .A1(n3244), .A2(n3023), .ZN(n3022) );
  NAND4_X1 U3985 ( .A1(n3247), .A2(n3227), .A3(n3024), .A4(n3248), .ZN(n4124)
         );
  OR2_X2 U3986 ( .A1(n3035), .A2(n5680), .ZN(n3027) );
  INV_X1 U3987 ( .A(n3032), .ZN(n3028) );
  OR2_X1 U3988 ( .A1(n3072), .A2(n3034), .ZN(n3033) );
  OAI21_X1 U3989 ( .B1(n2971), .B2(n3072), .A(n3029), .ZN(n3032) );
  INV_X1 U3990 ( .A(n3030), .ZN(n3029) );
  OAI22_X1 U3991 ( .A1(n5680), .A2(n2979), .B1(n5689), .B2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3030) );
  AND2_X1 U3992 ( .A1(n3035), .A2(n3031), .ZN(n5679) );
  AND2_X1 U3993 ( .A1(n3033), .A2(n2979), .ZN(n3031) );
  NAND3_X1 U3994 ( .A1(n3037), .A2(n4211), .A3(n3036), .ZN(n3035) );
  INV_X1 U3995 ( .A(n5716), .ZN(n3037) );
  NAND2_X1 U3996 ( .A1(n5670), .A2(n3092), .ZN(n3042) );
  NAND2_X1 U3998 ( .A1(n2975), .A2(n3054), .ZN(n3052) );
  NAND2_X1 U3999 ( .A1(n3056), .A2(n4885), .ZN(n3055) );
  NAND2_X1 U4000 ( .A1(n5226), .A2(n3061), .ZN(n4345) );
  NOR2_X2 U4001 ( .A1(n5404), .A2(n3063), .ZN(n5361) );
  INV_X2 U4002 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3068) );
  NAND2_X1 U4003 ( .A1(n3230), .A2(n4265), .ZN(n4263) );
  NAND3_X1 U4004 ( .A1(n3225), .A2(n4416), .A3(n3226), .ZN(n4229) );
  OR2_X2 U4006 ( .A1(n3071), .A2(n6196), .ZN(n3069) );
  INV_X1 U4007 ( .A(n5707), .ZN(n3073) );
  NAND2_X1 U4008 ( .A1(n3437), .A2(n3079), .ZN(n3078) );
  OAI211_X1 U4009 ( .C1(n3437), .C2(n3087), .A(n3086), .B(n3081), .ZN(n4176)
         );
  NAND2_X1 U4010 ( .A1(n3437), .A2(n3085), .ZN(n3081) );
  INV_X1 U4011 ( .A(n3086), .ZN(n3083) );
  NAND2_X1 U4012 ( .A1(n3096), .A2(n3095), .ZN(n3094) );
  NAND3_X1 U4013 ( .A1(n2957), .A2(n4703), .A3(n4978), .ZN(n4895) );
  NAND2_X1 U4014 ( .A1(n3507), .A2(n3506), .ZN(n4978) );
  OAI21_X1 U4016 ( .B1(n3266), .B2(n4263), .A(n4235), .ZN(n3274) );
  NAND2_X1 U4017 ( .A1(n3465), .A2(n3464), .ZN(n3498) );
  NAND2_X1 U4018 ( .A1(n5313), .A2(n5314), .ZN(n5174) );
  NAND2_X1 U4019 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  AND2_X1 U4020 ( .A1(n5157), .A2(n3105), .ZN(n4310) );
  NAND2_X1 U4021 ( .A1(n5157), .A2(n2984), .ZN(n3107) );
  NAND2_X1 U4022 ( .A1(n5157), .A2(n5158), .ZN(n4120) );
  NAND2_X1 U4023 ( .A1(n3371), .A2(n3370), .ZN(n4145) );
  INV_X1 U4024 ( .A(n5126), .ZN(n5129) );
  NAND2_X1 U4025 ( .A1(n5126), .A2(n5521), .ZN(n4422) );
  OAI21_X2 U4026 ( .B1(n5568), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4306), 
        .ZN(n4307) );
  INV_X1 U4027 ( .A(n6213), .ZN(n4156) );
  OAI21_X1 U4028 ( .B1(n4303), .B2(n4221), .A(n4220), .ZN(n4222) );
  INV_X1 U4029 ( .A(n3461), .ZN(n3465) );
  NOR2_X1 U4030 ( .A1(n5609), .A2(n5170), .ZN(n5173) );
  NAND2_X1 U4031 ( .A1(n5609), .A2(n4371), .ZN(n4374) );
  INV_X1 U4032 ( .A(n5521), .ZN(n5516) );
  INV_X1 U4033 ( .A(n5499), .ZN(n5521) );
  INV_X1 U4034 ( .A(READY_N), .ZN(n6591) );
  INV_X1 U4035 ( .A(n5873), .ZN(n6289) );
  OR2_X1 U4036 ( .A1(n4364), .A2(n6568), .ZN(n3108) );
  AND4_X1 U4037 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3109)
         );
  OR2_X1 U4038 ( .A1(n5172), .A2(n5171), .ZN(n3110) );
  OR2_X1 U4039 ( .A1(n5175), .A2(n5288), .ZN(n3112) );
  NAND3_X1 U4040 ( .A1(n4373), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n4372), .ZN(n3113) );
  INV_X1 U4041 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4449) );
  AND4_X1 U4042 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3114)
         );
  INV_X1 U4043 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4155) );
  AND2_X1 U4044 ( .A1(n4322), .A2(n4214), .ZN(n3115) );
  AND4_X1 U4045 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3116)
         );
  INV_X1 U4046 ( .A(n3573), .ZN(n3692) );
  NAND2_X1 U4047 ( .A1(n4447), .A2(n6442), .ZN(n5732) );
  INV_X2 U4048 ( .A(n5732), .ZN(n6217) );
  INV_X1 U4049 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6540) );
  AND2_X1 U4050 ( .A1(n4135), .A2(n4134), .ZN(n3117) );
  NAND2_X1 U4051 ( .A1(n4449), .A2(STATE_REG_1__SCAN_IN), .ZN(n6606) );
  OR2_X1 U4052 ( .A1(n4179), .A2(n6600), .ZN(n3118) );
  AND2_X1 U4053 ( .A1(n4429), .A2(n4430), .ZN(n3119) );
  NAND3_X1 U4054 ( .A1(n3538), .A2(n3537), .A3(n3536), .ZN(n3120) );
  AND2_X1 U4055 ( .A1(n4022), .A2(n4021), .ZN(n4979) );
  OR2_X1 U4056 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3121)
         );
  NOR2_X1 U4057 ( .A1(n5141), .A2(n2990), .ZN(n4305) );
  AND2_X1 U4058 ( .A1(n3237), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3238) );
  OR2_X1 U4059 ( .A1(n3434), .A2(n3433), .ZN(n4183) );
  OR2_X1 U4060 ( .A1(n3448), .A2(n3447), .ZN(n4182) );
  INV_X1 U4061 ( .A(n4735), .ZN(n3358) );
  AND2_X1 U4062 ( .A1(n3231), .A2(n3226), .ZN(n3243) );
  OR2_X1 U4063 ( .A1(n3786), .A2(n3785), .ZN(n3802) );
  AND4_X1 U4064 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3191)
         );
  INV_X1 U4065 ( .A(n4142), .ZN(n3361) );
  INV_X1 U4067 ( .A(n4896), .ZN(n3524) );
  AND2_X1 U4068 ( .A1(n3556), .A2(n3555), .ZN(n4430) );
  OR2_X1 U4069 ( .A1(n4089), .A2(n4085), .ZN(n4086) );
  INV_X1 U4070 ( .A(n4706), .ZN(n4004) );
  OAI211_X1 U4071 ( .C1(n4230), .C2(n3361), .A(n3360), .B(n3359), .ZN(n3369)
         );
  NAND2_X1 U4072 ( .A1(n4412), .A2(n4251), .ZN(n4513) );
  INV_X1 U4073 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5332) );
  INV_X1 U4074 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5391) );
  AND2_X1 U4075 ( .A1(n4058), .A2(n4057), .ZN(n5289) );
  OR3_X1 U4076 ( .A1(n4554), .A2(n4281), .A3(n4284), .ZN(n4282) );
  INV_X1 U4077 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4671) );
  XNOR2_X1 U4078 ( .A(n4487), .B(n4937), .ZN(n4580) );
  INV_X1 U4079 ( .A(n6387), .ZN(n5988) );
  INV_X1 U4080 ( .A(n5896), .ZN(n6394) );
  INV_X1 U4081 ( .A(n5445), .ZN(n4467) );
  OR2_X1 U4082 ( .A1(n5380), .A2(n4103), .ZN(n5237) );
  NAND2_X1 U4083 ( .A1(n6045), .A2(n4105), .ZN(n5380) );
  INV_X1 U4084 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4114) );
  OR3_X1 U4085 ( .A1(n6597), .A2(n6194), .A3(n3988), .ZN(n5441) );
  INV_X1 U4086 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5573) );
  NOR2_X2 U4087 ( .A1(n3026), .A2(n5034), .ZN(n3652) );
  INV_X1 U4088 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5415) );
  INV_X1 U4089 ( .A(n4881), .ZN(n4883) );
  NAND2_X1 U4090 ( .A1(n5577), .A2(n4304), .ZN(n5568) );
  OR2_X1 U4091 ( .A1(n5765), .A2(n4291), .ZN(n5149) );
  AND2_X1 U4092 ( .A1(n4049), .A2(n4048), .ZN(n5316) );
  INV_X1 U4093 ( .A(n4425), .ZN(n4030) );
  OR2_X1 U4094 ( .A1(n4276), .A2(n4662), .ZN(n5840) );
  NAND2_X1 U4095 ( .A1(n5884), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6443) );
  NOR2_X1 U4096 ( .A1(n5941), .A2(n6347), .ZN(n5910) );
  AND2_X1 U4097 ( .A1(n5039), .A2(n4989), .ZN(n6400) );
  INV_X1 U4098 ( .A(n4777), .ZN(n4936) );
  OR2_X1 U4099 ( .A1(n4743), .A2(n3990), .ZN(n6458) );
  OR2_X1 U4100 ( .A1(n4460), .A2(n4772), .ZN(n4466) );
  INV_X1 U4101 ( .A(n4312), .ZN(n6596) );
  INV_X1 U4102 ( .A(n5393), .ZN(n6093) );
  NAND2_X1 U4103 ( .A1(n5441), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4354) );
  INV_X1 U4104 ( .A(n4416), .ZN(n5164) );
  NOR2_X1 U4105 ( .A1(n5385), .A2(n5341), .ZN(n5371) );
  OR2_X1 U4106 ( .A1(n5554), .A2(n5555), .ZN(n5565) );
  NOR2_X1 U4107 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4614), .ZN(n4636) );
  INV_X1 U4108 ( .A(n6129), .ZN(n4561) );
  AND2_X1 U4109 ( .A1(n4662), .A2(n4698), .ZN(n4493) );
  OR2_X1 U4110 ( .A1(n4000), .A2(n4130), .ZN(n4245) );
  INV_X1 U4111 ( .A(n6184), .ZN(n6607) );
  OAI21_X1 U4112 ( .B1(n4499), .B2(n6591), .A(n4498), .ZN(n6179) );
  OR2_X1 U4113 ( .A1(n4242), .A2(n4264), .ZN(n4689) );
  OR2_X1 U4114 ( .A1(n5492), .A2(n5873), .ZN(n4397) );
  INV_X1 U4115 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6297) );
  OAI211_X1 U4116 ( .C1(n5908), .C2(n5910), .A(n6352), .B(n5907), .ZN(n5932)
         );
  OAI211_X1 U4117 ( .C1(n6442), .C2(n5906), .A(n4908), .B(n4944), .ZN(n4932)
         );
  OAI211_X1 U4118 ( .C1(n5086), .C2(n5089), .A(n6399), .B(n6387), .ZN(n5111)
         );
  NOR2_X2 U4119 ( .A1(n6307), .A2(n5979), .ZN(n6339) );
  OAI211_X1 U4120 ( .C1(n6354), .C2(n6353), .A(n6352), .B(n6351), .ZN(n6380)
         );
  OAI21_X1 U4121 ( .B1(n6354), .B2(n4947), .A(n4946), .ZN(n4970) );
  INV_X1 U4122 ( .A(n6402), .ZN(n6433) );
  AND2_X1 U4123 ( .A1(n4899), .A2(n3415), .ZN(n4777) );
  OAI211_X1 U4124 ( .C1(n6391), .C2(n6442), .A(n4781), .B(n4944), .ZN(n4805)
         );
  NOR2_X1 U4125 ( .A1(n4936), .A2(n6304), .ZN(n5975) );
  OAI211_X1 U4126 ( .C1(n6442), .C2(n5943), .A(n4854), .B(n4944), .ZN(n4877)
         );
  INV_X1 U4127 ( .A(n6471), .ZN(n6411) );
  OAI21_X1 U4128 ( .B1(n5990), .B2(n6447), .A(n5989), .ZN(n6021) );
  NOR2_X1 U4129 ( .A1(n5033), .A2(n6158), .ZN(n6468) );
  NOR2_X1 U4130 ( .A1(n5033), .A2(n6610), .ZN(n6506) );
  INV_X1 U4131 ( .A(n4995), .ZN(n5024) );
  INV_X1 U4132 ( .A(n5068), .ZN(n4843) );
  OAI211_X1 U4133 ( .C1(n6442), .C2(n4991), .A(n4812), .B(n4944), .ZN(n4839)
         );
  INV_X1 U4134 ( .A(n5038), .ZN(n5065) );
  INV_X1 U4135 ( .A(n6466), .ZN(n6361) );
  INV_X1 U4136 ( .A(n6499), .ZN(n6373) );
  AND2_X1 U4137 ( .A1(n3976), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6517) );
  INV_X1 U4138 ( .A(n6569), .ZN(n6570) );
  NAND2_X1 U4139 ( .A1(n4464), .A2(n4466), .ZN(n6597) );
  INV_X1 U4140 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6028) );
  INV_X1 U4141 ( .A(n6084), .ZN(n6097) );
  NAND2_X1 U4142 ( .A1(n5517), .A2(n4416), .ZN(n5499) );
  INV_X1 U4143 ( .A(n5565), .ZN(n5562) );
  OR2_X1 U4144 ( .A1(n4561), .A2(n6592), .ZN(n4560) );
  OR3_X1 U4145 ( .A1(n4500), .A2(n4493), .A3(n4492), .ZN(n6129) );
  INV_X1 U4146 ( .A(DATAI_0_), .ZN(n6154) );
  INV_X1 U4147 ( .A(DATAI_1_), .ZN(n6156) );
  INV_X1 U4148 ( .A(n6179), .ZN(n6130) );
  OR2_X1 U4149 ( .A1(n4500), .A2(n4698), .ZN(n6184) );
  INV_X1 U4150 ( .A(n4408), .ZN(n4409) );
  OAI21_X1 U4151 ( .B1(n5374), .B2(n5373), .A(n5372), .ZN(n5669) );
  NAND2_X1 U4152 ( .A1(n5727), .A2(n4546), .ZN(n6223) );
  OR2_X1 U4153 ( .A1(n4276), .A2(n4250), .ZN(n5873) );
  INV_X1 U4154 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6259) );
  OR2_X1 U4155 ( .A1(n4276), .A2(n4246), .ZN(n5882) );
  OR2_X1 U4156 ( .A1(n4618), .A2(n4990), .ZN(n6302) );
  INV_X1 U4157 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U4158 ( .A1(n4907), .A2(n4903), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5906), .ZN(n4935) );
  INV_X1 U4159 ( .A(n5084), .ZN(n5117) );
  OR2_X1 U4160 ( .A1(n6307), .A2(n6304), .ZN(n6383) );
  AOI22_X1 U4161 ( .A1(n4940), .A2(n4947), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6348), .ZN(n4973) );
  NAND2_X1 U4162 ( .A1(n4777), .A2(n4776), .ZN(n6438) );
  AOI22_X1 U4163 ( .A1(n4780), .A2(n4775), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6391), .ZN(n4808) );
  NAND2_X1 U4164 ( .A1(n6217), .A2(DATAI_21_), .ZN(n6487) );
  AOI22_X1 U4165 ( .A1(n4853), .A2(n4848), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5943), .ZN(n4880) );
  INV_X1 U4166 ( .A(n6461), .ZN(n5997) );
  INV_X1 U4167 ( .A(n6496), .ZN(n6017) );
  NAND2_X1 U4168 ( .A1(n6217), .A2(DATAI_19_), .ZN(n6478) );
  OR2_X1 U4169 ( .A1(n6444), .A2(n6304), .ZN(n6503) );
  OR2_X1 U4170 ( .A1(n4813), .A2(n4941), .ZN(n4995) );
  OR2_X1 U4171 ( .A1(n4813), .A2(n2955), .ZN(n5068) );
  NAND2_X1 U4172 ( .A1(n6217), .A2(DATAI_28_), .ZN(n6480) );
  NOR2_X1 U4173 ( .A1(n4311), .A2(n6028), .ZN(n4447) );
  INV_X1 U4174 ( .A(n6576), .ZN(n6522) );
  OR2_X1 U4175 ( .A1(n4098), .A2(STATE_REG_0__SCAN_IN), .ZN(n4492) );
  INV_X1 U4176 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6749) );
  INV_X1 U4177 ( .A(n6606), .ZN(n6546) );
  NAND2_X1 U4178 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6546), .ZN(n6569) );
  NAND2_X1 U4179 ( .A1(n4422), .A2(n4421), .ZN(U2829) );
  NAND2_X1 U4180 ( .A1(n4301), .A2(n4300), .ZN(U2987) );
  OAI21_X1 U4181 ( .B1(n5608), .B2(n5882), .A(n4385), .ZN(U2994) );
  INV_X1 U4182 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3122) );
  AND2_X2 U4183 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3122), .ZN(n3129)
         );
  AND2_X2 U4184 ( .A1(n3129), .A2(n4510), .ZN(n3326) );
  AOI22_X1 U4185 ( .A1(n3891), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3128) );
  INV_X1 U4186 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3123) );
  AND2_X2 U4187 ( .A1(n3123), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4522)
         );
  NOR2_X4 U4188 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4509) );
  AND2_X2 U4189 ( .A1(n3129), .A2(n4509), .ZN(n3341) );
  INV_X1 U4190 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3124) );
  AND2_X4 U4191 ( .A1(n3124), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4507)
         );
  AND2_X4 U4192 ( .A1(n4507), .A2(n3129), .ZN(n3889) );
  AND2_X2 U4193 ( .A1(n4522), .A2(n4579), .ZN(n3287) );
  AOI22_X1 U4194 ( .A1(n3889), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3126) );
  AND2_X2 U4195 ( .A1(n4582), .A2(n4509), .ZN(n3438) );
  AND2_X2 U4196 ( .A1(n4507), .A2(n4582), .ZN(n3342) );
  NOR2_X4 U4197 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4587) );
  AND2_X2 U4198 ( .A1(n4587), .A2(n4510), .ZN(n3293) );
  AOI22_X1 U4199 ( .A1(n3293), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3131) );
  AND2_X2 U4200 ( .A1(n4522), .A2(n4587), .ZN(n3349) );
  NAND2_X2 U4201 ( .A1(n3135), .A2(n3134), .ZN(n3224) );
  INV_X2 U4202 ( .A(n3224), .ZN(n3242) );
  AOI22_X1 U4203 ( .A1(n3889), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4204 ( .A1(n3342), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4205 ( .A1(n3438), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3137) );
  NAND4_X1 U4206 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3145)
         );
  AOI22_X1 U4207 ( .A1(n3847), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3899), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4208 ( .A1(n3349), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4209 ( .A1(n3891), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2956), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3140) );
  NAND4_X1 U4210 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n3144)
         );
  OR2_X2 U4211 ( .A1(n3145), .A2(n3144), .ZN(n3926) );
  NAND2_X2 U4212 ( .A1(n3242), .A2(n3926), .ZN(n3236) );
  AOI22_X1 U4213 ( .A1(n3292), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4214 ( .A1(n3342), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4215 ( .A1(n3293), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2950), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4216 ( .A1(n3294), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        INSTQUEUE_REG_2__3__SCAN_IN), .B2(n3349), .ZN(n3146) );
  AOI22_X1 U4217 ( .A1(n3891), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4218 ( .A1(n3847), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4219 ( .A1(n3889), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4220 ( .A1(n3438), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        INSTQUEUE_REG_12__3__SCAN_IN), .B2(n3899), .ZN(n3150) );
  AOI22_X1 U4221 ( .A1(n3292), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4222 ( .A1(n3342), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4223 ( .A1(n3438), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3899), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4224 ( .A1(n3891), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2950), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4225 ( .A1(n3349), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4226 ( .A1(n3847), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4227 ( .A1(n3889), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4228 ( .A1(n3326), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4229 ( .A1(n3114), .A2(n3162), .ZN(n3221) );
  AOI22_X1 U4230 ( .A1(n3847), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4231 ( .A1(n3891), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4232 ( .A1(n3889), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4233 ( .A1(n3438), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3899), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3163) );
  NAND4_X1 U4234 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3172)
         );
  AOI22_X1 U4235 ( .A1(n3342), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4236 ( .A1(n3292), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4237 ( .A1(n3293), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n2950), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4238 ( .A1(n3349), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U4239 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3171)
         );
  NAND3_X1 U4240 ( .A1(n3271), .A2(n4721), .A3(n4416), .ZN(n3223) );
  NAND2_X1 U4241 ( .A1(n3847), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3176)
         );
  NAND2_X1 U4242 ( .A1(n3341), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U4243 ( .A1(n3287), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3174)
         );
  NAND2_X1 U4244 ( .A1(n3889), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U4245 ( .A1(n3292), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U4246 ( .A1(n3314), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4247 ( .A1(n3342), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U4248 ( .A1(n2952), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3177)
         );
  NAND2_X1 U4249 ( .A1(n3438), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4250 ( .A1(n3326), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4251 ( .A1(n3891), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3182)
         );
  NAND2_X1 U4252 ( .A1(n3899), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3181)
         );
  NAND2_X1 U4253 ( .A1(n3349), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4254 ( .A1(n3294), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3187) );
  NAND2_X1 U4255 ( .A1(n3293), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4256 ( .A1(n2950), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3185)
         );
  MUX2_X1 U4257 ( .A(n3226), .B(n3926), .S(n3224), .Z(n3246) );
  AOI22_X1 U4258 ( .A1(n3891), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4259 ( .A1(n3847), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4260 ( .A1(n3889), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4261 ( .A1(n3438), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3899), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4262 ( .A1(n3342), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4263 ( .A1(n3292), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4264 ( .A1(n3293), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n2950), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4265 ( .A1(n3349), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4266 ( .A1(n3891), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3204)
         );
  NAND2_X1 U4267 ( .A1(n3342), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4268 ( .A1(n2952), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3202)
         );
  NAND2_X1 U4269 ( .A1(n3294), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4270 ( .A1(n3889), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4271 ( .A1(n3847), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4272 ( .A1(n3438), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4273 ( .A1(n3287), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4274 ( .A1(n3292), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4275 ( .A1(n3314), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4276 ( .A1(n3349), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4277 ( .A1(n2950), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3209)
         );
  NAND2_X1 U4278 ( .A1(n3341), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4279 ( .A1(n3326), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4280 ( .A1(n3899), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3214)
         );
  NAND2_X1 U4281 ( .A1(n3293), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3213) );
  AND4_X4 U4282 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n4735)
         );
  NAND2_X1 U4283 ( .A1(n3926), .A2(n3226), .ZN(n3249) );
  INV_X1 U4284 ( .A(n3249), .ZN(n3227) );
  NAND4_X1 U4285 ( .A1(n3271), .A2(n3227), .A3(n3250), .A4(n3221), .ZN(n3222)
         );
  OAI211_X1 U4286 ( .C1(n3223), .C2(n3246), .A(n4251), .B(n3222), .ZN(n3229)
         );
  NAND2_X1 U4287 ( .A1(n3231), .A2(n3224), .ZN(n3225) );
  AOI22_X1 U4288 ( .A1(n4229), .A2(n4499), .B1(n3227), .B2(n3991), .ZN(n3228)
         );
  NAND2_X1 U4289 ( .A1(n3229), .A2(n3228), .ZN(n3264) );
  INV_X1 U4290 ( .A(n3264), .ZN(n3235) );
  NAND2_X1 U4291 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4441) );
  OAI21_X1 U4292 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n4441), .ZN(n4098) );
  NAND2_X1 U4293 ( .A1(n3990), .A2(n4098), .ZN(n3245) );
  NAND2_X1 U4294 ( .A1(n3245), .A2(n3231), .ZN(n3233) );
  NAND2_X1 U4295 ( .A1(n3235), .A2(n3234), .ZN(n3256) );
  NAND2_X1 U4296 ( .A1(n3256), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4297 ( .A1(n3236), .A2(n3303), .ZN(n3259) );
  NAND2_X1 U4298 ( .A1(n3239), .A2(n3259), .ZN(n3283) );
  NAND2_X1 U4299 ( .A1(n3283), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4300 ( .A1(n6596), .A2(n6345), .ZN(n3241) );
  INV_X1 U4301 ( .A(n3976), .ZN(n4125) );
  NAND2_X1 U4302 ( .A1(n4125), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3240) );
  AND2_X1 U4303 ( .A1(n3242), .A2(n4416), .ZN(n3270) );
  NAND3_X1 U4304 ( .A1(n3243), .A2(n3098), .A3(n3270), .ZN(n4130) );
  INV_X1 U4305 ( .A(n4130), .ZN(n3244) );
  NAND2_X1 U4306 ( .A1(n3246), .A2(n4721), .ZN(n3248) );
  AND2_X1 U4307 ( .A1(n3271), .A2(n4416), .ZN(n3247) );
  INV_X1 U4308 ( .A(n4141), .ZN(n4725) );
  INV_X1 U4309 ( .A(n4513), .ZN(n3251) );
  NAND2_X1 U4310 ( .A1(n3251), .A2(n3250), .ZN(n4248) );
  NAND2_X1 U4311 ( .A1(n3252), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3281) );
  MUX2_X1 U4312 ( .A(n3976), .B(n4312), .S(n6390), .Z(n3258) );
  INV_X1 U4313 ( .A(n3258), .ZN(n3254) );
  NAND2_X1 U4314 ( .A1(n3256), .A2(n3255), .ZN(n3263) );
  INV_X1 U4315 ( .A(n3257), .ZN(n3261) );
  AND2_X1 U4316 ( .A1(n3259), .A2(n3258), .ZN(n3260) );
  NAND2_X1 U4317 ( .A1(n3236), .A2(n4247), .ZN(n3265) );
  NAND2_X1 U4318 ( .A1(n3265), .A2(n4141), .ZN(n3266) );
  INV_X1 U4319 ( .A(n5191), .ZN(n6514) );
  NOR2_X1 U4320 ( .A1(n6514), .A2(n6513), .ZN(n3267) );
  OAI211_X1 U4321 ( .C1(n4721), .C2(n4735), .A(n5445), .B(n3267), .ZN(n3268)
         );
  INV_X1 U4322 ( .A(n3268), .ZN(n3273) );
  NOR2_X1 U4323 ( .A1(n4141), .A2(n3221), .ZN(n3269) );
  NAND4_X1 U4324 ( .A1(n3270), .A2(n4735), .A3(n3269), .A4(n4247), .ZN(n4596)
         );
  NAND2_X1 U4325 ( .A1(n3271), .A2(n4499), .ZN(n3272) );
  NAND4_X1 U4326 ( .A1(n3274), .A2(n3273), .A3(n4596), .A4(n3272), .ZN(n3275)
         );
  INV_X1 U4327 ( .A(n3276), .ZN(n3337) );
  NAND2_X2 U4328 ( .A1(n3336), .A2(n3337), .ZN(n3339) );
  INV_X1 U4329 ( .A(n3339), .ZN(n3277) );
  NAND2_X1 U4330 ( .A1(n3307), .A2(n3277), .ZN(n3282) );
  INV_X1 U4331 ( .A(n3278), .ZN(n3279) );
  NOR2_X1 U4332 ( .A1(n3279), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3280)
         );
  OR2_X2 U4333 ( .A1(n3281), .A2(n3280), .ZN(n3308) );
  NAND2_X1 U4334 ( .A1(n3947), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6311) );
  MUX2_X1 U4335 ( .A(n6311), .B(n3947), .S(n6390), .Z(n3284) );
  NAND2_X1 U4336 ( .A1(n4671), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U4337 ( .A1(n3284), .A2(n4938), .ZN(n4996) );
  NAND2_X1 U4338 ( .A1(n4996), .A2(n6596), .ZN(n3285) );
  OAI21_X1 U4339 ( .B1(n3976), .B2(n3947), .A(n3285), .ZN(n3286) );
  NAND2_X1 U4340 ( .A1(n4525), .A2(n6513), .ZN(n3302) );
  AOI22_X1 U4341 ( .A1(n3897), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4342 ( .A1(n3776), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4343 ( .A1(n3696), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4344 ( .A1(n3871), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4345 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3300)
         );
  AOI22_X1 U4346 ( .A1(n3892), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4347 ( .A1(n3890), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4348 ( .A1(n2956), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4349 ( .A1(n3405), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4350 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  NAND2_X1 U4351 ( .A1(n4127), .A2(n4159), .ZN(n3301) );
  NAND2_X1 U4352 ( .A1(n4735), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3399) );
  INV_X1 U4353 ( .A(n3399), .ZN(n3304) );
  XNOR2_X2 U4354 ( .A(n3306), .B(n3305), .ZN(n3417) );
  NAND2_X1 U4355 ( .A1(n3308), .A2(n3307), .ZN(n3309) );
  XNOR2_X2 U4356 ( .A(n3309), .B(n3339), .ZN(n4511) );
  AOI22_X1 U4357 ( .A1(n3696), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4358 ( .A1(n3890), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4359 ( .A1(n3871), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4360 ( .A1(n4585), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3310) );
  NAND4_X1 U4361 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3320)
         );
  AOI22_X1 U4362 ( .A1(n3776), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4363 ( .A1(n3343), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4364 ( .A1(n3293), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4365 ( .A1(n3405), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3315) );
  NAND4_X1 U4366 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3319)
         );
  NAND2_X1 U4367 ( .A1(n4127), .A2(n4137), .ZN(n3321) );
  OAI21_X2 U4368 ( .B1(n4511), .B2(STATE2_REG_0__SCAN_IN), .A(n3321), .ZN(
        n3377) );
  AOI22_X1 U4369 ( .A1(n3897), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4370 ( .A1(n3890), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4371 ( .A1(n3892), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4372 ( .A1(n3776), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3322) );
  NAND4_X1 U4373 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3332)
         );
  AOI22_X1 U4374 ( .A1(n3696), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4375 ( .A1(n3871), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4377 ( .A1(n3293), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4378 ( .A1(n3558), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3327) );
  NAND4_X1 U4379 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3331)
         );
  INV_X1 U4380 ( .A(n4137), .ZN(n3333) );
  OR2_X1 U4381 ( .A1(n3333), .A2(n3399), .ZN(n3335) );
  NAND2_X1 U4382 ( .A1(n3303), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3334) );
  INV_X1 U4383 ( .A(n3336), .ZN(n3338) );
  NAND2_X1 U4384 ( .A1(n3338), .A2(n3276), .ZN(n3340) );
  NAND2_X1 U4385 ( .A1(n3340), .A2(n3339), .ZN(n3372) );
  AOI22_X1 U4386 ( .A1(n3696), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4387 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3890), .B1(n2952), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4388 ( .A1(n3871), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4389 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3558), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3345) );
  NAND4_X1 U4390 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3356)
         );
  AOI22_X1 U4391 ( .A1(n3897), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4392 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3892), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4393 ( .A1(n3776), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4394 ( .A1(n3326), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3351) );
  NAND4_X1 U4395 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3355)
         );
  XNOR2_X1 U4396 ( .A(n3361), .B(n4202), .ZN(n3357) );
  NAND2_X1 U4397 ( .A1(n3357), .A2(n4127), .ZN(n3367) );
  AOI21_X1 U4398 ( .B1(n3226), .B2(n4202), .A(n6513), .ZN(n3360) );
  NAND2_X1 U4399 ( .A1(n3303), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4400 ( .A1(n3362), .A2(n3369), .ZN(n3371) );
  NAND2_X1 U4401 ( .A1(n4127), .A2(n4202), .ZN(n3363) );
  NAND2_X1 U4402 ( .A1(n3377), .A2(n3378), .ZN(n3364) );
  INV_X1 U4403 ( .A(n3416), .ZN(n3366) );
  XNOR2_X1 U4404 ( .A(n3417), .B(n3366), .ZN(n4153) );
  AOI21_X1 U4405 ( .B1(n4153), .B2(n3652), .A(n3915), .ZN(n4638) );
  INV_X1 U4406 ( .A(n3367), .ZN(n3368) );
  AOI21_X1 U4407 ( .B1(n2955), .B2(n3242), .A(n5034), .ZN(n4544) );
  NAND2_X1 U4408 ( .A1(n3250), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3457) );
  INV_X1 U4409 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5201) );
  INV_X1 U4410 ( .A(n3652), .ZN(n3374) );
  OR2_X1 U4411 ( .A1(n3373), .A2(n3374), .ZN(n3376) );
  AOI22_X1 U4412 ( .A1(n3573), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n5034), .ZN(n3375) );
  OAI211_X1 U4413 ( .C1(n3457), .C2(n5201), .A(n3376), .B(n3375), .ZN(n4543)
         );
  MUX2_X1 U4414 ( .A(n3986), .B(n4544), .S(n4543), .Z(n4565) );
  NAND2_X1 U4415 ( .A1(n4136), .A2(n3652), .ZN(n3384) );
  AOI22_X1 U4416 ( .A1(n3573), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5034), .ZN(n3382) );
  INV_X1 U4417 ( .A(n3457), .ZN(n3380) );
  NAND2_X1 U4418 ( .A1(n3380), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3381) );
  AND2_X1 U4419 ( .A1(n3382), .A2(n3381), .ZN(n3383) );
  NAND2_X1 U4420 ( .A1(n3384), .A2(n3383), .ZN(n4564) );
  OAI21_X1 U4421 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3419), .ZN(n6222) );
  AOI22_X1 U4422 ( .A1(n3915), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3986), 
        .B2(n6222), .ZN(n3386) );
  NAND2_X1 U4423 ( .A1(n3743), .A2(EAX_REG_2__SCAN_IN), .ZN(n3385) );
  OAI211_X1 U4424 ( .C1(n3457), .C2(n3068), .A(n3386), .B(n3385), .ZN(n3388)
         );
  NAND2_X1 U4425 ( .A1(n4638), .A2(n3387), .ZN(n3389) );
  NAND2_X1 U4426 ( .A1(n4563), .A2(n2999), .ZN(n4640) );
  NAND2_X1 U4427 ( .A1(n3389), .A2(n4640), .ZN(n4639) );
  NAND2_X1 U4428 ( .A1(n3417), .A2(n3416), .ZN(n3414) );
  INV_X1 U4429 ( .A(n3390), .ZN(n3391) );
  NAND2_X1 U4430 ( .A1(n3392), .A2(n3391), .ZN(n4487) );
  NAND2_X1 U4431 ( .A1(n3393), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3397) );
  NAND2_X1 U4432 ( .A1(n6391), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U4433 ( .A1(n4802), .A2(n6312), .ZN(n3394) );
  NOR2_X1 U4434 ( .A1(n3976), .A2(n6312), .ZN(n3395) );
  AOI21_X1 U4435 ( .B1(n6344), .B2(n6596), .A(n3395), .ZN(n3396) );
  AOI22_X1 U4436 ( .A1(n3890), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4437 ( .A1(n3344), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4438 ( .A1(n4585), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4439 ( .A1(n3898), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3401) );
  NAND4_X1 U4440 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3411)
         );
  AOI22_X1 U4441 ( .A1(n3897), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4442 ( .A1(n3696), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4443 ( .A1(n3405), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4444 ( .A1(n3871), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3406) );
  NAND4_X1 U4445 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n3410)
         );
  AOI22_X1 U4446 ( .A1(n3969), .A2(n4169), .B1(n3303), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3412) );
  AOI21_X2 U4447 ( .B1(n4580), .B2(n6513), .A(n3413), .ZN(n3415) );
  NAND2_X1 U4448 ( .A1(n3414), .A2(n3415), .ZN(n3418) );
  INV_X1 U4449 ( .A(n3415), .ZN(n4709) );
  NAND3_X2 U4450 ( .A1(n3417), .A2(n4709), .A3(n3416), .ZN(n3461) );
  NAND2_X1 U4451 ( .A1(n3418), .A2(n3461), .ZN(n4165) );
  INV_X1 U4452 ( .A(n4165), .ZN(n4900) );
  INV_X1 U4453 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4584) );
  INV_X1 U4454 ( .A(n3419), .ZN(n3421) );
  INV_X1 U4455 ( .A(n3454), .ZN(n3420) );
  OAI21_X1 U4456 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3421), .A(n3420), 
        .ZN(n5450) );
  AOI22_X1 U4457 ( .A1(n3986), .A2(n5450), .B1(n3915), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4458 ( .A1(n3743), .A2(EAX_REG_3__SCAN_IN), .ZN(n3422) );
  OAI211_X1 U4459 ( .C1(n3457), .C2(n4584), .A(n3423), .B(n3422), .ZN(n3424)
         );
  AOI21_X1 U4460 ( .B1(n4900), .B2(n3652), .A(n3424), .ZN(n4702) );
  INV_X1 U4461 ( .A(n3461), .ZN(n3437) );
  AOI22_X1 U4462 ( .A1(n3696), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4463 ( .A1(n3776), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4464 ( .A1(n3344), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4465 ( .A1(n3816), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3425) );
  NAND4_X1 U4466 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3434)
         );
  AOI22_X1 U4467 ( .A1(n3890), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4468 ( .A1(n3897), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4469 ( .A1(n3871), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4470 ( .A1(n3405), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4471 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3433)
         );
  NAND2_X1 U4472 ( .A1(n3969), .A2(n4183), .ZN(n3436) );
  NAND2_X1 U4473 ( .A1(n3303), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4474 ( .A1(n3897), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4475 ( .A1(n3776), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4476 ( .A1(n3696), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3440) );
  INV_X1 U4477 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U4478 ( .A1(n3871), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3439) );
  NAND4_X1 U4479 ( .A1(n3442), .A2(n3441), .A3(n3440), .A4(n3439), .ZN(n3448)
         );
  AOI22_X1 U4480 ( .A1(n3892), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4481 ( .A1(n3890), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4482 ( .A1(n3900), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4483 ( .A1(n3405), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3443) );
  NAND4_X1 U4484 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n3447)
         );
  NAND2_X1 U4485 ( .A1(n3969), .A2(n4182), .ZN(n3450) );
  NAND2_X1 U4486 ( .A1(n3303), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U4487 ( .A1(n3450), .A2(n3449), .ZN(n3462) );
  NAND2_X1 U4488 ( .A1(n4176), .A2(n3652), .ZN(n3453) );
  NAND2_X1 U4489 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3454), .ZN(n3476)
         );
  XNOR2_X1 U4490 ( .A(n3476), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5433) );
  INV_X1 U4491 ( .A(n3915), .ZN(n3621) );
  INV_X1 U4492 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5431) );
  OAI22_X1 U4493 ( .A1(n5433), .A2(n3828), .B1(n3621), .B2(n5431), .ZN(n3451)
         );
  AOI21_X1 U4494 ( .B1(n3743), .B2(EAX_REG_5__SCAN_IN), .A(n3451), .ZN(n3452)
         );
  NAND2_X1 U4495 ( .A1(n3453), .A2(n3452), .ZN(n4881) );
  XNOR2_X1 U4496 ( .A(n3461), .B(n3463), .ZN(n4168) );
  NAND2_X1 U4497 ( .A1(n4168), .A2(n3652), .ZN(n3460) );
  OAI21_X1 U4498 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3454), .A(n3476), 
        .ZN(n6210) );
  OAI21_X1 U4499 ( .B1(n6028), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5034), 
        .ZN(n3456) );
  NAND2_X1 U4500 ( .A1(n3743), .A2(EAX_REG_4__SCAN_IN), .ZN(n3455) );
  OAI211_X1 U4501 ( .C1(n3457), .C2(n4491), .A(n3456), .B(n3455), .ZN(n3458)
         );
  OAI21_X1 U4502 ( .B1(n3828), .B2(n6210), .A(n3458), .ZN(n3459) );
  NAND2_X1 U4503 ( .A1(n3460), .A2(n3459), .ZN(n4749) );
  AOI22_X1 U4504 ( .A1(n3897), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4505 ( .A1(n3776), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4506 ( .A1(n3696), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4507 ( .A1(n3871), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4508 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3475)
         );
  AOI22_X1 U4509 ( .A1(n3892), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4510 ( .A1(n3890), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4511 ( .A1(n3900), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4512 ( .A1(n3405), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4513 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3474)
         );
  AOI22_X1 U4514 ( .A1(n3969), .A2(n4193), .B1(n3303), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U4515 ( .A1(n3498), .A2(n3499), .ZN(n4186) );
  NAND2_X1 U4516 ( .A1(n4186), .A2(n3652), .ZN(n3483) );
  INV_X1 U4517 ( .A(n3476), .ZN(n3477) );
  INV_X1 U4518 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3478) );
  NAND2_X1 U4519 ( .A1(n2992), .A2(n3478), .ZN(n3479) );
  NAND2_X1 U4520 ( .A1(n3504), .A2(n3479), .ZN(n6202) );
  INV_X1 U4521 ( .A(n6202), .ZN(n3481) );
  AOI22_X1 U4522 ( .A1(n3743), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n5034), .ZN(n3480) );
  MUX2_X1 U4523 ( .A(n3481), .B(n3480), .S(n3828), .Z(n3482) );
  NAND2_X1 U4524 ( .A1(n3483), .A2(n3482), .ZN(n4891) );
  AOI22_X1 U4525 ( .A1(n3776), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4526 ( .A1(n3344), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4527 ( .A1(n3815), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4528 ( .A1(n3900), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4529 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3493)
         );
  AOI22_X1 U4530 ( .A1(n3897), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4531 ( .A1(n3696), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4532 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3890), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4533 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3558), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4534 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3492)
         );
  OAI21_X1 U4535 ( .B1(n3493), .B2(n3492), .A(n3652), .ZN(n3497) );
  NAND2_X1 U4536 ( .A1(n3743), .A2(EAX_REG_8__SCAN_IN), .ZN(n3496) );
  XNOR2_X1 U4537 ( .A(n3508), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U4538 ( .A1(n6072), .A2(n3986), .ZN(n3495) );
  NAND2_X1 U4539 ( .A1(n3915), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3494)
         );
  NAND4_X1 U4540 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n5029)
         );
  NAND2_X1 U4541 ( .A1(n3969), .A2(n4202), .ZN(n3502) );
  NAND2_X1 U4542 ( .A1(n3303), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U4543 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  NAND2_X1 U4544 ( .A1(n4192), .A2(n3652), .ZN(n3507) );
  XNOR2_X1 U4545 ( .A(n3504), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5729) );
  OAI22_X1 U4546 ( .A1(n5729), .A2(n3828), .B1(n3621), .B2(n5726), .ZN(n3505)
         );
  AOI21_X1 U4547 ( .B1(n3743), .B2(EAX_REG_7__SCAN_IN), .A(n3505), .ZN(n3506)
         );
  XOR2_X1 U4548 ( .A(n5415), .B(n3525), .Z(n5712) );
  INV_X1 U4549 ( .A(n5712), .ZN(n3523) );
  AOI22_X1 U4550 ( .A1(n3897), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4551 ( .A1(n3890), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4552 ( .A1(n3815), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4553 ( .A1(n3816), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4554 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3518)
         );
  AOI22_X1 U4555 ( .A1(n3696), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4556 ( .A1(n3776), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4557 ( .A1(n3344), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4558 ( .A1(n3405), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4559 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3517)
         );
  OAI21_X1 U4560 ( .B1(n3518), .B2(n3517), .A(n3652), .ZN(n3521) );
  NAND2_X1 U4561 ( .A1(n3743), .A2(EAX_REG_9__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4562 ( .A1(n3915), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3519)
         );
  NAND3_X1 U4563 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3522) );
  AOI21_X1 U4564 ( .B1(n3523), .B2(n3986), .A(n3522), .ZN(n4896) );
  XNOR2_X1 U4565 ( .A(n3540), .B(n3007), .ZN(n6062) );
  OR2_X1 U4566 ( .A1(n6062), .A2(n3828), .ZN(n3538) );
  AOI22_X1 U4567 ( .A1(n3743), .A2(EAX_REG_10__SCAN_IN), .B1(n3915), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4568 ( .A1(n3871), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4569 ( .A1(n3897), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4570 ( .A1(n3892), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4571 ( .A1(n4585), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4572 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3535)
         );
  AOI22_X1 U4573 ( .A1(n3696), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4574 ( .A1(n3890), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4575 ( .A1(n3558), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4576 ( .A1(n3817), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3530) );
  NAND4_X1 U4577 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3534)
         );
  OAI21_X1 U4578 ( .B1(n3535), .B2(n3534), .A(n3652), .ZN(n3536) );
  AOI21_X1 U4579 ( .B1(n6648), .B2(n3541), .A(n2987), .ZN(n6187) );
  OR2_X1 U4580 ( .A1(n6187), .A2(n3828), .ZN(n3556) );
  AOI22_X1 U4581 ( .A1(n3897), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4582 ( .A1(n3696), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4583 ( .A1(n3344), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4584 ( .A1(n3898), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3542) );
  NAND4_X1 U4585 ( .A1(n3545), .A2(n3544), .A3(n3543), .A4(n3542), .ZN(n3551)
         );
  AOI22_X1 U4586 ( .A1(n3871), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4587 ( .A1(n3890), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4588 ( .A1(n4585), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4589 ( .A1(n3816), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3546) );
  NAND4_X1 U4590 ( .A1(n3549), .A2(n3548), .A3(n3547), .A4(n3546), .ZN(n3550)
         );
  OAI21_X1 U4591 ( .B1(n3551), .B2(n3550), .A(n3652), .ZN(n3554) );
  NAND2_X1 U4592 ( .A1(n3743), .A2(EAX_REG_11__SCAN_IN), .ZN(n3553) );
  NAND2_X1 U4593 ( .A1(n3915), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3552)
         );
  XNOR2_X1 U4594 ( .A(n2987), .B(n3009), .ZN(n5693) );
  AOI22_X1 U4595 ( .A1(n3743), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5034), .ZN(n3557) );
  MUX2_X1 U4596 ( .A(n5693), .B(n3557), .S(n3828), .Z(n3570) );
  AOI22_X1 U4597 ( .A1(n3696), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4598 ( .A1(n3344), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4599 ( .A1(n3815), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4600 ( .A1(n3776), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4601 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3568)
         );
  AOI22_X1 U4602 ( .A1(n3871), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4603 ( .A1(n3890), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4604 ( .A1(n4585), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4605 ( .A1(n3405), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4606 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3567)
         );
  OAI21_X1 U4607 ( .B1(n3568), .B2(n3567), .A(n3652), .ZN(n3569) );
  NAND2_X1 U4608 ( .A1(n3570), .A2(n3569), .ZN(n5401) );
  INV_X1 U4609 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4610 ( .A1(n3008), .A2(n3574), .ZN(n3572) );
  NAND2_X1 U4611 ( .A1(n3642), .A2(n3572), .ZN(n6055) );
  INV_X1 U4612 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5561) );
  OAI22_X1 U4613 ( .A1(n3692), .A2(n5561), .B1(n3574), .B2(n3621), .ZN(n3575)
         );
  AOI21_X1 U4614 ( .B1(n6055), .B2(n3986), .A(n3575), .ZN(n3576) );
  AOI22_X1 U4615 ( .A1(n3897), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4616 ( .A1(n3890), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4617 ( .A1(n3696), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4618 ( .A1(n3776), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4619 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3588)
         );
  AOI22_X1 U4620 ( .A1(n3344), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4621 ( .A1(n3871), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4622 ( .A1(n4585), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4623 ( .A1(n3816), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3583) );
  NAND4_X1 U4624 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3587)
         );
  OR2_X1 U4625 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  NAND2_X1 U4626 ( .A1(n5508), .A2(n5510), .ZN(n5509) );
  NAND2_X1 U4627 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3591) );
  NAND2_X1 U4628 ( .A1(n3609), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3674)
         );
  XNOR2_X1 U4629 ( .A(n3674), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5647)
         );
  NAND2_X1 U4630 ( .A1(n5647), .A2(n3986), .ZN(n3608) );
  NAND2_X1 U4631 ( .A1(n4247), .A2(n4416), .ZN(n3592) );
  AOI22_X1 U4632 ( .A1(n3897), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4633 ( .A1(n3776), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4634 ( .A1(n3696), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4635 ( .A1(n3871), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3593) );
  NAND4_X1 U4636 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3602)
         );
  AOI22_X1 U4637 ( .A1(n3892), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4638 ( .A1(n3890), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4639 ( .A1(n3900), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4640 ( .A1(n3405), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3597) );
  NAND4_X1 U4641 ( .A1(n3600), .A2(n3599), .A3(n3598), .A4(n3597), .ZN(n3601)
         );
  NOR2_X1 U4642 ( .A1(n3602), .A2(n3601), .ZN(n3606) );
  INV_X1 U4643 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3603) );
  AOI21_X1 U4644 ( .B1(n3603), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3604) );
  AOI21_X1 U4645 ( .B1(n3743), .B2(EAX_REG_17__SCAN_IN), .A(n3604), .ZN(n3605)
         );
  OAI21_X1 U4646 ( .B1(n3910), .B2(n3606), .A(n3605), .ZN(n3607) );
  NAND2_X1 U4647 ( .A1(n3608), .A2(n3607), .ZN(n5343) );
  INV_X1 U4648 ( .A(n3609), .ZN(n3610) );
  INV_X1 U4649 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U4650 ( .A(n3610), .B(n5358), .ZN(n5658) );
  NAND2_X1 U4651 ( .A1(n5658), .A2(n3986), .ZN(n3626) );
  AOI22_X1 U4652 ( .A1(n3871), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4653 ( .A1(n3890), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4654 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3776), .B1(n3900), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4655 ( .A1(n3892), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4656 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3620)
         );
  AOI22_X1 U4657 ( .A1(n3696), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4658 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3558), .B1(n3405), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4659 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4585), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4660 ( .A1(n3815), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4661 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3619)
         );
  OR2_X1 U4662 ( .A1(n3620), .A2(n3619), .ZN(n3624) );
  INV_X1 U4663 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3622) );
  OAI22_X1 U4664 ( .A1(n3692), .A2(n3622), .B1(n5358), .B2(n3621), .ZN(n3623)
         );
  AOI21_X1 U4665 ( .B1(n3884), .B2(n3624), .A(n3623), .ZN(n3625) );
  NAND2_X1 U4666 ( .A1(n3626), .A2(n3625), .ZN(n5357) );
  XNOR2_X1 U4667 ( .A(n3642), .B(n5391), .ZN(n5674) );
  NAND2_X1 U4668 ( .A1(n5674), .A2(n3986), .ZN(n3641) );
  AOI22_X1 U4669 ( .A1(n3890), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4670 ( .A1(n3696), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4671 ( .A1(n3871), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4672 ( .A1(n3558), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4673 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3636)
         );
  AOI22_X1 U4674 ( .A1(n3897), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4675 ( .A1(n3776), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4676 ( .A1(n3892), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4677 ( .A1(n3816), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3631) );
  NAND4_X1 U4678 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3635)
         );
  OAI21_X1 U4679 ( .B1(n3636), .B2(n3635), .A(n3652), .ZN(n3639) );
  NAND2_X1 U4680 ( .A1(n3743), .A2(EAX_REG_14__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4681 ( .A1(n3915), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3637)
         );
  AND3_X1 U4682 ( .A1(n3639), .A2(n3638), .A3(n3637), .ZN(n3640) );
  NAND2_X1 U4683 ( .A1(n3641), .A2(n3640), .ZN(n5386) );
  OR2_X1 U4684 ( .A1(n3642), .A2(n5391), .ZN(n3643) );
  INV_X1 U4685 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5377) );
  XNOR2_X1 U4686 ( .A(n3643), .B(n5377), .ZN(n5665) );
  NAND2_X1 U4687 ( .A1(n5665), .A2(n3986), .ZN(n3659) );
  AOI22_X1 U4688 ( .A1(n3776), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4689 ( .A1(n3890), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4690 ( .A1(n3815), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4691 ( .A1(n3405), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3644) );
  NAND4_X1 U4692 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3654)
         );
  AOI22_X1 U4693 ( .A1(n3897), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4694 ( .A1(n3696), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4695 ( .A1(n3892), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4696 ( .A1(n3900), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4697 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3653)
         );
  OAI21_X1 U4698 ( .B1(n3654), .B2(n3653), .A(n3652), .ZN(n3657) );
  NAND2_X1 U4699 ( .A1(n3743), .A2(EAX_REG_15__SCAN_IN), .ZN(n3656) );
  NAND2_X1 U4700 ( .A1(n3915), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3655)
         );
  AND3_X1 U4701 ( .A1(n3657), .A2(n3656), .A3(n3655), .ZN(n3658) );
  NAND2_X1 U4702 ( .A1(n3659), .A2(n3658), .ZN(n5373) );
  NAND3_X1 U4703 ( .A1(n5357), .A2(n5386), .A3(n5373), .ZN(n3660) );
  NOR2_X1 U4704 ( .A1(n5343), .A2(n3660), .ZN(n3661) );
  NAND2_X1 U4705 ( .A1(n5340), .A2(n3661), .ZN(n5329) );
  AOI22_X1 U4706 ( .A1(n3696), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4707 ( .A1(n3890), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4708 ( .A1(n4585), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4709 ( .A1(n3558), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4710 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4711 ( .A1(n3846), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4712 ( .A1(n3344), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4713 ( .A1(n3871), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4714 ( .A1(n3776), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4715 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NOR2_X1 U4716 ( .A1(n3671), .A2(n3670), .ZN(n3673) );
  AOI22_X1 U4717 ( .A1(n3573), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5034), .ZN(n3672) );
  OAI21_X1 U4718 ( .B1(n3910), .B2(n3673), .A(n3672), .ZN(n3678) );
  INV_X1 U4719 ( .A(n3674), .ZN(n3675) );
  NAND2_X1 U4720 ( .A1(n3676), .A2(n5332), .ZN(n3677) );
  NAND2_X1 U4721 ( .A1(n3709), .A2(n3677), .ZN(n5636) );
  MUX2_X1 U4722 ( .A(n3678), .B(n5636), .S(n3986), .Z(n5330) );
  INV_X1 U4723 ( .A(n5330), .ZN(n3679) );
  XNOR2_X1 U4724 ( .A(n3709), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5633)
         );
  AOI22_X1 U4725 ( .A1(n3897), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4726 ( .A1(n3776), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4727 ( .A1(n3696), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4728 ( .A1(n3871), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3680) );
  NAND4_X1 U4729 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3689)
         );
  AOI22_X1 U4730 ( .A1(n3892), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4731 ( .A1(n3890), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4732 ( .A1(n3900), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4733 ( .A1(n3405), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4734 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3688)
         );
  OR2_X1 U4735 ( .A1(n3689), .A2(n3688), .ZN(n3694) );
  INV_X1 U4736 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3691) );
  OAI21_X1 U4737 ( .B1(n6028), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5034), 
        .ZN(n3690) );
  OAI21_X1 U4738 ( .B1(n3692), .B2(n3691), .A(n3690), .ZN(n3693) );
  AOI21_X1 U4739 ( .B1(n3884), .B2(n3694), .A(n3693), .ZN(n3695) );
  AOI21_X1 U4740 ( .B1(n5633), .B2(n3986), .A(n3695), .ZN(n5314) );
  AOI22_X1 U4741 ( .A1(n3696), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4742 ( .A1(n3344), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4743 ( .A1(n3871), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4744 ( .A1(n3776), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4745 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3706)
         );
  AOI22_X1 U4746 ( .A1(n3890), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4747 ( .A1(n3897), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4748 ( .A1(n3405), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4749 ( .A1(n4585), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4750 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3705)
         );
  NOR2_X1 U4751 ( .A1(n3706), .A2(n3705), .ZN(n3708) );
  AOI22_X1 U4752 ( .A1(n3573), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5034), .ZN(n3707) );
  OAI21_X1 U4753 ( .B1(n3910), .B2(n3708), .A(n3707), .ZN(n3713) );
  NAND2_X1 U4754 ( .A1(n3711), .A2(n3710), .ZN(n3712) );
  NAND2_X1 U4755 ( .A1(n3773), .A2(n3712), .ZN(n5276) );
  MUX2_X1 U4756 ( .A(n3713), .B(n5276), .S(n3986), .Z(n3714) );
  INV_X1 U4757 ( .A(n3714), .ZN(n5175) );
  XNOR2_X1 U4758 ( .A(n3732), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5612)
         );
  AOI22_X1 U4759 ( .A1(n3897), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4760 ( .A1(n3892), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4761 ( .A1(n4585), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4762 ( .A1(n3816), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4763 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3724)
         );
  AOI22_X1 U4764 ( .A1(n3696), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4765 ( .A1(n3890), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4766 ( .A1(n3776), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4767 ( .A1(n3405), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4768 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3723)
         );
  OR2_X1 U4769 ( .A1(n3724), .A2(n3723), .ZN(n3727) );
  INV_X1 U4770 ( .A(EAX_REG_21__SCAN_IN), .ZN(n3725) );
  INV_X1 U4771 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5614) );
  OAI22_X1 U4772 ( .A1(n3692), .A2(n3725), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5614), .ZN(n3726) );
  AOI21_X1 U4773 ( .B1(n3884), .B2(n3727), .A(n3726), .ZN(n3728) );
  MUX2_X1 U4774 ( .A(n5612), .B(n3728), .S(n3828), .Z(n5288) );
  NAND2_X1 U4775 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  NAND2_X1 U4776 ( .A1(n3732), .A2(n3731), .ZN(n5621) );
  AOI22_X1 U4777 ( .A1(n3897), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4778 ( .A1(n3890), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4779 ( .A1(n3817), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4780 ( .A1(n3405), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4781 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3742)
         );
  AOI22_X1 U4782 ( .A1(n3696), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4783 ( .A1(n3344), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4784 ( .A1(n3776), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4785 ( .A1(n4585), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4786 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3741)
         );
  NOR2_X1 U4787 ( .A1(n3742), .A2(n3741), .ZN(n3746) );
  OAI21_X1 U4788 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6028), .A(n5034), 
        .ZN(n3745) );
  NAND2_X1 U4789 ( .A1(n3743), .A2(EAX_REG_20__SCAN_IN), .ZN(n3744) );
  OAI211_X1 U4790 ( .C1(n3910), .C2(n3746), .A(n3745), .B(n3744), .ZN(n3747)
         );
  OAI21_X1 U4791 ( .B1(n5621), .B2(n3828), .A(n3747), .ZN(n5301) );
  INV_X1 U4792 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3749) );
  XNOR2_X1 U4793 ( .A(n3773), .B(n3749), .ZN(n5266) );
  AOI22_X1 U4794 ( .A1(n3897), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4795 ( .A1(n3776), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4796 ( .A1(n3889), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4797 ( .A1(n3871), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4798 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4799 ( .A1(n3892), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4800 ( .A1(n3890), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4801 ( .A1(n3900), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4802 ( .A1(n3405), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4803 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  OR2_X1 U4804 ( .A1(n3759), .A2(n3758), .ZN(n3775) );
  AOI22_X1 U4805 ( .A1(n3897), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4806 ( .A1(n3776), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4807 ( .A1(n3889), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3761) );
  INV_X1 U4808 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U4809 ( .A1(n3871), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4810 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3769)
         );
  AOI22_X1 U4811 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3892), .B1(n3898), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4812 ( .A1(n3890), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4813 ( .A1(n3900), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4814 ( .A1(n3405), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4815 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  OR2_X1 U4816 ( .A1(n3769), .A2(n3768), .ZN(n3774) );
  XNOR2_X1 U4817 ( .A(n3775), .B(n3774), .ZN(n3771) );
  AOI22_X1 U4818 ( .A1(n3573), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5034), .ZN(n3770) );
  OAI21_X1 U4819 ( .B1(n3910), .B2(n3771), .A(n3770), .ZN(n3772) );
  MUX2_X1 U4820 ( .A(n5266), .B(n3772), .S(n3828), .Z(n4403) );
  XNOR2_X1 U4821 ( .A(n3806), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5601)
         );
  AOI22_X1 U4822 ( .A1(n3573), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n3915), .ZN(n3790) );
  AND2_X1 U4823 ( .A1(n3775), .A2(n3774), .ZN(n3801) );
  AOI22_X1 U4824 ( .A1(n3897), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4825 ( .A1(n3776), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4826 ( .A1(n3696), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4827 ( .A1(n3871), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4828 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3786)
         );
  AOI22_X1 U4829 ( .A1(n3892), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4830 ( .A1(n3890), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4831 ( .A1(n3900), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4832 ( .A1(n3405), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4833 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  NOR2_X1 U4834 ( .A1(n3801), .A2(n3802), .ZN(n3787) );
  AOI21_X1 U4835 ( .B1(n3801), .B2(n3802), .A(n3787), .ZN(n3788) );
  NAND2_X1 U4836 ( .A1(n3884), .A2(n3788), .ZN(n3789) );
  OAI211_X1 U4837 ( .C1(n5601), .C2(n3828), .A(n3790), .B(n3789), .ZN(n5258)
         );
  AOI22_X1 U4838 ( .A1(n3897), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4839 ( .A1(n3776), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4840 ( .A1(n3889), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4841 ( .A1(n3871), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4842 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4843 ( .A1(n3892), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4844 ( .A1(n3890), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4845 ( .A1(n3900), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4846 ( .A1(n3405), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4847 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  OR2_X1 U4848 ( .A1(n3800), .A2(n3799), .ZN(n3824) );
  XOR2_X1 U4849 ( .A(n3824), .B(n3825), .Z(n3805) );
  INV_X1 U4850 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3803) );
  OAI22_X1 U4851 ( .A1(n3692), .A2(n3803), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5595), .ZN(n3804) );
  AOI21_X1 U4852 ( .B1(n3884), .B2(n3805), .A(n3804), .ZN(n3807) );
  XNOR2_X1 U4853 ( .A(n2970), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5597)
         );
  MUX2_X1 U4854 ( .A(n3807), .B(n5597), .S(n3986), .Z(n5244) );
  INV_X1 U4855 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U4856 ( .A1(n3809), .A2(n3808), .ZN(n3810) );
  NAND2_X1 U4857 ( .A1(n3863), .A2(n3810), .ZN(n5589) );
  AOI22_X1 U4858 ( .A1(n3889), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4859 ( .A1(n3871), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4860 ( .A1(n3890), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4861 ( .A1(n3558), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4862 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3823)
         );
  AOI22_X1 U4863 ( .A1(n3846), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4864 ( .A1(n3344), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4865 ( .A1(n4585), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4866 ( .A1(n3900), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4867 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3822)
         );
  NOR2_X1 U4868 ( .A1(n3823), .A2(n3822), .ZN(n3831) );
  NAND2_X1 U4869 ( .A1(n3825), .A2(n3824), .ZN(n3830) );
  XNOR2_X1 U4870 ( .A(n3831), .B(n3830), .ZN(n3827) );
  AOI22_X1 U4871 ( .A1(n3573), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5034), .ZN(n3826) );
  OAI21_X1 U4872 ( .B1(n3827), .B2(n3910), .A(n3826), .ZN(n3829) );
  MUX2_X1 U4873 ( .A(n5589), .B(n3829), .S(n3828), .Z(n5233) );
  NOR2_X1 U4874 ( .A1(n3831), .A2(n3830), .ZN(n3860) );
  AOI22_X1 U4875 ( .A1(n3847), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4876 ( .A1(n3776), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4877 ( .A1(n3889), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4878 ( .A1(n3871), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4879 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3841)
         );
  AOI22_X1 U4880 ( .A1(n3892), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4881 ( .A1(n3890), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4882 ( .A1(n3900), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4883 ( .A1(n3405), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3836) );
  NAND4_X1 U4884 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3840)
         );
  OR2_X1 U4885 ( .A1(n3841), .A2(n3840), .ZN(n3859) );
  XOR2_X1 U4886 ( .A(n3860), .B(n3859), .Z(n3844) );
  INV_X1 U4887 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3842) );
  OAI22_X1 U4888 ( .A1(n3692), .A2(n3842), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5582), .ZN(n3843) );
  AOI21_X1 U4889 ( .B1(n3844), .B2(n3884), .A(n3843), .ZN(n3845) );
  XNOR2_X1 U4890 ( .A(n3863), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5580)
         );
  MUX2_X1 U4891 ( .A(n3845), .B(n5580), .S(n3986), .Z(n5223) );
  NOR2_X2 U4892 ( .A1(n5222), .A2(n5223), .ZN(n5157) );
  AOI22_X1 U4893 ( .A1(n3847), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4894 ( .A1(n3871), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4895 ( .A1(n3892), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4896 ( .A1(n3816), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4897 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3858)
         );
  AOI22_X1 U4898 ( .A1(n3890), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4899 ( .A1(n3889), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4900 ( .A1(n3891), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4901 ( .A1(n3405), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4902 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  NOR2_X1 U4903 ( .A1(n3858), .A2(n3857), .ZN(n3870) );
  NAND2_X1 U4904 ( .A1(n3860), .A2(n3859), .ZN(n3869) );
  XNOR2_X1 U4905 ( .A(n3870), .B(n3869), .ZN(n3862) );
  AOI22_X1 U4906 ( .A1(n3573), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5034), .ZN(n3861) );
  OAI21_X1 U4907 ( .B1(n3862), .B2(n3910), .A(n3861), .ZN(n3868) );
  INV_X1 U4908 ( .A(n3864), .ZN(n3866) );
  INV_X1 U4909 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3865) );
  NAND2_X1 U4910 ( .A1(n3866), .A2(n3865), .ZN(n3867) );
  NAND2_X1 U4911 ( .A1(n3912), .A2(n3867), .ZN(n5215) );
  MUX2_X1 U4912 ( .A(n3868), .B(n5215), .S(n3986), .Z(n5158) );
  NOR2_X1 U4913 ( .A1(n3870), .A2(n3869), .ZN(n3888) );
  AOI22_X1 U4914 ( .A1(n3897), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4915 ( .A1(n3891), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4585), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4916 ( .A1(n3889), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4917 ( .A1(n3871), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4918 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3881)
         );
  AOI22_X1 U4919 ( .A1(n3892), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3558), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4920 ( .A1(n3890), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4921 ( .A1(n3900), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3848), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4922 ( .A1(n3405), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4923 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3880)
         );
  OR2_X1 U4924 ( .A1(n3881), .A2(n3880), .ZN(n3887) );
  XOR2_X1 U4925 ( .A(n3888), .B(n3887), .Z(n3885) );
  INV_X1 U4926 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3882) );
  OAI22_X1 U4927 ( .A1(n3692), .A2(n3882), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5573), .ZN(n3883) );
  AOI21_X1 U4928 ( .B1(n3885), .B2(n3884), .A(n3883), .ZN(n3886) );
  XNOR2_X1 U4929 ( .A(n3912), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5571)
         );
  MUX2_X1 U4930 ( .A(n3886), .B(n5571), .S(n3986), .Z(n4121) );
  NAND2_X1 U4931 ( .A1(n3888), .A2(n3887), .ZN(n3908) );
  AOI22_X1 U4932 ( .A1(n3889), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4933 ( .A1(n3890), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3344), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4934 ( .A1(n3891), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4935 ( .A1(n3892), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4936 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3906)
         );
  AOI22_X1 U4937 ( .A1(n3897), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4938 ( .A1(n3558), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4939 ( .A1(n4585), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4940 ( .A1(n3816), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4941 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3905)
         );
  NOR2_X1 U4942 ( .A1(n3906), .A2(n3905), .ZN(n3907) );
  XNOR2_X1 U4943 ( .A(n3908), .B(n3907), .ZN(n3911) );
  AOI22_X1 U4944 ( .A1(n3573), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5034), .ZN(n3909) );
  OAI21_X1 U4945 ( .B1(n3911), .B2(n3910), .A(n3909), .ZN(n3914) );
  INV_X1 U4946 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3913) );
  XNOR2_X1 U4947 ( .A(n3918), .B(n3913), .ZN(n4361) );
  MUX2_X1 U4948 ( .A(n3914), .B(n4361), .S(n3986), .Z(n4308) );
  AOI22_X1 U4949 ( .A1(n3573), .A2(EAX_REG_31__SCAN_IN), .B1(n3915), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3916) );
  INV_X1 U4950 ( .A(n3935), .ZN(n3921) );
  XNOR2_X1 U4951 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3936) );
  XNOR2_X1 U4952 ( .A(n3921), .B(n3936), .ZN(n3982) );
  INV_X1 U4953 ( .A(n3982), .ZN(n3933) );
  AND2_X1 U4954 ( .A1(n5201), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3922)
         );
  NOR2_X1 U4955 ( .A1(n3935), .A2(n3922), .ZN(n3928) );
  NAND2_X1 U4956 ( .A1(n4264), .A2(n3928), .ZN(n3923) );
  NAND2_X1 U4957 ( .A1(n3923), .A2(n4230), .ZN(n3925) );
  NAND2_X1 U4958 ( .A1(n3231), .A2(n4230), .ZN(n3924) );
  NAND2_X1 U4959 ( .A1(n3924), .A2(n3990), .ZN(n3950) );
  NAND2_X1 U4960 ( .A1(n3925), .A2(n3950), .ZN(n3932) );
  NAND2_X1 U4961 ( .A1(n3969), .A2(n4235), .ZN(n3927) );
  NAND2_X1 U4962 ( .A1(n3927), .A2(n3926), .ZN(n3934) );
  AND2_X1 U4963 ( .A1(n3969), .A2(n3928), .ZN(n3929) );
  OAI211_X1 U4964 ( .C1(n3934), .C2(n3982), .A(n3929), .B(n3932), .ZN(n3930)
         );
  NAND2_X1 U4965 ( .A1(n3930), .A2(n3963), .ZN(n3931) );
  OAI21_X1 U4966 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n3943) );
  NAND3_X1 U4967 ( .A1(n3934), .A2(STATE2_REG_0__SCAN_IN), .A3(n3982), .ZN(
        n3942) );
  NAND2_X1 U4968 ( .A1(n3936), .A2(n3935), .ZN(n3938) );
  NAND2_X1 U4969 ( .A1(n4671), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3937) );
  NAND2_X1 U4970 ( .A1(n3938), .A2(n3937), .ZN(n3946) );
  XNOR2_X1 U4971 ( .A(n3947), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3944)
         );
  XNOR2_X1 U4972 ( .A(n3946), .B(n3944), .ZN(n3981) );
  INV_X1 U4973 ( .A(n3303), .ZN(n3958) );
  NAND2_X1 U4974 ( .A1(n3969), .A2(n3981), .ZN(n3939) );
  OAI211_X1 U4975 ( .C1(n3981), .C2(n3958), .A(n3939), .B(n3950), .ZN(n3940)
         );
  INV_X1 U4976 ( .A(n3940), .ZN(n3941) );
  AOI21_X1 U4977 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3962) );
  INV_X1 U4978 ( .A(n3944), .ZN(n3945) );
  NAND2_X1 U4979 ( .A1(n3946), .A2(n3945), .ZN(n3949) );
  NAND2_X1 U4980 ( .A1(n3947), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3948) );
  NAND2_X1 U4981 ( .A1(n3949), .A2(n3948), .ZN(n3955) );
  XNOR2_X1 U4982 ( .A(n6312), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3953)
         );
  XNOR2_X1 U4983 ( .A(n3955), .B(n3953), .ZN(n3983) );
  INV_X1 U4984 ( .A(n4201), .ZN(n4196) );
  INV_X1 U4985 ( .A(n3950), .ZN(n3951) );
  NAND3_X1 U4986 ( .A1(n3951), .A2(n3981), .A3(n3969), .ZN(n3952) );
  OAI21_X1 U4987 ( .B1(n3983), .B2(n4196), .A(n3952), .ZN(n3961) );
  INV_X1 U4988 ( .A(n3953), .ZN(n3954) );
  NAND2_X1 U4989 ( .A1(n3955), .A2(n3954), .ZN(n3957) );
  NAND2_X1 U4990 ( .A1(n6312), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3956) );
  NAND2_X1 U4991 ( .A1(n3957), .A2(n3956), .ZN(n3966) );
  INV_X1 U4992 ( .A(n3983), .ZN(n3959) );
  OAI21_X1 U4993 ( .B1(n3964), .B2(n3959), .A(n3958), .ZN(n3960) );
  OAI21_X1 U4994 ( .B1(n3962), .B2(n3961), .A(n3960), .ZN(n3972) );
  AOI22_X1 U4995 ( .A1(n3973), .A2(n3964), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6513), .ZN(n3971) );
  NAND2_X1 U4996 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4491), .ZN(n3967) );
  NAND2_X1 U4997 ( .A1(n3969), .A2(n3979), .ZN(n3970) );
  NAND3_X1 U4998 ( .A1(n3972), .A2(n3971), .A3(n3970), .ZN(n3975) );
  NAND2_X1 U4999 ( .A1(n3978), .A2(n4735), .ZN(n4684) );
  INV_X1 U5000 ( .A(n3979), .ZN(n3985) );
  NAND4_X1 U5001 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  NAND2_X1 U5002 ( .A1(n3985), .A2(n3984), .ZN(n4678) );
  NAND2_X1 U5003 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6601), .ZN(n4766) );
  INV_X1 U5004 ( .A(n4311), .ZN(n3987) );
  NAND2_X1 U5005 ( .A1(n3987), .A2(n3986), .ZN(n6518) );
  OAI21_X1 U5006 ( .B1(n4766), .B2(n6513), .A(n6518), .ZN(n3988) );
  NAND2_X1 U5007 ( .A1(n5166), .A2(n6087), .ZN(n4119) );
  OR2_X2 U5008 ( .A1(n3990), .A2(n4735), .ZN(n4000) );
  NAND2_X1 U5009 ( .A1(n4000), .A2(n3991), .ZN(n3992) );
  INV_X1 U5010 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3993) );
  INV_X1 U5011 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U5012 ( .A1(n3991), .A2(n5475), .ZN(n3994) );
  OAI21_X1 U5013 ( .B1(n4080), .B2(n5475), .A(n3994), .ZN(n4552) );
  MUX2_X1 U5014 ( .A(n4087), .B(n3991), .S(EBX_REG_2__SCAN_IN), .Z(n3998) );
  NOR2_X1 U5015 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3997)
         );
  NOR2_X1 U5016 ( .A1(n3998), .A2(n3997), .ZN(n4643) );
  NAND2_X1 U5017 ( .A1(n4644), .A2(n4643), .ZN(n4642) );
  INV_X1 U5018 ( .A(EBX_REG_3__SCAN_IN), .ZN(n3999) );
  NAND2_X1 U5019 ( .A1(n4068), .A2(n3999), .ZN(n4003) );
  INV_X1 U5020 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U5021 ( .A1(n4080), .A2(n6285), .ZN(n4001) );
  OAI211_X1 U5022 ( .C1(n4000), .C2(EBX_REG_3__SCAN_IN), .A(n4088), .B(n4001), 
        .ZN(n4002) );
  AND2_X1 U5023 ( .A1(n4003), .A2(n4002), .ZN(n4706) );
  INV_X1 U5024 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U5025 ( .A1(n4087), .A2(n6685), .ZN(n4008) );
  NAND2_X1 U5026 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4006)
         );
  OAI211_X1 U5027 ( .C1(n4000), .C2(EBX_REG_4__SCAN_IN), .A(n4006), .B(n4080), 
        .ZN(n4007) );
  NAND2_X1 U5028 ( .A1(n4008), .A2(n4007), .ZN(n4752) );
  INV_X1 U5029 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U5030 ( .A1(n4080), .A2(n6744), .ZN(n4009) );
  OAI211_X1 U5031 ( .C1(n4000), .C2(EBX_REG_5__SCAN_IN), .A(n4088), .B(n4009), 
        .ZN(n4010) );
  OAI21_X1 U5032 ( .B1(n4079), .B2(EBX_REG_5__SCAN_IN), .A(n4010), .ZN(n4885)
         );
  MUX2_X1 U5033 ( .A(n4087), .B(n3991), .S(EBX_REG_6__SCAN_IN), .Z(n4012) );
  NOR2_X1 U5034 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4011)
         );
  NOR2_X1 U5035 ( .A1(n4012), .A2(n4011), .ZN(n4974) );
  INV_X1 U5036 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U5037 ( .A1(n4068), .A2(n4013), .ZN(n4016) );
  INV_X1 U5038 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U5039 ( .B1(n3991), .B2(n6235), .A(n4080), .ZN(n4014) );
  OAI21_X1 U5040 ( .B1(EBX_REG_9__SCAN_IN), .B2(n4000), .A(n4014), .ZN(n4015)
         );
  AND2_X1 U5041 ( .A1(n4016), .A2(n4015), .ZN(n4986) );
  MUX2_X1 U5042 ( .A(n4087), .B(n3991), .S(EBX_REG_8__SCAN_IN), .Z(n4017) );
  INV_X1 U5043 ( .A(n4017), .ZN(n4018) );
  NAND2_X1 U5044 ( .A1(n4018), .A2(n3121), .ZN(n5122) );
  NOR2_X1 U5045 ( .A1(n4986), .A2(n5122), .ZN(n4023) );
  INV_X1 U5046 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U5047 ( .A1(n4068), .A2(n4019), .ZN(n4022) );
  NAND2_X1 U5048 ( .A1(n4080), .A2(n6259), .ZN(n4020) );
  OAI211_X1 U5049 ( .C1(n4000), .C2(EBX_REG_7__SCAN_IN), .A(n4088), .B(n4020), 
        .ZN(n4021) );
  MUX2_X1 U5050 ( .A(n4087), .B(n3991), .S(EBX_REG_10__SCAN_IN), .Z(n4025) );
  NOR2_X1 U5051 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4024)
         );
  NOR2_X1 U5052 ( .A1(n4025), .A2(n4024), .ZN(n5124) );
  NAND2_X1 U5053 ( .A1(n4985), .A2(n5124), .ZN(n4425) );
  INV_X1 U5054 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U5055 ( .A1(n4068), .A2(n5518), .ZN(n4028) );
  INV_X1 U5056 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U5057 ( .A1(n4080), .A2(n5685), .ZN(n4026) );
  OAI211_X1 U5058 ( .C1(n4000), .C2(EBX_REG_11__SCAN_IN), .A(n4088), .B(n4026), 
        .ZN(n4027) );
  INV_X1 U5059 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U5060 ( .A1(n4087), .A2(n5512), .ZN(n4033) );
  NAND2_X1 U5061 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4031) );
  OAI211_X1 U5062 ( .C1(n4000), .C2(EBX_REG_12__SCAN_IN), .A(n4031), .B(n4080), 
        .ZN(n4032) );
  NAND2_X1 U5063 ( .A1(n4033), .A2(n4032), .ZN(n5403) );
  INV_X1 U5064 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4034) );
  OAI21_X1 U5065 ( .B1(n3991), .B2(n4034), .A(n4080), .ZN(n4035) );
  OAI21_X1 U5066 ( .B1(EBX_REG_13__SCAN_IN), .B2(n4000), .A(n4035), .ZN(n4036)
         );
  OAI21_X1 U5067 ( .B1(n4079), .B2(EBX_REG_13__SCAN_IN), .A(n4036), .ZN(n5507)
         );
  MUX2_X1 U5068 ( .A(n4087), .B(n3991), .S(EBX_REG_14__SCAN_IN), .Z(n4037) );
  INV_X1 U5069 ( .A(n4037), .ZN(n4038) );
  OAI21_X1 U5070 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n4551), .A(n4038), 
        .ZN(n5388) );
  INV_X1 U5071 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U5072 ( .A1(n4087), .A2(n5503), .ZN(n4041) );
  NAND2_X1 U5073 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4039) );
  OAI211_X1 U5074 ( .C1(EBX_REG_16__SCAN_IN), .C2(n4000), .A(n4039), .B(n4080), 
        .ZN(n4040) );
  AND2_X1 U5075 ( .A1(n4041), .A2(n4040), .ZN(n5359) );
  NAND2_X1 U5076 ( .A1(n4080), .A2(n6750), .ZN(n4042) );
  OAI211_X1 U5077 ( .C1(n4000), .C2(EBX_REG_15__SCAN_IN), .A(n4088), .B(n4042), 
        .ZN(n4043) );
  OAI21_X1 U5078 ( .B1(n4079), .B2(EBX_REG_15__SCAN_IN), .A(n4043), .ZN(n5375)
         );
  NAND2_X1 U5079 ( .A1(n4080), .A2(n5803), .ZN(n4044) );
  OAI211_X1 U5080 ( .C1(n4000), .C2(EBX_REG_17__SCAN_IN), .A(n4088), .B(n4044), 
        .ZN(n4045) );
  OAI21_X1 U5081 ( .B1(n4079), .B2(EBX_REG_17__SCAN_IN), .A(n4045), .ZN(n5344)
         );
  AND2_X2 U5082 ( .A1(n5361), .A2(n5344), .ZN(n5345) );
  INV_X1 U5083 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U5084 ( .A1(n4087), .A2(n4046), .ZN(n4049) );
  NAND2_X1 U5085 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4047) );
  OAI211_X1 U5086 ( .C1(EBX_REG_19__SCAN_IN), .C2(n4000), .A(n4047), .B(n4080), 
        .ZN(n4048) );
  INV_X1 U5087 ( .A(n4551), .ZN(n4050) );
  INV_X1 U5088 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U5089 ( .A1(n4050), .A2(n5779), .ZN(n4051) );
  INV_X1 U5090 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U5091 ( .A1(n4567), .A2(n5501), .ZN(n4323) );
  OAI22_X1 U5092 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4000), .ZN(n5304) );
  NAND2_X1 U5093 ( .A1(n5303), .A2(n5304), .ZN(n4053) );
  NAND2_X1 U5094 ( .A1(n3991), .A2(EBX_REG_20__SCAN_IN), .ZN(n4052) );
  OAI211_X1 U5095 ( .C1(n5303), .C2(n3991), .A(n4053), .B(n4052), .ZN(n4054)
         );
  INV_X1 U5096 ( .A(EBX_REG_21__SCAN_IN), .ZN(n4055) );
  NAND2_X1 U5097 ( .A1(n4068), .A2(n4055), .ZN(n4058) );
  INV_X1 U5098 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U5099 ( .A1(n4080), .A2(n5169), .ZN(n4056) );
  OAI211_X1 U5100 ( .C1(n4000), .C2(EBX_REG_21__SCAN_IN), .A(n4088), .B(n4056), 
        .ZN(n4057) );
  MUX2_X1 U5101 ( .A(n4087), .B(n3991), .S(EBX_REG_22__SCAN_IN), .Z(n4060) );
  NOR2_X1 U5102 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4059)
         );
  NOR2_X1 U5103 ( .A1(n4060), .A2(n4059), .ZN(n5184) );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5105 ( .A1(n4080), .A2(n4369), .ZN(n4061) );
  OAI211_X1 U5106 ( .C1(n4000), .C2(EBX_REG_23__SCAN_IN), .A(n4088), .B(n4061), 
        .ZN(n4062) );
  OAI21_X1 U5107 ( .B1(n4079), .B2(EBX_REG_23__SCAN_IN), .A(n4062), .ZN(n4392)
         );
  NAND2_X1 U5108 ( .A1(n4391), .A2(n4392), .ZN(n4377) );
  INV_X1 U5109 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4063) );
  NAND2_X1 U5110 ( .A1(n4087), .A2(n4063), .ZN(n4066) );
  NAND2_X1 U5111 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4064) );
  OAI211_X1 U5112 ( .C1(EBX_REG_24__SCAN_IN), .C2(n4000), .A(n4064), .B(n4080), 
        .ZN(n4065) );
  NAND2_X1 U5113 ( .A1(n4066), .A2(n4065), .ZN(n4379) );
  INV_X1 U5114 ( .A(EBX_REG_25__SCAN_IN), .ZN(n4067) );
  NAND2_X1 U5115 ( .A1(n4068), .A2(n4067), .ZN(n4071) );
  INV_X1 U5116 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5142) );
  OAI21_X1 U5117 ( .B1(n3991), .B2(n5142), .A(n4080), .ZN(n4069) );
  OAI21_X1 U5118 ( .B1(EBX_REG_25__SCAN_IN), .B2(n4000), .A(n4069), .ZN(n4070)
         );
  INV_X1 U5119 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U5120 ( .A1(n4087), .A2(n6735), .ZN(n4075) );
  NAND2_X1 U5121 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4073) );
  OAI211_X1 U5122 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4000), .A(n4073), .B(n4080), 
        .ZN(n4074) );
  NAND2_X1 U5123 ( .A1(n4075), .A2(n4074), .ZN(n5235) );
  INV_X1 U5124 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4076) );
  NAND2_X1 U5125 ( .A1(n4080), .A2(n4076), .ZN(n4077) );
  OAI211_X1 U5126 ( .C1(n4000), .C2(EBX_REG_27__SCAN_IN), .A(n4088), .B(n4077), 
        .ZN(n4078) );
  OAI21_X1 U5127 ( .B1(n4079), .B2(EBX_REG_27__SCAN_IN), .A(n4078), .ZN(n5227)
         );
  INV_X1 U5128 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U5129 ( .A1(n4087), .A2(n5487), .ZN(n4083) );
  NAND2_X1 U5130 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4081) );
  OAI211_X1 U5131 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4000), .A(n4081), .B(n4080), 
        .ZN(n4082) );
  NAND2_X1 U5132 ( .A1(n4083), .A2(n4082), .ZN(n5147) );
  NOR2_X1 U5133 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4089)
         );
  INV_X1 U5134 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4084) );
  INV_X1 U5135 ( .A(n4087), .ZN(n4092) );
  MUX2_X1 U5136 ( .A(EBX_REG_29__SCAN_IN), .B(n4089), .S(n4088), .Z(n4090) );
  INV_X1 U5137 ( .A(n4090), .ZN(n4091) );
  OAI21_X1 U5138 ( .B1(EBX_REG_29__SCAN_IN), .B2(n4092), .A(n4091), .ZN(n5206)
         );
  AOI22_X1 U5139 ( .A1(n4551), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n4000), .ZN(n4347) );
  NAND2_X1 U5140 ( .A1(n5205), .A2(n4347), .ZN(n4093) );
  OAI22_X1 U5141 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4000), .ZN(n4094) );
  INV_X1 U5142 ( .A(n4094), .ZN(n4095) );
  NOR2_X1 U5143 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4112) );
  NAND2_X1 U5144 ( .A1(n4567), .A2(EBX_REG_31__SCAN_IN), .ZN(n4097) );
  OAI211_X1 U5145 ( .C1(n4686), .C2(n4235), .A(n4230), .B(n4112), .ZN(n4099)
         );
  INV_X1 U5146 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6529) );
  INV_X1 U5147 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6527) );
  NAND3_X1 U5148 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6094) );
  OR2_X1 U5149 ( .A1(n6527), .A2(n6094), .ZN(n5434) );
  NOR2_X1 U5150 ( .A1(n6529), .A2(n5434), .ZN(n5421) );
  INV_X1 U5151 ( .A(n5421), .ZN(n5422) );
  NOR2_X1 U5152 ( .A1(n6749), .A2(n5422), .ZN(n5420) );
  NAND3_X1 U5153 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n5420), .ZN(n5413) );
  NOR2_X2 U5154 ( .A1(n6095), .A2(n5413), .ZN(n6064) );
  NAND4_X1 U5155 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n6064), .ZN(n5409) );
  NOR2_X2 U5156 ( .A1(n6540), .A2(n5409), .ZN(n6045) );
  AND2_X1 U5157 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n4105) );
  AND3_X1 U5158 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U5159 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5308) );
  INV_X1 U5160 ( .A(n5308), .ZN(n4100) );
  AND2_X1 U5161 ( .A1(REIP_REG_20__SCAN_IN), .A2(n4100), .ZN(n4101) );
  NAND2_X1 U5162 ( .A1(n5324), .A2(n4101), .ZN(n5282) );
  NAND2_X1 U5163 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n4102) );
  NOR2_X1 U5164 ( .A1(n5282), .A2(n4102), .ZN(n5267) );
  NAND2_X1 U5165 ( .A1(n5267), .A2(REIP_REG_23__SCAN_IN), .ZN(n5255) );
  INV_X1 U5166 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6559) );
  OR2_X1 U5167 ( .A1(n5255), .A2(n6559), .ZN(n4103) );
  NAND2_X1 U5168 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n4108) );
  NOR2_X2 U5169 ( .A1(n5237), .A2(n4108), .ZN(n5230) );
  AND2_X1 U5170 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4111) );
  NAND2_X1 U5171 ( .A1(n5230), .A2(n4111), .ZN(n4353) );
  NOR2_X1 U5172 ( .A1(n4353), .A2(REIP_REG_29__SCAN_IN), .ZN(n5211) );
  INV_X1 U5173 ( .A(n5441), .ZN(n5466) );
  NAND3_X1 U5174 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n4104) );
  NOR3_X1 U5175 ( .A1(n5466), .A2(n5413), .A3(n4104), .ZN(n4423) );
  NAND2_X1 U5176 ( .A1(REIP_REG_12__SCAN_IN), .A2(n4423), .ZN(n5408) );
  INV_X1 U5177 ( .A(n4105), .ZN(n4106) );
  NAND2_X1 U5178 ( .A1(n6095), .A2(n5441), .ZN(n5479) );
  OAI21_X1 U5179 ( .B1(n5408), .B2(n4106), .A(n5479), .ZN(n5395) );
  NAND2_X1 U5180 ( .A1(n5479), .A2(n5255), .ZN(n4107) );
  NAND2_X1 U5181 ( .A1(n5395), .A2(n4107), .ZN(n5259) );
  INV_X1 U5182 ( .A(n4108), .ZN(n4109) );
  INV_X1 U5183 ( .A(n5479), .ZN(n4424) );
  AOI21_X1 U5184 ( .B1(REIP_REG_24__SCAN_IN), .B2(n4109), .A(n4424), .ZN(n4110) );
  NOR2_X1 U5185 ( .A1(n5259), .A2(n4110), .ZN(n5238) );
  OAI21_X1 U5186 ( .B1(n4111), .B2(n6095), .A(n5238), .ZN(n5218) );
  NOR2_X1 U5187 ( .A1(n5211), .A2(n5218), .ZN(n4364) );
  OAI21_X1 U5188 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6095), .A(n4364), .ZN(n4117) );
  INV_X1 U5189 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6709) );
  INV_X1 U5190 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6568) );
  NOR4_X1 U5191 ( .A1(n4353), .A2(REIP_REG_31__SCAN_IN), .A3(n6709), .A4(n6568), .ZN(n4116) );
  NAND2_X1 U5192 ( .A1(n4686), .A2(n4112), .ZN(n4697) );
  NAND2_X1 U5193 ( .A1(n4499), .A2(n4697), .ZN(n4113) );
  OR2_X1 U5194 ( .A1(n5446), .A2(n4113), .ZN(n4357) );
  INV_X1 U5195 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5203) );
  OAI22_X1 U5196 ( .A1(n6068), .A2(n4114), .B1(n4357), .B2(n5203), .ZN(n4115)
         );
  AOI211_X1 U5197 ( .C1(n4117), .C2(REIP_REG_31__SCAN_IN), .A(n4116), .B(n4115), .ZN(n4118) );
  AOI21_X1 U5198 ( .B1(n4120), .B2(n4121), .A(n4310), .ZN(n5575) );
  INV_X1 U5199 ( .A(n5575), .ZN(n5485) );
  NAND2_X1 U5200 ( .A1(n4663), .A2(n4735), .ZN(n4123) );
  NAND2_X1 U5201 ( .A1(n6771), .A2(n4123), .ZN(n4242) );
  INV_X1 U5202 ( .A(n4251), .ZN(n5428) );
  NOR2_X1 U5203 ( .A1(READY_N), .A2(n4678), .ZN(n4475) );
  NAND2_X1 U5204 ( .A1(n6517), .A2(n4475), .ZN(n4128) );
  NOR2_X1 U5205 ( .A1(n4416), .A2(n4125), .ZN(n4126) );
  NAND3_X1 U5206 ( .A1(n4127), .A2(n4126), .A3(n3026), .ZN(n4411) );
  OAI22_X1 U5207 ( .A1(n2953), .A2(n4128), .B1(n4513), .B2(n4411), .ZN(n4129)
         );
  INV_X1 U5208 ( .A(n4129), .ZN(n4131) );
  NAND2_X1 U5209 ( .A1(n3236), .A2(n4416), .ZN(n4132) );
  AOI22_X1 U5210 ( .A1(n5554), .A2(DATAI_29_), .B1(n5564), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n4135) );
  AND2_X1 U5211 ( .A1(n3231), .A2(n4416), .ZN(n4133) );
  NAND2_X1 U5212 ( .A1(n5555), .A2(DATAI_13_), .ZN(n4134) );
  OAI21_X1 U5213 ( .B1(n5485), .B2(n5567), .A(n3117), .ZN(U2862) );
  NAND2_X1 U5214 ( .A1(n4137), .A2(n4142), .ZN(n4161) );
  OAI21_X1 U5215 ( .B1(n4137), .B2(n4142), .A(n4161), .ZN(n4138) );
  OAI211_X1 U5216 ( .C1(n4138), .C2(n6600), .A(n3098), .B(n3926), .ZN(n4139)
         );
  INV_X1 U5217 ( .A(n4139), .ZN(n4140) );
  NAND2_X1 U5218 ( .A1(n4735), .A2(n4141), .ZN(n4150) );
  OAI21_X1 U5219 ( .B1(n6600), .B2(n4142), .A(n4150), .ZN(n4143) );
  INV_X1 U5220 ( .A(n4143), .ZN(n4144) );
  AND2_X1 U5221 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U5222 ( .A1(n4545), .A2(n6291), .ZN(n4148) );
  NAND2_X1 U5223 ( .A1(n4545), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4146)
         );
  NAND2_X1 U5224 ( .A1(n4146), .A2(n6297), .ZN(n4147) );
  AND2_X1 U5225 ( .A1(n4148), .A2(n4147), .ZN(n4569) );
  NAND2_X1 U5226 ( .A1(n4570), .A2(n4569), .ZN(n4149) );
  NAND2_X1 U5227 ( .A1(n6213), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4154)
         );
  XNOR2_X1 U5228 ( .A(n4161), .B(n4159), .ZN(n4151) );
  OAI21_X1 U5229 ( .B1(n4151), .B2(n6600), .A(n4150), .ZN(n4152) );
  AOI21_X2 U5230 ( .B1(n4153), .B2(n4201), .A(n4152), .ZN(n6215) );
  NAND2_X1 U5231 ( .A1(n4154), .A2(n6215), .ZN(n4158) );
  NAND2_X1 U5232 ( .A1(n4156), .A2(n4155), .ZN(n4157) );
  INV_X1 U5233 ( .A(n4159), .ZN(n4160) );
  NAND2_X1 U5234 ( .A1(n4161), .A2(n4160), .ZN(n4170) );
  INV_X1 U5235 ( .A(n4169), .ZN(n4162) );
  XNOR2_X1 U5236 ( .A(n4170), .B(n4162), .ZN(n4163) );
  NAND2_X1 U5237 ( .A1(n4163), .A2(n4499), .ZN(n4164) );
  OAI21_X2 U5238 ( .B1(n4165), .B2(n4196), .A(n4164), .ZN(n4166) );
  XNOR2_X1 U5239 ( .A(n4166), .B(n6285), .ZN(n4757) );
  NAND2_X1 U5240 ( .A1(n4755), .A2(n4757), .ZN(n4756) );
  NAND2_X1 U5241 ( .A1(n4166), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4167)
         );
  NAND2_X1 U5242 ( .A1(n4756), .A2(n4167), .ZN(n6204) );
  NAND2_X1 U5243 ( .A1(n4168), .A2(n4201), .ZN(n4173) );
  NAND2_X1 U5244 ( .A1(n4170), .A2(n4169), .ZN(n4185) );
  XNOR2_X1 U5245 ( .A(n4185), .B(n4183), .ZN(n4171) );
  NAND2_X1 U5246 ( .A1(n4171), .A2(n4499), .ZN(n4172) );
  NAND2_X1 U5247 ( .A1(n4173), .A2(n4172), .ZN(n4174) );
  INV_X1 U5248 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6277) );
  XNOR2_X1 U5249 ( .A(n4174), .B(n6277), .ZN(n6203) );
  NAND2_X1 U5250 ( .A1(n4174), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4175)
         );
  INV_X1 U5251 ( .A(n4185), .ZN(n4177) );
  NAND2_X1 U5252 ( .A1(n4177), .A2(n4183), .ZN(n4178) );
  XOR2_X1 U5253 ( .A(n4182), .B(n4178), .Z(n4179) );
  XOR2_X1 U5254 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .B(n4180), .Z(n5070) );
  INV_X1 U5255 ( .A(n4180), .ZN(n4181) );
  NAND2_X1 U5256 ( .A1(n4183), .A2(n4182), .ZN(n4184) );
  NOR2_X1 U5257 ( .A1(n4185), .A2(n4184), .ZN(n4194) );
  XNOR2_X1 U5258 ( .A(n4194), .B(n4193), .ZN(n4188) );
  NAND3_X1 U5259 ( .A1(n4200), .A2(n4201), .A3(n4186), .ZN(n4187) );
  OAI21_X1 U5260 ( .B1(n4188), .B2(n6600), .A(n4187), .ZN(n4189) );
  XOR2_X1 U5261 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .B(n4189), .Z(n6196) );
  INV_X1 U5262 ( .A(n4189), .ZN(n4190) );
  INV_X1 U5263 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6268) );
  INV_X1 U5264 ( .A(n4192), .ZN(n4197) );
  NAND2_X1 U5265 ( .A1(n4194), .A2(n4193), .ZN(n4205) );
  XOR2_X1 U5266 ( .A(n4202), .B(n4205), .Z(n4195) );
  XOR2_X1 U5267 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .B(n4198), .Z(n5723) );
  NAND2_X1 U5268 ( .A1(n4198), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4199)
         );
  NAND2_X1 U5269 ( .A1(n4499), .A2(n4202), .ZN(n4204) );
  AND2_X1 U5270 ( .A1(n4202), .A2(n4201), .ZN(n4203) );
  XOR2_X1 U5271 ( .A(n4206), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n5715) );
  INV_X1 U5272 ( .A(n4206), .ZN(n4207) );
  INV_X1 U5273 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6252) );
  INV_X4 U5274 ( .A(n5689), .ZN(n5686) );
  NAND2_X1 U5275 ( .A1(n5686), .A2(n6235), .ZN(n5705) );
  NOR2_X1 U5276 ( .A1(n5686), .A2(n6235), .ZN(n5707) );
  INV_X1 U5277 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U5278 ( .A1(n5685), .A2(n5684), .ZN(n4209) );
  OAI21_X1 U5279 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n4209), .A(n5689), 
        .ZN(n4211) );
  AOI21_X1 U5280 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5689), .ZN(n4210) );
  NOR2_X1 U5281 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5688)
         );
  NOR2_X1 U5282 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5672)
         );
  NOR2_X1 U5283 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4213) );
  NOR3_X1 U5284 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n4212) );
  AOI21_X1 U5285 ( .B1(n4213), .B2(n4212), .A(n5686), .ZN(n4215) );
  NAND2_X1 U5286 ( .A1(n5686), .A2(n6750), .ZN(n4322) );
  INV_X1 U5287 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U5288 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5780) );
  OAI21_X1 U5289 ( .B1(n5820), .B2(n5780), .A(n5686), .ZN(n4214) );
  NOR2_X1 U5290 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5626)
         );
  NAND2_X1 U5291 ( .A1(n5181), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U5292 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4370) );
  OAI21_X1 U5293 ( .B1(n4387), .B2(n4370), .A(n5686), .ZN(n4219) );
  NOR2_X1 U5294 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4381) );
  NOR2_X1 U5295 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5781) );
  NOR2_X1 U5296 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5180) );
  NAND3_X1 U5297 ( .A1(n4381), .A2(n5781), .A3(n5180), .ZN(n4216) );
  XNOR2_X1 U5298 ( .A(n5686), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5594)
         );
  NAND2_X1 U5299 ( .A1(n5141), .A2(n5594), .ZN(n4303) );
  INV_X1 U5300 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U5301 ( .A1(n5689), .A2(n6710), .ZN(n5587) );
  NOR3_X1 U5302 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4304) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5131) );
  INV_X1 U5304 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5737) );
  NAND3_X1 U5305 ( .A1(n4304), .A2(n5131), .A3(n5737), .ZN(n4221) );
  NAND2_X1 U5306 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4291) );
  NAND2_X1 U5307 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4292) );
  NAND3_X1 U5308 ( .A1(n4305), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4220) );
  XNOR2_X1 U5309 ( .A(n4222), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4340)
         );
  AOI21_X1 U5310 ( .B1(n3244), .B2(n6591), .A(n4735), .ZN(n4223) );
  NAND2_X1 U5311 ( .A1(n4680), .A2(n4223), .ZN(n4224) );
  OAI21_X1 U5312 ( .B1(n4686), .B2(n6600), .A(n4224), .ZN(n4226) );
  NAND2_X1 U5313 ( .A1(n4226), .A2(n4225), .ZN(n4240) );
  NAND2_X1 U5314 ( .A1(n4680), .A2(n4721), .ZN(n4228) );
  NOR2_X1 U5315 ( .A1(n4663), .A2(n3990), .ZN(n4270) );
  INV_X1 U5316 ( .A(n4270), .ZN(n4227) );
  NAND2_X1 U5317 ( .A1(n4228), .A2(n4227), .ZN(n4239) );
  NAND3_X1 U5318 ( .A1(n4229), .A2(n4230), .A3(n3236), .ZN(n4233) );
  INV_X1 U5319 ( .A(n3236), .ZN(n4231) );
  NAND2_X1 U5320 ( .A1(n4499), .A2(n4231), .ZN(n4232) );
  NAND2_X1 U5321 ( .A1(n4233), .A2(n4232), .ZN(n4259) );
  OR2_X1 U5322 ( .A1(n4242), .A2(n4259), .ZN(n4234) );
  NAND2_X1 U5323 ( .A1(n4684), .A2(n4234), .ZN(n4477) );
  NAND2_X1 U5324 ( .A1(n4235), .A2(n4492), .ZN(n4236) );
  NAND3_X1 U5325 ( .A1(n4236), .A2(n4475), .A3(n3221), .ZN(n4237) );
  NAND2_X1 U5326 ( .A1(n4477), .A2(n4237), .ZN(n4238) );
  AOI21_X1 U5327 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(n4241) );
  AND2_X1 U5328 ( .A1(n4527), .A2(n4689), .ZN(n4679) );
  INV_X1 U5329 ( .A(n4248), .ZN(n4243) );
  NAND2_X1 U5330 ( .A1(n4243), .A2(n4247), .ZN(n4244) );
  OAI21_X1 U5331 ( .B1(n4248), .B2(n4247), .A(n4698), .ZN(n4249) );
  INV_X1 U5332 ( .A(n4249), .ZN(n4250) );
  OAI21_X1 U5333 ( .B1(n4252), .B2(n3221), .A(n4251), .ZN(n4253) );
  OR2_X1 U5334 ( .A1(n3978), .A2(n4253), .ZN(n4262) );
  NAND2_X1 U5335 ( .A1(n4551), .A2(n4254), .ZN(n4256) );
  OAI21_X1 U5336 ( .B1(n4264), .B2(n4721), .A(n4467), .ZN(n4255) );
  NAND2_X1 U5337 ( .A1(n3250), .A2(n4735), .ZN(n4257) );
  NAND2_X1 U5338 ( .A1(n4257), .A2(n3221), .ZN(n4258) );
  NAND2_X1 U5339 ( .A1(n4271), .A2(n4258), .ZN(n4260) );
  NOR2_X1 U5340 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  NAND2_X1 U5341 ( .A1(n4262), .A2(n4261), .ZN(n4514) );
  INV_X1 U5342 ( .A(n4263), .ZN(n4267) );
  NAND2_X1 U5343 ( .A1(n4265), .A2(n4264), .ZN(n4266) );
  NAND2_X1 U5344 ( .A1(n4266), .A2(n3991), .ZN(n4512) );
  OAI21_X1 U5345 ( .B1(n4267), .B2(n4512), .A(n4596), .ZN(n4268) );
  NOR2_X1 U5346 ( .A1(n4514), .A2(n4268), .ZN(n4269) );
  NAND2_X1 U5347 ( .A1(n4271), .A2(n4270), .ZN(n4681) );
  NAND2_X1 U5348 ( .A1(n5813), .A2(n5867), .ZN(n5819) );
  AND2_X1 U5349 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4293) );
  INV_X1 U5350 ( .A(n5813), .ZN(n5870) );
  NAND2_X1 U5351 ( .A1(n5840), .A2(n4281), .ZN(n4573) );
  NAND2_X1 U5352 ( .A1(n5870), .A2(n4573), .ZN(n6296) );
  NAND2_X1 U5353 ( .A1(n5867), .A2(n6296), .ZN(n5875) );
  NOR2_X1 U5354 ( .A1(n6259), .A2(n6252), .ZN(n6247) );
  NAND3_X1 U5355 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6247), .ZN(n4273) );
  AOI21_X1 U5356 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6292) );
  NAND2_X1 U5357 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6273) );
  NOR2_X1 U5358 ( .A1(n6292), .A2(n6273), .ZN(n5072) );
  NAND2_X1 U5359 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5072), .ZN(n6263)
         );
  NOR2_X1 U5360 ( .A1(n6268), .A2(n6263), .ZN(n5868) );
  INV_X1 U5361 ( .A(n5868), .ZN(n5877) );
  OR2_X1 U5362 ( .A1(n4273), .A2(n5877), .ZN(n5811) );
  INV_X1 U5363 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4321) );
  NAND3_X1 U5364 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5844) );
  NOR2_X1 U5365 ( .A1(n4321), .A2(n5844), .ZN(n5810) );
  NAND3_X1 U5366 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5810), .ZN(n4274) );
  NOR2_X1 U5367 ( .A1(n5811), .A2(n4274), .ZN(n4327) );
  NAND2_X1 U5368 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U5369 ( .A1(n5780), .A2(n5782), .ZN(n4287) );
  NAND2_X1 U5370 ( .A1(n4327), .A2(n4287), .ZN(n4279) );
  NOR2_X1 U5371 ( .A1(n4155), .A2(n6297), .ZN(n5876) );
  INV_X1 U5372 ( .A(n5876), .ZN(n4272) );
  NOR2_X1 U5373 ( .A1(n4272), .A2(n6273), .ZN(n5073) );
  NAND3_X1 U5374 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5073), .ZN(n5871) );
  NOR2_X1 U5375 ( .A1(n5871), .A2(n4273), .ZN(n5814) );
  INV_X1 U5376 ( .A(n4274), .ZN(n4286) );
  AND2_X1 U5377 ( .A1(n5814), .A2(n4286), .ZN(n4275) );
  OR2_X1 U5378 ( .A1(n5813), .A2(n4275), .ZN(n4278) );
  OR2_X1 U5379 ( .A1(n4554), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4277)
         );
  NAND2_X1 U5380 ( .A1(n4276), .A2(n6211), .ZN(n4572) );
  NAND2_X1 U5381 ( .A1(n4278), .A2(n5866), .ZN(n4329) );
  AOI21_X1 U5382 ( .B1(n5819), .B2(n4279), .A(n4329), .ZN(n5179) );
  OAI21_X1 U5383 ( .B1(n5181), .B2(n5872), .A(n5179), .ZN(n4395) );
  AOI21_X1 U5384 ( .B1(n5875), .B2(n4370), .A(n4395), .ZN(n5754) );
  INV_X1 U5385 ( .A(n4291), .ZN(n4280) );
  NAND2_X1 U5386 ( .A1(n5754), .A2(n4280), .ZN(n5744) );
  NAND2_X1 U5387 ( .A1(n5754), .A2(n5872), .ZN(n5745) );
  OAI21_X1 U5388 ( .B1(n5744), .B2(n4292), .A(n5745), .ZN(n5738) );
  OAI21_X1 U5389 ( .B1(n5872), .B2(n4293), .A(n5738), .ZN(n4297) );
  INV_X1 U5390 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6573) );
  NOR2_X1 U5391 ( .A1(n6211), .A2(n6573), .ZN(n4337) );
  OR2_X1 U5392 ( .A1(n5867), .A2(n5811), .ZN(n4283) );
  INV_X1 U5393 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4281) );
  INV_X1 U5394 ( .A(n5814), .ZN(n4284) );
  NAND2_X1 U5395 ( .A1(n6231), .A2(n4286), .ZN(n5799) );
  INV_X1 U5396 ( .A(n4287), .ZN(n4288) );
  INV_X1 U5397 ( .A(n5181), .ZN(n4289) );
  NOR2_X1 U5398 ( .A1(n5773), .A2(n4289), .ZN(n4380) );
  INV_X1 U5399 ( .A(n4370), .ZN(n4290) );
  NAND2_X1 U5400 ( .A1(n4380), .A2(n4290), .ZN(n5765) );
  NOR2_X1 U5401 ( .A1(n5149), .A2(n4292), .ZN(n5734) );
  INV_X1 U5402 ( .A(n5734), .ZN(n4295) );
  INV_X1 U5403 ( .A(n4293), .ZN(n4294) );
  NOR3_X1 U5404 ( .A1(n4295), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4294), 
        .ZN(n4296) );
  AOI211_X1 U5405 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n4297), .A(n4337), .B(n4296), .ZN(n4298) );
  INV_X1 U5406 ( .A(n4299), .ZN(n4300) );
  NAND2_X1 U5407 ( .A1(n4305), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4306) );
  XNOR2_X1 U5408 ( .A(n4307), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5138)
         );
  NAND2_X1 U5409 ( .A1(n4312), .A2(n6593), .ZN(n4313) );
  NAND2_X1 U5410 ( .A1(n4313), .A2(n6513), .ZN(n4314) );
  NAND2_X1 U5411 ( .A1(n6513), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U5412 ( .A1(n6028), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U5413 ( .A1(n4316), .A2(n4315), .ZN(n4546) );
  NOR2_X1 U5414 ( .A1(n6211), .A2(n6568), .ZN(n5133) );
  AOI21_X1 U5415 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5133), 
        .ZN(n4317) );
  OAI21_X1 U5416 ( .B1(n4361), .B2(n6223), .A(n4317), .ZN(n4318) );
  AOI21_X1 U5417 ( .B1(n5126), .B2(n6217), .A(n4318), .ZN(n4319) );
  OAI21_X1 U5418 ( .B1(n5138), .B2(n6192), .A(n4319), .ZN(U2956) );
  NOR2_X1 U5419 ( .A1(n5686), .A2(n4321), .ZN(n5671) );
  XNOR2_X1 U5420 ( .A(n5686), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5663)
         );
  NOR2_X1 U5421 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5653)
         );
  NAND2_X1 U5422 ( .A1(n5635), .A2(n6294), .ZN(n4336) );
  INV_X1 U5423 ( .A(n4323), .ZN(n4324) );
  MUX2_X1 U5424 ( .A(n5303), .B(n4324), .S(n3991), .Z(n4325) );
  NAND2_X1 U5425 ( .A1(n5345), .A2(n4325), .ZN(n5317) );
  OR2_X1 U5426 ( .A1(n5345), .A2(n4325), .ZN(n4326) );
  NAND2_X1 U5427 ( .A1(n5317), .A2(n4326), .ZN(n5500) );
  AOI21_X1 U5428 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4327), .A(n5867), 
        .ZN(n4328) );
  NOR2_X1 U5429 ( .A1(n4329), .A2(n4328), .ZN(n5800) );
  INV_X1 U5430 ( .A(n6296), .ZN(n4330) );
  NAND2_X1 U5431 ( .A1(n5803), .A2(n4330), .ZN(n4331) );
  NAND2_X1 U5432 ( .A1(n5800), .A2(n4331), .ZN(n5778) );
  INV_X1 U5433 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6550) );
  NOR2_X1 U5434 ( .A1(n6211), .A2(n6550), .ZN(n5638) );
  NOR3_X1 U5435 ( .A1(n5799), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5803), 
        .ZN(n4332) );
  AOI211_X1 U5436 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5778), .A(n5638), .B(n4332), .ZN(n4333) );
  OAI21_X1 U5437 ( .B1(n5500), .B2(n5873), .A(n4333), .ZN(n4334) );
  INV_X1 U5438 ( .A(n4334), .ZN(n4335) );
  NAND2_X1 U5439 ( .A1(n4336), .A2(n4335), .ZN(U3000) );
  NAND2_X1 U5440 ( .A1(n5166), .A2(n6217), .ZN(n4343) );
  AOI21_X1 U5441 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4337), 
        .ZN(n4338) );
  OAI21_X1 U5442 ( .B1(n4356), .B2(n6223), .A(n4338), .ZN(n4339) );
  INV_X1 U5443 ( .A(n4339), .ZN(n4342) );
  OR2_X1 U5444 ( .A1(n4340), .A2(n6192), .ZN(n4341) );
  NAND3_X1 U5445 ( .A1(n4343), .A2(n4342), .A3(n4341), .ZN(U2955) );
  INV_X1 U5446 ( .A(n4347), .ZN(n4346) );
  OAI21_X1 U5447 ( .B1(n4350), .B2(n4345), .A(n4346), .ZN(n4351) );
  INV_X1 U5448 ( .A(n4345), .ZN(n4348) );
  OAI21_X1 U5449 ( .B1(n4348), .B2(n4088), .A(n4347), .ZN(n4349) );
  OAI22_X1 U5450 ( .A1(n4352), .A2(n4351), .B1(n4350), .B2(n4349), .ZN(n4417)
         );
  INV_X1 U5451 ( .A(n4417), .ZN(n5135) );
  NOR3_X1 U5452 ( .A1(n4353), .A2(REIP_REG_30__SCAN_IN), .A3(n6709), .ZN(n4363) );
  INV_X1 U5453 ( .A(n4354), .ZN(n4355) );
  OR2_X1 U5454 ( .A1(n4735), .A2(EBX_REG_31__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U5455 ( .A1(n5393), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6098), .ZN(n4360) );
  OAI21_X1 U5456 ( .B1(n6108), .B2(n4361), .A(n4360), .ZN(n4362) );
  AOI211_X1 U5457 ( .C1(n5135), .C2(n6082), .A(n4363), .B(n4362), .ZN(n4366)
         );
  NAND2_X1 U5458 ( .A1(n5126), .A2(n6087), .ZN(n4365) );
  NAND3_X1 U5459 ( .A1(n4366), .A2(n4365), .A3(n3108), .ZN(U2797) );
  NAND2_X1 U5460 ( .A1(n4369), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4368) );
  INV_X1 U5461 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U5462 ( .A1(n5689), .A2(n6628), .ZN(n5172) );
  INV_X1 U5463 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4382) );
  NAND4_X1 U5464 ( .A1(n5172), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n4382), .ZN(n4367) );
  INV_X1 U5465 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U5466 ( .A1(n5686), .A2(n6752), .ZN(n5625) );
  INV_X1 U5467 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5786) );
  XNOR2_X1 U5468 ( .A(n5686), .B(n5169), .ZN(n5611) );
  AOI21_X1 U5469 ( .B1(n4368), .B2(n4367), .A(n5609), .ZN(n4376) );
  NOR2_X1 U5470 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5171)
         );
  NAND2_X1 U5471 ( .A1(n5171), .A2(n4369), .ZN(n4373) );
  OAI21_X1 U5472 ( .B1(n4373), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n4370), 
        .ZN(n4371) );
  NAND3_X1 U5473 ( .A1(n5686), .A2(n5181), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5474 ( .A1(n4374), .A2(n3113), .ZN(n4375) );
  AOI21_X1 U5475 ( .B1(n4379), .B2(n4377), .A(n4378), .ZN(n5490) );
  NAND2_X1 U5476 ( .A1(n6194), .A2(REIP_REG_24__SCAN_IN), .ZN(n5602) );
  INV_X1 U5477 ( .A(n5602), .ZN(n4384) );
  INV_X1 U5478 ( .A(n4380), .ZN(n4393) );
  AOI211_X1 U5479 ( .C1(n4382), .C2(n4393), .A(n4381), .B(n5754), .ZN(n4383)
         );
  AOI211_X1 U5480 ( .C1(n5490), .C2(n6289), .A(n4384), .B(n4383), .ZN(n4385)
         );
  NOR2_X1 U5481 ( .A1(n5689), .A2(n4387), .ZN(n4388) );
  XNOR2_X1 U5482 ( .A(n4390), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4400)
         );
  NAND2_X1 U5483 ( .A1(n4400), .A2(n6294), .ZN(n4399) );
  OAI21_X1 U5484 ( .B1(n4391), .B2(n4392), .A(n4377), .ZN(n5492) );
  INV_X1 U5485 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6557) );
  NOR2_X1 U5486 ( .A1(n6211), .A2(n6557), .ZN(n4406) );
  NOR2_X1 U5487 ( .A1(n4393), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4394)
         );
  AOI211_X1 U5488 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n4395), .A(n4406), .B(n4394), .ZN(n4396) );
  NAND2_X1 U5489 ( .A1(n4399), .A2(n4398), .ZN(U2995) );
  NAND2_X1 U5490 ( .A1(n4400), .A2(n6219), .ZN(n4410) );
  NOR2_X1 U5491 ( .A1(n4402), .A2(n4403), .ZN(n4404) );
  NOR2_X1 U5492 ( .A1(n5266), .A2(n6223), .ZN(n4405) );
  AOI211_X1 U5493 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4406), 
        .B(n4405), .ZN(n4407) );
  NAND2_X1 U5494 ( .A1(n4410), .A2(n4409), .ZN(U2963) );
  INV_X1 U5495 ( .A(n4411), .ZN(n4413) );
  NAND3_X1 U5496 ( .A1(n4413), .A2(n4412), .A3(n4567), .ZN(n4414) );
  INV_X1 U5497 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4418) );
  OR2_X1 U5498 ( .A1(n5517), .A2(n4418), .ZN(n4419) );
  NAND2_X1 U5499 ( .A1(n5441), .A2(n4465), .ZN(n6084) );
  INV_X1 U5500 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6538) );
  NOR3_X1 U5501 ( .A1(n4424), .A2(n4423), .A3(n6538), .ZN(n4435) );
  OAI22_X1 U5502 ( .A1(n6093), .A2(n5518), .B1(n6648), .B2(n6068), .ZN(n4434)
         );
  NAND2_X1 U5503 ( .A1(n4425), .A2(n4426), .ZN(n4427) );
  NAND2_X1 U5504 ( .A1(n5404), .A2(n4427), .ZN(n5865) );
  NOR2_X1 U5505 ( .A1(n4428), .A2(n3119), .ZN(n6189) );
  NAND4_X1 U5506 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n6064), .A4(n6538), .ZN(n4431) );
  OAI211_X1 U5507 ( .C1(n5865), .C2(n6101), .A(n4432), .B(n4431), .ZN(n4433)
         );
  INV_X1 U5508 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4457) );
  INV_X1 U5509 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4450) );
  NOR2_X1 U5510 ( .A1(n4449), .A2(n4450), .ZN(n4442) );
  AND2_X1 U5511 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4451) );
  NAND2_X1 U5512 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4436) );
  OAI21_X1 U5513 ( .B1(n4442), .B2(n4451), .A(n4436), .ZN(n4437) );
  OAI211_X1 U5514 ( .C1(n6591), .C2(n4457), .A(n4437), .B(n4492), .ZN(U3182)
         );
  AOI221_X1 U5515 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6591), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4438) );
  AOI221_X1 U5516 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4438), .C2(HOLD), .A(n4449), .ZN(n4445) );
  AND2_X1 U5517 ( .A1(n4441), .A2(n4449), .ZN(n4440) );
  INV_X1 U5518 ( .A(NA_N), .ZN(n4443) );
  NAND2_X1 U5519 ( .A1(n4443), .A2(STATE_REG_2__SCAN_IN), .ZN(n4439) );
  AND2_X1 U5520 ( .A1(n4440), .A2(n4439), .ZN(n4452) );
  AOI22_X1 U5521 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4456) );
  INV_X1 U5522 ( .A(n4441), .ZN(n4455) );
  AOI21_X1 U5523 ( .B1(n4443), .B2(n4442), .A(n4455), .ZN(n4444) );
  OAI22_X1 U5524 ( .A1(n4445), .A2(n4452), .B1(n4456), .B2(n4444), .ZN(U3183)
         );
  NAND3_X1 U5525 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .A3(n6591), .ZN(n4446) );
  NAND2_X1 U5526 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4619), .ZN(n4700) );
  INV_X1 U5527 ( .A(n4700), .ZN(n4483) );
  AOI21_X1 U5528 ( .B1(n5034), .B2(n4446), .A(n4483), .ZN(n4448) );
  OR2_X1 U5529 ( .A1(n4448), .A2(n4447), .ZN(U3150) );
  OAI21_X1 U5530 ( .B1(n4451), .B2(n4450), .A(n6606), .ZN(n4454) );
  INV_X1 U5531 ( .A(n4452), .ZN(n4453) );
  OAI211_X1 U5532 ( .C1(n4456), .C2(n4455), .A(n4454), .B(n4453), .ZN(U3181)
         );
  INV_X1 U5533 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4459) );
  OAI21_X1 U5534 ( .B1(n4457), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4458) );
  OAI21_X1 U5535 ( .B1(n6546), .B2(n4459), .A(n6522), .ZN(U2789) );
  INV_X1 U5536 ( .A(n4680), .ZN(n4765) );
  AOI22_X1 U5537 ( .A1(n4765), .A2(n5428), .B1(n3977), .B2(n4460), .ZN(n4688)
         );
  INV_X1 U5538 ( .A(n4688), .ZN(n4461) );
  OAI21_X1 U5539 ( .B1(n4461), .B2(n4772), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4463) );
  NAND3_X1 U5540 ( .A1(n5191), .A2(STATE2_REG_0__SCAN_IN), .A3(n5034), .ZN(
        n4462) );
  NAND2_X1 U5541 ( .A1(n4463), .A2(n4462), .ZN(U2790) );
  NOR2_X1 U5542 ( .A1(n4498), .A2(n4465), .ZN(n4470) );
  INV_X1 U5543 ( .A(n4466), .ZN(n4472) );
  NOR2_X1 U5544 ( .A1(n4472), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4469) );
  NOR2_X1 U5545 ( .A1(n4467), .A2(n4499), .ZN(n4687) );
  INV_X1 U5546 ( .A(n4687), .ZN(n4468) );
  AOI22_X1 U5547 ( .A1(n4470), .A2(n4469), .B1(n6597), .B2(n4468), .ZN(U3474)
         );
  INV_X1 U5548 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4471) );
  OAI21_X1 U5549 ( .B1(n4472), .B2(n4471), .A(n4470), .ZN(U2788) );
  MUX2_X1 U5550 ( .A(n4681), .B(n4527), .S(n4680), .Z(n4482) );
  NAND2_X1 U5551 ( .A1(n4000), .A2(n4492), .ZN(n4473) );
  NAND2_X1 U5552 ( .A1(n4473), .A2(n6591), .ZN(n4474) );
  AOI21_X1 U5553 ( .B1(n4662), .B2(n4130), .A(n4474), .ZN(n4480) );
  INV_X1 U5554 ( .A(n4475), .ZN(n4478) );
  OR2_X1 U5555 ( .A1(n5445), .A2(n3221), .ZN(n4476) );
  OAI211_X1 U5556 ( .C1(n2953), .C2(n4478), .A(n4477), .B(n4476), .ZN(n4479)
         );
  AOI21_X1 U5557 ( .B1(n4680), .B2(n4480), .A(n4479), .ZN(n4481) );
  OR2_X1 U5558 ( .A1(n4666), .A2(n4772), .ZN(n4485) );
  NAND2_X1 U5559 ( .A1(n4483), .A2(FLUSH_REG_SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5560 ( .A1(n4485), .A2(n4484), .ZN(n4489) );
  NOR2_X1 U5561 ( .A1(n6733), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4486) );
  INV_X1 U5562 ( .A(n2953), .ZN(n4604) );
  INV_X1 U5563 ( .A(n4937), .ZN(n4989) );
  OR2_X1 U5564 ( .A1(n4487), .A2(n4989), .ZN(n4488) );
  XNOR2_X1 U5565 ( .A(n4488), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6090)
         );
  NAND4_X1 U5566 ( .A1(n4489), .A2(n4604), .A3(n5191), .A4(n6090), .ZN(n4490)
         );
  OAI21_X1 U5567 ( .B1(n5902), .B2(n4491), .A(n4490), .ZN(U3455) );
  INV_X1 U5568 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5569 ( .A1(n4561), .A2(EAX_REG_8__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4494) );
  OAI21_X1 U5570 ( .B1(n4560), .B2(n4495), .A(n4494), .ZN(U2915) );
  INV_X1 U5571 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4497) );
  AOI22_X1 U5572 ( .A1(n4561), .A2(EAX_REG_2__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4496) );
  OAI21_X1 U5573 ( .B1(n4560), .B2(n4497), .A(n4496), .ZN(U2921) );
  INV_X1 U5574 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6616) );
  INV_X1 U5575 ( .A(DATAI_8_), .ZN(n4501) );
  NOR2_X1 U5576 ( .A1(n6611), .A2(n4501), .ZN(n6139) );
  AOI21_X1 U5577 ( .B1(n6607), .B2(EAX_REG_8__SCAN_IN), .A(n6139), .ZN(n4502)
         );
  OAI21_X1 U5578 ( .B1(n6130), .B2(n6616), .A(n4502), .ZN(U2947) );
  INV_X1 U5579 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6737) );
  INV_X1 U5580 ( .A(DATAI_10_), .ZN(n4503) );
  NOR2_X1 U5581 ( .A1(n6611), .A2(n4503), .ZN(n6170) );
  AOI21_X1 U5582 ( .B1(n6607), .B2(EAX_REG_26__SCAN_IN), .A(n6170), .ZN(n4504)
         );
  OAI21_X1 U5583 ( .B1(n6737), .B2(n6130), .A(n4504), .ZN(U2934) );
  INV_X1 U5584 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6751) );
  INV_X1 U5585 ( .A(DATAI_11_), .ZN(n4505) );
  NOR2_X1 U5586 ( .A1(n6611), .A2(n4505), .ZN(n6144) );
  AOI21_X1 U5587 ( .B1(n6607), .B2(EAX_REG_11__SCAN_IN), .A(n6144), .ZN(n4506)
         );
  OAI21_X1 U5588 ( .B1(n6751), .B2(n6130), .A(n4506), .ZN(U2950) );
  INV_X1 U5589 ( .A(n4507), .ZN(n4520) );
  NAND2_X1 U5590 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5197) );
  INV_X1 U5591 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4508) );
  OAI22_X1 U5592 ( .A1(n6297), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4508), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4535) );
  NOR2_X1 U5593 ( .A1(n4509), .A2(n4510), .ZN(n4518) );
  NOR2_X1 U5594 ( .A1(n4662), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4517)
         );
  NAND4_X1 U5595 ( .A1(n2953), .A2(n4130), .A3(n4513), .A4(n4512), .ZN(n4515)
         );
  NOR2_X1 U5596 ( .A1(n4515), .A2(n4514), .ZN(n4664) );
  NOR2_X1 U5597 ( .A1(n4511), .A2(n4664), .ZN(n4516) );
  AOI211_X1 U5598 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4516), .ZN(n4667)
         );
  OAI222_X1 U5599 ( .A1(n5899), .A2(n4520), .B1(n5197), .B2(n4535), .C1(n6514), 
        .C2(n4667), .ZN(n4521) );
  NAND2_X1 U5600 ( .A1(n4521), .A2(n5902), .ZN(n4524) );
  INV_X1 U5601 ( .A(n5899), .ZN(n5196) );
  AOI22_X1 U5602 ( .A1(n5200), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n4522), .B2(n5196), .ZN(n4523) );
  NAND2_X1 U5603 ( .A1(n4524), .A2(n4523), .ZN(U3460) );
  INV_X1 U5604 ( .A(n4510), .ZN(n4537) );
  AOI21_X1 U5605 ( .B1(n5196), .B2(n4537), .A(n5200), .ZN(n4542) );
  INV_X1 U5606 ( .A(n4664), .ZN(n4581) );
  XNOR2_X1 U5607 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U5608 ( .A1(n4527), .A2(n4681), .ZN(n4590) );
  XNOR2_X1 U5609 ( .A(n4510), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4528)
         );
  NAND2_X1 U5610 ( .A1(n4590), .A2(n4528), .ZN(n4532) );
  INV_X1 U5611 ( .A(n4596), .ZN(n4530) );
  INV_X1 U5612 ( .A(n4528), .ZN(n4529) );
  NAND2_X1 U5613 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  OAI211_X1 U5614 ( .C1(n4533), .C2(n4662), .A(n4532), .B(n4531), .ZN(n4534)
         );
  AOI21_X1 U5615 ( .B1(n4526), .B2(n4581), .A(n4534), .ZN(n4602) );
  INV_X1 U5616 ( .A(n4602), .ZN(n4540) );
  INV_X1 U5617 ( .A(n4535), .ZN(n4536) );
  NOR2_X1 U5618 ( .A1(n5197), .A2(n4536), .ZN(n4539) );
  NOR3_X1 U5619 ( .A1(n5899), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4537), 
        .ZN(n4538) );
  AOI211_X1 U5620 ( .C1(n4540), .C2(n5191), .A(n4539), .B(n4538), .ZN(n4541)
         );
  OAI22_X1 U5621 ( .A1(n4542), .A2(n3068), .B1(n5200), .B2(n4541), .ZN(U3459)
         );
  XNOR2_X1 U5622 ( .A(n4544), .B(n4543), .ZN(n5482) );
  XOR2_X1 U5623 ( .A(n4545), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4550) );
  NAND2_X1 U5624 ( .A1(n4550), .A2(n6219), .ZN(n4549) );
  OR2_X1 U5625 ( .A1(n6212), .A2(n4546), .ZN(n4547) );
  AOI22_X1 U5626 ( .A1(n4547), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6194), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4548) );
  OAI211_X1 U5627 ( .C1(n5482), .C2(n5732), .A(n4549), .B(n4548), .ZN(U2986)
         );
  INV_X1 U5628 ( .A(n4550), .ZN(n4559) );
  NOR2_X1 U5629 ( .A1(n4551), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4553)
         );
  OR2_X1 U5630 ( .A1(n4553), .A2(n4552), .ZN(n5476) );
  INV_X1 U5631 ( .A(n5476), .ZN(n4557) );
  INV_X1 U5632 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U5633 ( .A1(n5867), .A2(n4554), .ZN(n5842) );
  NAND2_X1 U5634 ( .A1(n4281), .A2(n5842), .ZN(n4571) );
  OAI21_X1 U5635 ( .B1(n6211), .B2(n6585), .A(n4571), .ZN(n4556) );
  AOI21_X1 U5636 ( .B1(n5840), .B2(n4572), .A(n4281), .ZN(n4555) );
  AOI211_X1 U5637 ( .C1(n4557), .C2(n6289), .A(n4556), .B(n4555), .ZN(n4558)
         );
  OAI21_X1 U5638 ( .B1(n4559), .B2(n5882), .A(n4558), .ZN(U3018) );
  AOI222_X1 U5639 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6592), .B1(n6127), .B2(
        DATAO_REG_11__SCAN_IN), .C1(EAX_REG_11__SCAN_IN), .C2(n4561), .ZN(
        n4562) );
  INV_X1 U5640 ( .A(n4562), .ZN(U2912) );
  OAI21_X1 U5641 ( .B1(n4565), .B2(n4564), .A(n4563), .ZN(n5474) );
  XNOR2_X1 U5642 ( .A(n4566), .B(n4567), .ZN(n5465) );
  AOI22_X1 U5643 ( .A1(n5514), .A2(n5465), .B1(n5504), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4568) );
  OAI21_X1 U5644 ( .B1(n5474), .B2(n5516), .A(n4568), .ZN(U2858) );
  OAI222_X1 U5645 ( .A1(n5476), .A2(n5519), .B1(n5517), .B2(n5475), .C1(n5516), 
        .C2(n5482), .ZN(U2859) );
  XNOR2_X1 U5646 ( .A(n4570), .B(n4569), .ZN(n4627) );
  INV_X1 U5647 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U5648 ( .A1(n6211), .A2(n6578), .ZN(n4577) );
  NAND2_X1 U5649 ( .A1(n4572), .A2(n4571), .ZN(n4575) );
  AND2_X1 U5650 ( .A1(n5819), .A2(n4573), .ZN(n4574) );
  MUX2_X1 U5651 ( .A(n4575), .B(n4574), .S(n6297), .Z(n4576) );
  AOI211_X1 U5652 ( .C1(n6289), .C2(n5465), .A(n4577), .B(n4576), .ZN(n4578)
         );
  OAI21_X1 U5653 ( .B1(n4627), .B2(n5882), .A(n4578), .ZN(U3017) );
  INV_X1 U5654 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6126) );
  OAI222_X1 U5655 ( .A1(n5474), .A2(n5567), .B1(n5562), .B2(n6156), .C1(n5560), 
        .C2(n6126), .ZN(U2890) );
  INV_X1 U5656 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6030) );
  NAND2_X1 U5657 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6030), .ZN(n4611) );
  INV_X1 U5658 ( .A(n4579), .ZN(n4610) );
  NAND2_X1 U5659 ( .A1(n6347), .A2(n4581), .ZN(n4599) );
  INV_X1 U5660 ( .A(n4582), .ZN(n4583) );
  OAI21_X1 U5661 ( .B1(n4510), .B2(n4584), .A(n4583), .ZN(n4586) );
  NOR2_X1 U5662 ( .A1(n4586), .A2(n4585), .ZN(n5900) );
  MUX2_X1 U5663 ( .A(n4587), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4510), 
        .Z(n4588) );
  NOR2_X1 U5664 ( .A1(n4588), .A2(n4579), .ZN(n4589) );
  NAND2_X1 U5665 ( .A1(n4590), .A2(n4589), .ZN(n4595) );
  NAND2_X1 U5666 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4592) );
  INV_X1 U5667 ( .A(n4592), .ZN(n4591) );
  MUX2_X1 U5668 ( .A(n4592), .B(n4591), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4593) );
  OR2_X1 U5669 ( .A1(n4662), .A2(n4593), .ZN(n4594) );
  OAI211_X1 U5670 ( .C1(n5900), .C2(n4596), .A(n4595), .B(n4594), .ZN(n4597)
         );
  INV_X1 U5671 ( .A(n4597), .ZN(n4598) );
  NAND2_X1 U5672 ( .A1(n4599), .A2(n4598), .ZN(n5898) );
  INV_X1 U5673 ( .A(n4666), .ZN(n4601) );
  AND2_X1 U5674 ( .A1(n4666), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4600)
         );
  AOI21_X1 U5675 ( .B1(n5898), .B2(n4601), .A(n4600), .ZN(n4674) );
  INV_X1 U5676 ( .A(n4674), .ZN(n4675) );
  MUX2_X1 U5677 ( .A(n4602), .B(n3068), .S(n4666), .Z(n4673) );
  INV_X1 U5678 ( .A(n4673), .ZN(n4603) );
  NAND3_X1 U5679 ( .A1(n4675), .A2(n5194), .A3(n4603), .ZN(n4609) );
  NAND3_X1 U5680 ( .A1(n6090), .A2(n4604), .A3(n5194), .ZN(n4608) );
  NAND2_X1 U5681 ( .A1(n4666), .A2(n5194), .ZN(n4605) );
  NAND2_X1 U5682 ( .A1(n4605), .A2(n4611), .ZN(n4606) );
  NAND2_X1 U5683 ( .A1(n4606), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4607) );
  OAI211_X1 U5684 ( .C1(n4611), .C2(n4610), .A(n4609), .B(n4612), .ZN(n4692)
         );
  NAND2_X1 U5685 ( .A1(n4612), .A2(n4509), .ZN(n4613) );
  NAND2_X1 U5686 ( .A1(n4692), .A2(n4613), .ZN(n4620) );
  AOI21_X1 U5687 ( .B1(n4620), .B2(n6030), .A(n4700), .ZN(n4618) );
  INV_X1 U5688 ( .A(n6601), .ZN(n4615) );
  NAND2_X1 U5689 ( .A1(n4615), .A2(n4614), .ZN(n4616) );
  INV_X1 U5690 ( .A(n5033), .ZN(n4990) );
  AND2_X1 U5691 ( .A1(n4620), .A2(n4619), .ZN(n4768) );
  AND2_X1 U5692 ( .A1(n6733), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5895) );
  OAI22_X1 U5693 ( .A1(n2955), .A2(n6593), .B1(n5895), .B2(n3373), .ZN(n4621)
         );
  OAI21_X1 U5694 ( .B1(n4768), .B2(n4621), .A(n6302), .ZN(n4622) );
  OAI21_X1 U5695 ( .B1(n6302), .B2(n6390), .A(n4622), .ZN(U3465) );
  INV_X1 U5696 ( .A(n5474), .ZN(n4625) );
  INV_X1 U5697 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U5698 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6194), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4623) );
  OAI21_X1 U5699 ( .B1(n6223), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4623), 
        .ZN(n4624) );
  AOI21_X1 U5700 ( .B1(n4625), .B2(n6217), .A(n4624), .ZN(n4626) );
  OAI21_X1 U5701 ( .B1(n4627), .B2(n6192), .A(n4626), .ZN(U2985) );
  AOI222_X1 U5702 ( .A1(EAX_REG_30__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_30__SCAN_IN), .C1(n6592), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4628) );
  INV_X1 U5703 ( .A(n4628), .ZN(U2893) );
  AOI222_X1 U5704 ( .A1(EAX_REG_16__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_16__SCAN_IN), .C1(n4636), .C2(UWORD_REG_0__SCAN_IN), .ZN(
        n4629) );
  INV_X1 U5705 ( .A(n4629), .ZN(U2907) );
  AOI222_X1 U5706 ( .A1(EAX_REG_23__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_23__SCAN_IN), .C1(n4636), .C2(UWORD_REG_7__SCAN_IN), .ZN(
        n4630) );
  INV_X1 U5707 ( .A(n4630), .ZN(U2900) );
  AOI222_X1 U5708 ( .A1(EAX_REG_24__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_24__SCAN_IN), .C1(n4636), .C2(UWORD_REG_8__SCAN_IN), .ZN(
        n4631) );
  INV_X1 U5709 ( .A(n4631), .ZN(U2899) );
  AOI222_X1 U5710 ( .A1(EAX_REG_25__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_25__SCAN_IN), .C1(n4636), .C2(UWORD_REG_9__SCAN_IN), .ZN(
        n4632) );
  INV_X1 U5711 ( .A(n4632), .ZN(U2898) );
  AOI222_X1 U5712 ( .A1(EAX_REG_22__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_22__SCAN_IN), .C1(n6592), .C2(UWORD_REG_6__SCAN_IN), .ZN(
        n4633) );
  INV_X1 U5713 ( .A(n4633), .ZN(U2901) );
  AOI222_X1 U5714 ( .A1(EAX_REG_27__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n4636), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4634) );
  INV_X1 U5715 ( .A(n4634), .ZN(U2896) );
  AOI222_X1 U5716 ( .A1(EAX_REG_28__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_28__SCAN_IN), .C1(n6592), .C2(UWORD_REG_12__SCAN_IN), .ZN(
        n4635) );
  INV_X1 U5717 ( .A(n4635), .ZN(U2895) );
  AOI222_X1 U5718 ( .A1(EAX_REG_29__SCAN_IN), .A2(n4660), .B1(n6127), .B2(
        DATAO_REG_29__SCAN_IN), .C1(n4636), .C2(UWORD_REG_13__SCAN_IN), .ZN(
        n4637) );
  INV_X1 U5719 ( .A(n4637), .ZN(U2894) );
  INV_X1 U5720 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6731) );
  OAI222_X1 U5721 ( .A1(n5567), .A2(n5482), .B1(n5560), .B2(n6731), .C1(n6154), 
        .C2(n5562), .ZN(U2891) );
  INV_X1 U5722 ( .A(n4638), .ZN(n4641) );
  OAI21_X1 U5723 ( .B1(n4641), .B2(n4640), .A(n4639), .ZN(n6216) );
  OR2_X1 U5724 ( .A1(n4644), .A2(n4643), .ZN(n4645) );
  AND2_X1 U5725 ( .A1(n4642), .A2(n4645), .ZN(n6288) );
  AOI22_X1 U5726 ( .A1(n5514), .A2(n6288), .B1(n5504), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4646) );
  OAI21_X1 U5727 ( .B1(n6216), .B2(n5499), .A(n4646), .ZN(U2857) );
  AOI22_X1 U5728 ( .A1(n5565), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n5564), .ZN(n4647) );
  OAI21_X1 U5729 ( .B1(n6216), .B2(n5567), .A(n4647), .ZN(U2889) );
  AOI222_X1 U5730 ( .A1(n6127), .A2(DATAO_REG_20__SCAN_IN), .B1(n4660), .B2(
        EAX_REG_20__SCAN_IN), .C1(n6592), .C2(UWORD_REG_4__SCAN_IN), .ZN(n4648) );
  INV_X1 U5731 ( .A(n4648), .ZN(U2903) );
  INV_X1 U5732 ( .A(n4660), .ZN(n4659) );
  INV_X1 U5733 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5734 ( .A1(n6127), .A2(DATAO_REG_18__SCAN_IN), .ZN(n4650) );
  NAND2_X1 U5735 ( .A1(n6592), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4649) );
  OAI211_X1 U5736 ( .C1(n4659), .C2(n4651), .A(n4650), .B(n4649), .ZN(U2905)
         );
  NAND2_X1 U5737 ( .A1(n6127), .A2(DATAO_REG_19__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U5738 ( .A1(n6592), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4652) );
  OAI211_X1 U5739 ( .C1(n4659), .C2(n3691), .A(n4653), .B(n4652), .ZN(U2904)
         );
  NAND2_X1 U5740 ( .A1(n6127), .A2(DATAO_REG_21__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U5741 ( .A1(n6592), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4654) );
  OAI211_X1 U5742 ( .C1(n4659), .C2(n3725), .A(n4655), .B(n4654), .ZN(U2902)
         );
  INV_X1 U5743 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4658) );
  NAND2_X1 U5744 ( .A1(n6127), .A2(DATAO_REG_17__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5745 ( .A1(n6592), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4656) );
  OAI211_X1 U5746 ( .C1(n4659), .C2(n4658), .A(n4657), .B(n4656), .ZN(U2906)
         );
  AOI222_X1 U5747 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6592), .B1(n6127), .B2(
        DATAO_REG_26__SCAN_IN), .C1(EAX_REG_26__SCAN_IN), .C2(n4660), .ZN(
        n4661) );
  INV_X1 U5748 ( .A(n4661), .ZN(U2897) );
  INV_X1 U5749 ( .A(n4662), .ZN(n5192) );
  OAI22_X1 U5750 ( .A1(n3373), .A2(n4664), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4663), .ZN(n5193) );
  AOI211_X1 U5751 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n5192), .A(n6390), .B(n5193), .ZN(n4665) );
  INV_X1 U5752 ( .A(n4665), .ZN(n4670) );
  OAI22_X1 U5753 ( .A1(n4667), .A2(n4666), .B1(n4665), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5754 ( .A1(n4673), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4668) );
  OAI211_X1 U5755 ( .C1(n4671), .C2(n4670), .A(n4669), .B(n4668), .ZN(n4672)
         );
  OAI21_X1 U5756 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4673), .A(n4672), 
        .ZN(n4677) );
  NAND2_X1 U5757 ( .A1(n4674), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5758 ( .A1(n4677), .A2(n4676), .B1(n6312), .B2(n4675), .ZN(n4694)
         );
  INV_X1 U5759 ( .A(n4678), .ZN(n4685) );
  AND2_X1 U5760 ( .A1(n4679), .A2(n3977), .ZN(n4682) );
  MUX2_X1 U5761 ( .A(n4682), .B(n4681), .S(n4680), .Z(n4683) );
  OAI21_X1 U5762 ( .B1(n4685), .B2(n4684), .A(n4683), .ZN(n6590) );
  OAI21_X1 U5763 ( .B1(n4687), .B2(n4686), .A(n6591), .ZN(n6598) );
  NAND2_X1 U5764 ( .A1(n4688), .A2(n6598), .ZN(n6029) );
  NOR2_X1 U5765 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n4690) );
  OAI21_X1 U5766 ( .B1(n6029), .B2(n4690), .A(n4689), .ZN(n4691) );
  NOR3_X1 U5767 ( .A1(n4692), .A2(n6590), .A3(n4691), .ZN(n4693) );
  OAI21_X1 U5768 ( .B1(n4694), .B2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n4693), 
        .ZN(n4762) );
  NAND2_X1 U5769 ( .A1(n4762), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U5770 ( .A1(n6592), .A2(READY_N), .ZN(n4695) );
  NAND2_X1 U5771 ( .A1(n4772), .A2(n4695), .ZN(n4763) );
  OAI211_X1 U5772 ( .C1(n4698), .C2(n4697), .A(n4696), .B(n4763), .ZN(n6515)
         );
  INV_X1 U5773 ( .A(n6515), .ZN(n4699) );
  OAI21_X1 U5774 ( .B1(n4699), .B2(n6513), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4701) );
  NAND2_X1 U5775 ( .A1(n4701), .A2(n4700), .ZN(U3453) );
  AND2_X1 U5776 ( .A1(n4639), .A2(n4702), .ZN(n4704) );
  OR2_X1 U5777 ( .A1(n4704), .A2(n4703), .ZN(n5455) );
  NAND2_X1 U5778 ( .A1(n4642), .A2(n4706), .ZN(n4707) );
  AND2_X1 U5779 ( .A1(n4705), .A2(n4707), .ZN(n6279) );
  AOI22_X1 U5780 ( .A1(n5514), .A2(n6279), .B1(n5504), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4708) );
  OAI21_X1 U5781 ( .B1(n5455), .B2(n5516), .A(n4708), .ZN(U2856) );
  INV_X1 U5782 ( .A(DATAI_3_), .ZN(n6160) );
  INV_X1 U5783 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6124) );
  OAI222_X1 U5784 ( .A1(n5455), .A2(n5567), .B1(n5562), .B2(n6160), .C1(n5560), 
        .C2(n6124), .ZN(U2888) );
  AND2_X1 U5785 ( .A1(n5884), .A2(n4709), .ZN(n4710) );
  NAND2_X1 U5786 ( .A1(n4899), .A2(n4710), .ZN(n4711) );
  NAND2_X1 U5787 ( .A1(n6217), .A2(DATAI_29_), .ZN(n6492) );
  AND2_X1 U5788 ( .A1(n4711), .A2(n6217), .ZN(n4713) );
  INV_X1 U5789 ( .A(n4511), .ZN(n4846) );
  INV_X1 U5790 ( .A(n4744), .ZN(n4712) );
  AOI21_X1 U5791 ( .B1(n4847), .B2(n5039), .A(n4712), .ZN(n4716) );
  OAI21_X1 U5792 ( .B1(n4713), .B2(n6394), .A(n4716), .ZN(n4714) );
  NAND2_X1 U5793 ( .A1(n4742), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4720)
         );
  INV_X1 U5794 ( .A(n6487), .ZN(n6370) );
  NOR2_X1 U5795 ( .A1(n6304), .A2(n3415), .ZN(n4715) );
  INV_X1 U5796 ( .A(n4716), .ZN(n4717) );
  AOI22_X1 U5797 ( .A1(n4717), .A2(n6442), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5032), .ZN(n4745) );
  INV_X1 U5798 ( .A(DATAI_5_), .ZN(n6164) );
  OAI22_X1 U5799 ( .A1(n4745), .A2(n6013), .B1(n4744), .B2(n6486), .ZN(n4718)
         );
  AOI21_X1 U5800 ( .B1(n6370), .B2(n5936), .A(n4718), .ZN(n4719) );
  OAI211_X1 U5801 ( .C1(n5038), .C2(n6492), .A(n4720), .B(n4719), .ZN(U3145)
         );
  NAND2_X1 U5802 ( .A1(n6217), .A2(DATAI_26_), .ZN(n6471) );
  NAND2_X1 U5803 ( .A1(n4742), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4724)
         );
  INV_X1 U5804 ( .A(DATAI_2_), .ZN(n6158) );
  OAI22_X1 U5805 ( .A1(n4745), .A2(n6001), .B1(n4744), .B2(n6465), .ZN(n4722)
         );
  AOI21_X1 U5806 ( .B1(n6361), .B2(n5936), .A(n4722), .ZN(n4723) );
  OAI211_X1 U5807 ( .C1(n5038), .C2(n6471), .A(n4724), .B(n4723), .ZN(U3142)
         );
  NAND2_X1 U5808 ( .A1(n6217), .A2(DATAI_27_), .ZN(n6473) );
  NAND2_X1 U5809 ( .A1(n4742), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4728)
         );
  INV_X1 U5810 ( .A(n6478), .ZN(n6364) );
  OR2_X1 U5811 ( .A1(n4743), .A2(n4725), .ZN(n6472) );
  OAI22_X1 U5812 ( .A1(n4745), .A2(n6005), .B1(n4744), .B2(n6472), .ZN(n4726)
         );
  AOI21_X1 U5813 ( .B1(n6364), .B2(n5936), .A(n4726), .ZN(n4727) );
  OAI211_X1 U5814 ( .C1(n5038), .C2(n6473), .A(n4728), .B(n4727), .ZN(U3143)
         );
  NAND2_X1 U5815 ( .A1(n6217), .A2(DATAI_31_), .ZN(n6511) );
  NAND2_X1 U5816 ( .A1(n4742), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4731)
         );
  INV_X1 U5817 ( .A(n6502), .ZN(n6379) );
  INV_X1 U5818 ( .A(DATAI_7_), .ZN(n6610) );
  OAI22_X1 U5819 ( .A1(n4745), .A2(n6024), .B1(n4744), .B2(n6501), .ZN(n4729)
         );
  AOI21_X1 U5820 ( .B1(n6379), .B2(n5936), .A(n4729), .ZN(n4730) );
  OAI211_X1 U5821 ( .C1(n5038), .C2(n6511), .A(n4731), .B(n4730), .ZN(U3147)
         );
  NAND2_X1 U5822 ( .A1(n6217), .A2(DATAI_25_), .ZN(n6464) );
  NAND2_X1 U5823 ( .A1(n4742), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4734)
         );
  INV_X1 U5824 ( .A(n6459), .ZN(n6358) );
  OAI22_X1 U5825 ( .A1(n4745), .A2(n5997), .B1(n4744), .B2(n6458), .ZN(n4732)
         );
  AOI21_X1 U5826 ( .B1(n6358), .B2(n5936), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5827 ( .C1(n5038), .C2(n6464), .A(n4734), .B(n4733), .ZN(U3141)
         );
  NAND2_X1 U5828 ( .A1(n6217), .A2(DATAI_24_), .ZN(n6440) );
  NAND2_X1 U5829 ( .A1(n4742), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4738)
         );
  INV_X1 U5830 ( .A(n6457), .ZN(n6355) );
  OR2_X1 U5831 ( .A1(n4743), .A2(n4735), .ZN(n6439) );
  OAI22_X1 U5832 ( .A1(n4745), .A2(n5993), .B1(n4744), .B2(n6439), .ZN(n4736)
         );
  AOI21_X1 U5833 ( .B1(n6355), .B2(n5936), .A(n4736), .ZN(n4737) );
  OAI211_X1 U5834 ( .C1(n5038), .C2(n6440), .A(n4738), .B(n4737), .ZN(U3140)
         );
  NAND2_X1 U5835 ( .A1(n6217), .A2(DATAI_30_), .ZN(n6494) );
  NAND2_X1 U5836 ( .A1(n4742), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4741)
         );
  INV_X1 U5837 ( .A(DATAI_6_), .ZN(n6166) );
  OAI22_X1 U5838 ( .A1(n4745), .A2(n6017), .B1(n4744), .B2(n6493), .ZN(n4739)
         );
  AOI21_X1 U5839 ( .B1(n6373), .B2(n5936), .A(n4739), .ZN(n4740) );
  OAI211_X1 U5840 ( .C1(n5038), .C2(n6494), .A(n4741), .B(n4740), .ZN(U3146)
         );
  NAND2_X1 U5841 ( .A1(n4742), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4748)
         );
  INV_X1 U5842 ( .A(n6485), .ZN(n6367) );
  INV_X1 U5843 ( .A(DATAI_4_), .ZN(n6162) );
  OAI22_X1 U5844 ( .A1(n4745), .A2(n6009), .B1(n4744), .B2(n6479), .ZN(n4746)
         );
  AOI21_X1 U5845 ( .B1(n6367), .B2(n5936), .A(n4746), .ZN(n4747) );
  OAI211_X1 U5846 ( .C1(n5038), .C2(n6480), .A(n4748), .B(n4747), .ZN(U3144)
         );
  NAND2_X1 U5847 ( .A1(n4703), .A2(n4749), .ZN(n4882) );
  OR2_X1 U5848 ( .A1(n4703), .A2(n4749), .ZN(n4750) );
  INV_X1 U5849 ( .A(n6207), .ZN(n4754) );
  AOI21_X1 U5850 ( .B1(n4752), .B2(n4705), .A(n4751), .ZN(n6271) );
  AOI22_X1 U5851 ( .A1(n6271), .A2(n5514), .B1(n5504), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4753) );
  OAI21_X1 U5852 ( .B1(n4754), .B2(n5499), .A(n4753), .ZN(U2855) );
  INV_X1 U5853 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6122) );
  OAI222_X1 U5854 ( .A1(n4754), .A2(n5567), .B1(n5562), .B2(n6162), .C1(n6122), 
        .C2(n5560), .ZN(U2887) );
  OAI21_X1 U5855 ( .B1(n4755), .B2(n4757), .A(n4756), .ZN(n4758) );
  INV_X1 U5856 ( .A(n4758), .ZN(n6281) );
  NAND2_X1 U5857 ( .A1(n6281), .A2(n6219), .ZN(n4761) );
  INV_X1 U5858 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U5859 ( .A1(n6211), .A2(n5444), .ZN(n6278) );
  NOR2_X1 U5860 ( .A1(n6223), .A2(n5450), .ZN(n4759) );
  AOI211_X1 U5861 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6278), 
        .B(n4759), .ZN(n4760) );
  OAI211_X1 U5862 ( .C1(n5732), .C2(n5455), .A(n4761), .B(n4760), .ZN(U2983)
         );
  INV_X1 U5863 ( .A(n4762), .ZN(n4773) );
  INV_X1 U5864 ( .A(n4763), .ZN(n4764) );
  OAI21_X1 U5865 ( .B1(n4765), .B2(n4766), .A(n4764), .ZN(n4770) );
  OAI21_X1 U5866 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6591), .A(n6515), .ZN(
        n6512) );
  INV_X1 U5867 ( .A(n4766), .ZN(n4767) );
  NOR3_X1 U5868 ( .A1(n6512), .A2(n4768), .A3(n4767), .ZN(n4769) );
  MUX2_X1 U5869 ( .A(n4770), .B(n4769), .S(STATE2_REG_0__SCAN_IN), .Z(n4771)
         );
  OAI21_X1 U5870 ( .B1(n4773), .B2(n4772), .A(n4771), .ZN(U3148) );
  NOR2_X1 U5871 ( .A1(n4936), .A2(n6443), .ZN(n5893) );
  NOR2_X1 U5872 ( .A1(n5893), .A2(n6593), .ZN(n4780) );
  INV_X1 U5873 ( .A(n4802), .ZN(n4774) );
  AOI21_X1 U5874 ( .B1(n6400), .B2(n6446), .A(n4774), .ZN(n4779) );
  INV_X1 U5875 ( .A(n4779), .ZN(n4775) );
  INV_X1 U5876 ( .A(n6473), .ZN(n6415) );
  NAND2_X1 U5877 ( .A1(n5884), .A2(n2955), .ZN(n5979) );
  INV_X1 U5878 ( .A(n5979), .ZN(n4776) );
  OAI22_X1 U5879 ( .A1(n4803), .A2(n6478), .B1(n4802), .B2(n6472), .ZN(n4778)
         );
  AOI21_X1 U5880 ( .B1(n6415), .B2(n6393), .A(n4778), .ZN(n4783) );
  NAND2_X1 U5881 ( .A1(n4780), .A2(n4779), .ZN(n4781) );
  NAND2_X1 U5882 ( .A1(n4805), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4782) );
  OAI211_X1 U5883 ( .C1(n4808), .C2(n6005), .A(n4783), .B(n4782), .ZN(U3079)
         );
  INV_X1 U5884 ( .A(n6492), .ZN(n6423) );
  OAI22_X1 U5885 ( .A1(n4803), .A2(n6487), .B1(n4802), .B2(n6486), .ZN(n4784)
         );
  AOI21_X1 U5886 ( .B1(n6423), .B2(n6393), .A(n4784), .ZN(n4786) );
  NAND2_X1 U5887 ( .A1(n4805), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4785) );
  OAI211_X1 U5888 ( .C1(n4808), .C2(n6013), .A(n4786), .B(n4785), .ZN(U3081)
         );
  INV_X1 U5889 ( .A(n6494), .ZN(n6427) );
  OAI22_X1 U5890 ( .A1(n4803), .A2(n6499), .B1(n4802), .B2(n6493), .ZN(n4787)
         );
  AOI21_X1 U5891 ( .B1(n6427), .B2(n6393), .A(n4787), .ZN(n4789) );
  NAND2_X1 U5892 ( .A1(n4805), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4788) );
  OAI211_X1 U5893 ( .C1(n4808), .C2(n6017), .A(n4789), .B(n4788), .ZN(U3082)
         );
  OAI22_X1 U5894 ( .A1(n4803), .A2(n6457), .B1(n4802), .B2(n6439), .ZN(n4790)
         );
  AOI21_X1 U5895 ( .B1(n6403), .B2(n6393), .A(n4790), .ZN(n4792) );
  NAND2_X1 U5896 ( .A1(n4805), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4791) );
  OAI211_X1 U5897 ( .C1(n4808), .C2(n5993), .A(n4792), .B(n4791), .ZN(U3076)
         );
  INV_X1 U5898 ( .A(n6464), .ZN(n6407) );
  OAI22_X1 U5899 ( .A1(n4803), .A2(n6459), .B1(n4802), .B2(n6458), .ZN(n4793)
         );
  AOI21_X1 U5900 ( .B1(n6407), .B2(n6393), .A(n4793), .ZN(n4795) );
  NAND2_X1 U5901 ( .A1(n4805), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4794) );
  OAI211_X1 U5902 ( .C1(n4808), .C2(n5997), .A(n4795), .B(n4794), .ZN(U3077)
         );
  OAI22_X1 U5903 ( .A1(n4803), .A2(n6466), .B1(n4802), .B2(n6465), .ZN(n4796)
         );
  AOI21_X1 U5904 ( .B1(n6411), .B2(n6393), .A(n4796), .ZN(n4798) );
  NAND2_X1 U5905 ( .A1(n4805), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4797) );
  OAI211_X1 U5906 ( .C1(n4808), .C2(n6001), .A(n4798), .B(n4797), .ZN(U3078)
         );
  OAI22_X1 U5907 ( .A1(n4803), .A2(n6485), .B1(n4802), .B2(n6479), .ZN(n4799)
         );
  AOI21_X1 U5908 ( .B1(n6419), .B2(n6393), .A(n4799), .ZN(n4801) );
  NAND2_X1 U5909 ( .A1(n4805), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4800) );
  OAI211_X1 U5910 ( .C1(n4808), .C2(n6009), .A(n4801), .B(n4800), .ZN(U3080)
         );
  OAI22_X1 U5911 ( .A1(n4803), .A2(n6502), .B1(n4802), .B2(n6501), .ZN(n4804)
         );
  AOI21_X1 U5912 ( .B1(n6434), .B2(n6393), .A(n4804), .ZN(n4807) );
  NAND2_X1 U5913 ( .A1(n4805), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4806) );
  OAI211_X1 U5914 ( .C1(n4808), .C2(n6024), .A(n4807), .B(n4806), .ZN(U3083)
         );
  NOR2_X1 U5915 ( .A1(n5884), .A2(n3415), .ZN(n4809) );
  NAND2_X1 U5916 ( .A1(n4899), .A2(n4809), .ZN(n4813) );
  NOR2_X1 U5917 ( .A1(n4938), .A2(n6312), .ZN(n4991) );
  NOR2_X1 U5918 ( .A1(n4813), .A2(n6028), .ZN(n5891) );
  INV_X1 U5919 ( .A(n5891), .ZN(n4811) );
  NAND2_X1 U5920 ( .A1(n4526), .A2(n4511), .ZN(n6346) );
  INV_X1 U5921 ( .A(n6346), .ZN(n4998) );
  INV_X1 U5922 ( .A(n4991), .ZN(n4810) );
  NOR2_X1 U5923 ( .A1(n4810), .A2(n6390), .ZN(n4817) );
  AOI21_X1 U5924 ( .B1(n4847), .B2(n4998), .A(n4817), .ZN(n4815) );
  NAND3_X1 U5925 ( .A1(n4811), .A2(n6442), .A3(n4815), .ZN(n4812) );
  NAND2_X1 U5926 ( .A1(n4839), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4820)
         );
  NAND2_X1 U5927 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4814) );
  OAI22_X1 U5928 ( .A1(n4815), .A2(n6593), .B1(n4814), .B2(n4938), .ZN(n4816)
         );
  INV_X1 U5929 ( .A(n4817), .ZN(n4840) );
  OAI22_X1 U5930 ( .A1(n4841), .A2(n6024), .B1(n6501), .B2(n4840), .ZN(n4818)
         );
  AOI21_X1 U5931 ( .B1(n6379), .B2(n4843), .A(n4818), .ZN(n4819) );
  OAI211_X1 U5932 ( .C1(n4995), .C2(n6511), .A(n4820), .B(n4819), .ZN(U3131)
         );
  NAND2_X1 U5933 ( .A1(n4839), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4823)
         );
  OAI22_X1 U5934 ( .A1(n4841), .A2(n6005), .B1(n6472), .B2(n4840), .ZN(n4821)
         );
  AOI21_X1 U5935 ( .B1(n6364), .B2(n4843), .A(n4821), .ZN(n4822) );
  OAI211_X1 U5936 ( .C1(n4995), .C2(n6473), .A(n4823), .B(n4822), .ZN(U3127)
         );
  NAND2_X1 U5937 ( .A1(n4839), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4826)
         );
  OAI22_X1 U5938 ( .A1(n4841), .A2(n5997), .B1(n6458), .B2(n4840), .ZN(n4824)
         );
  AOI21_X1 U5939 ( .B1(n6358), .B2(n4843), .A(n4824), .ZN(n4825) );
  OAI211_X1 U5940 ( .C1(n4995), .C2(n6464), .A(n4826), .B(n4825), .ZN(U3125)
         );
  NAND2_X1 U5941 ( .A1(n4839), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4829)
         );
  OAI22_X1 U5942 ( .A1(n4841), .A2(n6017), .B1(n6493), .B2(n4840), .ZN(n4827)
         );
  AOI21_X1 U5943 ( .B1(n6373), .B2(n4843), .A(n4827), .ZN(n4828) );
  OAI211_X1 U5944 ( .C1(n4995), .C2(n6494), .A(n4829), .B(n4828), .ZN(U3130)
         );
  NAND2_X1 U5945 ( .A1(n4839), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4832)
         );
  OAI22_X1 U5946 ( .A1(n4841), .A2(n6009), .B1(n6479), .B2(n4840), .ZN(n4830)
         );
  AOI21_X1 U5947 ( .B1(n6367), .B2(n4843), .A(n4830), .ZN(n4831) );
  OAI211_X1 U5948 ( .C1(n4995), .C2(n6480), .A(n4832), .B(n4831), .ZN(U3128)
         );
  NAND2_X1 U5949 ( .A1(n4839), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4835)
         );
  OAI22_X1 U5950 ( .A1(n4841), .A2(n6001), .B1(n6465), .B2(n4840), .ZN(n4833)
         );
  AOI21_X1 U5951 ( .B1(n6361), .B2(n4843), .A(n4833), .ZN(n4834) );
  OAI211_X1 U5952 ( .C1(n4995), .C2(n6471), .A(n4835), .B(n4834), .ZN(U3126)
         );
  NAND2_X1 U5953 ( .A1(n4839), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4838)
         );
  OAI22_X1 U5954 ( .A1(n4841), .A2(n5993), .B1(n6439), .B2(n4840), .ZN(n4836)
         );
  AOI21_X1 U5955 ( .B1(n6355), .B2(n4843), .A(n4836), .ZN(n4837) );
  OAI211_X1 U5956 ( .C1(n4995), .C2(n6440), .A(n4838), .B(n4837), .ZN(U3124)
         );
  NAND2_X1 U5957 ( .A1(n4839), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4845)
         );
  OAI22_X1 U5958 ( .A1(n4841), .A2(n6013), .B1(n6486), .B2(n4840), .ZN(n4842)
         );
  AOI21_X1 U5959 ( .B1(n6370), .B2(n4843), .A(n4842), .ZN(n4844) );
  OAI211_X1 U5960 ( .C1(n4995), .C2(n6492), .A(n4845), .B(n4844), .ZN(U3129)
         );
  INV_X1 U5961 ( .A(n4899), .ZN(n5887) );
  OAI21_X1 U5962 ( .B1(n4849), .B2(n6593), .A(n5896), .ZN(n4853) );
  INV_X1 U5963 ( .A(n5941), .ZN(n5948) );
  NOR2_X1 U5964 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4901) );
  AND2_X1 U5965 ( .A1(n4901), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5943)
         );
  AND2_X1 U5966 ( .A1(n5943), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4850)
         );
  AOI21_X1 U5967 ( .B1(n4847), .B2(n5948), .A(n4850), .ZN(n4852) );
  INV_X1 U5968 ( .A(n4852), .ZN(n4848) );
  AND2_X1 U5969 ( .A1(n4849), .A2(n2955), .ZN(n5940) );
  INV_X1 U5970 ( .A(n4850), .ZN(n4875) );
  OAI22_X1 U5971 ( .A1(n5984), .A2(n6457), .B1(n6439), .B2(n4875), .ZN(n4851)
         );
  AOI21_X1 U5972 ( .B1(n6403), .B2(n5940), .A(n4851), .ZN(n4856) );
  NAND2_X1 U5973 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  NAND2_X1 U5974 ( .A1(n4877), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4855) );
  OAI211_X1 U5975 ( .C1(n4880), .C2(n5993), .A(n4856), .B(n4855), .ZN(U3092)
         );
  OAI22_X1 U5976 ( .A1(n5984), .A2(n6459), .B1(n6458), .B2(n4875), .ZN(n4857)
         );
  AOI21_X1 U5977 ( .B1(n6407), .B2(n5940), .A(n4857), .ZN(n4859) );
  NAND2_X1 U5978 ( .A1(n4877), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4858) );
  OAI211_X1 U5979 ( .C1(n4880), .C2(n5997), .A(n4859), .B(n4858), .ZN(U3093)
         );
  OAI22_X1 U5980 ( .A1(n5984), .A2(n6502), .B1(n6501), .B2(n4875), .ZN(n4860)
         );
  AOI21_X1 U5981 ( .B1(n6434), .B2(n5940), .A(n4860), .ZN(n4862) );
  NAND2_X1 U5982 ( .A1(n4877), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4861) );
  OAI211_X1 U5983 ( .C1(n4880), .C2(n6024), .A(n4862), .B(n4861), .ZN(U3099)
         );
  OAI22_X1 U5984 ( .A1(n5984), .A2(n6466), .B1(n6465), .B2(n4875), .ZN(n4863)
         );
  AOI21_X1 U5985 ( .B1(n6411), .B2(n5940), .A(n4863), .ZN(n4865) );
  NAND2_X1 U5986 ( .A1(n4877), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4864) );
  OAI211_X1 U5987 ( .C1(n4880), .C2(n6001), .A(n4865), .B(n4864), .ZN(U3094)
         );
  OAI22_X1 U5988 ( .A1(n5984), .A2(n6487), .B1(n6486), .B2(n4875), .ZN(n4866)
         );
  AOI21_X1 U5989 ( .B1(n6423), .B2(n5940), .A(n4866), .ZN(n4868) );
  NAND2_X1 U5990 ( .A1(n4877), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4867) );
  OAI211_X1 U5991 ( .C1(n4880), .C2(n6013), .A(n4868), .B(n4867), .ZN(U3097)
         );
  OAI22_X1 U5992 ( .A1(n5984), .A2(n6499), .B1(n6493), .B2(n4875), .ZN(n4869)
         );
  AOI21_X1 U5993 ( .B1(n6427), .B2(n5940), .A(n4869), .ZN(n4871) );
  NAND2_X1 U5994 ( .A1(n4877), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4870) );
  OAI211_X1 U5995 ( .C1(n4880), .C2(n6017), .A(n4871), .B(n4870), .ZN(U3098)
         );
  OAI22_X1 U5996 ( .A1(n5984), .A2(n6485), .B1(n6479), .B2(n4875), .ZN(n4872)
         );
  AOI21_X1 U5997 ( .B1(n6419), .B2(n5940), .A(n4872), .ZN(n4874) );
  NAND2_X1 U5998 ( .A1(n4877), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4873) );
  OAI211_X1 U5999 ( .C1(n4880), .C2(n6009), .A(n4874), .B(n4873), .ZN(U3096)
         );
  OAI22_X1 U6000 ( .A1(n5984), .A2(n6478), .B1(n6472), .B2(n4875), .ZN(n4876)
         );
  AOI21_X1 U6001 ( .B1(n6415), .B2(n5940), .A(n4876), .ZN(n4879) );
  NAND2_X1 U6002 ( .A1(n4877), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4878) );
  OAI211_X1 U6003 ( .C1(n4880), .C2(n6005), .A(n4879), .B(n4878), .ZN(U3095)
         );
  AOI21_X1 U6004 ( .B1(n4883), .B2(n4882), .A(n4892), .ZN(n5429) );
  NOR2_X1 U6005 ( .A1(n4751), .A2(n4885), .ZN(n4886) );
  OR2_X1 U6006 ( .A1(n4884), .A2(n4886), .ZN(n5430) );
  INV_X1 U6007 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4887) );
  OAI22_X1 U6008 ( .A1(n5430), .A2(n5519), .B1(n4887), .B2(n5517), .ZN(n4888)
         );
  AOI21_X1 U6009 ( .B1(n5429), .B2(n5521), .A(n4888), .ZN(n4889) );
  INV_X1 U6010 ( .A(n4889), .ZN(U2854) );
  INV_X1 U6011 ( .A(n5429), .ZN(n4890) );
  INV_X1 U6012 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6120) );
  OAI222_X1 U6013 ( .A1(n4890), .A2(n5567), .B1(n5562), .B2(n6164), .C1(n5560), 
        .C2(n6120), .ZN(U2886) );
  NAND2_X1 U6014 ( .A1(n4892), .A2(n4891), .ZN(n5028) );
  OAI21_X1 U6015 ( .B1(n4892), .B2(n4891), .A(n5028), .ZN(n6081) );
  AOI22_X1 U6016 ( .A1(n5565), .A2(DATAI_6_), .B1(EAX_REG_6__SCAN_IN), .B2(
        n5564), .ZN(n4893) );
  OAI21_X1 U6017 ( .B1(n6081), .B2(n5567), .A(n4893), .ZN(U2885) );
  NAND2_X1 U6018 ( .A1(n4895), .A2(n4896), .ZN(n4897) );
  NAND2_X1 U6019 ( .A1(n4894), .A2(n4897), .ZN(n5709) );
  AOI22_X1 U6020 ( .A1(n5565), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5564), .ZN(n4898) );
  OAI21_X1 U6021 ( .B1(n5709), .B2(n5567), .A(n4898), .ZN(U2882) );
  OAI21_X1 U6022 ( .B1(n4904), .B2(n6593), .A(n5896), .ZN(n4907) );
  AND2_X1 U6023 ( .A1(n4901), .A2(n6312), .ZN(n5906) );
  NAND2_X1 U6024 ( .A1(n5906), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4929) );
  INV_X1 U6025 ( .A(n4929), .ZN(n4902) );
  AOI21_X1 U6026 ( .B1(n5910), .B2(n6446), .A(n4902), .ZN(n4906) );
  INV_X1 U6027 ( .A(n4906), .ZN(n4903) );
  NAND2_X1 U6028 ( .A1(n4904), .A2(n2955), .ZN(n5939) );
  OAI22_X1 U6029 ( .A1(n5117), .A2(n6502), .B1(n6501), .B2(n4929), .ZN(n4905)
         );
  AOI21_X1 U6030 ( .B1(n6434), .B2(n4931), .A(n4905), .ZN(n4910) );
  NAND2_X1 U6031 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  NAND2_X1 U6032 ( .A1(n4932), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4909) );
  OAI211_X1 U6033 ( .C1(n4935), .C2(n6024), .A(n4910), .B(n4909), .ZN(U3035)
         );
  OAI22_X1 U6034 ( .A1(n5117), .A2(n6457), .B1(n6439), .B2(n4929), .ZN(n4911)
         );
  AOI21_X1 U6035 ( .B1(n6403), .B2(n4931), .A(n4911), .ZN(n4913) );
  NAND2_X1 U6036 ( .A1(n4932), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4912) );
  OAI211_X1 U6037 ( .C1(n4935), .C2(n5993), .A(n4913), .B(n4912), .ZN(U3028)
         );
  OAI22_X1 U6038 ( .A1(n5117), .A2(n6466), .B1(n6465), .B2(n4929), .ZN(n4914)
         );
  AOI21_X1 U6039 ( .B1(n6411), .B2(n4931), .A(n4914), .ZN(n4916) );
  NAND2_X1 U6040 ( .A1(n4932), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4915) );
  OAI211_X1 U6041 ( .C1(n4935), .C2(n6001), .A(n4916), .B(n4915), .ZN(U3030)
         );
  OAI22_X1 U6042 ( .A1(n5117), .A2(n6499), .B1(n6493), .B2(n4929), .ZN(n4917)
         );
  AOI21_X1 U6043 ( .B1(n6427), .B2(n4931), .A(n4917), .ZN(n4919) );
  NAND2_X1 U6044 ( .A1(n4932), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4918) );
  OAI211_X1 U6045 ( .C1(n4935), .C2(n6017), .A(n4919), .B(n4918), .ZN(U3034)
         );
  OAI22_X1 U6046 ( .A1(n5117), .A2(n6485), .B1(n6479), .B2(n4929), .ZN(n4920)
         );
  AOI21_X1 U6047 ( .B1(n6419), .B2(n4931), .A(n4920), .ZN(n4922) );
  NAND2_X1 U6048 ( .A1(n4932), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4921) );
  OAI211_X1 U6049 ( .C1(n4935), .C2(n6009), .A(n4922), .B(n4921), .ZN(U3032)
         );
  OAI22_X1 U6050 ( .A1(n5117), .A2(n6487), .B1(n6486), .B2(n4929), .ZN(n4923)
         );
  AOI21_X1 U6051 ( .B1(n6423), .B2(n4931), .A(n4923), .ZN(n4925) );
  NAND2_X1 U6052 ( .A1(n4932), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4924) );
  OAI211_X1 U6053 ( .C1(n4935), .C2(n6013), .A(n4925), .B(n4924), .ZN(U3033)
         );
  OAI22_X1 U6054 ( .A1(n5117), .A2(n6478), .B1(n6472), .B2(n4929), .ZN(n4926)
         );
  AOI21_X1 U6055 ( .B1(n6415), .B2(n4931), .A(n4926), .ZN(n4928) );
  NAND2_X1 U6056 ( .A1(n4932), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4927) );
  OAI211_X1 U6057 ( .C1(n4935), .C2(n6005), .A(n4928), .B(n4927), .ZN(U3031)
         );
  OAI22_X1 U6058 ( .A1(n5117), .A2(n6459), .B1(n6458), .B2(n4929), .ZN(n4930)
         );
  AOI21_X1 U6059 ( .B1(n6407), .B2(n4931), .A(n4930), .ZN(n4934) );
  NAND2_X1 U6060 ( .A1(n4932), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4933) );
  OAI211_X1 U6061 ( .C1(n4935), .C2(n5997), .A(n4934), .B(n4933), .ZN(U3029)
         );
  INV_X1 U6062 ( .A(n6354), .ZN(n4940) );
  OR2_X1 U6063 ( .A1(n6346), .A2(n4937), .ZN(n6349) );
  OR2_X1 U6064 ( .A1(n6349), .A2(n3373), .ZN(n4939) );
  NOR2_X1 U6065 ( .A1(n4938), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6348)
         );
  NAND2_X1 U6066 ( .A1(n6348), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6067 ( .A1(n4939), .A2(n4968), .ZN(n4947) );
  NOR2_X2 U6068 ( .A1(n4942), .A2(n4941), .ZN(n6378) );
  OR2_X1 U6069 ( .A1(n4942), .A2(n2955), .ZN(n6402) );
  OAI22_X1 U6070 ( .A1(n6402), .A2(n6459), .B1(n6458), .B2(n4968), .ZN(n4943)
         );
  AOI21_X1 U6071 ( .B1(n6407), .B2(n6378), .A(n4943), .ZN(n4949) );
  INV_X1 U6072 ( .A(n6348), .ZN(n4945) );
  INV_X1 U6073 ( .A(n4944), .ZN(n6310) );
  AOI21_X1 U6074 ( .B1(n6593), .B2(n4945), .A(n6310), .ZN(n4946) );
  NAND2_X1 U6075 ( .A1(n4970), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4948) );
  OAI211_X1 U6076 ( .C1(n4973), .C2(n5997), .A(n4949), .B(n4948), .ZN(U3061)
         );
  OAI22_X1 U6077 ( .A1(n6402), .A2(n6466), .B1(n6465), .B2(n4968), .ZN(n4950)
         );
  AOI21_X1 U6078 ( .B1(n6411), .B2(n6378), .A(n4950), .ZN(n4952) );
  NAND2_X1 U6079 ( .A1(n4970), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4951) );
  OAI211_X1 U6080 ( .C1(n4973), .C2(n6001), .A(n4952), .B(n4951), .ZN(U3062)
         );
  OAI22_X1 U6081 ( .A1(n6402), .A2(n6485), .B1(n6479), .B2(n4968), .ZN(n4953)
         );
  AOI21_X1 U6082 ( .B1(n6419), .B2(n6378), .A(n4953), .ZN(n4955) );
  NAND2_X1 U6083 ( .A1(n4970), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4954) );
  OAI211_X1 U6084 ( .C1(n4973), .C2(n6009), .A(n4955), .B(n4954), .ZN(U3064)
         );
  OAI22_X1 U6085 ( .A1(n6402), .A2(n6502), .B1(n6501), .B2(n4968), .ZN(n4956)
         );
  AOI21_X1 U6086 ( .B1(n6434), .B2(n6378), .A(n4956), .ZN(n4958) );
  NAND2_X1 U6087 ( .A1(n4970), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4957) );
  OAI211_X1 U6088 ( .C1(n4973), .C2(n6024), .A(n4958), .B(n4957), .ZN(U3067)
         );
  OAI22_X1 U6089 ( .A1(n6402), .A2(n6457), .B1(n6439), .B2(n4968), .ZN(n4959)
         );
  AOI21_X1 U6090 ( .B1(n6403), .B2(n6378), .A(n4959), .ZN(n4961) );
  NAND2_X1 U6091 ( .A1(n4970), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4960) );
  OAI211_X1 U6092 ( .C1(n4973), .C2(n5993), .A(n4961), .B(n4960), .ZN(U3060)
         );
  OAI22_X1 U6093 ( .A1(n6402), .A2(n6499), .B1(n6493), .B2(n4968), .ZN(n4962)
         );
  AOI21_X1 U6094 ( .B1(n6427), .B2(n6378), .A(n4962), .ZN(n4964) );
  NAND2_X1 U6095 ( .A1(n4970), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4963) );
  OAI211_X1 U6096 ( .C1(n4973), .C2(n6017), .A(n4964), .B(n4963), .ZN(U3066)
         );
  OAI22_X1 U6097 ( .A1(n6402), .A2(n6478), .B1(n6472), .B2(n4968), .ZN(n4965)
         );
  AOI21_X1 U6098 ( .B1(n6415), .B2(n6378), .A(n4965), .ZN(n4967) );
  NAND2_X1 U6099 ( .A1(n4970), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4966) );
  OAI211_X1 U6100 ( .C1(n4973), .C2(n6005), .A(n4967), .B(n4966), .ZN(U3063)
         );
  OAI22_X1 U6101 ( .A1(n6402), .A2(n6487), .B1(n6486), .B2(n4968), .ZN(n4969)
         );
  AOI21_X1 U6102 ( .B1(n6423), .B2(n6378), .A(n4969), .ZN(n4972) );
  NAND2_X1 U6103 ( .A1(n4970), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4971) );
  OAI211_X1 U6104 ( .C1(n4973), .C2(n6013), .A(n4972), .B(n4971), .ZN(U3065)
         );
  INV_X1 U6105 ( .A(n4974), .ZN(n4976) );
  INV_X1 U6106 ( .A(n4884), .ZN(n4975) );
  INV_X1 U6107 ( .A(n4980), .ZN(n4982) );
  AOI21_X1 U6108 ( .B1(n4976), .B2(n4975), .A(n4982), .ZN(n6262) );
  INV_X1 U6109 ( .A(n6262), .ZN(n4977) );
  INV_X1 U6110 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6741) );
  OAI222_X1 U6111 ( .A1(n4977), .A2(n5519), .B1(n5517), .B2(n6741), .C1(n5516), 
        .C2(n6081), .ZN(U2853) );
  INV_X1 U6112 ( .A(n4978), .ZN(n5027) );
  XNOR2_X1 U6113 ( .A(n5028), .B(n5027), .ZN(n5733) );
  INV_X1 U6114 ( .A(n4979), .ZN(n4981) );
  OR2_X1 U6115 ( .A1(n4980), .A2(n4979), .ZN(n5121) );
  OAI21_X1 U6116 ( .B1(n4982), .B2(n4981), .A(n5121), .ZN(n5419) );
  INV_X1 U6117 ( .A(n5419), .ZN(n6254) );
  AOI22_X1 U6118 ( .A1(n6254), .A2(n5514), .B1(n5504), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4983) );
  OAI21_X1 U6119 ( .B1(n5733), .B2(n5499), .A(n4983), .ZN(U2852) );
  AOI22_X1 U6120 ( .A1(n5565), .A2(DATAI_7_), .B1(EAX_REG_7__SCAN_IN), .B2(
        n5564), .ZN(n4984) );
  OAI21_X1 U6121 ( .B1(n5733), .B2(n5567), .A(n4984), .ZN(U2884) );
  INV_X1 U6122 ( .A(n4985), .ZN(n4988) );
  OR2_X1 U6123 ( .A1(n5121), .A2(n5122), .ZN(n5119) );
  NAND2_X1 U6124 ( .A1(n5119), .A2(n4986), .ZN(n4987) );
  NAND2_X1 U6125 ( .A1(n4988), .A2(n4987), .ZN(n5874) );
  OAI222_X1 U6126 ( .A1(n5874), .A2(n5519), .B1(n5517), .B2(n4013), .C1(n5516), 
        .C2(n5709), .ZN(U2850) );
  AOI21_X1 U6127 ( .B1(n6503), .B2(n4995), .A(n6028), .ZN(n4994) );
  OAI21_X1 U6128 ( .B1(n6346), .B2(n4989), .A(n6442), .ZN(n4993) );
  INV_X1 U6129 ( .A(n6344), .ZN(n4997) );
  INV_X1 U6130 ( .A(n6345), .ZN(n5088) );
  OAI21_X1 U6131 ( .B1(n5034), .B2(n5088), .A(n4990), .ZN(n5905) );
  AOI21_X1 U6132 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4997), .A(n5905), .ZN(
        n5945) );
  NAND2_X1 U6133 ( .A1(n4991), .A2(n6390), .ZN(n5021) );
  AOI21_X1 U6134 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5021), .A(n6396), .ZN(
        n4992) );
  NAND2_X1 U6135 ( .A1(n5020), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5001)
         );
  NOR2_X1 U6136 ( .A1(n6384), .A2(n6593), .ZN(n5949) );
  NAND2_X1 U6137 ( .A1(n4996), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6387) );
  NOR2_X1 U6138 ( .A1(n4997), .A2(n6345), .ZN(n5947) );
  AOI22_X1 U6139 ( .A1(n5949), .A2(n4998), .B1(n5988), .B2(n5947), .ZN(n5022)
         );
  OAI22_X1 U6140 ( .A1(n5022), .A2(n6024), .B1(n6501), .B2(n5021), .ZN(n4999)
         );
  AOI21_X1 U6141 ( .B1(n5024), .B2(n6379), .A(n4999), .ZN(n5000) );
  OAI211_X1 U6142 ( .C1(n6503), .C2(n6511), .A(n5001), .B(n5000), .ZN(U3123)
         );
  NAND2_X1 U6143 ( .A1(n5020), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5004)
         );
  OAI22_X1 U6144 ( .A1(n5022), .A2(n6001), .B1(n6465), .B2(n5021), .ZN(n5002)
         );
  AOI21_X1 U6145 ( .B1(n5024), .B2(n6361), .A(n5002), .ZN(n5003) );
  OAI211_X1 U6146 ( .C1(n6503), .C2(n6471), .A(n5004), .B(n5003), .ZN(U3118)
         );
  NAND2_X1 U6147 ( .A1(n5020), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5007)
         );
  OAI22_X1 U6148 ( .A1(n5022), .A2(n5997), .B1(n6458), .B2(n5021), .ZN(n5005)
         );
  AOI21_X1 U6149 ( .B1(n5024), .B2(n6358), .A(n5005), .ZN(n5006) );
  OAI211_X1 U6150 ( .C1(n6503), .C2(n6464), .A(n5007), .B(n5006), .ZN(U3117)
         );
  NAND2_X1 U6151 ( .A1(n5020), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5010)
         );
  OAI22_X1 U6152 ( .A1(n5022), .A2(n6005), .B1(n6472), .B2(n5021), .ZN(n5008)
         );
  AOI21_X1 U6153 ( .B1(n5024), .B2(n6364), .A(n5008), .ZN(n5009) );
  OAI211_X1 U6154 ( .C1(n6503), .C2(n6473), .A(n5010), .B(n5009), .ZN(U3119)
         );
  NAND2_X1 U6155 ( .A1(n5020), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5013)
         );
  OAI22_X1 U6156 ( .A1(n5022), .A2(n6009), .B1(n6479), .B2(n5021), .ZN(n5011)
         );
  AOI21_X1 U6157 ( .B1(n5024), .B2(n6367), .A(n5011), .ZN(n5012) );
  OAI211_X1 U6158 ( .C1(n6503), .C2(n6480), .A(n5013), .B(n5012), .ZN(U3120)
         );
  NAND2_X1 U6159 ( .A1(n5020), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5016)
         );
  OAI22_X1 U6160 ( .A1(n5022), .A2(n6013), .B1(n6486), .B2(n5021), .ZN(n5014)
         );
  AOI21_X1 U6161 ( .B1(n5024), .B2(n6370), .A(n5014), .ZN(n5015) );
  OAI211_X1 U6162 ( .C1(n6503), .C2(n6492), .A(n5016), .B(n5015), .ZN(U3121)
         );
  NAND2_X1 U6163 ( .A1(n5020), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5019)
         );
  OAI22_X1 U6164 ( .A1(n5022), .A2(n6017), .B1(n6493), .B2(n5021), .ZN(n5017)
         );
  AOI21_X1 U6165 ( .B1(n5024), .B2(n6373), .A(n5017), .ZN(n5018) );
  OAI211_X1 U6166 ( .C1(n6503), .C2(n6494), .A(n5019), .B(n5018), .ZN(U3122)
         );
  NAND2_X1 U6167 ( .A1(n5020), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5026)
         );
  OAI22_X1 U6168 ( .A1(n5022), .A2(n5993), .B1(n6439), .B2(n5021), .ZN(n5023)
         );
  AOI21_X1 U6169 ( .B1(n5024), .B2(n6355), .A(n5023), .ZN(n5025) );
  OAI211_X1 U6170 ( .C1(n6503), .C2(n6440), .A(n5026), .B(n5025), .ZN(U3116)
         );
  NOR2_X1 U6171 ( .A1(n5028), .A2(n5027), .ZN(n5030) );
  OAI21_X1 U6172 ( .B1(n5030), .B2(n5029), .A(n4895), .ZN(n6071) );
  AOI22_X1 U6173 ( .A1(n5565), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5564), .ZN(n5031) );
  OAI21_X1 U6174 ( .B1(n6071), .B2(n5567), .A(n5031), .ZN(U2883) );
  AOI21_X1 U6175 ( .B1(n5068), .B2(n5038), .A(n6028), .ZN(n5037) );
  INV_X1 U6176 ( .A(n5039), .ZN(n6388) );
  OAI21_X1 U6177 ( .B1(n6388), .B2(n6384), .A(n6442), .ZN(n5036) );
  NAND2_X1 U6178 ( .A1(n5032), .A2(n6390), .ZN(n5062) );
  AOI21_X1 U6179 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5088), .A(n5033), .ZN(
        n6399) );
  OAI21_X1 U6180 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5034), .A(n6399), 
        .ZN(n5987) );
  AOI211_X1 U6181 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5062), .A(n6396), .B(
        n5987), .ZN(n5035) );
  NAND2_X1 U6182 ( .A1(n5061), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5042)
         );
  NOR2_X1 U6183 ( .A1(n5088), .A2(n6312), .ZN(n5983) );
  AOI22_X1 U6184 ( .A1(n5949), .A2(n5039), .B1(n5988), .B2(n5983), .ZN(n5063)
         );
  OAI22_X1 U6185 ( .A1(n5063), .A2(n5997), .B1(n6458), .B2(n5062), .ZN(n5040)
         );
  AOI21_X1 U6186 ( .B1(n5065), .B2(n6358), .A(n5040), .ZN(n5041) );
  OAI211_X1 U6187 ( .C1(n5068), .C2(n6464), .A(n5042), .B(n5041), .ZN(U3133)
         );
  NAND2_X1 U6188 ( .A1(n5061), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5045)
         );
  OAI22_X1 U6189 ( .A1(n5063), .A2(n6009), .B1(n6479), .B2(n5062), .ZN(n5043)
         );
  AOI21_X1 U6190 ( .B1(n5065), .B2(n6367), .A(n5043), .ZN(n5044) );
  OAI211_X1 U6191 ( .C1(n5068), .C2(n6480), .A(n5045), .B(n5044), .ZN(U3136)
         );
  NAND2_X1 U6192 ( .A1(n5061), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5048)
         );
  OAI22_X1 U6193 ( .A1(n5063), .A2(n6005), .B1(n6472), .B2(n5062), .ZN(n5046)
         );
  AOI21_X1 U6194 ( .B1(n5065), .B2(n6364), .A(n5046), .ZN(n5047) );
  OAI211_X1 U6195 ( .C1(n5068), .C2(n6473), .A(n5048), .B(n5047), .ZN(U3135)
         );
  NAND2_X1 U6196 ( .A1(n5061), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5051)
         );
  OAI22_X1 U6197 ( .A1(n5063), .A2(n6001), .B1(n6465), .B2(n5062), .ZN(n5049)
         );
  AOI21_X1 U6198 ( .B1(n5065), .B2(n6361), .A(n5049), .ZN(n5050) );
  OAI211_X1 U6199 ( .C1(n5068), .C2(n6471), .A(n5051), .B(n5050), .ZN(U3134)
         );
  NAND2_X1 U6200 ( .A1(n5061), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5054)
         );
  OAI22_X1 U6201 ( .A1(n5063), .A2(n6024), .B1(n6501), .B2(n5062), .ZN(n5052)
         );
  AOI21_X1 U6202 ( .B1(n5065), .B2(n6379), .A(n5052), .ZN(n5053) );
  OAI211_X1 U6203 ( .C1(n5068), .C2(n6511), .A(n5054), .B(n5053), .ZN(U3139)
         );
  NAND2_X1 U6204 ( .A1(n5061), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5057)
         );
  OAI22_X1 U6205 ( .A1(n5063), .A2(n6017), .B1(n6493), .B2(n5062), .ZN(n5055)
         );
  AOI21_X1 U6206 ( .B1(n5065), .B2(n6373), .A(n5055), .ZN(n5056) );
  OAI211_X1 U6207 ( .C1(n5068), .C2(n6494), .A(n5057), .B(n5056), .ZN(U3138)
         );
  NAND2_X1 U6208 ( .A1(n5061), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5060)
         );
  OAI22_X1 U6209 ( .A1(n5063), .A2(n6013), .B1(n6486), .B2(n5062), .ZN(n5058)
         );
  AOI21_X1 U6210 ( .B1(n5065), .B2(n6370), .A(n5058), .ZN(n5059) );
  OAI211_X1 U6211 ( .C1(n5068), .C2(n6492), .A(n5060), .B(n5059), .ZN(U3137)
         );
  NAND2_X1 U6212 ( .A1(n5061), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5067)
         );
  OAI22_X1 U6213 ( .A1(n5063), .A2(n5993), .B1(n6439), .B2(n5062), .ZN(n5064)
         );
  AOI21_X1 U6214 ( .B1(n5065), .B2(n6355), .A(n5064), .ZN(n5066) );
  OAI211_X1 U6215 ( .C1(n5068), .C2(n6440), .A(n5067), .B(n5066), .ZN(U3132)
         );
  OAI21_X1 U6216 ( .B1(n5071), .B2(n5070), .A(n5069), .ZN(n5083) );
  INV_X1 U6217 ( .A(n5430), .ZN(n5077) );
  NOR2_X1 U6218 ( .A1(n6211), .A2(n6529), .ZN(n5080) );
  OAI21_X1 U6219 ( .B1(n5876), .B2(n5813), .A(n5866), .ZN(n6295) );
  AOI21_X1 U6220 ( .B1(n6263), .B2(n5819), .A(n6295), .ZN(n6269) );
  AOI21_X1 U6221 ( .B1(n6290), .B2(n5072), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n5075) );
  NAND2_X1 U6222 ( .A1(n5073), .A2(n6744), .ZN(n5074) );
  OAI22_X1 U6223 ( .A1(n6269), .A2(n5075), .B1(n6296), .B2(n5074), .ZN(n5076)
         );
  AOI211_X1 U6224 ( .C1(n6289), .C2(n5077), .A(n5080), .B(n5076), .ZN(n5078)
         );
  OAI21_X1 U6225 ( .B1(n5882), .B2(n5083), .A(n5078), .ZN(U3013) );
  NAND2_X1 U6226 ( .A1(n5429), .A2(n6217), .ZN(n5082) );
  NOR2_X1 U6227 ( .A1(n5727), .A2(n5431), .ZN(n5079) );
  AOI211_X1 U6228 ( .C1(n6188), .C2(n5433), .A(n5080), .B(n5079), .ZN(n5081)
         );
  OAI211_X1 U6229 ( .C1(n5083), .C2(n6192), .A(n5082), .B(n5081), .ZN(U2981)
         );
  OAI21_X1 U6230 ( .B1(n5084), .B2(n6339), .A(n5896), .ZN(n5085) );
  OR2_X1 U6231 ( .A1(n4526), .A2(n4511), .ZN(n5981) );
  AOI21_X1 U6232 ( .B1(n5085), .B2(n5087), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5086) );
  OR2_X1 U6233 ( .A1(n6311), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6314)
         );
  NOR2_X1 U6234 ( .A1(n6314), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5089)
         );
  NAND2_X1 U6235 ( .A1(n5111), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5092) );
  INV_X1 U6236 ( .A(n5087), .ZN(n6309) );
  NOR2_X1 U6237 ( .A1(n5088), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6385)
         );
  AOI22_X1 U6238 ( .A1(n6309), .A2(n6442), .B1(n6396), .B2(n6385), .ZN(n5113)
         );
  INV_X1 U6239 ( .A(n5089), .ZN(n5112) );
  OAI22_X1 U6240 ( .A1(n5113), .A2(n6024), .B1(n6501), .B2(n5112), .ZN(n5090)
         );
  AOI21_X1 U6241 ( .B1(n6339), .B2(n6379), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6242 ( .C1(n5117), .C2(n6511), .A(n5092), .B(n5091), .ZN(U3043)
         );
  NAND2_X1 U6243 ( .A1(n5111), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5095) );
  OAI22_X1 U6244 ( .A1(n5113), .A2(n6009), .B1(n6479), .B2(n5112), .ZN(n5093)
         );
  AOI21_X1 U6245 ( .B1(n6339), .B2(n6367), .A(n5093), .ZN(n5094) );
  OAI211_X1 U6246 ( .C1(n5117), .C2(n6480), .A(n5095), .B(n5094), .ZN(U3040)
         );
  NAND2_X1 U6247 ( .A1(n5111), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5098) );
  OAI22_X1 U6248 ( .A1(n5113), .A2(n5997), .B1(n6458), .B2(n5112), .ZN(n5096)
         );
  AOI21_X1 U6249 ( .B1(n6339), .B2(n6358), .A(n5096), .ZN(n5097) );
  OAI211_X1 U6250 ( .C1(n5117), .C2(n6464), .A(n5098), .B(n5097), .ZN(U3037)
         );
  NAND2_X1 U6251 ( .A1(n5111), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5101) );
  OAI22_X1 U6252 ( .A1(n5113), .A2(n5993), .B1(n6439), .B2(n5112), .ZN(n5099)
         );
  AOI21_X1 U6253 ( .B1(n6339), .B2(n6355), .A(n5099), .ZN(n5100) );
  OAI211_X1 U6254 ( .C1(n5117), .C2(n6440), .A(n5101), .B(n5100), .ZN(U3036)
         );
  NAND2_X1 U6255 ( .A1(n5111), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5104) );
  OAI22_X1 U6256 ( .A1(n5113), .A2(n6005), .B1(n6472), .B2(n5112), .ZN(n5102)
         );
  AOI21_X1 U6257 ( .B1(n6339), .B2(n6364), .A(n5102), .ZN(n5103) );
  OAI211_X1 U6258 ( .C1(n5117), .C2(n6473), .A(n5104), .B(n5103), .ZN(U3039)
         );
  NAND2_X1 U6259 ( .A1(n5111), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5107) );
  OAI22_X1 U6260 ( .A1(n5113), .A2(n6017), .B1(n6493), .B2(n5112), .ZN(n5105)
         );
  AOI21_X1 U6261 ( .B1(n6339), .B2(n6373), .A(n5105), .ZN(n5106) );
  OAI211_X1 U6262 ( .C1(n5117), .C2(n6494), .A(n5107), .B(n5106), .ZN(U3042)
         );
  NAND2_X1 U6263 ( .A1(n5111), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5110) );
  OAI22_X1 U6264 ( .A1(n5113), .A2(n6001), .B1(n6465), .B2(n5112), .ZN(n5108)
         );
  AOI21_X1 U6265 ( .B1(n6339), .B2(n6361), .A(n5108), .ZN(n5109) );
  OAI211_X1 U6266 ( .C1(n5117), .C2(n6471), .A(n5110), .B(n5109), .ZN(U3038)
         );
  NAND2_X1 U6267 ( .A1(n5111), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5116) );
  OAI22_X1 U6268 ( .A1(n5113), .A2(n6013), .B1(n6486), .B2(n5112), .ZN(n5114)
         );
  AOI21_X1 U6269 ( .B1(n6339), .B2(n6370), .A(n5114), .ZN(n5115) );
  OAI211_X1 U6270 ( .C1(n5117), .C2(n6492), .A(n5116), .B(n5115), .ZN(U3041)
         );
  OAI21_X1 U6271 ( .B1(n3539), .B2(n3120), .A(n4429), .ZN(n6060) );
  AOI22_X1 U6272 ( .A1(n5565), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5564), .ZN(n5118) );
  OAI21_X1 U6273 ( .B1(n6060), .B2(n5567), .A(n5118), .ZN(U2881) );
  INV_X1 U6274 ( .A(n5119), .ZN(n5120) );
  AOI21_X1 U6275 ( .B1(n5122), .B2(n5121), .A(n5120), .ZN(n6246) );
  INV_X1 U6276 ( .A(n6246), .ZN(n5123) );
  INV_X1 U6277 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6742) );
  OAI222_X1 U6278 ( .A1(n5123), .A2(n5519), .B1(n5517), .B2(n6742), .C1(n5516), 
        .C2(n6071), .ZN(U2851) );
  OAI21_X1 U6279 ( .B1(n4985), .B2(n5124), .A(n4425), .ZN(n6236) );
  INV_X1 U6280 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5125) );
  OAI222_X1 U6281 ( .A1(n6236), .A2(n5519), .B1(n5125), .B2(n5517), .C1(n6060), 
        .C2(n5516), .ZN(U2849) );
  AOI22_X1 U6282 ( .A1(n5554), .A2(DATAI_30_), .B1(n5564), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6283 ( .A1(n5555), .A2(DATAI_14_), .ZN(n5127) );
  OAI211_X1 U6284 ( .C1(n5129), .C2(n5567), .A(n5128), .B(n5127), .ZN(U2861)
         );
  NOR2_X1 U6285 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5134)
         );
  INV_X1 U6286 ( .A(n5745), .ZN(n5130) );
  AOI211_X1 U6287 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5738), .A(n5131), .B(n5130), .ZN(n5132) );
  AOI211_X1 U6288 ( .C1(n5734), .C2(n5134), .A(n5133), .B(n5132), .ZN(n5137)
         );
  NAND2_X1 U6289 ( .A1(n5135), .A2(n6289), .ZN(n5136) );
  OAI211_X1 U6290 ( .C1(n5138), .C2(n5882), .A(n5137), .B(n5136), .ZN(U2988)
         );
  INV_X1 U6291 ( .A(n5577), .ZN(n5140) );
  NAND2_X1 U6292 ( .A1(n5140), .A2(n5139), .ZN(n5144) );
  INV_X1 U6293 ( .A(n5587), .ZN(n5143) );
  NAND3_X1 U6294 ( .A1(n5141), .A2(n5143), .A3(n5142), .ZN(n5578) );
  XNOR2_X1 U6295 ( .A(n5145), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5163)
         );
  NAND2_X1 U6296 ( .A1(n5146), .A2(n5147), .ZN(n5148) );
  NAND2_X1 U6297 ( .A1(n4345), .A2(n5148), .ZN(n5486) );
  INV_X1 U6298 ( .A(n5486), .ZN(n5155) );
  NOR2_X1 U6299 ( .A1(n5149), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5749)
         );
  AOI21_X1 U6300 ( .B1(n5745), .B2(n5744), .A(n5749), .ZN(n5153) );
  INV_X1 U6301 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6302 ( .A1(n6194), .A2(REIP_REG_28__SCAN_IN), .ZN(n5160) );
  INV_X1 U6303 ( .A(n5149), .ZN(n5150) );
  NAND3_X1 U6304 ( .A1(n5150), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5152), .ZN(n5151) );
  OAI211_X1 U6305 ( .C1(n5153), .C2(n5152), .A(n5160), .B(n5151), .ZN(n5154)
         );
  AOI21_X1 U6306 ( .B1(n5155), .B2(n6289), .A(n5154), .ZN(n5156) );
  OAI21_X1 U6307 ( .B1(n5163), .B2(n5882), .A(n5156), .ZN(U2990) );
  NAND2_X1 U6308 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5159)
         );
  OAI211_X1 U6309 ( .C1(n5215), .C2(n6223), .A(n5160), .B(n5159), .ZN(n5161)
         );
  OAI21_X1 U6310 ( .B1(n5163), .B2(n6192), .A(n5162), .ZN(U2958) );
  AND2_X1 U6311 ( .A1(n5560), .A2(n5164), .ZN(n5165) );
  NAND2_X1 U6312 ( .A1(n5166), .A2(n5165), .ZN(n5168) );
  AOI22_X1 U6313 ( .A1(n5554), .A2(DATAI_31_), .B1(n5564), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6314 ( .A1(n5168), .A2(n5167), .ZN(U2860) );
  AOI21_X1 U6315 ( .B1(n5175), .B2(n5286), .A(n4402), .ZN(n5274) );
  INV_X1 U6316 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6555) );
  NOR2_X1 U6317 ( .A1(n6211), .A2(n6555), .ZN(n5183) );
  AOI21_X1 U6318 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5183), 
        .ZN(n5176) );
  OAI21_X1 U6319 ( .B1(n5276), .B2(n6223), .A(n5176), .ZN(n5177) );
  AOI21_X1 U6320 ( .B1(n5274), .B2(n6217), .A(n5177), .ZN(n5178) );
  OAI21_X1 U6321 ( .B1(n5190), .B2(n6192), .A(n5178), .ZN(U2964) );
  INV_X1 U6322 ( .A(n5179), .ZN(n5770) );
  NOR3_X1 U6323 ( .A1(n5773), .A2(n5181), .A3(n5180), .ZN(n5182) );
  AOI211_X1 U6324 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5770), .A(n5183), .B(n5182), .ZN(n5189) );
  INV_X1 U6325 ( .A(n5184), .ZN(n5187) );
  INV_X1 U6326 ( .A(n5185), .ZN(n5186) );
  AOI21_X1 U6327 ( .B1(n5187), .B2(n5186), .A(n4391), .ZN(n5494) );
  NAND2_X1 U6328 ( .A1(n5494), .A2(n6289), .ZN(n5188) );
  OAI211_X1 U6329 ( .C1(n5190), .C2(n5882), .A(n5189), .B(n5188), .ZN(U2996)
         );
  AOI21_X1 U6330 ( .B1(n5192), .B2(n5191), .A(n5200), .ZN(n5202) );
  INV_X1 U6331 ( .A(n5193), .ZN(n5195) );
  OAI21_X1 U6332 ( .B1(n5195), .B2(STATE2_REG_3__SCAN_IN), .A(n5194), .ZN(
        n5198) );
  AOI22_X1 U6333 ( .A1(n5198), .A2(n5197), .B1(n5196), .B2(n5201), .ZN(n5199)
         );
  OAI22_X1 U6334 ( .A1(n5202), .A2(n5201), .B1(n5200), .B2(n5199), .ZN(U3461)
         );
  OAI22_X1 U6335 ( .A1(n5204), .A2(n5519), .B1(n5203), .B2(n5517), .ZN(U2828)
         );
  AOI21_X1 U6336 ( .B1(n4345), .B2(n5206), .A(n5205), .ZN(n5740) );
  INV_X1 U6337 ( .A(n5571), .ZN(n5209) );
  NAND2_X1 U6338 ( .A1(n5218), .A2(REIP_REG_29__SCAN_IN), .ZN(n5208) );
  AOI22_X1 U6339 ( .A1(n5393), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6098), .ZN(n5207) );
  OAI211_X1 U6340 ( .C1(n6108), .C2(n5209), .A(n5208), .B(n5207), .ZN(n5210)
         );
  AOI211_X1 U6341 ( .C1(n5740), .C2(n6082), .A(n5211), .B(n5210), .ZN(n5212)
         );
  OAI21_X1 U6342 ( .B1(n5485), .B2(n6059), .A(n5212), .ZN(U2798) );
  AOI22_X1 U6343 ( .A1(n5393), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6098), .ZN(n5214) );
  OAI21_X1 U6344 ( .B1(n6108), .B2(n5215), .A(n5214), .ZN(n5217) );
  NOR2_X1 U6345 ( .A1(n5486), .A2(n6101), .ZN(n5216) );
  AOI211_X1 U6346 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5218), .A(n5217), .B(n5216), .ZN(n5221) );
  INV_X1 U6347 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5219) );
  NAND3_X1 U6348 ( .A1(n5230), .A2(REIP_REG_27__SCAN_IN), .A3(n5219), .ZN(
        n5220) );
  OAI211_X1 U6349 ( .C1(n5213), .C2(n6059), .A(n5221), .B(n5220), .ZN(U2799)
         );
  AOI21_X1 U6350 ( .B1(n5223), .B2(n5222), .A(n5157), .ZN(n5584) );
  INV_X1 U6351 ( .A(n5584), .ZN(n5527) );
  INV_X1 U6352 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6566) );
  AOI22_X1 U6353 ( .A1(n5393), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6098), .ZN(n5225) );
  NAND2_X1 U6354 ( .A1(n6073), .A2(n5580), .ZN(n5224) );
  OAI211_X1 U6355 ( .C1(n5238), .C2(n6566), .A(n5225), .B(n5224), .ZN(n5229)
         );
  OAI21_X1 U6356 ( .B1(n5234), .B2(n5227), .A(n5146), .ZN(n5743) );
  NOR2_X1 U6357 ( .A1(n5743), .A2(n6101), .ZN(n5228) );
  AOI211_X1 U6358 ( .C1(n5230), .C2(n6566), .A(n5229), .B(n5228), .ZN(n5231)
         );
  OAI21_X1 U6359 ( .B1(n5527), .B2(n6059), .A(n5231), .ZN(U2800) );
  OAI21_X1 U6360 ( .B1(n5232), .B2(n5233), .A(n5222), .ZN(n5593) );
  AOI21_X1 U6361 ( .B1(n5235), .B2(n5246), .A(n5234), .ZN(n5488) );
  AOI22_X1 U6362 ( .A1(n5393), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6098), .ZN(n5236) );
  OAI21_X1 U6363 ( .B1(n6108), .B2(n5589), .A(n5236), .ZN(n5241) );
  INV_X1 U6364 ( .A(n5237), .ZN(n5254) );
  AOI21_X1 U6365 ( .B1(n5254), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5239) );
  NOR2_X1 U6366 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  AOI211_X1 U6367 ( .C1(n5488), .C2(n6082), .A(n5241), .B(n5240), .ZN(n5242)
         );
  OAI21_X1 U6368 ( .B1(n5593), .B2(n6059), .A(n5242), .ZN(U2801) );
  AOI21_X1 U6369 ( .B1(n5244), .B2(n5243), .A(n5232), .ZN(n5245) );
  INV_X1 U6370 ( .A(n5245), .ZN(n5600) );
  INV_X1 U6371 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6561) );
  INV_X1 U6372 ( .A(n5597), .ZN(n5252) );
  INV_X1 U6373 ( .A(n5246), .ZN(n5247) );
  AOI21_X1 U6374 ( .B1(n5249), .B2(n5248), .A(n5247), .ZN(n5767) );
  NAND2_X1 U6375 ( .A1(n5767), .A2(n6082), .ZN(n5251) );
  AOI22_X1 U6376 ( .A1(n5393), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6098), .ZN(n5250) );
  OAI211_X1 U6377 ( .C1(n6108), .C2(n5252), .A(n5251), .B(n5250), .ZN(n5253)
         );
  AOI21_X1 U6378 ( .B1(n5254), .B2(n6561), .A(n5253), .ZN(n5257) );
  NOR3_X1 U6379 ( .A1(n5380), .A2(REIP_REG_24__SCAN_IN), .A3(n5255), .ZN(n5262) );
  OAI21_X1 U6380 ( .B1(n5262), .B2(n5259), .A(REIP_REG_25__SCAN_IN), .ZN(n5256) );
  OAI211_X1 U6381 ( .C1(n5600), .C2(n6059), .A(n5257), .B(n5256), .ZN(U2802)
         );
  XOR2_X1 U6382 ( .A(n5258), .B(n4401), .Z(n5606) );
  INV_X1 U6383 ( .A(n5606), .ZN(n5534) );
  INV_X1 U6384 ( .A(n5259), .ZN(n5268) );
  AOI22_X1 U6385 ( .A1(n5393), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6098), .ZN(n5261) );
  NAND2_X1 U6386 ( .A1(n6073), .A2(n5601), .ZN(n5260) );
  OAI211_X1 U6387 ( .C1(n5268), .C2(n6559), .A(n5261), .B(n5260), .ZN(n5263)
         );
  AOI211_X1 U6388 ( .C1(n5490), .C2(n6082), .A(n5263), .B(n5262), .ZN(n5264)
         );
  OAI21_X1 U6389 ( .B1(n5534), .B2(n6059), .A(n5264), .ZN(U2803) );
  INV_X1 U6390 ( .A(n5492), .ZN(n5272) );
  AOI22_X1 U6391 ( .A1(n5393), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6098), .ZN(n5265) );
  OAI21_X1 U6392 ( .B1(n6108), .B2(n5266), .A(n5265), .ZN(n5271) );
  INV_X1 U6393 ( .A(n5380), .ZN(n5369) );
  AOI21_X1 U6394 ( .B1(n5369), .B2(n5267), .A(REIP_REG_23__SCAN_IN), .ZN(n5269) );
  NOR2_X1 U6395 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  AOI211_X1 U6396 ( .C1(n6082), .C2(n5272), .A(n5271), .B(n5270), .ZN(n5273)
         );
  OAI21_X1 U6397 ( .B1(n5537), .B2(n6059), .A(n5273), .ZN(U2804) );
  INV_X1 U6398 ( .A(n5274), .ZN(n5540) );
  AOI22_X1 U6399 ( .A1(n5393), .A2(EBX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6098), .ZN(n5275) );
  OAI21_X1 U6400 ( .B1(n6108), .B2(n5276), .A(n5275), .ZN(n5278) );
  INV_X1 U6401 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5279) );
  NOR4_X1 U6402 ( .A1(n5380), .A2(REIP_REG_22__SCAN_IN), .A3(n5282), .A4(n5279), .ZN(n5277) );
  AOI211_X1 U6403 ( .C1(n6082), .C2(n5494), .A(n5278), .B(n5277), .ZN(n5285)
         );
  INV_X1 U6404 ( .A(n5282), .ZN(n5280) );
  NAND2_X1 U6405 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NOR2_X1 U6406 ( .A1(n5380), .A2(n5281), .ZN(n5296) );
  NAND2_X1 U6407 ( .A1(n5479), .A2(n5282), .ZN(n5283) );
  NAND2_X1 U6408 ( .A1(n5395), .A2(n5283), .ZN(n5309) );
  OAI21_X1 U6409 ( .B1(n5296), .B2(n5309), .A(REIP_REG_22__SCAN_IN), .ZN(n5284) );
  OAI211_X1 U6410 ( .C1(n5540), .C2(n6059), .A(n5285), .B(n5284), .ZN(U2805)
         );
  INV_X1 U6411 ( .A(n5286), .ZN(n5287) );
  AOI21_X1 U6412 ( .B1(n5288), .B2(n5299), .A(n5287), .ZN(n5616) );
  INV_X1 U6413 ( .A(n5616), .ZN(n5543) );
  AND2_X1 U6414 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  NOR2_X1 U6415 ( .A1(n5185), .A2(n5291), .ZN(n5775) );
  AND2_X1 U6416 ( .A1(n5309), .A2(REIP_REG_21__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6417 ( .A1(n6073), .A2(n5612), .ZN(n5293) );
  AOI22_X1 U6418 ( .A1(n5393), .A2(EBX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6098), .ZN(n5292) );
  NAND2_X1 U6419 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  AOI211_X1 U6420 ( .C1(n5775), .C2(n6082), .A(n5295), .B(n5294), .ZN(n5298)
         );
  INV_X1 U6421 ( .A(n5296), .ZN(n5297) );
  OAI211_X1 U6422 ( .C1(n5543), .C2(n6059), .A(n5298), .B(n5297), .ZN(U2806)
         );
  INV_X1 U6423 ( .A(n5299), .ZN(n5300) );
  AOI21_X1 U6424 ( .B1(n5301), .B2(n5174), .A(n5300), .ZN(n5623) );
  INV_X1 U6425 ( .A(n5623), .ZN(n5546) );
  MUX2_X1 U6426 ( .A(n5303), .B(n3991), .S(n5302), .Z(n5305) );
  XNOR2_X1 U6427 ( .A(n5305), .B(n5304), .ZN(n5788) );
  AOI22_X1 U6428 ( .A1(n5393), .A2(EBX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6098), .ZN(n5306) );
  OAI21_X1 U6429 ( .B1(n6108), .B2(n5621), .A(n5306), .ZN(n5307) );
  AOI21_X1 U6430 ( .B1(n5788), .B2(n6082), .A(n5307), .ZN(n5312) );
  NAND2_X1 U6431 ( .A1(n5369), .A2(n5324), .ZN(n5323) );
  NOR2_X1 U6432 ( .A1(n5323), .A2(n5308), .ZN(n5310) );
  OAI21_X1 U6433 ( .B1(n5310), .B2(REIP_REG_20__SCAN_IN), .A(n5309), .ZN(n5311) );
  OAI211_X1 U6434 ( .C1(n5546), .C2(n6059), .A(n5312), .B(n5311), .ZN(U2807)
         );
  OR2_X1 U6435 ( .A1(n5313), .A2(n5314), .ZN(n5315) );
  NAND2_X1 U6436 ( .A1(n5174), .A2(n5315), .ZN(n5630) );
  XNOR2_X1 U6437 ( .A(n5317), .B(n5316), .ZN(n5796) );
  INV_X1 U6438 ( .A(n5633), .ZN(n5320) );
  INV_X1 U6439 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5629) );
  OAI21_X1 U6440 ( .B1(n6068), .B2(n5629), .A(n6084), .ZN(n5318) );
  AOI21_X1 U6441 ( .B1(EBX_REG_19__SCAN_IN), .B2(n5393), .A(n5318), .ZN(n5319)
         );
  OAI21_X1 U6442 ( .B1(n6108), .B2(n5320), .A(n5319), .ZN(n5322) );
  NOR3_X1 U6443 ( .A1(n5323), .A2(REIP_REG_19__SCAN_IN), .A3(n6550), .ZN(n5321) );
  AOI211_X1 U6444 ( .C1(n5796), .C2(n6082), .A(n5322), .B(n5321), .ZN(n5328)
         );
  NOR2_X1 U6445 ( .A1(n5323), .A2(REIP_REG_18__SCAN_IN), .ZN(n5338) );
  INV_X1 U6446 ( .A(n5324), .ZN(n5325) );
  NAND2_X1 U6447 ( .A1(n5479), .A2(n5325), .ZN(n5326) );
  NAND2_X1 U6448 ( .A1(n5395), .A2(n5326), .ZN(n5352) );
  OAI21_X1 U6449 ( .B1(n5338), .B2(n5352), .A(REIP_REG_19__SCAN_IN), .ZN(n5327) );
  OAI211_X1 U6450 ( .C1(n5630), .C2(n6059), .A(n5328), .B(n5327), .ZN(U2808)
         );
  INV_X1 U6451 ( .A(n5329), .ZN(n5342) );
  INV_X1 U6452 ( .A(n5500), .ZN(n5334) );
  NAND2_X1 U6453 ( .A1(n5393), .A2(EBX_REG_18__SCAN_IN), .ZN(n5331) );
  OAI211_X1 U6454 ( .C1(n6068), .C2(n5332), .A(n5331), .B(n6084), .ZN(n5333)
         );
  AOI21_X1 U6455 ( .B1(n5334), .B2(n6082), .A(n5333), .ZN(n5336) );
  NAND2_X1 U6456 ( .A1(n5352), .A2(REIP_REG_18__SCAN_IN), .ZN(n5335) );
  OAI211_X1 U6457 ( .C1(n6108), .C2(n5636), .A(n5336), .B(n5335), .ZN(n5337)
         );
  NOR2_X1 U6458 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  OAI21_X1 U6459 ( .B1(n5641), .B2(n6059), .A(n5339), .ZN(U2809) );
  NAND2_X1 U6460 ( .A1(n5340), .A2(n5386), .ZN(n5385) );
  INV_X1 U6461 ( .A(n5373), .ZN(n5341) );
  NAND2_X1 U6462 ( .A1(n5371), .A2(n5357), .ZN(n5356) );
  AOI21_X1 U6463 ( .B1(n5356), .B2(n5343), .A(n5342), .ZN(n5651) );
  INV_X1 U6464 ( .A(n5651), .ZN(n5553) );
  INV_X1 U6465 ( .A(n5344), .ZN(n5347) );
  INV_X1 U6466 ( .A(n5361), .ZN(n5346) );
  AOI21_X1 U6467 ( .B1(n5347), .B2(n5346), .A(n5345), .ZN(n5805) );
  INV_X1 U6468 ( .A(n5805), .ZN(n5350) );
  AOI21_X1 U6469 ( .B1(n6098), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6097), 
        .ZN(n5349) );
  NAND2_X1 U6470 ( .A1(n5393), .A2(EBX_REG_17__SCAN_IN), .ZN(n5348) );
  OAI211_X1 U6471 ( .C1(n5350), .C2(n6101), .A(n5349), .B(n5348), .ZN(n5351)
         );
  AOI21_X1 U6472 ( .B1(n5647), .B2(n6073), .A(n5351), .ZN(n5355) );
  INV_X1 U6473 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6547) );
  INV_X1 U6474 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6543) );
  NOR3_X1 U6475 ( .A1(n5380), .A2(n6547), .A3(n6543), .ZN(n5353) );
  OAI21_X1 U6476 ( .B1(n5353), .B2(REIP_REG_17__SCAN_IN), .A(n5352), .ZN(n5354) );
  OAI211_X1 U6477 ( .C1(n5553), .C2(n6059), .A(n5355), .B(n5354), .ZN(U2810)
         );
  OAI21_X1 U6478 ( .B1(n5371), .B2(n5357), .A(n5356), .ZN(n5656) );
  XOR2_X1 U6479 ( .A(REIP_REG_16__SCAN_IN), .B(REIP_REG_15__SCAN_IN), .Z(n5368) );
  NOR2_X1 U6480 ( .A1(n5395), .A2(n6547), .ZN(n5367) );
  OAI21_X1 U6481 ( .B1(n6068), .B2(n5358), .A(n6084), .ZN(n5364) );
  INV_X1 U6482 ( .A(n5389), .ZN(n5360) );
  AOI21_X1 U6483 ( .B1(n5360), .B2(n5375), .A(n5359), .ZN(n5362) );
  OR2_X1 U6484 ( .A1(n5362), .A2(n5361), .ZN(n5809) );
  NOR2_X1 U6485 ( .A1(n5809), .A2(n6101), .ZN(n5363) );
  AOI211_X1 U6486 ( .C1(EBX_REG_16__SCAN_IN), .C2(n5393), .A(n5364), .B(n5363), 
        .ZN(n5365) );
  OAI21_X1 U6487 ( .B1(n5658), .B2(n6108), .A(n5365), .ZN(n5366) );
  AOI211_X1 U6488 ( .C1(n5369), .C2(n5368), .A(n5367), .B(n5366), .ZN(n5370)
         );
  OAI21_X1 U6489 ( .B1(n5656), .B2(n6059), .A(n5370), .ZN(U2811) );
  INV_X1 U6490 ( .A(n5385), .ZN(n5374) );
  INV_X1 U6491 ( .A(n5371), .ZN(n5372) );
  INV_X1 U6492 ( .A(n5395), .ZN(n5383) );
  XNOR2_X1 U6493 ( .A(n5389), .B(n5375), .ZN(n5835) );
  NAND2_X1 U6494 ( .A1(n5393), .A2(EBX_REG_15__SCAN_IN), .ZN(n5376) );
  OAI211_X1 U6495 ( .C1(n6068), .C2(n5377), .A(n5376), .B(n6084), .ZN(n5378)
         );
  AOI21_X1 U6496 ( .B1(n5835), .B2(n6082), .A(n5378), .ZN(n5379) );
  OAI21_X1 U6497 ( .B1(n6108), .B2(n5665), .A(n5379), .ZN(n5382) );
  NOR2_X1 U6498 ( .A1(n5380), .A2(REIP_REG_15__SCAN_IN), .ZN(n5381) );
  AOI211_X1 U6499 ( .C1(n5383), .C2(REIP_REG_15__SCAN_IN), .A(n5382), .B(n5381), .ZN(n5384) );
  OAI21_X1 U6500 ( .B1(n5669), .B2(n6059), .A(n5384), .ZN(U2812) );
  OAI21_X1 U6501 ( .B1(n5340), .B2(n5386), .A(n5385), .ZN(n5678) );
  INV_X1 U6502 ( .A(n5674), .ZN(n5399) );
  INV_X1 U6503 ( .A(n5387), .ZN(n5390) );
  OAI21_X1 U6504 ( .B1(n5390), .B2(n3064), .A(n5389), .ZN(n5850) );
  OAI21_X1 U6505 ( .B1(n6068), .B2(n5391), .A(n6084), .ZN(n5392) );
  AOI21_X1 U6506 ( .B1(EBX_REG_14__SCAN_IN), .B2(n5393), .A(n5392), .ZN(n5394)
         );
  OAI21_X1 U6507 ( .B1(n5850), .B2(n6101), .A(n5394), .ZN(n5398) );
  AOI21_X1 U6508 ( .B1(n6045), .B2(REIP_REG_13__SCAN_IN), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5396) );
  NOR2_X1 U6509 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  AOI211_X1 U6510 ( .C1(n6073), .C2(n5399), .A(n5398), .B(n5397), .ZN(n5400)
         );
  OAI21_X1 U6511 ( .B1(n6059), .B2(n5678), .A(n5400), .ZN(U2813) );
  XNOR2_X1 U6512 ( .A(n4428), .B(n5401), .ZN(n5696) );
  AND2_X1 U6513 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NOR2_X1 U6514 ( .A1(n5402), .A2(n5405), .ZN(n6225) );
  NAND2_X1 U6515 ( .A1(n6225), .A2(n6082), .ZN(n5407) );
  AOI21_X1 U6516 ( .B1(n6098), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6097), 
        .ZN(n5406) );
  OAI211_X1 U6517 ( .C1(n5512), .C2(n6093), .A(n5407), .B(n5406), .ZN(n5411)
         );
  NAND2_X1 U6518 ( .A1(n5479), .A2(n5408), .ZN(n6048) );
  AOI21_X1 U6519 ( .B1(n6540), .B2(n5409), .A(n6048), .ZN(n5410) );
  AOI211_X1 U6520 ( .C1(n6073), .C2(n5693), .A(n5411), .B(n5410), .ZN(n5412)
         );
  OAI21_X1 U6521 ( .B1(n5696), .B2(n6059), .A(n5412), .ZN(U2815) );
  OAI21_X1 U6522 ( .B1(n5466), .B2(n5413), .A(n5479), .ZN(n6079) );
  INV_X1 U6523 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6535) );
  OAI22_X1 U6524 ( .A1(n6079), .A2(n6535), .B1(n6101), .B2(n5874), .ZN(n5417)
         );
  AOI22_X1 U6525 ( .A1(n6064), .A2(n6535), .B1(n5393), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5414) );
  OAI211_X1 U6526 ( .C1(n6068), .C2(n5415), .A(n5414), .B(n6084), .ZN(n5416)
         );
  AOI211_X1 U6527 ( .C1(n5712), .C2(n6073), .A(n5417), .B(n5416), .ZN(n5418)
         );
  OAI21_X1 U6528 ( .B1(n6059), .B2(n5709), .A(n5418), .ZN(U2818) );
  OAI22_X1 U6529 ( .A1(n6101), .A2(n5419), .B1(n6093), .B2(n4019), .ZN(n5426)
         );
  INV_X1 U6531 ( .A(n6095), .ZN(n5469) );
  AND2_X1 U6532 ( .A1(n5469), .A2(n5420), .ZN(n6067) );
  INV_X1 U6533 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U6534 ( .B1(n6095), .B2(n5421), .A(n5441), .ZN(n6080) );
  NOR3_X1 U6535 ( .A1(n6095), .A2(REIP_REG_6__SCAN_IN), .A3(n5422), .ZN(n6086)
         );
  OAI33_X1 U6536 ( .A1(1'b0), .A2(n6067), .A3(REIP_REG_7__SCAN_IN), .B1(n6533), 
        .B2(n6080), .B3(n6086), .ZN(n5424) );
  OAI211_X1 U6537 ( .C1(n6068), .C2(n5726), .A(n5424), .B(n6084), .ZN(n5425)
         );
  AOI211_X1 U6538 ( .C1(n6073), .C2(n5729), .A(n5426), .B(n5425), .ZN(n5427)
         );
  OAI21_X1 U6539 ( .B1(n5733), .B2(n6059), .A(n5427), .ZN(U2820) );
  OAI21_X1 U6540 ( .B1(n5428), .B2(n5446), .A(n6059), .ZN(n6105) );
  NAND2_X1 U6541 ( .A1(n6105), .A2(n5429), .ZN(n5439) );
  OAI22_X1 U6542 ( .A1(n5431), .A2(n6068), .B1(n6101), .B2(n5430), .ZN(n5432)
         );
  AOI211_X1 U6543 ( .C1(n5393), .C2(EBX_REG_5__SCAN_IN), .A(n5432), .B(n6097), 
        .ZN(n5438) );
  NAND2_X1 U6544 ( .A1(n6073), .A2(n5433), .ZN(n5437) );
  OAI21_X1 U6545 ( .B1(n6095), .B2(n5434), .A(n6529), .ZN(n5435) );
  NAND2_X1 U6546 ( .A1(n6080), .A2(n5435), .ZN(n5436) );
  NAND4_X1 U6547 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(U2822)
         );
  INV_X1 U6548 ( .A(n6105), .ZN(n5483) );
  INV_X1 U6549 ( .A(n6094), .ZN(n5440) );
  OAI21_X1 U6550 ( .B1(n6095), .B2(n5440), .A(n5441), .ZN(n6104) );
  NAND2_X1 U6551 ( .A1(n5441), .A2(REIP_REG_1__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6552 ( .A1(n5479), .A2(n5442), .ZN(n5443) );
  NAND2_X1 U6553 ( .A1(n5443), .A2(REIP_REG_2__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6554 ( .A1(n5462), .A2(n5444), .ZN(n5453) );
  NAND2_X1 U6555 ( .A1(n5393), .A2(EBX_REG_3__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6556 ( .A1(n6082), .A2(n6279), .ZN(n5448) );
  NOR2_X1 U6557 ( .A1(n5446), .A2(n5445), .ZN(n5464) );
  AOI22_X1 U6558 ( .A1(n5464), .A2(n6347), .B1(n6098), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5447) );
  NAND3_X1 U6559 ( .A1(n5449), .A2(n5448), .A3(n5447), .ZN(n5452) );
  NOR2_X1 U6560 ( .A1(n6108), .A2(n5450), .ZN(n5451) );
  AOI211_X1 U6561 ( .C1(n6104), .C2(n5453), .A(n5452), .B(n5451), .ZN(n5454)
         );
  OAI21_X1 U6562 ( .B1(n5483), .B2(n5455), .A(n5454), .ZN(U2824) );
  INV_X1 U6563 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6524) );
  OAI21_X1 U6564 ( .B1(n6095), .B2(n6578), .A(n6524), .ZN(n5461) );
  NAND2_X1 U6565 ( .A1(n5393), .A2(EBX_REG_2__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6566 ( .A1(n6082), .A2(n6288), .ZN(n5457) );
  AOI22_X1 U6567 ( .A1(n5464), .A2(n4526), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6098), .ZN(n5456) );
  NAND3_X1 U6568 ( .A1(n5458), .A2(n5457), .A3(n5456), .ZN(n5460) );
  NOR2_X1 U6569 ( .A1(n6108), .A2(n6222), .ZN(n5459) );
  AOI211_X1 U6570 ( .C1(n5462), .C2(n5461), .A(n5460), .B(n5459), .ZN(n5463)
         );
  OAI21_X1 U6571 ( .B1(n5483), .B2(n6216), .A(n5463), .ZN(U2825) );
  INV_X1 U6572 ( .A(n5464), .ZN(n6092) );
  AOI22_X1 U6573 ( .A1(n5466), .A2(REIP_REG_1__SCAN_IN), .B1(n6082), .B2(n5465), .ZN(n5467) );
  OAI21_X1 U6574 ( .B1(n6068), .B2(n6745), .A(n5467), .ZN(n5468) );
  AOI21_X1 U6575 ( .B1(n5469), .B2(n6578), .A(n5468), .ZN(n5470) );
  OAI21_X1 U6576 ( .B1(n4511), .B2(n6092), .A(n5470), .ZN(n5472) );
  NOR2_X1 U6577 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5471)
         );
  AOI211_X1 U6578 ( .C1(EBX_REG_1__SCAN_IN), .C2(n5393), .A(n5472), .B(n5471), 
        .ZN(n5473) );
  OAI21_X1 U6579 ( .B1(n5483), .B2(n5474), .A(n5473), .ZN(U2826) );
  NOR2_X1 U6580 ( .A1(n6093), .A2(n5475), .ZN(n5478) );
  OAI22_X1 U6581 ( .A1(n6101), .A2(n5476), .B1(n3373), .B2(n6092), .ZN(n5477)
         );
  AOI211_X1 U6582 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5479), .A(n5478), .B(n5477), 
        .ZN(n5481) );
  OAI21_X1 U6583 ( .B1(n6073), .B2(n6098), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5480) );
  OAI211_X1 U6584 ( .C1(n5483), .C2(n5482), .A(n5481), .B(n5480), .ZN(U2827)
         );
  AOI22_X1 U6585 ( .A1(n5740), .A2(n5514), .B1(n5504), .B2(EBX_REG_29__SCAN_IN), .ZN(n5484) );
  OAI21_X1 U6586 ( .B1(n5485), .B2(n5499), .A(n5484), .ZN(U2830) );
  OAI222_X1 U6587 ( .A1(n5487), .A2(n5517), .B1(n5519), .B2(n5486), .C1(n5213), 
        .C2(n5516), .ZN(U2831) );
  INV_X1 U6588 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6736) );
  OAI222_X1 U6589 ( .A1(n6736), .A2(n5517), .B1(n5519), .B2(n5743), .C1(n5527), 
        .C2(n5499), .ZN(U2832) );
  INV_X1 U6590 ( .A(n5488), .ZN(n5760) );
  OAI222_X1 U6591 ( .A1(n6735), .A2(n5517), .B1(n5519), .B2(n5760), .C1(n5593), 
        .C2(n5499), .ZN(U2833) );
  AOI22_X1 U6592 ( .A1(n5767), .A2(n5514), .B1(n5504), .B2(EBX_REG_25__SCAN_IN), .ZN(n5489) );
  OAI21_X1 U6593 ( .B1(n5600), .B2(n5499), .A(n5489), .ZN(U2834) );
  AOI22_X1 U6594 ( .A1(n5490), .A2(n5514), .B1(n5504), .B2(EBX_REG_24__SCAN_IN), .ZN(n5491) );
  OAI21_X1 U6595 ( .B1(n5534), .B2(n5499), .A(n5491), .ZN(U2835) );
  INV_X1 U6596 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5493) );
  OAI222_X1 U6597 ( .A1(n5493), .A2(n5517), .B1(n5519), .B2(n5492), .C1(n5537), 
        .C2(n5516), .ZN(U2836) );
  AOI22_X1 U6598 ( .A1(n5494), .A2(n5514), .B1(n5504), .B2(EBX_REG_22__SCAN_IN), .ZN(n5495) );
  OAI21_X1 U6599 ( .B1(n5540), .B2(n5499), .A(n5495), .ZN(U2837) );
  AOI22_X1 U6600 ( .A1(n5775), .A2(n5514), .B1(n5504), .B2(EBX_REG_21__SCAN_IN), .ZN(n5496) );
  OAI21_X1 U6601 ( .B1(n5543), .B2(n5499), .A(n5496), .ZN(U2838) );
  AOI22_X1 U6602 ( .A1(n5788), .A2(n5514), .B1(EBX_REG_20__SCAN_IN), .B2(n5504), .ZN(n5497) );
  OAI21_X1 U6603 ( .B1(n5546), .B2(n5499), .A(n5497), .ZN(U2839) );
  AOI22_X1 U6604 ( .A1(n5796), .A2(n5514), .B1(n5504), .B2(EBX_REG_19__SCAN_IN), .ZN(n5498) );
  OAI21_X1 U6605 ( .B1(n5630), .B2(n5499), .A(n5498), .ZN(U2840) );
  OAI222_X1 U6606 ( .A1(n5501), .A2(n5517), .B1(n5519), .B2(n5500), .C1(n5641), 
        .C2(n5516), .ZN(U2841) );
  AOI22_X1 U6607 ( .A1(n5805), .A2(n5514), .B1(n5504), .B2(EBX_REG_17__SCAN_IN), .ZN(n5502) );
  OAI21_X1 U6608 ( .B1(n5553), .B2(n5516), .A(n5502), .ZN(U2842) );
  OAI222_X1 U6609 ( .A1(n5809), .A2(n5519), .B1(n5503), .B2(n5517), .C1(n5656), 
        .C2(n5516), .ZN(U2843) );
  AOI22_X1 U6610 ( .A1(n5835), .A2(n5514), .B1(n5504), .B2(EBX_REG_15__SCAN_IN), .ZN(n5505) );
  OAI21_X1 U6611 ( .B1(n5669), .B2(n5516), .A(n5505), .ZN(U2844) );
  INV_X1 U6612 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5506) );
  OAI222_X1 U6613 ( .A1(n5850), .A2(n5519), .B1(n5506), .B2(n5517), .C1(n5678), 
        .C2(n5516), .ZN(U2845) );
  OAI21_X1 U6614 ( .B1(n5402), .B2(n5507), .A(n5387), .ZN(n6051) );
  INV_X1 U6615 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5511) );
  OAI21_X1 U6616 ( .B1(n5508), .B2(n5510), .A(n5509), .ZN(n6044) );
  OAI222_X1 U6617 ( .A1(n6051), .A2(n5519), .B1(n5517), .B2(n5511), .C1(n5516), 
        .C2(n6044), .ZN(U2846) );
  NOR2_X1 U6618 ( .A1(n5517), .A2(n5512), .ZN(n5513) );
  AOI21_X1 U6619 ( .B1(n6225), .B2(n5514), .A(n5513), .ZN(n5515) );
  OAI21_X1 U6620 ( .B1(n5696), .B2(n5516), .A(n5515), .ZN(U2847) );
  OAI22_X1 U6621 ( .A1(n5865), .A2(n5519), .B1(n5518), .B2(n5517), .ZN(n5520)
         );
  AOI21_X1 U6622 ( .B1(n6189), .B2(n5521), .A(n5520), .ZN(n5522) );
  INV_X1 U6623 ( .A(n5522), .ZN(U2848) );
  AOI22_X1 U6624 ( .A1(n5554), .A2(DATAI_28_), .B1(n5564), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6625 ( .A1(n5555), .A2(DATAI_12_), .ZN(n5523) );
  OAI211_X1 U6626 ( .C1(n5213), .C2(n5567), .A(n5524), .B(n5523), .ZN(U2863)
         );
  AOI22_X1 U6627 ( .A1(n5554), .A2(DATAI_27_), .B1(n5564), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6628 ( .A1(n5555), .A2(DATAI_11_), .ZN(n5525) );
  OAI211_X1 U6629 ( .C1(n5527), .C2(n5567), .A(n5526), .B(n5525), .ZN(U2864)
         );
  AOI22_X1 U6630 ( .A1(n5554), .A2(DATAI_26_), .B1(n5564), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6631 ( .A1(n5555), .A2(DATAI_10_), .ZN(n5528) );
  OAI211_X1 U6632 ( .C1(n5593), .C2(n5567), .A(n5529), .B(n5528), .ZN(U2865)
         );
  AOI22_X1 U6633 ( .A1(n5554), .A2(DATAI_25_), .B1(n5564), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6634 ( .A1(n5555), .A2(DATAI_9_), .ZN(n5530) );
  OAI211_X1 U6635 ( .C1(n5600), .C2(n5567), .A(n5531), .B(n5530), .ZN(U2866)
         );
  AOI22_X1 U6636 ( .A1(n5554), .A2(DATAI_24_), .B1(n5564), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U6637 ( .A1(n5555), .A2(DATAI_8_), .ZN(n5532) );
  OAI211_X1 U6638 ( .C1(n5534), .C2(n5567), .A(n5533), .B(n5532), .ZN(U2867)
         );
  AOI22_X1 U6639 ( .A1(n5554), .A2(DATAI_23_), .B1(n5564), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U6640 ( .A1(n5555), .A2(DATAI_7_), .ZN(n5535) );
  OAI211_X1 U6641 ( .C1(n5537), .C2(n5567), .A(n5536), .B(n5535), .ZN(U2868)
         );
  AOI22_X1 U6642 ( .A1(n5554), .A2(DATAI_22_), .B1(n5564), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U6643 ( .A1(n5555), .A2(DATAI_6_), .ZN(n5538) );
  OAI211_X1 U6644 ( .C1(n5540), .C2(n5567), .A(n5539), .B(n5538), .ZN(U2869)
         );
  AOI22_X1 U6645 ( .A1(n5554), .A2(DATAI_21_), .B1(n5564), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U6646 ( .A1(n5555), .A2(DATAI_5_), .ZN(n5541) );
  OAI211_X1 U6647 ( .C1(n5543), .C2(n5567), .A(n5542), .B(n5541), .ZN(U2870)
         );
  AOI22_X1 U6648 ( .A1(n5554), .A2(DATAI_20_), .B1(n5564), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6649 ( .A1(n5555), .A2(DATAI_4_), .ZN(n5544) );
  OAI211_X1 U6650 ( .C1(n5546), .C2(n5567), .A(n5545), .B(n5544), .ZN(U2871)
         );
  AOI22_X1 U6651 ( .A1(n5554), .A2(DATAI_19_), .B1(n5564), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6652 ( .A1(n5555), .A2(DATAI_3_), .ZN(n5547) );
  OAI211_X1 U6653 ( .C1(n5630), .C2(n5567), .A(n5548), .B(n5547), .ZN(U2872)
         );
  AOI22_X1 U6654 ( .A1(n5554), .A2(DATAI_18_), .B1(n5564), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6655 ( .A1(n5555), .A2(DATAI_2_), .ZN(n5549) );
  OAI211_X1 U6656 ( .C1(n5641), .C2(n5567), .A(n5550), .B(n5549), .ZN(U2873)
         );
  AOI22_X1 U6657 ( .A1(n5554), .A2(DATAI_17_), .B1(n5564), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6658 ( .A1(n5555), .A2(DATAI_1_), .ZN(n5551) );
  OAI211_X1 U6659 ( .C1(n5553), .C2(n5567), .A(n5552), .B(n5551), .ZN(U2874)
         );
  AOI22_X1 U6660 ( .A1(n5554), .A2(DATAI_16_), .B1(n5564), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U6661 ( .A1(n5555), .A2(DATAI_0_), .ZN(n5556) );
  OAI211_X1 U6662 ( .C1(n5656), .C2(n5567), .A(n5557), .B(n5556), .ZN(U2875)
         );
  AOI22_X1 U6663 ( .A1(n5565), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5564), .ZN(n5558) );
  OAI21_X1 U6664 ( .B1(n5669), .B2(n5567), .A(n5558), .ZN(U2876) );
  AOI22_X1 U6665 ( .A1(n5565), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5564), .ZN(n5559) );
  OAI21_X1 U6666 ( .B1(n5678), .B2(n5567), .A(n5559), .ZN(U2877) );
  INV_X1 U6667 ( .A(DATAI_13_), .ZN(n6149) );
  OAI222_X1 U6668 ( .A1(n6044), .A2(n5567), .B1(n6149), .B2(n5562), .C1(n5561), 
        .C2(n5560), .ZN(U2878) );
  AOI22_X1 U6669 ( .A1(n5565), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5564), .ZN(n5563) );
  OAI21_X1 U6670 ( .B1(n5696), .B2(n5567), .A(n5563), .ZN(U2879) );
  AOI22_X1 U6671 ( .A1(n5565), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5564), .ZN(n5566) );
  OAI21_X1 U6672 ( .B1(n3014), .B2(n5567), .A(n5566), .ZN(U2880) );
  INV_X1 U6673 ( .A(n4305), .ZN(n5569) );
  NAND2_X1 U6674 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  XNOR2_X1 U6675 ( .A(n5570), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5742)
         );
  NAND2_X1 U6676 ( .A1(n5571), .A2(n6188), .ZN(n5572) );
  NAND2_X1 U6677 ( .A1(n6194), .A2(REIP_REG_29__SCAN_IN), .ZN(n5735) );
  OAI211_X1 U6678 ( .C1(n5727), .C2(n5573), .A(n5572), .B(n5735), .ZN(n5574)
         );
  AOI21_X1 U6679 ( .B1(n5575), .B2(n6217), .A(n5574), .ZN(n5576) );
  OAI21_X1 U6680 ( .B1(n5742), .B2(n6192), .A(n5576), .ZN(U2957) );
  NAND2_X1 U6681 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5586) );
  OAI21_X1 U6682 ( .B1(n5577), .B2(n5586), .A(n5578), .ZN(n5579) );
  XNOR2_X1 U6683 ( .A(n5579), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5752)
         );
  NAND2_X1 U6684 ( .A1(n5580), .A2(n6188), .ZN(n5581) );
  NAND2_X1 U6685 ( .A1(n6194), .A2(REIP_REG_27__SCAN_IN), .ZN(n5746) );
  OAI211_X1 U6686 ( .C1(n5727), .C2(n5582), .A(n5581), .B(n5746), .ZN(n5583)
         );
  AOI21_X1 U6687 ( .B1(n5584), .B2(n6217), .A(n5583), .ZN(n5585) );
  OAI21_X1 U6688 ( .B1(n5752), .B2(n6192), .A(n5585), .ZN(U2959) );
  NAND2_X1 U6689 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  XNOR2_X1 U6690 ( .A(n5577), .B(n5588), .ZN(n5753) );
  NAND2_X1 U6691 ( .A1(n5753), .A2(n6219), .ZN(n5592) );
  AND2_X1 U6692 ( .A1(n6194), .A2(REIP_REG_26__SCAN_IN), .ZN(n5757) );
  NOR2_X1 U6693 ( .A1(n5589), .A2(n6223), .ZN(n5590) );
  AOI211_X1 U6694 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5757), 
        .B(n5590), .ZN(n5591) );
  OAI211_X1 U6695 ( .C1(n5732), .C2(n5593), .A(n5592), .B(n5591), .ZN(U2960)
         );
  OAI21_X1 U6696 ( .B1(n5141), .B2(n5594), .A(n4303), .ZN(n5761) );
  NAND2_X1 U6697 ( .A1(n5761), .A2(n6219), .ZN(n5599) );
  NAND2_X1 U6698 ( .A1(n6194), .A2(REIP_REG_25__SCAN_IN), .ZN(n5763) );
  OAI21_X1 U6699 ( .B1(n5727), .B2(n5595), .A(n5763), .ZN(n5596) );
  AOI21_X1 U6700 ( .B1(n5597), .B2(n6188), .A(n5596), .ZN(n5598) );
  OAI211_X1 U6701 ( .C1(n5732), .C2(n5600), .A(n5599), .B(n5598), .ZN(U2961)
         );
  NAND2_X1 U6702 ( .A1(n5601), .A2(n6188), .ZN(n5603) );
  OAI211_X1 U6703 ( .C1(n5727), .C2(n5604), .A(n5603), .B(n5602), .ZN(n5605)
         );
  AOI21_X1 U6704 ( .B1(n5606), .B2(n6217), .A(n5605), .ZN(n5607) );
  OAI21_X1 U6705 ( .B1(n5608), .B2(n6192), .A(n5607), .ZN(U2962) );
  AOI21_X1 U6706 ( .B1(n5611), .B2(n5610), .A(n5609), .ZN(n5777) );
  NAND2_X1 U6707 ( .A1(n5612), .A2(n6188), .ZN(n5613) );
  NAND2_X1 U6708 ( .A1(n6194), .A2(REIP_REG_21__SCAN_IN), .ZN(n5771) );
  OAI211_X1 U6709 ( .C1(n5727), .C2(n5614), .A(n5613), .B(n5771), .ZN(n5615)
         );
  AOI21_X1 U6710 ( .B1(n5616), .B2(n6217), .A(n5615), .ZN(n5617) );
  OAI21_X1 U6711 ( .B1(n5777), .B2(n6192), .A(n5617), .ZN(U2965) );
  XNOR2_X1 U6712 ( .A(n5689), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5619)
         );
  XNOR2_X1 U6713 ( .A(n5618), .B(n5619), .ZN(n5790) );
  NAND2_X1 U6714 ( .A1(n6194), .A2(REIP_REG_20__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U6715 ( .A1(n6212), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5620)
         );
  OAI211_X1 U6716 ( .C1(n5621), .C2(n6223), .A(n5785), .B(n5620), .ZN(n5622)
         );
  AOI21_X1 U6717 ( .B1(n5623), .B2(n6217), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6718 ( .B1(n5790), .B2(n6192), .A(n5624), .ZN(U2966) );
  NOR2_X1 U6719 ( .A1(n5626), .A2(n5625), .ZN(n5628) );
  XOR2_X1 U6720 ( .A(n5628), .B(n5627), .Z(n5798) );
  NAND2_X1 U6721 ( .A1(n6194), .A2(REIP_REG_19__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U6722 ( .B1(n5727), .B2(n5629), .A(n5793), .ZN(n5632) );
  NOR2_X1 U6723 ( .A1(n5630), .A2(n5732), .ZN(n5631) );
  AOI211_X1 U6724 ( .C1(n6188), .C2(n5633), .A(n5632), .B(n5631), .ZN(n5634)
         );
  OAI21_X1 U6725 ( .B1(n5798), .B2(n6192), .A(n5634), .ZN(U2967) );
  NAND2_X1 U6726 ( .A1(n5635), .A2(n6219), .ZN(n5640) );
  NOR2_X1 U6727 ( .A1(n6223), .A2(n5636), .ZN(n5637) );
  AOI211_X1 U6728 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5638), 
        .B(n5637), .ZN(n5639) );
  OAI211_X1 U6729 ( .C1(n5732), .C2(n5641), .A(n5640), .B(n5639), .ZN(U2968)
         );
  OAI21_X1 U6730 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5686), .A(n2983), 
        .ZN(n5642) );
  OAI21_X1 U6731 ( .B1(n5653), .B2(n5803), .A(n5642), .ZN(n5646) );
  INV_X1 U6732 ( .A(n5643), .ZN(n5644) );
  AOI21_X1 U6733 ( .B1(n5646), .B2(n5645), .A(n5644), .ZN(n5808) );
  INV_X1 U6734 ( .A(n5647), .ZN(n5649) );
  INV_X1 U6735 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6545) );
  NOR2_X1 U6736 ( .A1(n6211), .A2(n6545), .ZN(n5802) );
  AOI21_X1 U6737 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n5802), 
        .ZN(n5648) );
  OAI21_X1 U6738 ( .B1(n5649), .B2(n6223), .A(n5648), .ZN(n5650) );
  AOI21_X1 U6739 ( .B1(n5651), .B2(n6217), .A(n5650), .ZN(n5652) );
  OAI21_X1 U6740 ( .B1(n5808), .B2(n6192), .A(n5652), .ZN(U2969) );
  AOI21_X1 U6741 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5686), .A(n5653), 
        .ZN(n5654) );
  XNOR2_X1 U6742 ( .A(n5655), .B(n5654), .ZN(n5828) );
  INV_X1 U6743 ( .A(n5656), .ZN(n5660) );
  NOR2_X1 U6744 ( .A1(n6211), .A2(n6547), .ZN(n5824) );
  AOI21_X1 U6745 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5824), 
        .ZN(n5657) );
  OAI21_X1 U6746 ( .B1(n5658), .B2(n6223), .A(n5657), .ZN(n5659) );
  AOI21_X1 U6747 ( .B1(n5660), .B2(n6217), .A(n5659), .ZN(n5661) );
  OAI21_X1 U6748 ( .B1(n5828), .B2(n6192), .A(n5661), .ZN(U2970) );
  OAI21_X1 U6749 ( .B1(n5664), .B2(n5663), .A(n2949), .ZN(n5829) );
  NAND2_X1 U6750 ( .A1(n5829), .A2(n6219), .ZN(n5668) );
  NOR2_X1 U6751 ( .A1(n6211), .A2(n6543), .ZN(n5830) );
  NOR2_X1 U6752 ( .A1(n6223), .A2(n5665), .ZN(n5666) );
  AOI211_X1 U6753 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5830), 
        .B(n5666), .ZN(n5667) );
  OAI211_X1 U6754 ( .C1(n5732), .C2(n5669), .A(n5668), .B(n5667), .ZN(U2971)
         );
  NOR2_X1 U6755 ( .A1(n5672), .A2(n5671), .ZN(n5673) );
  XNOR2_X1 U6756 ( .A(n5670), .B(n5673), .ZN(n5838) );
  NAND2_X1 U6757 ( .A1(n5838), .A2(n6219), .ZN(n5677) );
  INV_X1 U6758 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6542) );
  NOR2_X1 U6759 ( .A1(n6211), .A2(n6542), .ZN(n5846) );
  NOR2_X1 U6760 ( .A1(n6223), .A2(n5674), .ZN(n5675) );
  AOI211_X1 U6761 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5846), 
        .B(n5675), .ZN(n5676) );
  OAI211_X1 U6762 ( .C1(n5732), .C2(n5678), .A(n5677), .B(n5676), .ZN(U2972)
         );
  XNOR2_X1 U6763 ( .A(n5679), .B(n5680), .ZN(n5851) );
  NAND2_X1 U6764 ( .A1(n5851), .A2(n6219), .ZN(n5683) );
  INV_X1 U6765 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6047) );
  NOR2_X1 U6766 ( .A1(n6211), .A2(n6047), .ZN(n5855) );
  NOR2_X1 U6767 ( .A1(n6223), .A2(n6055), .ZN(n5681) );
  AOI211_X1 U6768 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5855), 
        .B(n5681), .ZN(n5682) );
  OAI211_X1 U6769 ( .C1(n5732), .C2(n6044), .A(n5683), .B(n5682), .ZN(U2973)
         );
  NOR2_X1 U6770 ( .A1(n5686), .A2(n5684), .ZN(n5697) );
  NAND2_X1 U6771 ( .A1(n5686), .A2(n5684), .ZN(n5698) );
  NAND2_X1 U6772 ( .A1(n2963), .A2(n5698), .ZN(n5860) );
  AOI21_X1 U6773 ( .B1(n5686), .B2(n5685), .A(n5860), .ZN(n5687) );
  AOI211_X1 U6774 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5689), .A(n5697), .B(n5687), .ZN(n5691) );
  AOI21_X1 U6775 ( .B1(n5689), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5688), 
        .ZN(n5690) );
  XNOR2_X1 U6776 ( .A(n5691), .B(n5690), .ZN(n6230) );
  NAND2_X1 U6777 ( .A1(n6230), .A2(n6219), .ZN(n5695) );
  NOR2_X1 U6778 ( .A1(n6211), .A2(n6540), .ZN(n6224) );
  NOR2_X1 U6779 ( .A1(n5727), .A2(n3009), .ZN(n5692) );
  AOI211_X1 U6780 ( .C1(n6188), .C2(n5693), .A(n6224), .B(n5692), .ZN(n5694)
         );
  OAI211_X1 U6781 ( .C1(n5696), .C2(n5732), .A(n5695), .B(n5694), .ZN(U2974)
         );
  INV_X1 U6782 ( .A(n5697), .ZN(n5859) );
  NAND2_X1 U6783 ( .A1(n5859), .A2(n5698), .ZN(n5699) );
  XNOR2_X1 U6784 ( .A(n2963), .B(n5699), .ZN(n6240) );
  NAND2_X1 U6785 ( .A1(n6240), .A2(n6219), .ZN(n5703) );
  INV_X1 U6786 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5700) );
  NOR2_X1 U6787 ( .A1(n6211), .A2(n5700), .ZN(n6237) );
  NOR2_X1 U6788 ( .A1(n5727), .A2(n3007), .ZN(n5701) );
  AOI211_X1 U6789 ( .C1(n6188), .C2(n6062), .A(n6237), .B(n5701), .ZN(n5702)
         );
  OAI211_X1 U6790 ( .C1(n5732), .C2(n6060), .A(n5703), .B(n5702), .ZN(U2976)
         );
  INV_X1 U6791 ( .A(n5705), .ZN(n5706) );
  NOR2_X1 U6792 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  XNOR2_X1 U6793 ( .A(n5704), .B(n5708), .ZN(n5883) );
  NAND2_X1 U6794 ( .A1(n6194), .A2(REIP_REG_9__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U6795 ( .B1(n5727), .B2(n5415), .A(n5878), .ZN(n5711) );
  NOR2_X1 U6796 ( .A1(n5709), .A2(n5732), .ZN(n5710) );
  AOI211_X1 U6797 ( .C1(n6188), .C2(n5712), .A(n5711), .B(n5710), .ZN(n5713)
         );
  OAI21_X1 U6798 ( .B1(n5883), .B2(n6192), .A(n5713), .ZN(U2977) );
  OAI21_X1 U6799 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5717) );
  INV_X1 U6800 ( .A(n5717), .ZN(n6249) );
  NAND2_X1 U6801 ( .A1(n6249), .A2(n6219), .ZN(n5721) );
  INV_X1 U6802 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5718) );
  NOR2_X1 U6803 ( .A1(n6211), .A2(n5718), .ZN(n6245) );
  NOR2_X1 U6804 ( .A1(n6223), .A2(n6072), .ZN(n5719) );
  AOI211_X1 U6805 ( .C1(n6212), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6245), 
        .B(n5719), .ZN(n5720) );
  OAI211_X1 U6806 ( .C1(n5732), .C2(n6071), .A(n5721), .B(n5720), .ZN(U2978)
         );
  OAI21_X1 U6807 ( .B1(n5724), .B2(n5723), .A(n5722), .ZN(n5725) );
  INV_X1 U6808 ( .A(n5725), .ZN(n6256) );
  NAND2_X1 U6809 ( .A1(n6256), .A2(n6219), .ZN(n5731) );
  NOR2_X1 U6810 ( .A1(n6211), .A2(n6533), .ZN(n6253) );
  NOR2_X1 U6811 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  AOI211_X1 U6812 ( .C1(n6188), .C2(n5729), .A(n6253), .B(n5728), .ZN(n5730)
         );
  OAI211_X1 U6813 ( .C1(n5733), .C2(n5732), .A(n5731), .B(n5730), .ZN(U2979)
         );
  NAND2_X1 U6814 ( .A1(n5734), .A2(n5737), .ZN(n5736) );
  OAI211_X1 U6815 ( .C1(n5738), .C2(n5737), .A(n5736), .B(n5735), .ZN(n5739)
         );
  AOI21_X1 U6816 ( .B1(n5740), .B2(n6289), .A(n5739), .ZN(n5741) );
  OAI21_X1 U6817 ( .B1(n5742), .B2(n5882), .A(n5741), .ZN(U2989) );
  INV_X1 U6818 ( .A(n5743), .ZN(n5750) );
  NAND3_X1 U6819 ( .A1(n5745), .A2(n5744), .A3(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U6820 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  AOI211_X1 U6821 ( .C1(n5750), .C2(n6289), .A(n5749), .B(n5748), .ZN(n5751)
         );
  OAI21_X1 U6822 ( .B1(n5752), .B2(n5882), .A(n5751), .ZN(U2991) );
  NAND2_X1 U6823 ( .A1(n5753), .A2(n6294), .ZN(n5759) );
  INV_X1 U6824 ( .A(n5754), .ZN(n5762) );
  XNOR2_X1 U6825 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5755) );
  NOR2_X1 U6826 ( .A1(n5765), .A2(n5755), .ZN(n5756) );
  AOI211_X1 U6827 ( .C1(n5762), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5757), .B(n5756), .ZN(n5758) );
  OAI211_X1 U6828 ( .C1(n5873), .C2(n5760), .A(n5759), .B(n5758), .ZN(U2992)
         );
  INV_X1 U6829 ( .A(n5761), .ZN(n5769) );
  NAND2_X1 U6830 ( .A1(n5762), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U6831 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5765), .A(n5764), .B(n5763), .ZN(n5766) );
  AOI21_X1 U6832 ( .B1(n5767), .B2(n6289), .A(n5766), .ZN(n5768) );
  OAI21_X1 U6833 ( .B1(n5769), .B2(n5882), .A(n5768), .ZN(U2993) );
  NAND2_X1 U6834 ( .A1(n5770), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5772) );
  OAI211_X1 U6835 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5773), .A(n5772), .B(n5771), .ZN(n5774) );
  AOI21_X1 U6836 ( .B1(n5775), .B2(n6289), .A(n5774), .ZN(n5776) );
  OAI21_X1 U6837 ( .B1(n5777), .B2(n5882), .A(n5776), .ZN(U2997) );
  AOI21_X1 U6838 ( .B1(n5779), .B2(n5819), .A(n5778), .ZN(n5794) );
  NOR2_X1 U6839 ( .A1(n5799), .A2(n5780), .ZN(n5791) );
  INV_X1 U6840 ( .A(n5781), .ZN(n5783) );
  NAND3_X1 U6841 ( .A1(n5791), .A2(n5783), .A3(n5782), .ZN(n5784) );
  OAI211_X1 U6842 ( .C1(n5794), .C2(n5786), .A(n5785), .B(n5784), .ZN(n5787)
         );
  AOI21_X1 U6843 ( .B1(n5788), .B2(n6289), .A(n5787), .ZN(n5789) );
  OAI21_X1 U6844 ( .B1(n5790), .B2(n5882), .A(n5789), .ZN(U2998) );
  NAND2_X1 U6845 ( .A1(n5791), .A2(n6752), .ZN(n5792) );
  OAI211_X1 U6846 ( .C1(n5794), .C2(n6752), .A(n5793), .B(n5792), .ZN(n5795)
         );
  AOI21_X1 U6847 ( .B1(n5796), .B2(n6289), .A(n5795), .ZN(n5797) );
  OAI21_X1 U6848 ( .B1(n5798), .B2(n5882), .A(n5797), .ZN(U2999) );
  INV_X1 U6849 ( .A(n5799), .ZN(n5804) );
  NOR2_X1 U6850 ( .A1(n5800), .A2(n5803), .ZN(n5801) );
  AOI211_X1 U6851 ( .C1(n5804), .C2(n5803), .A(n5802), .B(n5801), .ZN(n5807)
         );
  NAND2_X1 U6852 ( .A1(n5805), .A2(n6289), .ZN(n5806) );
  OAI211_X1 U6853 ( .C1(n5808), .C2(n5882), .A(n5807), .B(n5806), .ZN(U3001)
         );
  NOR2_X1 U6854 ( .A1(n5809), .A2(n5873), .ZN(n5826) );
  AND2_X1 U6855 ( .A1(n6231), .A2(n5810), .ZN(n5821) );
  NAND2_X1 U6856 ( .A1(n5821), .A2(n6750), .ZN(n5832) );
  INV_X1 U6857 ( .A(n5810), .ZN(n5818) );
  INV_X1 U6858 ( .A(n5811), .ZN(n5812) );
  OR2_X1 U6859 ( .A1(n5867), .A2(n5812), .ZN(n5817) );
  OAI21_X1 U6860 ( .B1(n5814), .B2(n5813), .A(n5866), .ZN(n5815) );
  INV_X1 U6861 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U6862 ( .A1(n5817), .A2(n5816), .ZN(n6226) );
  AOI21_X1 U6863 ( .B1(n5819), .B2(n5818), .A(n6226), .ZN(n5833) );
  AOI21_X1 U6864 ( .B1(n5832), .B2(n5833), .A(n5820), .ZN(n5825) );
  INV_X1 U6865 ( .A(n5821), .ZN(n5822) );
  NOR3_X1 U6866 ( .A1(n5822), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6750), 
        .ZN(n5823) );
  NOR4_X1 U6867 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n5827)
         );
  OAI21_X1 U6868 ( .B1(n5828), .B2(n5882), .A(n5827), .ZN(U3002) );
  INV_X1 U6869 ( .A(n5829), .ZN(n5837) );
  INV_X1 U6870 ( .A(n5830), .ZN(n5831) );
  OAI211_X1 U6871 ( .C1(n5833), .C2(n6750), .A(n5832), .B(n5831), .ZN(n5834)
         );
  AOI21_X1 U6872 ( .B1(n5835), .B2(n6289), .A(n5834), .ZN(n5836) );
  OAI21_X1 U6873 ( .B1(n5837), .B2(n5882), .A(n5836), .ZN(U3003) );
  NAND2_X1 U6874 ( .A1(n5838), .A2(n6294), .ZN(n5849) );
  NAND2_X1 U6875 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5853) );
  INV_X1 U6876 ( .A(n5844), .ZN(n5839) );
  NOR2_X1 U6877 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  AOI211_X1 U6878 ( .C1(n5853), .C2(n5842), .A(n5841), .B(n6226), .ZN(n5852)
         );
  OAI21_X1 U6879 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5843), .A(n5852), 
        .ZN(n5847) );
  INV_X1 U6880 ( .A(n6231), .ZN(n6228) );
  NOR3_X1 U6881 ( .A1(n6228), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n5844), 
        .ZN(n5845) );
  AOI211_X1 U6882 ( .C1(n5847), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5846), .B(n5845), .ZN(n5848) );
  OAI211_X1 U6883 ( .C1(n5873), .C2(n5850), .A(n5849), .B(n5848), .ZN(U3004)
         );
  NAND2_X1 U6884 ( .A1(n5851), .A2(n6294), .ZN(n5858) );
  INV_X1 U6885 ( .A(n5852), .ZN(n5856) );
  NOR3_X1 U6886 ( .A1(n6228), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5853), 
        .ZN(n5854) );
  AOI211_X1 U6887 ( .C1(INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n5856), .A(n5855), .B(n5854), .ZN(n5857) );
  OAI211_X1 U6888 ( .C1(n5873), .C2(n6051), .A(n5858), .B(n5857), .ZN(U3005)
         );
  NAND2_X1 U6889 ( .A1(n5860), .A2(n5859), .ZN(n5862) );
  XNOR2_X1 U6890 ( .A(n5686), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5861)
         );
  XNOR2_X1 U6891 ( .A(n5862), .B(n5861), .ZN(n6193) );
  OAI22_X1 U6892 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6228), .B1(n6193), .B2(n5882), .ZN(n5863) );
  NOR2_X1 U6893 ( .A1(n6211), .A2(n6538), .ZN(n6186) );
  AOI211_X1 U6894 ( .C1(n6226), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5863), .B(n6186), .ZN(n5864) );
  OAI21_X1 U6895 ( .B1(n5865), .B2(n5873), .A(n5864), .ZN(U3007) );
  OAI21_X1 U6896 ( .B1(n5868), .B2(n5867), .A(n5866), .ZN(n5869) );
  AOI21_X1 U6897 ( .B1(n5871), .B2(n5870), .A(n5869), .ZN(n6260) );
  OAI21_X1 U6898 ( .B1(n5872), .B2(n6247), .A(n6260), .ZN(n6239) );
  NOR2_X1 U6899 ( .A1(n5874), .A2(n5873), .ZN(n5880) );
  OAI21_X1 U6900 ( .B1(n5876), .B2(n6290), .A(n5875), .ZN(n6280) );
  NOR2_X1 U6901 ( .A1(n5877), .A2(n6280), .ZN(n6255) );
  NAND2_X1 U6902 ( .A1(n6247), .A2(n6255), .ZN(n6244) );
  OAI21_X1 U6903 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6244), .A(n5878), 
        .ZN(n5879) );
  AOI211_X1 U6904 ( .C1(n6239), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5880), 
        .B(n5879), .ZN(n5881) );
  OAI21_X1 U6905 ( .B1(n5883), .B2(n5882), .A(n5881), .ZN(U3009) );
  OAI211_X1 U6906 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5884), .A(n6443), .B(
        n6442), .ZN(n5885) );
  OAI21_X1 U6907 ( .B1(n5895), .B2(n4511), .A(n5885), .ZN(n5886) );
  MUX2_X1 U6908 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5886), .S(n6302), 
        .Z(U3464) );
  XNOR2_X1 U6909 ( .A(n5887), .B(n6443), .ZN(n5889) );
  INV_X1 U6910 ( .A(n4526), .ZN(n5888) );
  OAI22_X1 U6911 ( .A1(n5889), .A2(n6593), .B1(n5895), .B2(n5888), .ZN(n5890)
         );
  MUX2_X1 U6912 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5890), .S(n6302), 
        .Z(U3463) );
  INV_X1 U6913 ( .A(n6444), .ZN(n5892) );
  NOR3_X1 U6914 ( .A1(n5893), .A2(n5892), .A3(n5891), .ZN(n5894) );
  OAI222_X1 U6915 ( .A1(n4165), .A2(n5896), .B1(n6384), .B2(n5895), .C1(n6593), 
        .C2(n5894), .ZN(n5897) );
  MUX2_X1 U6916 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5897), .S(n6302), 
        .Z(U3462) );
  INV_X1 U6917 ( .A(n5898), .ZN(n5901) );
  OAI22_X1 U6918 ( .A1(n5901), .A2(n6514), .B1(n5900), .B2(n5899), .ZN(n5903)
         );
  MUX2_X1 U6919 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5903), .S(n5902), 
        .Z(U3456) );
  NOR2_X1 U6920 ( .A1(n5936), .A2(n6593), .ZN(n5904) );
  AOI21_X1 U6921 ( .B1(n5939), .B2(n5904), .A(n6394), .ZN(n5908) );
  AOI21_X1 U6922 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6344), .A(n5905), .ZN(
        n6352) );
  NAND2_X1 U6923 ( .A1(n5906), .A2(n6390), .ZN(n5933) );
  AOI21_X1 U6924 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5933), .A(n5988), .ZN(
        n5907) );
  NAND2_X1 U6925 ( .A1(n5932), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5913) );
  NOR2_X1 U6926 ( .A1(n6344), .A2(n6345), .ZN(n5909) );
  AOI22_X1 U6927 ( .A1(n5910), .A2(n6442), .B1(n6396), .B2(n5909), .ZN(n5934)
         );
  OAI22_X1 U6928 ( .A1(n5934), .A2(n5993), .B1(n6439), .B2(n5933), .ZN(n5911)
         );
  AOI21_X1 U6929 ( .B1(n5936), .B2(n6403), .A(n5911), .ZN(n5912) );
  OAI211_X1 U6930 ( .C1(n5939), .C2(n6457), .A(n5913), .B(n5912), .ZN(U3020)
         );
  NAND2_X1 U6931 ( .A1(n5932), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5916) );
  OAI22_X1 U6932 ( .A1(n5934), .A2(n5997), .B1(n6458), .B2(n5933), .ZN(n5914)
         );
  AOI21_X1 U6933 ( .B1(n5936), .B2(n6407), .A(n5914), .ZN(n5915) );
  OAI211_X1 U6934 ( .C1(n5939), .C2(n6459), .A(n5916), .B(n5915), .ZN(U3021)
         );
  NAND2_X1 U6935 ( .A1(n5932), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5919) );
  OAI22_X1 U6936 ( .A1(n5934), .A2(n6001), .B1(n6465), .B2(n5933), .ZN(n5917)
         );
  AOI21_X1 U6937 ( .B1(n5936), .B2(n6411), .A(n5917), .ZN(n5918) );
  OAI211_X1 U6938 ( .C1(n5939), .C2(n6466), .A(n5919), .B(n5918), .ZN(U3022)
         );
  NAND2_X1 U6939 ( .A1(n5932), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5922) );
  OAI22_X1 U6940 ( .A1(n5934), .A2(n6005), .B1(n6472), .B2(n5933), .ZN(n5920)
         );
  AOI21_X1 U6941 ( .B1(n5936), .B2(n6415), .A(n5920), .ZN(n5921) );
  OAI211_X1 U6942 ( .C1(n5939), .C2(n6478), .A(n5922), .B(n5921), .ZN(U3023)
         );
  NAND2_X1 U6943 ( .A1(n5932), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5925) );
  OAI22_X1 U6944 ( .A1(n5934), .A2(n6009), .B1(n6479), .B2(n5933), .ZN(n5923)
         );
  AOI21_X1 U6945 ( .B1(n5936), .B2(n6419), .A(n5923), .ZN(n5924) );
  OAI211_X1 U6946 ( .C1(n5939), .C2(n6485), .A(n5925), .B(n5924), .ZN(U3024)
         );
  NAND2_X1 U6947 ( .A1(n5932), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5928) );
  OAI22_X1 U6948 ( .A1(n5934), .A2(n6013), .B1(n6486), .B2(n5933), .ZN(n5926)
         );
  AOI21_X1 U6949 ( .B1(n5936), .B2(n6423), .A(n5926), .ZN(n5927) );
  OAI211_X1 U6950 ( .C1(n5939), .C2(n6487), .A(n5928), .B(n5927), .ZN(U3025)
         );
  NAND2_X1 U6951 ( .A1(n5932), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5931) );
  OAI22_X1 U6952 ( .A1(n5934), .A2(n6017), .B1(n6493), .B2(n5933), .ZN(n5929)
         );
  AOI21_X1 U6953 ( .B1(n5936), .B2(n6427), .A(n5929), .ZN(n5930) );
  OAI211_X1 U6954 ( .C1(n5939), .C2(n6499), .A(n5931), .B(n5930), .ZN(U3026)
         );
  NAND2_X1 U6955 ( .A1(n5932), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5938) );
  OAI22_X1 U6956 ( .A1(n5934), .A2(n6024), .B1(n6501), .B2(n5933), .ZN(n5935)
         );
  AOI21_X1 U6957 ( .B1(n5936), .B2(n6434), .A(n5935), .ZN(n5937) );
  OAI211_X1 U6958 ( .C1(n5939), .C2(n6502), .A(n5938), .B(n5937), .ZN(U3027)
         );
  NOR3_X1 U6959 ( .A1(n5940), .A2(n5975), .A3(n6593), .ZN(n5942) );
  OAI22_X1 U6960 ( .A1(n5942), .A2(n6394), .B1(n6384), .B2(n5941), .ZN(n5946)
         );
  NAND2_X1 U6961 ( .A1(n5943), .A2(n6390), .ZN(n5972) );
  AOI21_X1 U6962 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5972), .A(n5988), .ZN(
        n5944) );
  NAND3_X1 U6963 ( .A1(n5946), .A2(n5945), .A3(n5944), .ZN(n5971) );
  NAND2_X1 U6964 ( .A1(n5971), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5952) );
  AOI22_X1 U6965 ( .A1(n5949), .A2(n5948), .B1(n6396), .B2(n5947), .ZN(n5973)
         );
  OAI22_X1 U6966 ( .A1(n5973), .A2(n5993), .B1(n6439), .B2(n5972), .ZN(n5950)
         );
  AOI21_X1 U6967 ( .B1(n5975), .B2(n6403), .A(n5950), .ZN(n5951) );
  OAI211_X1 U6968 ( .C1(n5978), .C2(n6457), .A(n5952), .B(n5951), .ZN(U3084)
         );
  NAND2_X1 U6969 ( .A1(n5971), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5955) );
  OAI22_X1 U6970 ( .A1(n5973), .A2(n5997), .B1(n6458), .B2(n5972), .ZN(n5953)
         );
  AOI21_X1 U6971 ( .B1(n5975), .B2(n6407), .A(n5953), .ZN(n5954) );
  OAI211_X1 U6972 ( .C1(n5978), .C2(n6459), .A(n5955), .B(n5954), .ZN(U3085)
         );
  NAND2_X1 U6973 ( .A1(n5971), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5958) );
  OAI22_X1 U6974 ( .A1(n5973), .A2(n6001), .B1(n6465), .B2(n5972), .ZN(n5956)
         );
  AOI21_X1 U6975 ( .B1(n5975), .B2(n6411), .A(n5956), .ZN(n5957) );
  OAI211_X1 U6976 ( .C1(n5978), .C2(n6466), .A(n5958), .B(n5957), .ZN(U3086)
         );
  NAND2_X1 U6977 ( .A1(n5971), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5961) );
  OAI22_X1 U6978 ( .A1(n5973), .A2(n6005), .B1(n6472), .B2(n5972), .ZN(n5959)
         );
  AOI21_X1 U6979 ( .B1(n5975), .B2(n6415), .A(n5959), .ZN(n5960) );
  OAI211_X1 U6980 ( .C1(n5978), .C2(n6478), .A(n5961), .B(n5960), .ZN(U3087)
         );
  NAND2_X1 U6981 ( .A1(n5971), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5964) );
  OAI22_X1 U6982 ( .A1(n5973), .A2(n6009), .B1(n6479), .B2(n5972), .ZN(n5962)
         );
  AOI21_X1 U6983 ( .B1(n5975), .B2(n6419), .A(n5962), .ZN(n5963) );
  OAI211_X1 U6984 ( .C1(n5978), .C2(n6485), .A(n5964), .B(n5963), .ZN(U3088)
         );
  NAND2_X1 U6985 ( .A1(n5971), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5967) );
  OAI22_X1 U6986 ( .A1(n5973), .A2(n6013), .B1(n6486), .B2(n5972), .ZN(n5965)
         );
  AOI21_X1 U6987 ( .B1(n5975), .B2(n6423), .A(n5965), .ZN(n5966) );
  OAI211_X1 U6988 ( .C1(n5978), .C2(n6487), .A(n5967), .B(n5966), .ZN(U3089)
         );
  NAND2_X1 U6989 ( .A1(n5971), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5970) );
  OAI22_X1 U6990 ( .A1(n5973), .A2(n6017), .B1(n6493), .B2(n5972), .ZN(n5968)
         );
  AOI21_X1 U6991 ( .B1(n5975), .B2(n6427), .A(n5968), .ZN(n5969) );
  OAI211_X1 U6992 ( .C1(n5978), .C2(n6499), .A(n5970), .B(n5969), .ZN(U3090)
         );
  NAND2_X1 U6993 ( .A1(n5971), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5977) );
  OAI22_X1 U6994 ( .A1(n5973), .A2(n6024), .B1(n6501), .B2(n5972), .ZN(n5974)
         );
  AOI21_X1 U6995 ( .B1(n5975), .B2(n6434), .A(n5974), .ZN(n5976) );
  OAI211_X1 U6996 ( .C1(n5978), .C2(n6502), .A(n5977), .B(n5976), .ZN(U3091)
         );
  AOI21_X1 U6997 ( .B1(n5984), .B2(n6510), .A(n6028), .ZN(n5980) );
  NOR2_X1 U6998 ( .A1(n5980), .A2(n6593), .ZN(n5986) );
  INV_X1 U6999 ( .A(n5981), .ZN(n5982) );
  NOR2_X1 U7000 ( .A1(n6311), .A2(n6312), .ZN(n6450) );
  NAND2_X1 U7001 ( .A1(n6450), .A2(n6390), .ZN(n6018) );
  OAI22_X1 U7002 ( .A1(n6510), .A2(n6457), .B1(n6018), .B2(n6439), .ZN(n5985)
         );
  AOI21_X1 U7003 ( .B1(n6020), .B2(n6403), .A(n5985), .ZN(n5992) );
  INV_X1 U7004 ( .A(n5986), .ZN(n5990) );
  AOI211_X1 U7005 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6018), .A(n5988), .B(
        n5987), .ZN(n5989) );
  NAND2_X1 U7006 ( .A1(n6021), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5991)
         );
  OAI211_X1 U7007 ( .C1(n6025), .C2(n5993), .A(n5992), .B(n5991), .ZN(U3100)
         );
  OAI22_X1 U7008 ( .A1(n6510), .A2(n6459), .B1(n6018), .B2(n6458), .ZN(n5994)
         );
  AOI21_X1 U7009 ( .B1(n6020), .B2(n6407), .A(n5994), .ZN(n5996) );
  NAND2_X1 U7010 ( .A1(n6021), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5995)
         );
  OAI211_X1 U7011 ( .C1(n6025), .C2(n5997), .A(n5996), .B(n5995), .ZN(U3101)
         );
  OAI22_X1 U7012 ( .A1(n6510), .A2(n6466), .B1(n6018), .B2(n6465), .ZN(n5998)
         );
  AOI21_X1 U7013 ( .B1(n6020), .B2(n6411), .A(n5998), .ZN(n6000) );
  NAND2_X1 U7014 ( .A1(n6021), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5999)
         );
  OAI211_X1 U7015 ( .C1(n6025), .C2(n6001), .A(n6000), .B(n5999), .ZN(U3102)
         );
  OAI22_X1 U7016 ( .A1(n6510), .A2(n6478), .B1(n6018), .B2(n6472), .ZN(n6002)
         );
  AOI21_X1 U7017 ( .B1(n6020), .B2(n6415), .A(n6002), .ZN(n6004) );
  NAND2_X1 U7018 ( .A1(n6021), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6003)
         );
  OAI211_X1 U7019 ( .C1(n6025), .C2(n6005), .A(n6004), .B(n6003), .ZN(U3103)
         );
  OAI22_X1 U7020 ( .A1(n6510), .A2(n6485), .B1(n6018), .B2(n6479), .ZN(n6006)
         );
  AOI21_X1 U7021 ( .B1(n6020), .B2(n6419), .A(n6006), .ZN(n6008) );
  NAND2_X1 U7022 ( .A1(n6021), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6007)
         );
  OAI211_X1 U7023 ( .C1(n6025), .C2(n6009), .A(n6008), .B(n6007), .ZN(U3104)
         );
  OAI22_X1 U7024 ( .A1(n6510), .A2(n6487), .B1(n6018), .B2(n6486), .ZN(n6010)
         );
  AOI21_X1 U7025 ( .B1(n6020), .B2(n6423), .A(n6010), .ZN(n6012) );
  NAND2_X1 U7026 ( .A1(n6021), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6011)
         );
  OAI211_X1 U7027 ( .C1(n6025), .C2(n6013), .A(n6012), .B(n6011), .ZN(U3105)
         );
  OAI22_X1 U7028 ( .A1(n6510), .A2(n6499), .B1(n6018), .B2(n6493), .ZN(n6014)
         );
  AOI21_X1 U7029 ( .B1(n6020), .B2(n6427), .A(n6014), .ZN(n6016) );
  NAND2_X1 U7030 ( .A1(n6021), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6015)
         );
  OAI211_X1 U7031 ( .C1(n6025), .C2(n6017), .A(n6016), .B(n6015), .ZN(U3106)
         );
  OAI22_X1 U7032 ( .A1(n6510), .A2(n6502), .B1(n6018), .B2(n6501), .ZN(n6019)
         );
  AOI21_X1 U7033 ( .B1(n6020), .B2(n6434), .A(n6019), .ZN(n6023) );
  NAND2_X1 U7034 ( .A1(n6021), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6022)
         );
  OAI211_X1 U7035 ( .C1(n6025), .C2(n6024), .A(n6023), .B(n6022), .ZN(U3107)
         );
  AND2_X1 U7036 ( .A1(n6127), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7037 ( .A(n6546), .ZN(n6588) );
  NOR2_X1 U7038 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6027) );
  OAI21_X1 U7039 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6027), .A(n6606), .ZN(n6026)
         );
  OAI21_X1 U7040 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6588), .A(n6026), .ZN(
        U2791) );
  OAI21_X1 U7041 ( .B1(BS16_N), .B2(n6027), .A(n6576), .ZN(n6575) );
  OAI21_X1 U7042 ( .B1(n6576), .B2(n6028), .A(n6575), .ZN(U2792) );
  AND2_X1 U7043 ( .A1(n6029), .A2(n6517), .ZN(n6589) );
  OAI21_X1 U7044 ( .B1(n6589), .B2(n6030), .A(n6192), .ZN(U2793) );
  NOR4_X1 U7045 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6040)
         );
  NOR4_X1 U7046 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6039) );
  NOR4_X1 U7047 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6031) );
  INV_X1 U7048 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6673) );
  INV_X1 U7049 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6627) );
  NAND3_X1 U7050 ( .A1(n6031), .A2(n6673), .A3(n6627), .ZN(n6037) );
  NOR4_X1 U7051 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6035) );
  NOR4_X1 U7052 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6034) );
  NOR4_X1 U7053 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6033) );
  NOR4_X1 U7054 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n6032) );
  NAND4_X1 U7055 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n6036)
         );
  AOI211_X1 U7056 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6037), .B(n6036), .ZN(n6038) );
  NAND3_X1 U7057 ( .A1(n6040), .A2(n6039), .A3(n6038), .ZN(n6584) );
  NOR2_X1 U7058 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6584), .ZN(n6586) );
  INV_X1 U7059 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U7060 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6577) );
  NAND3_X1 U7061 ( .A1(n6585), .A2(n6651), .A3(n6577), .ZN(n6043) );
  INV_X1 U7062 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6041) );
  AOI22_X1 U7063 ( .A1(n6586), .A2(n6043), .B1(n6584), .B2(n6041), .ZN(U2794)
         );
  AOI22_X1 U7064 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6584), .B1(n6586), 
        .B2(n6651), .ZN(n6042) );
  OAI21_X1 U7065 ( .B1(n6584), .B2(n6043), .A(n6042), .ZN(U2795) );
  INV_X1 U7066 ( .A(n6044), .ZN(n6053) );
  AOI22_X1 U7067 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6098), .B1(n6045), 
        .B2(n6047), .ZN(n6046) );
  OAI211_X1 U7068 ( .C1(n6048), .C2(n6047), .A(n6084), .B(n6046), .ZN(n6049)
         );
  AOI21_X1 U7069 ( .B1(n5393), .B2(EBX_REG_13__SCAN_IN), .A(n6049), .ZN(n6050)
         );
  OAI21_X1 U7070 ( .B1(n6051), .B2(n6101), .A(n6050), .ZN(n6052) );
  AOI21_X1 U7071 ( .B1(n6053), .B2(n6087), .A(n6052), .ZN(n6054) );
  OAI21_X1 U7072 ( .B1(n6055), .B2(n6108), .A(n6054), .ZN(U2814) );
  OAI21_X1 U7073 ( .B1(n6068), .B2(n3007), .A(n6084), .ZN(n6057) );
  NOR2_X1 U7074 ( .A1(n6236), .A2(n6101), .ZN(n6056) );
  AOI211_X1 U7075 ( .C1(EBX_REG_10__SCAN_IN), .C2(n5393), .A(n6057), .B(n6056), 
        .ZN(n6058) );
  OAI21_X1 U7076 ( .B1(n6060), .B2(n6059), .A(n6058), .ZN(n6061) );
  AOI21_X1 U7077 ( .B1(n6062), .B2(n6073), .A(n6061), .ZN(n6066) );
  NAND2_X1 U7078 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6063) );
  OAI211_X1 U7079 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n6064), .B(n6063), .ZN(n6065) );
  OAI211_X1 U7080 ( .C1(n6079), .C2(n5700), .A(n6066), .B(n6065), .ZN(U2817)
         );
  AOI21_X1 U7081 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6067), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6078) );
  INV_X1 U7082 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6069) );
  OAI22_X1 U7083 ( .A1(n6093), .A2(n6742), .B1(n6069), .B2(n6068), .ZN(n6070)
         );
  AOI211_X1 U7084 ( .C1(n6082), .C2(n6246), .A(n6097), .B(n6070), .ZN(n6077)
         );
  INV_X1 U7085 ( .A(n6071), .ZN(n6075) );
  INV_X1 U7086 ( .A(n6072), .ZN(n6074) );
  AOI22_X1 U7087 ( .A1(n6075), .A2(n6087), .B1(n6074), .B2(n6073), .ZN(n6076)
         );
  OAI211_X1 U7088 ( .C1(n6079), .C2(n6078), .A(n6077), .B(n6076), .ZN(U2819)
         );
  AOI22_X1 U7089 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6080), .B1(n5393), .B2(
        EBX_REG_6__SCAN_IN), .ZN(n6089) );
  INV_X1 U7090 ( .A(n6081), .ZN(n6199) );
  AOI22_X1 U7091 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6098), .B1(n6082), 
        .B2(n6262), .ZN(n6083) );
  NAND2_X1 U7092 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  AOI211_X1 U7093 ( .C1(n6199), .C2(n6087), .A(n6086), .B(n6085), .ZN(n6088)
         );
  OAI211_X1 U7094 ( .C1(n6202), .C2(n6108), .A(n6089), .B(n6088), .ZN(U2821)
         );
  INV_X1 U7095 ( .A(n6090), .ZN(n6091) );
  OAI22_X1 U7096 ( .A1(n6093), .A2(n6685), .B1(n6092), .B2(n6091), .ZN(n6103)
         );
  INV_X1 U7097 ( .A(n6271), .ZN(n6100) );
  NOR3_X1 U7098 ( .A1(n6095), .A2(n6094), .A3(REIP_REG_4__SCAN_IN), .ZN(n6096)
         );
  AOI211_X1 U7099 ( .C1(n6098), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6097), 
        .B(n6096), .ZN(n6099) );
  OAI21_X1 U7100 ( .B1(n6101), .B2(n6100), .A(n6099), .ZN(n6102) );
  AOI211_X1 U7101 ( .C1(n6104), .C2(REIP_REG_4__SCAN_IN), .A(n6103), .B(n6102), 
        .ZN(n6107) );
  NAND2_X1 U7102 ( .A1(n6105), .A2(n6207), .ZN(n6106) );
  OAI211_X1 U7103 ( .C1(n6108), .C2(n6210), .A(n6107), .B(n6106), .ZN(U2823)
         );
  INV_X1 U7104 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6185) );
  AOI22_X1 U7105 ( .A1(n6127), .A2(DATAO_REG_15__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7106 ( .B1(n6185), .B2(n6129), .A(n6109), .ZN(U2908) );
  INV_X1 U7107 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6181) );
  AOI22_X1 U7108 ( .A1(n6127), .A2(DATAO_REG_14__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7109 ( .B1(n6181), .B2(n6129), .A(n6110), .ZN(U2909) );
  AOI22_X1 U7110 ( .A1(n6127), .A2(DATAO_REG_13__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7111 ( .B1(n5561), .B2(n6129), .A(n6111), .ZN(U2910) );
  INV_X1 U7112 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6175) );
  AOI22_X1 U7113 ( .A1(n6127), .A2(DATAO_REG_12__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7114 ( .B1(n6175), .B2(n6129), .A(n6112), .ZN(U2911) );
  INV_X1 U7115 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6172) );
  AOI22_X1 U7116 ( .A1(n6127), .A2(DATAO_REG_10__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7117 ( .B1(n6172), .B2(n6129), .A(n6113), .ZN(U2913) );
  INV_X1 U7118 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6169) );
  AOI22_X1 U7119 ( .A1(n6127), .A2(DATAO_REG_9__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7120 ( .B1(n6169), .B2(n6129), .A(n6114), .ZN(U2914) );
  INV_X1 U7121 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6116) );
  AOI22_X1 U7122 ( .A1(n6127), .A2(DATAO_REG_7__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7123 ( .B1(n6116), .B2(n6129), .A(n6115), .ZN(U2916) );
  INV_X1 U7124 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6118) );
  AOI22_X1 U7125 ( .A1(n6127), .A2(DATAO_REG_6__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7126 ( .B1(n6118), .B2(n6129), .A(n6117), .ZN(U2917) );
  AOI22_X1 U7127 ( .A1(n6127), .A2(DATAO_REG_5__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7128 ( .B1(n6120), .B2(n6129), .A(n6119), .ZN(U2918) );
  AOI22_X1 U7129 ( .A1(n6127), .A2(DATAO_REG_4__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7130 ( .B1(n6122), .B2(n6129), .A(n6121), .ZN(U2919) );
  AOI22_X1 U7131 ( .A1(n6127), .A2(DATAO_REG_3__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7132 ( .B1(n6124), .B2(n6129), .A(n6123), .ZN(U2920) );
  AOI22_X1 U7133 ( .A1(n6127), .A2(DATAO_REG_1__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7134 ( .B1(n6126), .B2(n6129), .A(n6125), .ZN(U2922) );
  AOI22_X1 U7135 ( .A1(n6127), .A2(DATAO_REG_0__SCAN_IN), .B1(n6592), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U7136 ( .B1(n6731), .B2(n6129), .A(n6128), .ZN(U2923) );
  AOI22_X1 U7137 ( .A1(n6608), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6607), .ZN(n6131) );
  OAI21_X1 U7138 ( .B1(n6611), .B2(n6154), .A(n6131), .ZN(U2924) );
  AOI22_X1 U7139 ( .A1(n6608), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6607), .ZN(n6132) );
  OAI21_X1 U7140 ( .B1(n6611), .B2(n6156), .A(n6132), .ZN(U2925) );
  AOI22_X1 U7141 ( .A1(n6608), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6607), .ZN(n6133) );
  OAI21_X1 U7142 ( .B1(n6611), .B2(n6158), .A(n6133), .ZN(U2926) );
  AOI22_X1 U7143 ( .A1(n6608), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6607), .ZN(n6134) );
  OAI21_X1 U7144 ( .B1(n6611), .B2(n6160), .A(n6134), .ZN(U2927) );
  AOI22_X1 U7145 ( .A1(n6608), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6607), .ZN(n6135) );
  OAI21_X1 U7146 ( .B1(n6611), .B2(n6162), .A(n6135), .ZN(U2928) );
  AOI22_X1 U7147 ( .A1(n6608), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6607), .ZN(n6136) );
  OAI21_X1 U7148 ( .B1(n6611), .B2(n6164), .A(n6136), .ZN(U2929) );
  AOI22_X1 U7149 ( .A1(n6608), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6607), .ZN(n6137) );
  OAI21_X1 U7150 ( .B1(n6611), .B2(n6166), .A(n6137), .ZN(U2930) );
  AOI22_X1 U7151 ( .A1(n6608), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6607), .ZN(n6138) );
  OAI21_X1 U7152 ( .B1(n6611), .B2(n6610), .A(n6138), .ZN(U2931) );
  INV_X1 U7153 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6141) );
  AOI21_X1 U7154 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6608), .A(n6139), .ZN(n6140) );
  OAI21_X1 U7155 ( .B1(n6141), .B2(n6184), .A(n6140), .ZN(U2932) );
  INV_X1 U7156 ( .A(DATAI_9_), .ZN(n6142) );
  NOR2_X1 U7157 ( .A1(n6611), .A2(n6142), .ZN(n6167) );
  AOI21_X1 U7158 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6608), .A(n6167), .ZN(n6143) );
  OAI21_X1 U7159 ( .B1(n3803), .B2(n6184), .A(n6143), .ZN(U2933) );
  AOI21_X1 U7160 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6608), .A(n6144), .ZN(
        n6145) );
  OAI21_X1 U7161 ( .B1(n3842), .B2(n6184), .A(n6145), .ZN(U2935) );
  INV_X1 U7162 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6148) );
  INV_X1 U7163 ( .A(DATAI_12_), .ZN(n6146) );
  NOR2_X1 U7164 ( .A1(n6611), .A2(n6146), .ZN(n6173) );
  AOI21_X1 U7165 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6608), .A(n6173), .ZN(
        n6147) );
  OAI21_X1 U7166 ( .B1(n6148), .B2(n6184), .A(n6147), .ZN(U2936) );
  NOR2_X1 U7167 ( .A1(n6611), .A2(n6149), .ZN(n6176) );
  AOI21_X1 U7168 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6608), .A(n6176), .ZN(
        n6150) );
  OAI21_X1 U7169 ( .B1(n3882), .B2(n6184), .A(n6150), .ZN(U2937) );
  INV_X1 U7170 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6656) );
  INV_X1 U7171 ( .A(DATAI_14_), .ZN(n6151) );
  NOR2_X1 U7172 ( .A1(n6611), .A2(n6151), .ZN(n6178) );
  AOI21_X1 U7173 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6608), .A(n6178), .ZN(
        n6152) );
  OAI21_X1 U7174 ( .B1(n6656), .B2(n6184), .A(n6152), .ZN(U2938) );
  AOI22_X1 U7175 ( .A1(n6608), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6607), .ZN(n6153) );
  OAI21_X1 U7176 ( .B1(n6611), .B2(n6154), .A(n6153), .ZN(U2939) );
  AOI22_X1 U7177 ( .A1(n6608), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6607), .ZN(n6155) );
  OAI21_X1 U7178 ( .B1(n6611), .B2(n6156), .A(n6155), .ZN(U2940) );
  AOI22_X1 U7179 ( .A1(n6608), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6607), .ZN(n6157) );
  OAI21_X1 U7180 ( .B1(n6611), .B2(n6158), .A(n6157), .ZN(U2941) );
  AOI22_X1 U7181 ( .A1(n6608), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6607), .ZN(n6159) );
  OAI21_X1 U7182 ( .B1(n6611), .B2(n6160), .A(n6159), .ZN(U2942) );
  AOI22_X1 U7183 ( .A1(n6608), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6607), .ZN(n6161) );
  OAI21_X1 U7184 ( .B1(n6611), .B2(n6162), .A(n6161), .ZN(U2943) );
  AOI22_X1 U7185 ( .A1(n6608), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6607), .ZN(n6163) );
  OAI21_X1 U7186 ( .B1(n6611), .B2(n6164), .A(n6163), .ZN(U2944) );
  AOI22_X1 U7187 ( .A1(n6608), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6607), .ZN(n6165) );
  OAI21_X1 U7188 ( .B1(n6611), .B2(n6166), .A(n6165), .ZN(U2945) );
  AOI21_X1 U7189 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6179), .A(n6167), .ZN(n6168) );
  OAI21_X1 U7190 ( .B1(n6169), .B2(n6184), .A(n6168), .ZN(U2948) );
  AOI21_X1 U7191 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6179), .A(n6170), .ZN(
        n6171) );
  OAI21_X1 U7192 ( .B1(n6172), .B2(n6184), .A(n6171), .ZN(U2949) );
  AOI21_X1 U7193 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6179), .A(n6173), .ZN(
        n6174) );
  OAI21_X1 U7194 ( .B1(n6175), .B2(n6184), .A(n6174), .ZN(U2951) );
  AOI21_X1 U7195 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6179), .A(n6176), .ZN(
        n6177) );
  OAI21_X1 U7196 ( .B1(n5561), .B2(n6184), .A(n6177), .ZN(U2952) );
  AOI21_X1 U7197 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6179), .A(n6178), .ZN(
        n6180) );
  OAI21_X1 U7198 ( .B1(n6181), .B2(n6184), .A(n6180), .ZN(U2953) );
  INV_X1 U7199 ( .A(n6611), .ZN(n6182) );
  AOI22_X1 U7200 ( .A1(n6608), .A2(LWORD_REG_15__SCAN_IN), .B1(n6182), .B2(
        DATAI_15_), .ZN(n6183) );
  OAI21_X1 U7201 ( .B1(n6185), .B2(n6184), .A(n6183), .ZN(U2954) );
  AOI21_X1 U7202 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6186), 
        .ZN(n6191) );
  AOI22_X1 U7203 ( .A1(n6189), .A2(n6217), .B1(n6188), .B2(n6187), .ZN(n6190)
         );
  OAI211_X1 U7204 ( .C1(n6193), .C2(n6192), .A(n6191), .B(n6190), .ZN(U2975)
         );
  AND2_X1 U7205 ( .A1(n6194), .A2(REIP_REG_6__SCAN_IN), .ZN(n6261) );
  AOI21_X1 U7206 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6261), 
        .ZN(n6201) );
  OAI21_X1 U7207 ( .B1(n6197), .B2(n6196), .A(n6195), .ZN(n6198) );
  INV_X1 U7208 ( .A(n6198), .ZN(n6265) );
  AOI22_X1 U7209 ( .A1(n6265), .A2(n6219), .B1(n6217), .B2(n6199), .ZN(n6200)
         );
  OAI211_X1 U7210 ( .C1(n6223), .C2(n6202), .A(n6201), .B(n6200), .ZN(U2980)
         );
  NOR2_X1 U7211 ( .A1(n6211), .A2(n6527), .ZN(n6270) );
  AOI21_X1 U7212 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6270), 
        .ZN(n6209) );
  OR2_X1 U7213 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  AND2_X1 U7214 ( .A1(n6206), .A2(n6205), .ZN(n6272) );
  AOI22_X1 U7215 ( .A1(n6219), .A2(n6272), .B1(n6207), .B2(n6217), .ZN(n6208)
         );
  OAI211_X1 U7216 ( .C1(n6223), .C2(n6210), .A(n6209), .B(n6208), .ZN(U2982)
         );
  NOR2_X1 U7217 ( .A1(n6211), .A2(n6524), .ZN(n6287) );
  AOI21_X1 U7218 ( .B1(n6212), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6287), 
        .ZN(n6221) );
  XOR2_X1 U7219 ( .A(n6213), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6214) );
  XNOR2_X1 U7220 ( .A(n6215), .B(n6214), .ZN(n6293) );
  INV_X1 U7221 ( .A(n6216), .ZN(n6218) );
  AOI22_X1 U7222 ( .A1(n6293), .A2(n6219), .B1(n6218), .B2(n6217), .ZN(n6220)
         );
  OAI211_X1 U7223 ( .C1(n6223), .C2(n6222), .A(n6221), .B(n6220), .ZN(U2984)
         );
  AOI21_X1 U7224 ( .B1(n6225), .B2(n6289), .A(n6224), .ZN(n6234) );
  INV_X1 U7225 ( .A(n6226), .ZN(n6227) );
  OAI21_X1 U7226 ( .B1(n6228), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n6227), 
        .ZN(n6229) );
  AOI22_X1 U7227 ( .A1(n6230), .A2(n6294), .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6229), .ZN(n6233) );
  INV_X1 U7228 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6653) );
  NAND3_X1 U7229 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6653), .A3(n6231), .ZN(n6232) );
  NAND3_X1 U7230 ( .A1(n6234), .A2(n6233), .A3(n6232), .ZN(U3006) );
  AOI22_X1 U7231 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5684), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6235), .ZN(n6243) );
  INV_X1 U7232 ( .A(n6236), .ZN(n6238) );
  AOI21_X1 U7233 ( .B1(n6238), .B2(n6289), .A(n6237), .ZN(n6242) );
  AOI22_X1 U7234 ( .A1(n6240), .A2(n6294), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6239), .ZN(n6241) );
  OAI211_X1 U7235 ( .C1(n6244), .C2(n6243), .A(n6242), .B(n6241), .ZN(U3008)
         );
  AOI21_X1 U7236 ( .B1(n6246), .B2(n6289), .A(n6245), .ZN(n6251) );
  AOI21_X1 U7237 ( .B1(n6259), .B2(n6252), .A(n6247), .ZN(n6248) );
  AOI22_X1 U7238 ( .A1(n6249), .A2(n6294), .B1(n6255), .B2(n6248), .ZN(n6250)
         );
  OAI211_X1 U7239 ( .C1(n6260), .C2(n6252), .A(n6251), .B(n6250), .ZN(U3010)
         );
  AOI21_X1 U7240 ( .B1(n6254), .B2(n6289), .A(n6253), .ZN(n6258) );
  AOI22_X1 U7241 ( .A1(n6256), .A2(n6294), .B1(n6255), .B2(n6259), .ZN(n6257)
         );
  OAI211_X1 U7242 ( .C1(n6260), .C2(n6259), .A(n6258), .B(n6257), .ZN(U3011)
         );
  AOI21_X1 U7243 ( .B1(n6262), .B2(n6289), .A(n6261), .ZN(n6267) );
  NOR3_X1 U7244 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6263), .A3(n6280), 
        .ZN(n6264) );
  AOI21_X1 U7245 ( .B1(n6265), .B2(n6294), .A(n6264), .ZN(n6266) );
  OAI211_X1 U7246 ( .C1(n6269), .C2(n6268), .A(n6267), .B(n6266), .ZN(U3012)
         );
  AOI21_X1 U7247 ( .B1(n6290), .B2(n6292), .A(n6295), .ZN(n6286) );
  AOI21_X1 U7248 ( .B1(n6289), .B2(n6271), .A(n6270), .ZN(n6276) );
  AOI211_X1 U7249 ( .C1(n6285), .C2(n6277), .A(n6292), .B(n6280), .ZN(n6274)
         );
  AOI22_X1 U7250 ( .A1(n6274), .A2(n6273), .B1(n6294), .B2(n6272), .ZN(n6275)
         );
  OAI211_X1 U7251 ( .C1(n6286), .C2(n6277), .A(n6276), .B(n6275), .ZN(U3014)
         );
  AOI21_X1 U7252 ( .B1(n6289), .B2(n6279), .A(n6278), .ZN(n6284) );
  NOR2_X1 U7253 ( .A1(n6292), .A2(n6280), .ZN(n6282) );
  AOI22_X1 U7254 ( .A1(n6282), .A2(n6285), .B1(n6281), .B2(n6294), .ZN(n6283)
         );
  OAI211_X1 U7255 ( .C1(n6286), .C2(n6285), .A(n6284), .B(n6283), .ZN(U3015)
         );
  AOI21_X1 U7256 ( .B1(n6289), .B2(n6288), .A(n6287), .ZN(n6301) );
  OAI221_X1 U7257 ( .B1(n6292), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .C1(n6292), .C2(n6291), .A(n6290), .ZN(n6300) );
  AOI22_X1 U7258 ( .A1(n6295), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6294), 
        .B2(n6293), .ZN(n6299) );
  OR3_X1 U7259 ( .A1(n6297), .A2(n6296), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6298) );
  NAND4_X1 U7260 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(U3016)
         );
  NOR2_X1 U7261 ( .A1(n6303), .A2(n6302), .ZN(U3019) );
  INV_X1 U7262 ( .A(n6314), .ZN(n6305) );
  NAND2_X1 U7263 ( .A1(n6305), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6337) );
  NOR2_X1 U7264 ( .A1(n6439), .A2(n6337), .ZN(n6306) );
  AOI21_X1 U7265 ( .B1(n6339), .B2(n6403), .A(n6306), .ZN(n6318) );
  OAI21_X1 U7266 ( .B1(n6307), .B2(n6443), .A(n6442), .ZN(n6316) );
  INV_X1 U7267 ( .A(n6337), .ZN(n6308) );
  AOI21_X1 U7268 ( .B1(n6309), .B2(n6446), .A(n6308), .ZN(n6315) );
  INV_X1 U7269 ( .A(n6315), .ZN(n6313) );
  AOI21_X1 U7270 ( .B1(n6311), .B2(n6593), .A(n6310), .ZN(n6448) );
  OAI211_X1 U7271 ( .C1(n6316), .C2(n6313), .A(n6448), .B(n6312), .ZN(n6341)
         );
  OAI22_X1 U7272 ( .A1(n6316), .A2(n6315), .B1(n5034), .B2(n6314), .ZN(n6340)
         );
  AOI22_X1 U7273 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6341), .B1(n6454), 
        .B2(n6340), .ZN(n6317) );
  OAI211_X1 U7274 ( .C1(n6457), .C2(n6383), .A(n6318), .B(n6317), .ZN(U3044)
         );
  NOR2_X1 U7275 ( .A1(n6458), .A2(n6337), .ZN(n6319) );
  AOI21_X1 U7276 ( .B1(n6339), .B2(n6407), .A(n6319), .ZN(n6321) );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6341), .B1(n6461), 
        .B2(n6340), .ZN(n6320) );
  OAI211_X1 U7278 ( .C1(n6459), .C2(n6383), .A(n6321), .B(n6320), .ZN(U3045)
         );
  NOR2_X1 U7279 ( .A1(n6465), .A2(n6337), .ZN(n6322) );
  AOI21_X1 U7280 ( .B1(n6339), .B2(n6411), .A(n6322), .ZN(n6324) );
  AOI22_X1 U7281 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6341), .B1(n6468), 
        .B2(n6340), .ZN(n6323) );
  OAI211_X1 U7282 ( .C1(n6466), .C2(n6383), .A(n6324), .B(n6323), .ZN(U3046)
         );
  NOR2_X1 U7283 ( .A1(n6472), .A2(n6337), .ZN(n6325) );
  AOI21_X1 U7284 ( .B1(n6339), .B2(n6415), .A(n6325), .ZN(n6327) );
  AOI22_X1 U7285 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6341), .B1(n6475), 
        .B2(n6340), .ZN(n6326) );
  OAI211_X1 U7286 ( .C1(n6478), .C2(n6383), .A(n6327), .B(n6326), .ZN(U3047)
         );
  NOR2_X1 U7287 ( .A1(n6479), .A2(n6337), .ZN(n6328) );
  AOI21_X1 U7288 ( .B1(n6339), .B2(n6419), .A(n6328), .ZN(n6330) );
  AOI22_X1 U7289 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6341), .B1(n6482), 
        .B2(n6340), .ZN(n6329) );
  OAI211_X1 U7290 ( .C1(n6485), .C2(n6383), .A(n6330), .B(n6329), .ZN(U3048)
         );
  NOR2_X1 U7291 ( .A1(n6486), .A2(n6337), .ZN(n6331) );
  AOI21_X1 U7292 ( .B1(n6339), .B2(n6423), .A(n6331), .ZN(n6333) );
  AOI22_X1 U7293 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6341), .B1(n6489), 
        .B2(n6340), .ZN(n6332) );
  OAI211_X1 U7294 ( .C1(n6487), .C2(n6383), .A(n6333), .B(n6332), .ZN(U3049)
         );
  NOR2_X1 U7295 ( .A1(n6493), .A2(n6337), .ZN(n6334) );
  AOI21_X1 U7296 ( .B1(n6339), .B2(n6427), .A(n6334), .ZN(n6336) );
  AOI22_X1 U7297 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6341), .B1(n6496), 
        .B2(n6340), .ZN(n6335) );
  OAI211_X1 U7298 ( .C1(n6499), .C2(n6383), .A(n6336), .B(n6335), .ZN(U3050)
         );
  NOR2_X1 U7299 ( .A1(n6501), .A2(n6337), .ZN(n6338) );
  AOI21_X1 U7300 ( .B1(n6339), .B2(n6434), .A(n6338), .ZN(n6343) );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6341), .B1(n6506), 
        .B2(n6340), .ZN(n6342) );
  OAI211_X1 U7302 ( .C1(n6502), .C2(n6383), .A(n6343), .B(n6342), .ZN(U3051)
         );
  OAI33_X1 U7303 ( .A1(n6347), .A2(n6346), .A3(n6593), .B1(n6345), .B2(n6387), 
        .B3(n6344), .ZN(n6377) );
  INV_X1 U7304 ( .A(n6439), .ZN(n6392) );
  NAND2_X1 U7305 ( .A1(n6348), .A2(n6390), .ZN(n6350) );
  INV_X1 U7306 ( .A(n6350), .ZN(n6376) );
  AOI22_X1 U7307 ( .A1(n6377), .A2(n6454), .B1(n6392), .B2(n6376), .ZN(n6357)
         );
  OAI21_X1 U7308 ( .B1(n6383), .B2(n6394), .A(n6349), .ZN(n6353) );
  AOI21_X1 U7309 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6350), .A(n6396), .ZN(
        n6351) );
  AOI22_X1 U7310 ( .A1(n6380), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6355), 
        .B2(n6378), .ZN(n6356) );
  OAI211_X1 U7311 ( .C1(n6440), .C2(n6383), .A(n6357), .B(n6356), .ZN(U3052)
         );
  INV_X1 U7312 ( .A(n6458), .ZN(n6406) );
  AOI22_X1 U7313 ( .A1(n6377), .A2(n6461), .B1(n6406), .B2(n6376), .ZN(n6360)
         );
  AOI22_X1 U7314 ( .A1(n6380), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6358), 
        .B2(n6378), .ZN(n6359) );
  OAI211_X1 U7315 ( .C1(n6464), .C2(n6383), .A(n6360), .B(n6359), .ZN(U3053)
         );
  INV_X1 U7316 ( .A(n6465), .ZN(n6410) );
  AOI22_X1 U7317 ( .A1(n2994), .A2(n6468), .B1(n6410), .B2(n6376), .ZN(n6363)
         );
  AOI22_X1 U7318 ( .A1(n6380), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6361), 
        .B2(n6378), .ZN(n6362) );
  OAI211_X1 U7319 ( .C1(n6471), .C2(n6383), .A(n6363), .B(n6362), .ZN(U3054)
         );
  INV_X1 U7320 ( .A(n6472), .ZN(n6414) );
  AOI22_X1 U7321 ( .A1(n6377), .A2(n6475), .B1(n6414), .B2(n6376), .ZN(n6366)
         );
  AOI22_X1 U7322 ( .A1(n6380), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6364), 
        .B2(n6378), .ZN(n6365) );
  OAI211_X1 U7323 ( .C1(n6473), .C2(n6383), .A(n6366), .B(n6365), .ZN(U3055)
         );
  INV_X1 U7324 ( .A(n6479), .ZN(n6418) );
  AOI22_X1 U7325 ( .A1(n2994), .A2(n6482), .B1(n6418), .B2(n6376), .ZN(n6369)
         );
  AOI22_X1 U7326 ( .A1(n6380), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6367), 
        .B2(n6378), .ZN(n6368) );
  OAI211_X1 U7327 ( .C1(n6480), .C2(n6383), .A(n6369), .B(n6368), .ZN(U3056)
         );
  INV_X1 U7328 ( .A(n6486), .ZN(n6422) );
  AOI22_X1 U7329 ( .A1(n2994), .A2(n6489), .B1(n6422), .B2(n6376), .ZN(n6372)
         );
  AOI22_X1 U7330 ( .A1(n6380), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6370), 
        .B2(n6378), .ZN(n6371) );
  OAI211_X1 U7331 ( .C1(n6492), .C2(n6383), .A(n6372), .B(n6371), .ZN(U3057)
         );
  INV_X1 U7332 ( .A(n6493), .ZN(n6426) );
  AOI22_X1 U7333 ( .A1(n6377), .A2(n6496), .B1(n6426), .B2(n6376), .ZN(n6375)
         );
  AOI22_X1 U7334 ( .A1(n6380), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6373), 
        .B2(n6378), .ZN(n6374) );
  OAI211_X1 U7335 ( .C1(n6494), .C2(n6383), .A(n6375), .B(n6374), .ZN(U3058)
         );
  INV_X1 U7336 ( .A(n6501), .ZN(n6431) );
  AOI22_X1 U7337 ( .A1(n2994), .A2(n6506), .B1(n6431), .B2(n6376), .ZN(n6382)
         );
  AOI22_X1 U7338 ( .A1(n6380), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6379), 
        .B2(n6378), .ZN(n6381) );
  OAI211_X1 U7339 ( .C1(n6511), .C2(n6383), .A(n6382), .B(n6381), .ZN(U3059)
         );
  NAND2_X1 U7340 ( .A1(n6384), .A2(n6442), .ZN(n6389) );
  INV_X1 U7341 ( .A(n6385), .ZN(n6386) );
  OAI22_X1 U7342 ( .A1(n6389), .A2(n6388), .B1(n6387), .B2(n6386), .ZN(n6432)
         );
  NAND2_X1 U7343 ( .A1(n6391), .A2(n6390), .ZN(n6397) );
  INV_X1 U7344 ( .A(n6397), .ZN(n6430) );
  AOI22_X1 U7345 ( .A1(n6432), .A2(n6454), .B1(n6392), .B2(n6430), .ZN(n6405)
         );
  NOR2_X1 U7346 ( .A1(n6393), .A2(n6593), .ZN(n6395) );
  AOI21_X1 U7347 ( .B1(n6395), .B2(n6402), .A(n6394), .ZN(n6401) );
  AOI211_X1 U7348 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6397), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6396), .ZN(n6398) );
  AOI22_X1 U7349 ( .A1(n6435), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6403), 
        .B2(n6433), .ZN(n6404) );
  OAI211_X1 U7350 ( .C1(n6457), .C2(n6438), .A(n6405), .B(n6404), .ZN(U3068)
         );
  AOI22_X1 U7351 ( .A1(n6432), .A2(n6461), .B1(n6406), .B2(n6430), .ZN(n6409)
         );
  AOI22_X1 U7352 ( .A1(n6435), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6407), 
        .B2(n6433), .ZN(n6408) );
  OAI211_X1 U7353 ( .C1(n6459), .C2(n6438), .A(n6409), .B(n6408), .ZN(U3069)
         );
  AOI22_X1 U7354 ( .A1(n6432), .A2(n6468), .B1(n6410), .B2(n6430), .ZN(n6413)
         );
  AOI22_X1 U7355 ( .A1(n6435), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6411), 
        .B2(n6433), .ZN(n6412) );
  OAI211_X1 U7356 ( .C1(n6466), .C2(n6438), .A(n6413), .B(n6412), .ZN(U3070)
         );
  AOI22_X1 U7357 ( .A1(n6432), .A2(n6475), .B1(n6414), .B2(n6430), .ZN(n6417)
         );
  AOI22_X1 U7358 ( .A1(n6435), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6415), 
        .B2(n6433), .ZN(n6416) );
  OAI211_X1 U7359 ( .C1(n6478), .C2(n6438), .A(n6417), .B(n6416), .ZN(U3071)
         );
  AOI22_X1 U7360 ( .A1(n6432), .A2(n6482), .B1(n6418), .B2(n6430), .ZN(n6421)
         );
  AOI22_X1 U7361 ( .A1(n6435), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6419), 
        .B2(n6433), .ZN(n6420) );
  OAI211_X1 U7362 ( .C1(n6485), .C2(n6438), .A(n6421), .B(n6420), .ZN(U3072)
         );
  AOI22_X1 U7363 ( .A1(n6432), .A2(n6489), .B1(n6422), .B2(n6430), .ZN(n6425)
         );
  AOI22_X1 U7364 ( .A1(n6435), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6423), 
        .B2(n6433), .ZN(n6424) );
  OAI211_X1 U7365 ( .C1(n6487), .C2(n6438), .A(n6425), .B(n6424), .ZN(U3073)
         );
  AOI22_X1 U7366 ( .A1(n6432), .A2(n6496), .B1(n6426), .B2(n6430), .ZN(n6429)
         );
  AOI22_X1 U7367 ( .A1(n6435), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6427), 
        .B2(n6433), .ZN(n6428) );
  OAI211_X1 U7368 ( .C1(n6499), .C2(n6438), .A(n6429), .B(n6428), .ZN(U3074)
         );
  AOI22_X1 U7369 ( .A1(n6432), .A2(n6506), .B1(n6431), .B2(n6430), .ZN(n6437)
         );
  AOI22_X1 U7370 ( .A1(n6435), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6434), 
        .B2(n6433), .ZN(n6436) );
  OAI211_X1 U7371 ( .C1(n6502), .C2(n6438), .A(n6437), .B(n6436), .ZN(U3075)
         );
  NAND2_X1 U7372 ( .A1(n6450), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6500) );
  OAI22_X1 U7373 ( .A1(n6510), .A2(n6440), .B1(n6439), .B2(n6500), .ZN(n6441)
         );
  INV_X1 U7374 ( .A(n6441), .ZN(n6456) );
  OAI21_X1 U7375 ( .B1(n6444), .B2(n6443), .A(n6442), .ZN(n6453) );
  INV_X1 U7376 ( .A(n6500), .ZN(n6445) );
  AOI21_X1 U7377 ( .B1(n6447), .B2(n6446), .A(n6445), .ZN(n6452) );
  INV_X1 U7378 ( .A(n6452), .ZN(n6449) );
  OAI211_X1 U7379 ( .C1(n6453), .C2(n6449), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6448), .ZN(n6507) );
  INV_X1 U7380 ( .A(n6450), .ZN(n6451) );
  OAI22_X1 U7381 ( .A1(n6453), .A2(n6452), .B1(n5034), .B2(n6451), .ZN(n6505)
         );
  AOI22_X1 U7382 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6507), .B1(n6454), 
        .B2(n6505), .ZN(n6455) );
  OAI211_X1 U7383 ( .C1(n6457), .C2(n6503), .A(n6456), .B(n6455), .ZN(U3108)
         );
  OAI22_X1 U7384 ( .A1(n6503), .A2(n6459), .B1(n6458), .B2(n6500), .ZN(n6460)
         );
  INV_X1 U7385 ( .A(n6460), .ZN(n6463) );
  AOI22_X1 U7386 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6507), .B1(n6461), 
        .B2(n6505), .ZN(n6462) );
  OAI211_X1 U7387 ( .C1(n6464), .C2(n6510), .A(n6463), .B(n6462), .ZN(U3109)
         );
  OAI22_X1 U7388 ( .A1(n6503), .A2(n6466), .B1(n6465), .B2(n6500), .ZN(n6467)
         );
  INV_X1 U7389 ( .A(n6467), .ZN(n6470) );
  AOI22_X1 U7390 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6507), .B1(n6468), 
        .B2(n6505), .ZN(n6469) );
  OAI211_X1 U7391 ( .C1(n6471), .C2(n6510), .A(n6470), .B(n6469), .ZN(U3110)
         );
  OAI22_X1 U7392 ( .A1(n6510), .A2(n6473), .B1(n6472), .B2(n6500), .ZN(n6474)
         );
  INV_X1 U7393 ( .A(n6474), .ZN(n6477) );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6507), .B1(n6475), 
        .B2(n6505), .ZN(n6476) );
  OAI211_X1 U7395 ( .C1(n6478), .C2(n6503), .A(n6477), .B(n6476), .ZN(U3111)
         );
  OAI22_X1 U7396 ( .A1(n6510), .A2(n6480), .B1(n6479), .B2(n6500), .ZN(n6481)
         );
  INV_X1 U7397 ( .A(n6481), .ZN(n6484) );
  AOI22_X1 U7398 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6507), .B1(n6482), 
        .B2(n6505), .ZN(n6483) );
  OAI211_X1 U7399 ( .C1(n6485), .C2(n6503), .A(n6484), .B(n6483), .ZN(U3112)
         );
  OAI22_X1 U7400 ( .A1(n6503), .A2(n6487), .B1(n6486), .B2(n6500), .ZN(n6488)
         );
  INV_X1 U7401 ( .A(n6488), .ZN(n6491) );
  AOI22_X1 U7402 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6507), .B1(n6489), 
        .B2(n6505), .ZN(n6490) );
  OAI211_X1 U7403 ( .C1(n6492), .C2(n6510), .A(n6491), .B(n6490), .ZN(U3113)
         );
  OAI22_X1 U7404 ( .A1(n6510), .A2(n6494), .B1(n6493), .B2(n6500), .ZN(n6495)
         );
  INV_X1 U7405 ( .A(n6495), .ZN(n6498) );
  AOI22_X1 U7406 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6507), .B1(n6496), 
        .B2(n6505), .ZN(n6497) );
  OAI211_X1 U7407 ( .C1(n6499), .C2(n6503), .A(n6498), .B(n6497), .ZN(U3114)
         );
  OAI22_X1 U7408 ( .A1(n6503), .A2(n6502), .B1(n6501), .B2(n6500), .ZN(n6504)
         );
  INV_X1 U7409 ( .A(n6504), .ZN(n6509) );
  AOI22_X1 U7410 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6507), .B1(n6506), 
        .B2(n6505), .ZN(n6508) );
  OAI211_X1 U7411 ( .C1(n6511), .C2(n6510), .A(n6509), .B(n6508), .ZN(U3115)
         );
  OAI211_X1 U7412 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6512), .ZN(n6521) );
  NOR3_X1 U7413 ( .A1(n6514), .A2(READY_N), .A3(n6513), .ZN(n6516) );
  OAI21_X1 U7414 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6519) );
  AND2_X1 U7415 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NAND2_X1 U7416 ( .A1(n6521), .A2(n6520), .ZN(U3149) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6522), .ZN(U3151) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6522), .ZN(U3152) );
  NOR2_X1 U7419 ( .A1(n6576), .A2(n6673), .ZN(U3153) );
  NOR2_X1 U7420 ( .A1(n6576), .A2(n6627), .ZN(U3154) );
  INV_X1 U7421 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U7422 ( .A1(n6576), .A2(n6753), .ZN(U3155) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6522), .ZN(U3156) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6522), .ZN(U3157) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6522), .ZN(U3158) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6522), .ZN(U3159) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6522), .ZN(U3160) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6522), .ZN(U3161) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6522), .ZN(U3162) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6522), .ZN(U3163) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6522), .ZN(U3164) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6522), .ZN(U3165) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6522), .ZN(U3166) );
  AND2_X1 U7434 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6522), .ZN(U3167) );
  AND2_X1 U7435 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6522), .ZN(U3168) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6522), .ZN(U3169) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6522), .ZN(U3170) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6522), .ZN(U3171) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6522), .ZN(U3172) );
  AND2_X1 U7440 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6522), .ZN(U3173) );
  AND2_X1 U7441 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6522), .ZN(U3174) );
  AND2_X1 U7442 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6522), .ZN(U3175) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6522), .ZN(U3176) );
  AND2_X1 U7444 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6522), .ZN(U3177) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6522), .ZN(U3178) );
  AND2_X1 U7446 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6522), .ZN(U3179) );
  AND2_X1 U7447 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6522), .ZN(U3180) );
  NOR2_X1 U7448 ( .A1(n6606), .A2(STATE_REG_2__SCAN_IN), .ZN(n6564) );
  INV_X1 U7449 ( .A(n6564), .ZN(n6572) );
  AOI22_X1 U7450 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6588), .ZN(n6523) );
  OAI21_X1 U7451 ( .B1(n6524), .B2(n6572), .A(n6523), .ZN(U3184) );
  AOI222_X1 U7452 ( .A1(n6570), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6606), .C1(REIP_REG_3__SCAN_IN), .C2(
        n6564), .ZN(n6525) );
  INV_X1 U7453 ( .A(n6525), .ZN(U3185) );
  AOI22_X1 U7454 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6588), .ZN(n6526) );
  OAI21_X1 U7455 ( .B1(n6527), .B2(n6572), .A(n6526), .ZN(U3186) );
  AOI22_X1 U7456 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6588), .ZN(n6528) );
  OAI21_X1 U7457 ( .B1(n6529), .B2(n6572), .A(n6528), .ZN(U3187) );
  AOI22_X1 U7458 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6606), .ZN(n6530) );
  OAI21_X1 U7459 ( .B1(n6749), .B2(n6572), .A(n6530), .ZN(U3188) );
  AOI22_X1 U7460 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6606), .ZN(n6531) );
  OAI21_X1 U7461 ( .B1(n6533), .B2(n6572), .A(n6531), .ZN(U3189) );
  AOI22_X1 U7462 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6606), .ZN(n6532) );
  OAI21_X1 U7463 ( .B1(n6533), .B2(n6569), .A(n6532), .ZN(U3190) );
  AOI22_X1 U7464 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6606), .ZN(n6534) );
  OAI21_X1 U7465 ( .B1(n6535), .B2(n6572), .A(n6534), .ZN(U3191) );
  INV_X1 U7466 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6679) );
  OAI222_X1 U7467 ( .A1(n6569), .A2(n6535), .B1(n6679), .B2(n6546), .C1(n5700), 
        .C2(n6572), .ZN(U3192) );
  AOI22_X1 U7468 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6606), .ZN(n6536) );
  OAI21_X1 U7469 ( .B1(n5700), .B2(n6569), .A(n6536), .ZN(U3193) );
  AOI22_X1 U7470 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6606), .ZN(n6537) );
  OAI21_X1 U7471 ( .B1(n6538), .B2(n6569), .A(n6537), .ZN(U3194) );
  AOI22_X1 U7472 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6606), .ZN(n6539) );
  OAI21_X1 U7473 ( .B1(n6540), .B2(n6569), .A(n6539), .ZN(U3195) );
  AOI22_X1 U7474 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6606), .ZN(n6541) );
  OAI21_X1 U7475 ( .B1(n6542), .B2(n6572), .A(n6541), .ZN(U3196) );
  INV_X1 U7476 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6655) );
  OAI222_X1 U7477 ( .A1(n6572), .A2(n6543), .B1(n6655), .B2(n6546), .C1(n6542), 
        .C2(n6569), .ZN(U3197) );
  AOI22_X1 U7478 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6606), .ZN(n6544) );
  OAI21_X1 U7479 ( .B1(n6547), .B2(n6572), .A(n6544), .ZN(U3198) );
  INV_X1 U7480 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6631) );
  OAI222_X1 U7481 ( .A1(n6569), .A2(n6547), .B1(n6631), .B2(n6546), .C1(n6545), 
        .C2(n6572), .ZN(U3199) );
  AOI22_X1 U7482 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6588), .ZN(n6548) );
  OAI21_X1 U7483 ( .B1(n6550), .B2(n6572), .A(n6548), .ZN(U3200) );
  AOI22_X1 U7484 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6588), .ZN(n6549) );
  OAI21_X1 U7485 ( .B1(n6550), .B2(n6569), .A(n6549), .ZN(U3201) );
  INV_X1 U7486 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6553) );
  AOI22_X1 U7487 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6588), .ZN(n6551) );
  OAI21_X1 U7488 ( .B1(n6553), .B2(n6572), .A(n6551), .ZN(U3202) );
  AOI22_X1 U7489 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6588), .ZN(n6552) );
  OAI21_X1 U7490 ( .B1(n6553), .B2(n6569), .A(n6552), .ZN(U3203) );
  AOI22_X1 U7491 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6588), .ZN(n6554) );
  OAI21_X1 U7492 ( .B1(n6555), .B2(n6572), .A(n6554), .ZN(U3204) );
  AOI22_X1 U7493 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6588), .ZN(n6556) );
  OAI21_X1 U7494 ( .B1(n6557), .B2(n6572), .A(n6556), .ZN(U3205) );
  AOI22_X1 U7495 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6588), .ZN(n6558) );
  OAI21_X1 U7496 ( .B1(n6559), .B2(n6572), .A(n6558), .ZN(U3206) );
  AOI22_X1 U7497 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6588), .ZN(n6560) );
  OAI21_X1 U7498 ( .B1(n6561), .B2(n6572), .A(n6560), .ZN(U3207) );
  INV_X1 U7499 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U7500 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6588), .ZN(n6562) );
  OAI21_X1 U7501 ( .B1(n6665), .B2(n6572), .A(n6562), .ZN(U3208) );
  AOI22_X1 U7502 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6588), .ZN(n6563) );
  OAI21_X1 U7503 ( .B1(n6665), .B2(n6569), .A(n6563), .ZN(U3209) );
  AOI22_X1 U7504 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6564), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6588), .ZN(n6565) );
  OAI21_X1 U7505 ( .B1(n6566), .B2(n6569), .A(n6565), .ZN(U3210) );
  AOI22_X1 U7506 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6588), .ZN(n6567) );
  OAI21_X1 U7507 ( .B1(n6709), .B2(n6572), .A(n6567), .ZN(U3211) );
  INV_X1 U7508 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U7509 ( .A1(n6569), .A2(n6709), .B1(n6641), .B2(n6546), .C1(n6568), 
        .C2(n6572), .ZN(U3212) );
  AOI22_X1 U7510 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6570), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6588), .ZN(n6571) );
  OAI21_X1 U7511 ( .B1(n6573), .B2(n6572), .A(n6571), .ZN(U3213) );
  MUX2_X1 U7512 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6606), .Z(U3445) );
  MUX2_X1 U7513 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6606), .Z(U3446) );
  MUX2_X1 U7514 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6606), .Z(U3447) );
  MUX2_X1 U7515 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6606), .Z(U3448) );
  OAI21_X1 U7516 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6576), .A(n6575), .ZN(
        n6574) );
  INV_X1 U7517 ( .A(n6574), .ZN(U3451) );
  OAI21_X1 U7518 ( .B1(n6576), .B2(n6651), .A(n6575), .ZN(U3452) );
  OAI211_X1 U7519 ( .C1(n6577), .C2(n6585), .A(n6651), .B(n6586), .ZN(n6582)
         );
  INV_X1 U7520 ( .A(n6584), .ZN(n6580) );
  OAI21_X1 U7521 ( .B1(n6585), .B2(n6578), .A(n6580), .ZN(n6579) );
  OAI21_X1 U7522 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6580), .A(n6579), .ZN(
        n6581) );
  NAND2_X1 U7523 ( .A1(n6582), .A2(n6581), .ZN(U3468) );
  INV_X1 U7524 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6583) );
  AOI22_X1 U7525 ( .A1(n6586), .A2(n6585), .B1(n6584), .B2(n6583), .ZN(U3469)
         );
  NAND2_X1 U7526 ( .A1(n6588), .A2(W_R_N_REG_SCAN_IN), .ZN(n6587) );
  OAI21_X1 U7527 ( .B1(n6588), .B2(READREQUEST_REG_SCAN_IN), .A(n6587), .ZN(
        U3470) );
  MUX2_X1 U7528 ( .A(MORE_REG_SCAN_IN), .B(n6590), .S(n6589), .Z(U3471) );
  NAND2_X1 U7529 ( .A1(n6592), .A2(n6591), .ZN(n6594) );
  NAND2_X1 U7530 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  NOR3_X1 U7531 ( .A1(n6597), .A2(n6596), .A3(n6595), .ZN(n6605) );
  INV_X1 U7532 ( .A(n6598), .ZN(n6599) );
  OAI211_X1 U7533 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6600), .A(n6599), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6602) );
  AOI21_X1 U7534 ( .B1(n6602), .B2(STATE2_REG_0__SCAN_IN), .A(n6601), .ZN(
        n6604) );
  NAND2_X1 U7535 ( .A1(n6605), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6603) );
  OAI21_X1 U7536 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(U3472) );
  MUX2_X1 U7537 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6606), .Z(U3473) );
  AOI22_X1 U7538 ( .A1(n6608), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6607), .ZN(n6609) );
  OAI21_X1 U7539 ( .B1(n6611), .B2(n6610), .A(n6609), .ZN(n6770) );
  INV_X1 U7540 ( .A(DATAI_27_), .ZN(n6614) );
  INV_X1 U7541 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6613) );
  AOI22_X1 U7542 ( .A1(n6614), .A2(keyinput7), .B1(n6613), .B2(keyinput46), 
        .ZN(n6612) );
  OAI221_X1 U7543 ( .B1(n6614), .B2(keyinput7), .C1(n6613), .C2(keyinput46), 
        .A(n6612), .ZN(n6625) );
  INV_X1 U7544 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6617) );
  AOI22_X1 U7545 ( .A1(n6617), .A2(keyinput22), .B1(keyinput16), .B2(n6616), 
        .ZN(n6615) );
  OAI221_X1 U7546 ( .B1(n6617), .B2(keyinput22), .C1(n6616), .C2(keyinput16), 
        .A(n6615), .ZN(n6624) );
  INV_X1 U7547 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6619) );
  AOI22_X1 U7548 ( .A1(n6619), .A2(keyinput45), .B1(keyinput58), .B2(n6750), 
        .ZN(n6618) );
  OAI221_X1 U7549 ( .B1(n6619), .B2(keyinput45), .C1(n6750), .C2(keyinput58), 
        .A(n6618), .ZN(n6623) );
  XNOR2_X1 U7550 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput29), .ZN(n6621)
         );
  XNOR2_X1 U7551 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .B(keyinput38), .ZN(n6620) );
  NAND2_X1 U7552 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  NOR4_X1 U7553 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6768)
         );
  AOI22_X1 U7554 ( .A1(n6628), .A2(keyinput8), .B1(keyinput21), .B2(n6627), 
        .ZN(n6626) );
  OAI221_X1 U7555 ( .B1(n6628), .B2(keyinput8), .C1(n6627), .C2(keyinput21), 
        .A(n6626), .ZN(n6638) );
  INV_X1 U7556 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6630) );
  AOI22_X1 U7557 ( .A1(n6631), .A2(keyinput44), .B1(n6630), .B2(keyinput1), 
        .ZN(n6629) );
  OAI221_X1 U7558 ( .B1(n6631), .B2(keyinput44), .C1(n6630), .C2(keyinput1), 
        .A(n6629), .ZN(n6637) );
  XNOR2_X1 U7559 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(keyinput49), .ZN(
        n6634) );
  XNOR2_X1 U7560 ( .A(STATE2_REG_3__SCAN_IN), .B(keyinput31), .ZN(n6633) );
  XNOR2_X1 U7561 ( .A(keyinput15), .B(EAX_REG_16__SCAN_IN), .ZN(n6632) );
  NAND3_X1 U7562 ( .A1(n6634), .A2(n6633), .A3(n6632), .ZN(n6636) );
  XNOR2_X1 U7563 ( .A(n6737), .B(keyinput9), .ZN(n6635) );
  NOR4_X1 U7564 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6767)
         );
  INV_X1 U7565 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7566 ( .A1(n6743), .A2(keyinput60), .B1(keyinput28), .B2(n6752), 
        .ZN(n6639) );
  OAI221_X1 U7567 ( .B1(n6743), .B2(keyinput60), .C1(n6752), .C2(keyinput28), 
        .A(n6639), .ZN(n6724) );
  INV_X1 U7568 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6642) );
  AOI22_X1 U7569 ( .A1(n6642), .A2(keyinput25), .B1(keyinput57), .B2(n6641), 
        .ZN(n6640) );
  OAI221_X1 U7570 ( .B1(n6642), .B2(keyinput25), .C1(n6641), .C2(keyinput57), 
        .A(n6640), .ZN(n6723) );
  INV_X1 U7571 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6644) );
  OAI22_X1 U7572 ( .A1(n6644), .A2(keyinput39), .B1(n6749), .B2(keyinput62), 
        .ZN(n6643) );
  AOI221_X1 U7573 ( .B1(n6644), .B2(keyinput39), .C1(keyinput62), .C2(n6749), 
        .A(n6643), .ZN(n6663) );
  INV_X1 U7574 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6646) );
  OAI22_X1 U7575 ( .A1(n4495), .A2(keyinput30), .B1(n6646), .B2(keyinput5), 
        .ZN(n6645) );
  AOI221_X1 U7576 ( .B1(n4495), .B2(keyinput30), .C1(keyinput5), .C2(n6646), 
        .A(n6645), .ZN(n6662) );
  INV_X1 U7577 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7578 ( .A1(n6649), .A2(keyinput13), .B1(n6648), .B2(keyinput42), 
        .ZN(n6647) );
  OAI221_X1 U7579 ( .B1(n6649), .B2(keyinput13), .C1(n6648), .C2(keyinput42), 
        .A(n6647), .ZN(n6660) );
  AOI22_X1 U7580 ( .A1(n6651), .A2(keyinput27), .B1(keyinput33), .B2(n6751), 
        .ZN(n6650) );
  OAI221_X1 U7581 ( .B1(n6651), .B2(keyinput27), .C1(n6751), .C2(keyinput33), 
        .A(n6650), .ZN(n6659) );
  AOI22_X1 U7582 ( .A1(n6653), .A2(keyinput2), .B1(keyinput10), .B2(n6753), 
        .ZN(n6652) );
  OAI221_X1 U7583 ( .B1(n6653), .B2(keyinput2), .C1(n6753), .C2(keyinput10), 
        .A(n6652), .ZN(n6658) );
  AOI22_X1 U7584 ( .A1(n6656), .A2(keyinput61), .B1(keyinput53), .B2(n6655), 
        .ZN(n6654) );
  OAI221_X1 U7585 ( .B1(n6656), .B2(keyinput61), .C1(n6655), .C2(keyinput53), 
        .A(n6654), .ZN(n6657) );
  NOR4_X1 U7586 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6661)
         );
  NAND3_X1 U7587 ( .A1(n6663), .A2(n6662), .A3(n6661), .ZN(n6722) );
  INV_X1 U7588 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U7589 ( .A1(n6666), .A2(keyinput47), .B1(keyinput50), .B2(n6665), 
        .ZN(n6664) );
  OAI221_X1 U7590 ( .B1(n6666), .B2(keyinput47), .C1(n6665), .C2(keyinput50), 
        .A(n6664), .ZN(n6677) );
  INV_X1 U7591 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7592 ( .A1(n6668), .A2(keyinput20), .B1(n6744), .B2(keyinput4), 
        .ZN(n6667) );
  OAI221_X1 U7593 ( .B1(n6668), .B2(keyinput20), .C1(n6744), .C2(keyinput4), 
        .A(n6667), .ZN(n6676) );
  INV_X1 U7594 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7595 ( .A1(n6671), .A2(keyinput55), .B1(n6670), .B2(keyinput26), 
        .ZN(n6669) );
  OAI221_X1 U7596 ( .B1(n6671), .B2(keyinput55), .C1(n6670), .C2(keyinput26), 
        .A(n6669), .ZN(n6675) );
  AOI22_X1 U7597 ( .A1(n4497), .A2(keyinput40), .B1(keyinput41), .B2(n6673), 
        .ZN(n6672) );
  OAI221_X1 U7598 ( .B1(n4497), .B2(keyinput40), .C1(n6673), .C2(keyinput41), 
        .A(n6672), .ZN(n6674) );
  NOR4_X1 U7599 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6720)
         );
  INV_X1 U7600 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6680) );
  AOI22_X1 U7601 ( .A1(n6680), .A2(keyinput43), .B1(keyinput34), .B2(n6679), 
        .ZN(n6678) );
  OAI221_X1 U7602 ( .B1(n6680), .B2(keyinput43), .C1(n6679), .C2(keyinput34), 
        .A(n6678), .ZN(n6691) );
  INV_X1 U7603 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6682) );
  AOI22_X1 U7604 ( .A1(n6682), .A2(keyinput63), .B1(keyinput11), .B2(n6742), 
        .ZN(n6681) );
  OAI221_X1 U7605 ( .B1(n6682), .B2(keyinput63), .C1(n6742), .C2(keyinput11), 
        .A(n6681), .ZN(n6690) );
  INV_X1 U7606 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U7607 ( .A1(n6685), .A2(keyinput0), .B1(keyinput56), .B2(n6684), 
        .ZN(n6683) );
  OAI221_X1 U7608 ( .B1(n6685), .B2(keyinput0), .C1(n6684), .C2(keyinput56), 
        .A(n6683), .ZN(n6689) );
  XOR2_X1 U7609 ( .A(n6741), .B(keyinput24), .Z(n6687) );
  XNOR2_X1 U7610 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .B(keyinput14), .ZN(n6686)
         );
  NAND2_X1 U7611 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  NOR4_X1 U7612 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6719)
         );
  AOI22_X1 U7613 ( .A1(n6735), .A2(keyinput52), .B1(n6725), .B2(keyinput32), 
        .ZN(n6692) );
  OAI221_X1 U7614 ( .B1(n6735), .B2(keyinput52), .C1(n6725), .C2(keyinput32), 
        .A(n6692), .ZN(n6702) );
  INV_X1 U7615 ( .A(DATAI_26_), .ZN(n6694) );
  AOI22_X1 U7616 ( .A1(n6745), .A2(keyinput48), .B1(keyinput17), .B2(n6694), 
        .ZN(n6693) );
  OAI221_X1 U7617 ( .B1(n6745), .B2(keyinput48), .C1(n6694), .C2(keyinput17), 
        .A(n6693), .ZN(n6701) );
  INV_X1 U7618 ( .A(DATAI_23_), .ZN(n6696) );
  AOI22_X1 U7619 ( .A1(n6696), .A2(keyinput6), .B1(n6730), .B2(keyinput51), 
        .ZN(n6695) );
  OAI221_X1 U7620 ( .B1(n6696), .B2(keyinput6), .C1(n6730), .C2(keyinput51), 
        .A(n6695), .ZN(n6700) );
  XNOR2_X1 U7621 ( .A(EBX_REG_27__SCAN_IN), .B(keyinput37), .ZN(n6698) );
  XNOR2_X1 U7622 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput35), .ZN(n6697) );
  NAND2_X1 U7623 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  NOR4_X1 U7624 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n6718)
         );
  INV_X1 U7625 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6705) );
  INV_X1 U7626 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U7627 ( .A1(n6705), .A2(keyinput59), .B1(keyinput23), .B2(n6704), 
        .ZN(n6703) );
  OAI221_X1 U7628 ( .B1(n6705), .B2(keyinput59), .C1(n6704), .C2(keyinput23), 
        .A(n6703), .ZN(n6716) );
  INV_X1 U7629 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U7630 ( .A1(n6731), .A2(keyinput54), .B1(n6707), .B2(keyinput18), 
        .ZN(n6706) );
  OAI221_X1 U7631 ( .B1(n6731), .B2(keyinput54), .C1(n6707), .C2(keyinput18), 
        .A(n6706), .ZN(n6715) );
  AOI22_X1 U7632 ( .A1(n6710), .A2(keyinput36), .B1(keyinput12), .B2(n6709), 
        .ZN(n6708) );
  OAI221_X1 U7633 ( .B1(n6710), .B2(keyinput36), .C1(n6709), .C2(keyinput12), 
        .A(n6708), .ZN(n6714) );
  XNOR2_X1 U7634 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .B(keyinput3), .ZN(n6712)
         );
  XNOR2_X1 U7635 ( .A(keyinput19), .B(EAX_REG_22__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U7636 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  NOR4_X1 U7637 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6717)
         );
  NAND4_X1 U7638 ( .A1(n6720), .A2(n6719), .A3(n6718), .A4(n6717), .ZN(n6721)
         );
  NOR4_X1 U7639 ( .A1(n6724), .A2(n6723), .A3(n6722), .A4(n6721), .ZN(n6766)
         );
  NOR4_X1 U7640 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        INSTQUEUE_REG_10__6__SCAN_IN), .A3(INSTQUEUE_REG_2__6__SCAN_IN), .A4(
        INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6764) );
  NAND3_X1 U7641 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6725), .ZN(n6727) );
  NAND4_X1 U7642 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(
        INSTQUEUE_REG_1__4__SCAN_IN), .A3(INSTQUEUE_REG_2__4__SCAN_IN), .A4(
        INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6726) );
  NOR4_X1 U7643 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n6727), .A3(n6726), 
        .A4(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6729) );
  INV_X1 U7644 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6728) );
  AND4_X1 U7645 ( .A1(n6729), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .A3(
        INSTQUEUE_REG_9__1__SCAN_IN), .A4(n6728), .ZN(n6763) );
  INV_X1 U7646 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6734) );
  AND4_X1 U7647 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        EAX_REG_22__SCAN_IN), .A3(n6731), .A4(n6730), .ZN(n6732) );
  AND4_X1 U7648 ( .A1(n6734), .A2(n6733), .A3(EAX_REG_23__SCAN_IN), .A4(n6732), 
        .ZN(n6740) );
  AND4_X1 U7649 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        EAX_REG_16__SCAN_IN), .A3(ADDRESS_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6739) );
  AND4_X1 U7650 ( .A1(n6736), .A2(n6735), .A3(REIP_REG_29__SCAN_IN), .A4(
        DATAI_23_), .ZN(n6738) );
  AND4_X1 U7651 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6762)
         );
  NAND4_X1 U7652 ( .A1(EBX_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_29__SCAN_IN), 
        .A3(n6742), .A4(n6741), .ZN(n6760) );
  NOR3_X1 U7653 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(
        INSTQUEUE_REG_11__7__SCAN_IN), .A3(n6743), .ZN(n6748) );
  NOR4_X1 U7654 ( .A1(UWORD_REG_4__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        DATAO_REG_2__SCAN_IN), .A4(n6744), .ZN(n6747) );
  NOR4_X1 U7655 ( .A1(ADDRESS_REG_1__SCAN_IN), .A2(DATAI_26_), .A3(
        ADDRESS_REG_8__SCAN_IN), .A4(n6745), .ZN(n6746) );
  NAND4_X1 U7656 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6748), .A3(n6747), 
        .A4(n6746), .ZN(n6759) );
  NAND4_X1 U7657 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        DATAO_REG_8__SCAN_IN), .A3(UWORD_REG_0__SCAN_IN), .A4(n6749), .ZN(
        n6758) );
  NOR3_X1 U7658 ( .A1(DATAI_27_), .A2(ADDRESS_REG_28__SCAN_IN), .A3(n6750), 
        .ZN(n6756) );
  NOR4_X1 U7659 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(CODEFETCH_REG_SCAN_IN), 
        .A3(n6752), .A4(n6751), .ZN(n6755) );
  NOR4_X1 U7660 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        EAX_REG_30__SCAN_IN), .A3(ADDRESS_REG_13__SCAN_IN), .A4(n6753), .ZN(
        n6754) );
  NAND4_X1 U7661 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6756), .A3(n6755), .A4(
        n6754), .ZN(n6757) );
  NOR4_X1 U7662 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6761)
         );
  NAND4_X1 U7663 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6765)
         );
  NAND4_X1 U7664 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6769)
         );
  XNOR2_X1 U7665 ( .A(n6770), .B(n6769), .ZN(U2946) );
  CLKBUF_X1 U3432 ( .A(n3558), .Z(n3898) );
  CLKBUF_X1 U3435 ( .A(n2950), .Z(n3350) );
  CLKBUF_X1 U3441 ( .A(n3350), .Z(n3848) );
  NAND2_X1 U3518 ( .A1(n3465), .A2(n2974), .ZN(n4200) );
  CLKBUF_X1 U3997 ( .A(n3232), .Z(n4235) );
  CLKBUF_X1 U4005 ( .A(n3358), .Z(n4230) );
  CLKBUF_X1 U4015 ( .A(n4145), .Z(n2955) );
  AND3_X1 U4066 ( .A1(n3230), .A2(n4265), .A3(n3098), .ZN(n6771) );
endmodule

