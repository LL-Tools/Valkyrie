

module b15_C_gen_AntiSAT_k_256_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3152, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3192, n3194,
         n3195, n3196, n3197, n3198, n3199, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000;

  AND2_X1 U3600 ( .A1(n4565), .A2(n3241), .ZN(n4630) );
  AND2_X1 U3601 ( .A1(n3753), .A2(n3408), .ZN(n3776) );
  CLKBUF_X2 U3602 ( .A(n3396), .Z(n3507) );
  CLKBUF_X2 U3603 ( .A(n3617), .Z(n3190) );
  CLKBUF_X2 U3604 ( .A(n3612), .Z(n3154) );
  CLKBUF_X2 U3605 ( .A(n3581), .Z(n3192) );
  AND2_X1 U3607 ( .A1(n3303), .A2(n3315), .ZN(n3187) );
  INV_X1 U3608 ( .A(n3513), .ZN(n3204) );
  AND2_X2 U3610 ( .A1(n3304), .A2(n4604), .ZN(n3611) );
  AND2_X2 U3611 ( .A1(n3304), .A2(n4587), .ZN(n3617) );
  AND2_X2 U3612 ( .A1(n3229), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3304)
         );
  INV_X1 U3613 ( .A(n3512), .ZN(n3156) );
  BUF_X1 U3614 ( .A(n3581), .Z(n3195) );
  INV_X2 U3615 ( .A(n4294), .ZN(n3152) );
  INV_X2 U3616 ( .A(n4511), .ZN(n4468) );
  INV_X1 U3618 ( .A(n3727), .ZN(n5194) );
  NOR2_X1 U3620 ( .A1(n4996), .A2(n3222), .ZN(n5015) );
  AND2_X2 U3621 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U3622 ( .A1(n3591), .A2(n3592), .ZN(n3656) );
  OR2_X1 U3623 ( .A1(n5233), .A2(n5088), .ZN(n4483) );
  AND2_X1 U3624 ( .A1(n3234), .A2(n3232), .ZN(n3207) );
  OAI21_X1 U3625 ( .B1(n4995), .B2(n4997), .A(n4996), .ZN(n5353) );
  NAND2_X2 U3627 ( .A1(n4588), .A2(n4535), .ZN(n3169) );
  INV_X1 U3628 ( .A(n3610), .ZN(n3158) );
  NAND2_X1 U3629 ( .A1(n4701), .A2(n4700), .ZN(n4699) );
  AOI21_X1 U3630 ( .B1(n5368), .B2(n5367), .A(n5366), .ZN(n5430) );
  NAND2_X2 U3631 ( .A1(n5123), .A2(n3741), .ZN(n5185) );
  NOR3_X1 U3632 ( .A1(n5194), .A2(n4416), .A3(n5409), .ZN(n3747) );
  OR2_X1 U3633 ( .A1(n4477), .A2(n3247), .ZN(n3246) );
  CLKBUF_X2 U3634 ( .A(n5740), .Z(n5791) );
  NAND2_X1 U3635 ( .A1(n3207), .A2(n4844), .ZN(n4850) );
  NAND2_X1 U3636 ( .A1(n3506), .A2(n3505), .ZN(n3562) );
  NAND2_X1 U3637 ( .A1(n3447), .A2(n3446), .ZN(n3567) );
  CLKBUF_X2 U3638 ( .A(n4304), .Z(n3184) );
  NAND2_X1 U3639 ( .A1(n4660), .A2(n3534), .ZN(n4977) );
  INV_X2 U3640 ( .A(n3445), .ZN(n3534) );
  CLKBUF_X2 U3641 ( .A(n3171), .Z(n4216) );
  INV_X2 U3642 ( .A(n3158), .ZN(n3203) );
  CLKBUF_X2 U3644 ( .A(n3398), .Z(n4236) );
  AND2_X2 U3645 ( .A1(n4587), .A2(n4535), .ZN(n3581) );
  OR2_X1 U3646 ( .A1(n4440), .A2(n5878), .ZN(n4267) );
  NAND2_X1 U3647 ( .A1(n5111), .A2(n5110), .ZN(n5367) );
  AND2_X1 U3648 ( .A1(n3209), .A2(n3746), .ZN(n5342) );
  NAND2_X1 U3649 ( .A1(n4263), .A2(n3292), .ZN(n4416) );
  AOI211_X1 U3650 ( .C1(n5349), .C2(n5626), .A(n5001), .B(n5000), .ZN(n5002)
         );
  XNOR2_X1 U3651 ( .A(n4257), .B(n4256), .ZN(n5092) );
  XNOR2_X1 U3652 ( .A(n5015), .B(n4466), .ZN(n5339) );
  NOR2_X1 U3653 ( .A1(n5030), .A2(n5031), .ZN(n4995) );
  AND2_X1 U3654 ( .A1(n4483), .A2(n3296), .ZN(n4484) );
  AOI211_X1 U3655 ( .C1(n5256), .C2(n5601), .A(n5255), .B(n5254), .ZN(n5258)
         );
  CLKBUF_X1 U3656 ( .A(n5814), .Z(n3179) );
  AOI21_X1 U3657 ( .B1(n4429), .B2(n4475), .A(n4481), .ZN(n4432) );
  AOI21_X1 U3658 ( .B1(n3260), .B2(n3262), .A(n3259), .ZN(n3258) );
  NOR2_X1 U3659 ( .A1(n4474), .A2(n4428), .ZN(n4477) );
  AND2_X1 U3660 ( .A1(n4918), .A2(n3271), .ZN(n3270) );
  AND2_X1 U3661 ( .A1(n3180), .A2(n3181), .ZN(n3165) );
  AND2_X1 U3662 ( .A1(n3181), .A2(n5829), .ZN(n3164) );
  NAND2_X1 U3663 ( .A1(n3868), .A2(n3867), .ZN(n4781) );
  OR2_X1 U3664 ( .A1(n5835), .A2(n3182), .ZN(n3181) );
  NAND2_X2 U3665 ( .A1(n3711), .A2(n3720), .ZN(n3727) );
  NAND3_X1 U3666 ( .A1(n4624), .A2(n4561), .A3(n4696), .ZN(n4642) );
  AND2_X1 U3667 ( .A1(n4623), .A2(n4632), .ZN(n4624) );
  NAND2_X1 U3668 ( .A1(n3697), .A2(n3696), .ZN(n3711) );
  OR2_X1 U3669 ( .A1(n3848), .A2(n3847), .ZN(n4563) );
  NOR2_X1 U3671 ( .A1(n4636), .A2(n3659), .ZN(n3660) );
  OR2_X1 U3672 ( .A1(n3591), .A2(n3592), .ZN(n3593) );
  NAND2_X2 U3673 ( .A1(n5674), .A2(n3435), .ZN(n5086) );
  AND2_X1 U3675 ( .A1(n3173), .A2(n3174), .ZN(n3255) );
  CLKBUF_X1 U3676 ( .A(n4586), .Z(n6362) );
  OR2_X1 U3677 ( .A1(n4652), .A2(n4979), .ZN(n5237) );
  XNOR2_X1 U3678 ( .A(n3562), .B(n3563), .ZN(n3553) );
  NAND2_X1 U3679 ( .A1(n3494), .A2(n3493), .ZN(n6282) );
  CLKBUF_X1 U3680 ( .A(n3834), .Z(n6482) );
  NAND2_X1 U3681 ( .A1(n3566), .A2(n3464), .ZN(n3834) );
  AND2_X2 U3682 ( .A1(n3566), .A2(n3464), .ZN(n3159) );
  AOI21_X1 U3683 ( .B1(n3602), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3570), 
        .ZN(n3573) );
  NOR2_X1 U3684 ( .A1(n4302), .A2(n3461), .ZN(n3463) );
  XNOR2_X1 U3685 ( .A(n3214), .B(n4553), .ZN(n5642) );
  AND2_X1 U3686 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  NAND2_X1 U3687 ( .A1(n3530), .A2(n3529), .ZN(n4287) );
  OR3_X1 U3688 ( .A1(n3779), .A2(n3778), .A3(n3777), .ZN(n3780) );
  NOR2_X1 U3689 ( .A1(n4648), .A2(n4288), .ZN(n4327) );
  AND2_X1 U3690 ( .A1(n4529), .A2(n3436), .ZN(n3459) );
  AND2_X1 U3691 ( .A1(n4403), .A2(n4294), .ZN(n4555) );
  NAND2_X1 U3692 ( .A1(n3227), .A2(n3535), .ZN(n4648) );
  NAND2_X1 U3693 ( .A1(n3776), .A2(n3749), .ZN(n3797) );
  NAND2_X1 U3694 ( .A1(n3609), .A2(n3608), .ZN(n3804) );
  NAND2_X2 U3695 ( .A1(n4671), .A2(n3445), .ZN(n4403) );
  INV_X1 U3696 ( .A(n4297), .ZN(n3809) );
  NAND2_X1 U3697 ( .A1(n3532), .A2(n3450), .ZN(n4297) );
  AND2_X1 U3698 ( .A1(n4660), .A2(n3445), .ZN(n3496) );
  INV_X1 U3699 ( .A(n3532), .ZN(n4671) );
  OR2_X1 U3700 ( .A1(n3474), .A2(n3473), .ZN(n3554) );
  OR2_X1 U3701 ( .A1(n3486), .A2(n3485), .ZN(n3719) );
  AND2_X1 U3702 ( .A1(n3445), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3753) );
  INV_X1 U3703 ( .A(n3450), .ZN(n4295) );
  AND4_X1 U3704 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3330)
         );
  NAND2_X2 U3705 ( .A1(n3379), .A2(n3378), .ZN(n3435) );
  NAND4_X2 U3706 ( .A1(n3349), .A2(n3350), .A3(n3347), .A4(n3348), .ZN(n3531)
         );
  AND4_X2 U3707 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3450)
         );
  AND4_X1 U3708 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3403)
         );
  AND4_X1 U3709 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3405)
         );
  AND4_X1 U3710 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n3213)
         );
  AND4_X1 U3711 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3368)
         );
  AND4_X1 U3712 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3349)
         );
  AND4_X1 U3713 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3431)
         );
  AND4_X1 U3714 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3347)
         );
  AND4_X1 U3715 ( .A1(n3421), .A2(n3420), .A3(n3419), .A4(n3418), .ZN(n3432)
         );
  AND4_X1 U3716 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3379)
         );
  AND4_X1 U3717 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3310)
         );
  CLKBUF_X1 U3718 ( .A(n6572), .Z(n6577) );
  AND4_X1 U3719 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3404)
         );
  AND4_X1 U3720 ( .A1(n3385), .A2(n3384), .A3(n3383), .A4(n3382), .ZN(n3406)
         );
  INV_X1 U3721 ( .A(n3170), .ZN(n3171) );
  NAND2_X2 U3722 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6998), .ZN(n6575) );
  AND2_X1 U3723 ( .A1(n3318), .A2(n3316), .ZN(n3178) );
  AND4_X1 U3724 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(n3378)
         );
  AND4_X1 U3725 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3350)
         );
  AND4_X1 U3726 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3367)
         );
  AND4_X1 U3727 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3369)
         );
  AND4_X1 U3728 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3430)
         );
  AND4_X1 U3729 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3348)
         );
  AND4_X1 U3730 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3433)
         );
  BUF_X2 U3731 ( .A(n3581), .Z(n3196) );
  AND2_X2 U3732 ( .A1(n6599), .A2(n4613), .ZN(n4833) );
  BUF_X2 U3734 ( .A(n3611), .Z(n3475) );
  BUF_X2 U3735 ( .A(n3417), .Z(n3869) );
  INV_X4 U3736 ( .A(n3169), .ZN(n3157) );
  NOR2_X1 U3737 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6596), .ZN(n4254) );
  CLKBUF_X1 U3738 ( .A(n6405), .Z(n6603) );
  INV_X1 U3739 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3298) );
  INV_X2 U3740 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6251) );
  AND2_X2 U3741 ( .A1(n4587), .A2(n4534), .ZN(n3417) );
  NAND2_X1 U3742 ( .A1(n3832), .A2(n3831), .ZN(n4508) );
  BUF_X2 U3743 ( .A(n3381), .Z(n4187) );
  INV_X2 U3744 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3229) );
  AND4_X1 U3745 ( .A1(n3308), .A2(n3306), .A3(n3307), .A4(n3305), .ZN(n3309)
         );
  AOI22_X1 U3746 ( .A1(n3198), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3306) );
  XNOR2_X1 U3747 ( .A(n3681), .B(n3682), .ZN(n3852) );
  XNOR2_X1 U3748 ( .A(n3711), .B(n3710), .ZN(n3860) );
  NAND2_X1 U3749 ( .A1(n3434), .A2(n3534), .ZN(n3160) );
  NAND2_X1 U3750 ( .A1(n5035), .A2(n5037), .ZN(n3161) );
  OR2_X2 U3751 ( .A1(n3161), .A2(n3162), .ZN(n4996) );
  OR2_X1 U3752 ( .A1(n3163), .A2(n5031), .ZN(n3162) );
  INV_X1 U3753 ( .A(n4997), .ZN(n3163) );
  INV_X1 U3754 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3166) );
  AND2_X1 U3755 ( .A1(n3303), .A2(n3315), .ZN(n3397) );
  INV_X1 U3756 ( .A(n3156), .ZN(n3167) );
  NAND2_X1 U3757 ( .A1(n3184), .A2(n3532), .ZN(n3168) );
  INV_X1 U3758 ( .A(n3156), .ZN(n3199) );
  INV_X1 U3759 ( .A(n3391), .ZN(n3170) );
  OR2_X2 U3760 ( .A1(n3462), .A2(n3463), .ZN(n3172) );
  AND2_X4 U3761 ( .A1(n3297), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4588)
         );
  NAND2_X1 U3762 ( .A1(n4527), .A2(n3176), .ZN(n3173) );
  OR2_X1 U3763 ( .A1(n3175), .A2(n3551), .ZN(n3174) );
  INV_X1 U3764 ( .A(n3563), .ZN(n3175) );
  AND2_X1 U3765 ( .A1(n6599), .A2(n3563), .ZN(n3176) );
  NAND2_X1 U3766 ( .A1(n4527), .A2(n6599), .ZN(n3177) );
  XNOR2_X2 U3767 ( .A(n3549), .B(n3548), .ZN(n4527) );
  AND3_X2 U3768 ( .A1(n3178), .A2(n3317), .A3(n3319), .ZN(n3320) );
  AND2_X2 U3769 ( .A1(n4588), .A2(n3303), .ZN(n3610) );
  AND2_X2 U3770 ( .A1(n4534), .A2(n4588), .ZN(n3512) );
  NOR2_X2 U3771 ( .A1(n5269), .A2(n4455), .ZN(n5263) );
  NOR2_X2 U3772 ( .A1(n6562), .A2(n5552), .ZN(n5537) );
  AOI21_X1 U3773 ( .B1(n4441), .B2(n3536), .A(n4327), .ZN(n3537) );
  NOR2_X2 U3774 ( .A1(n5605), .A2(n5606), .ZN(n4644) );
  NOR2_X2 U3775 ( .A1(n4510), .A2(n3214), .ZN(n4565) );
  NOR3_X4 U3776 ( .A1(n5450), .A2(n5449), .A3(n3237), .ZN(n5059) );
  NAND2_X1 U3777 ( .A1(n4699), .A2(n3183), .ZN(n3180) );
  INV_X1 U3778 ( .A(n3680), .ZN(n3182) );
  AND2_X1 U3779 ( .A1(n3655), .A2(n3680), .ZN(n3183) );
  NAND2_X1 U3780 ( .A1(n5820), .A2(n3718), .ZN(n5814) );
  AND2_X4 U3781 ( .A1(n3656), .A2(n3593), .ZN(n4634) );
  AND2_X2 U3782 ( .A1(n3543), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3303)
         );
  NAND2_X2 U3783 ( .A1(n3850), .A2(n3849), .ZN(n4561) );
  AND2_X1 U3784 ( .A1(n4263), .A2(n3263), .ZN(n5343) );
  NOR2_X2 U3785 ( .A1(n5367), .A2(n5368), .ZN(n5366) );
  INV_X2 U3786 ( .A(n3409), .ZN(n4686) );
  NAND2_X2 U3787 ( .A1(n5064), .A2(n5066), .ZN(n5005) );
  XNOR2_X1 U3788 ( .A(n3553), .B(n3564), .ZN(n4618) );
  NOR2_X2 U3790 ( .A1(n4642), .A2(n4643), .ZN(n4780) );
  NOR2_X2 U3791 ( .A1(n4521), .A2(n4516), .ZN(n4421) );
  AOI21_X2 U3792 ( .B1(n3567), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3449), 
        .ZN(n3462) );
  AND2_X2 U3793 ( .A1(n4274), .A2(n4660), .ZN(n4521) );
  AND2_X2 U3794 ( .A1(n3527), .A2(n3526), .ZN(n4274) );
  OAI22_X2 U3795 ( .A1(n5185), .A2(n5184), .B1(n5194), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5176) );
  NAND2_X2 U3796 ( .A1(n3266), .A2(n3265), .ZN(n4263) );
  BUF_X2 U3797 ( .A(n4618), .Z(n3185) );
  AOI21_X1 U3798 ( .B1(n3440), .B2(n3409), .A(n3408), .ZN(n3525) );
  INV_X2 U3799 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3297) );
  AND2_X1 U3800 ( .A1(n3303), .A2(n3315), .ZN(n3186) );
  AND2_X1 U3801 ( .A1(n3304), .A2(n4588), .ZN(n3188) );
  NAND2_X4 U3802 ( .A1(n3321), .A2(n3320), .ZN(n3438) );
  NOR2_X4 U3803 ( .A1(n4847), .A2(n4854), .ZN(n3955) );
  OAI21_X2 U3804 ( .B1(n4201), .B2(n4202), .A(n5014), .ZN(n5097) );
  OAI21_X2 U3805 ( .B1(n4887), .B2(n3269), .A(n3267), .ZN(n5207) );
  OAI21_X2 U3806 ( .B1(n5796), .B2(n3731), .A(n3730), .ZN(n4887) );
  AND2_X4 U3807 ( .A1(n4534), .A2(n3315), .ZN(n3189) );
  INV_X2 U3808 ( .A(n3169), .ZN(n3197) );
  INV_X2 U3809 ( .A(n3169), .ZN(n3198) );
  AND2_X1 U3810 ( .A1(n3304), .A2(n4588), .ZN(n3612) );
  OAI21_X2 U3814 ( .B1(n5129), .B2(n3737), .A(n3736), .ZN(n5195) );
  OAI21_X2 U3815 ( .B1(n5207), .B2(n3735), .A(n3734), .ZN(n5129) );
  AND2_X2 U3816 ( .A1(n4933), .A2(n3225), .ZN(n5064) );
  NOR2_X4 U3817 ( .A1(n4906), .A2(n5131), .ZN(n4933) );
  INV_X1 U3818 ( .A(n3513), .ZN(n3205) );
  INV_X1 U3819 ( .A(n3476), .ZN(n3206) );
  AOI22_X1 U3820 ( .A1(n3612), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U3821 ( .A1(n3673), .A2(n3672), .ZN(n3682) );
  NAND2_X1 U3822 ( .A1(n3683), .A2(n3682), .ZN(n3699) );
  INV_X1 U3823 ( .A(n3681), .ZN(n3683) );
  AND2_X1 U3824 ( .A1(n3695), .A2(n3694), .ZN(n3698) );
  OR2_X1 U3825 ( .A1(n4427), .A2(n3289), .ZN(n4428) );
  NAND2_X1 U3826 ( .A1(n5185), .A2(n3745), .ZN(n3266) );
  OR2_X1 U3827 ( .A1(n4403), .A2(n4468), .ZN(n4394) );
  NAND2_X1 U3828 ( .A1(n3152), .A2(n3216), .ZN(n3240) );
  NAND2_X1 U3829 ( .A1(n3534), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3609) );
  INV_X1 U3830 ( .A(n5003), .ZN(n3238) );
  INV_X1 U3831 ( .A(n5004), .ZN(n3239) );
  OR3_X1 U3832 ( .A1(n4652), .A2(READY_N), .A3(n4651), .ZN(n5713) );
  AOI22_X1 U3833 ( .A1(n4253), .A2(n5336), .B1(n4252), .B2(n4251), .ZN(n4465)
         );
  NAND2_X1 U3834 ( .A1(n5343), .A2(n5139), .ZN(n5227) );
  OR2_X1 U3835 ( .A1(n4423), .A2(n4307), .ZN(n4919) );
  OR2_X1 U3836 ( .A1(n4419), .A2(n3752), .ZN(n6495) );
  AND2_X1 U3837 ( .A1(n3808), .A2(n3442), .ZN(n3443) );
  AND2_X1 U3838 ( .A1(n3809), .A2(n3441), .ZN(n3442) );
  NAND2_X1 U3839 ( .A1(n3634), .A2(n3660), .ZN(n3681) );
  INV_X1 U3840 ( .A(n3776), .ZN(n3794) );
  INV_X1 U3841 ( .A(n3719), .ZN(n3722) );
  NAND2_X1 U3842 ( .A1(n3452), .A2(n3410), .ZN(n3526) );
  AOI22_X1 U3843 ( .A1(n3437), .A2(n3440), .B1(n3435), .B2(n4295), .ZN(n3410)
         );
  NAND2_X1 U3844 ( .A1(n4202), .A2(n3273), .ZN(n3272) );
  INV_X1 U3845 ( .A(n5020), .ZN(n3273) );
  NAND2_X1 U3846 ( .A1(n5052), .A2(n3283), .ZN(n3282) );
  INV_X1 U3847 ( .A(n5007), .ZN(n3283) );
  NAND2_X1 U3848 ( .A1(n3940), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3959)
         );
  OR2_X1 U3849 ( .A1(n3275), .A2(n3278), .ZN(n3274) );
  INV_X1 U3850 ( .A(n4849), .ZN(n3278) );
  OR2_X1 U3851 ( .A1(n3276), .A2(n4843), .ZN(n3275) );
  AND2_X1 U3852 ( .A1(n3827), .A2(EAX_REG_7__SCAN_IN), .ZN(n3866) );
  NOR2_X2 U3853 ( .A1(n3409), .A2(n6251), .ZN(n3981) );
  INV_X1 U3854 ( .A(n5029), .ZN(n3245) );
  INV_X1 U3855 ( .A(n3698), .ZN(n3696) );
  INV_X1 U3856 ( .A(n3699), .ZN(n3697) );
  NAND2_X1 U3857 ( .A1(n4888), .A2(n4889), .ZN(n3271) );
  NOR2_X1 U3858 ( .A1(n3495), .A2(n3408), .ZN(n4304) );
  INV_X1 U3859 ( .A(n3726), .ZN(n3262) );
  INV_X1 U3860 ( .A(n3261), .ZN(n3260) );
  OAI21_X1 U3861 ( .B1(n5813), .B2(n3262), .A(n5804), .ZN(n3261) );
  NOR2_X1 U3862 ( .A1(n4783), .A2(n3236), .ZN(n3235) );
  INV_X1 U3863 ( .A(n4776), .ZN(n3236) );
  INV_X1 U3864 ( .A(n4784), .ZN(n3234) );
  INV_X1 U3865 ( .A(n3551), .ZN(n3252) );
  NAND2_X1 U3866 ( .A1(n3588), .A2(n3550), .ZN(n3253) );
  NOR2_X1 U3867 ( .A1(n4533), .A2(n4308), .ZN(n4579) );
  OAI21_X1 U3868 ( .B1(n4614), .B2(n4613), .A(n6510), .ZN(n4659) );
  INV_X1 U3869 ( .A(n5073), .ZN(n3237) );
  NAND2_X1 U3870 ( .A1(n4480), .A2(n3249), .ZN(n5233) );
  NAND2_X1 U3871 ( .A1(n4479), .A2(n4478), .ZN(n4480) );
  NAND2_X1 U3872 ( .A1(n3246), .A2(n4473), .ZN(n3249) );
  NAND2_X1 U3873 ( .A1(n5050), .A2(n3244), .ZN(n5023) );
  AND2_X1 U3874 ( .A1(n3210), .A2(n4991), .ZN(n3244) );
  AND2_X1 U3875 ( .A1(n5354), .A2(n3221), .ZN(n3265) );
  NOR2_X2 U3876 ( .A1(n4851), .A2(n4850), .ZN(n4856) );
  INV_X1 U3877 ( .A(n5910), .ZN(n5197) );
  NAND2_X1 U3878 ( .A1(n3179), .A2(n5813), .ZN(n5812) );
  NAND2_X1 U3879 ( .A1(n4644), .A2(n4645), .ZN(n4784) );
  AND2_X1 U3880 ( .A1(n4566), .A2(n3242), .ZN(n3241) );
  INV_X1 U3881 ( .A(n4631), .ZN(n3242) );
  AND2_X1 U3882 ( .A1(n4293), .A2(n4292), .ZN(n4423) );
  OAI21_X1 U3883 ( .B1(n6282), .B2(n3495), .A(n3498), .ZN(n5871) );
  NAND2_X2 U3884 ( .A1(n3806), .A2(n3805), .ZN(n4978) );
  NAND2_X1 U3885 ( .A1(n3803), .A2(n3802), .ZN(n3806) );
  AND2_X1 U3886 ( .A1(n3155), .A2(n6282), .ZN(n6210) );
  NAND2_X1 U3887 ( .A1(n6599), .A2(n4659), .ZN(n4761) );
  NOR2_X1 U3888 ( .A1(n4445), .A2(n4487), .ZN(n5592) );
  INV_X1 U3889 ( .A(n4488), .ZN(n4445) );
  INV_X1 U3890 ( .A(n5644), .ZN(n5658) );
  AND2_X1 U3891 ( .A1(n5090), .A2(n4657), .ZN(n5684) );
  AND2_X1 U3892 ( .A1(n5090), .A2(n4655), .ZN(n5688) );
  NAND2_X1 U3893 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  NAND2_X1 U3894 ( .A1(n5227), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5228) );
  INV_X1 U3895 ( .A(n4465), .ZN(n4466) );
  OR2_X1 U3896 ( .A1(n4652), .A2(n6495), .ZN(n5878) );
  INV_X1 U3897 ( .A(n3211), .ZN(n3231) );
  INV_X1 U3898 ( .A(n5233), .ZN(n5244) );
  AND2_X1 U3899 ( .A1(n6502), .A2(n6501), .ZN(n6520) );
  NAND2_X1 U3900 ( .A1(n3646), .A2(n3645), .ZN(n3658) );
  OR2_X1 U3901 ( .A1(n3693), .A2(n3692), .ZN(n3712) );
  OR2_X1 U3902 ( .A1(n3671), .A2(n3670), .ZN(n3700) );
  AOI21_X1 U3903 ( .B1(n4468), .B2(n4512), .A(n3152), .ZN(n4332) );
  NAND2_X1 U3904 ( .A1(n3538), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3545) );
  AOI21_X1 U3905 ( .B1(n5224), .B2(n6493), .A(n3792), .ZN(n3800) );
  NOR2_X1 U3906 ( .A1(n3791), .A2(n3790), .ZN(n3792) );
  AND2_X1 U3907 ( .A1(n3794), .A2(n3786), .ZN(n3787) );
  AOI22_X1 U3908 ( .A1(n3188), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U3909 ( .A1(n3512), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U3910 ( .A1(n3610), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3611), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U3911 ( .A1(n3196), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3300) );
  OR2_X1 U3912 ( .A1(n3623), .A2(n3622), .ZN(n3648) );
  OR2_X1 U3913 ( .A1(n3519), .A2(n3518), .ZN(n3555) );
  AOI22_X1 U3914 ( .A1(n3610), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U3915 ( .A1(n3617), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U3916 ( .A1(n3512), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U3917 ( .A1(n3157), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3372) );
  OR2_X1 U3918 ( .A1(n4138), .A2(n4137), .ZN(n4152) );
  INV_X1 U3919 ( .A(n5069), .ZN(n3279) );
  NOR2_X1 U3920 ( .A1(n3281), .A2(n5389), .ZN(n3280) );
  INV_X1 U3921 ( .A(n4935), .ZN(n3281) );
  NAND2_X1 U3922 ( .A1(n3277), .A2(n4839), .ZN(n3276) );
  NOR2_X1 U3923 ( .A1(n4294), .A2(n3248), .ZN(n3247) );
  NAND2_X1 U3924 ( .A1(n4468), .A2(n4294), .ZN(n4402) );
  INV_X1 U3925 ( .A(n4402), .ZN(n4407) );
  NAND2_X1 U3926 ( .A1(n3172), .A2(n3565), .ZN(n3575) );
  INV_X1 U3927 ( .A(n3797), .ZN(n3801) );
  OR2_X1 U3928 ( .A1(n6139), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3603)
         );
  AND2_X1 U3929 ( .A1(n4585), .A2(n4584), .ZN(n6489) );
  INV_X1 U3930 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5532) );
  NOR2_X1 U3931 ( .A1(n3926), .A2(n3925), .ZN(n3940) );
  INV_X1 U3932 ( .A(n5611), .ZN(n5630) );
  NAND2_X1 U3933 ( .A1(n4856), .A2(n4855), .ZN(n4883) );
  NAND2_X1 U3934 ( .A1(n4686), .A2(n3438), .ZN(n4654) );
  AND2_X1 U3935 ( .A1(n4504), .A2(n4986), .ZN(n5692) );
  NAND2_X1 U3936 ( .A1(n5793), .A2(n4503), .ZN(n4504) );
  OR2_X1 U3937 ( .A1(n4652), .A2(n6478), .ZN(n4503) );
  XNOR2_X1 U3938 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .B(n4260), .ZN(n4488)
         );
  NOR2_X1 U3939 ( .A1(n4214), .A2(n4213), .ZN(n4215) );
  AOI22_X1 U3940 ( .A1(n4253), .A2(n4489), .B1(n4200), .B2(n4199), .ZN(n4202)
         );
  NOR2_X1 U3941 ( .A1(n4167), .A2(n4993), .ZN(n4168) );
  NAND2_X1 U3942 ( .A1(n4168), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4214)
         );
  AOI22_X1 U3943 ( .A1(n4253), .A2(n5349), .B1(n4166), .B2(n4165), .ZN(n4997)
         );
  NOR2_X1 U3944 ( .A1(n4135), .A2(n4134), .ZN(n4136) );
  NAND2_X1 U3945 ( .A1(n4136), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4167)
         );
  OR2_X1 U3946 ( .A1(n5274), .A2(n4232), .ZN(n4133) );
  NOR2_X1 U3947 ( .A1(n4089), .A2(n4088), .ZN(n4090) );
  NAND2_X1 U3948 ( .A1(n4090), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4135)
         );
  AND2_X1 U3949 ( .A1(n4253), .A2(n5362), .ZN(n4085) );
  NOR2_X1 U3950 ( .A1(n4058), .A2(n5303), .ZN(n4059) );
  NOR2_X1 U3951 ( .A1(n4031), .A2(n4030), .ZN(n4032) );
  NAND2_X1 U3952 ( .A1(n4032), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4058)
         );
  AND2_X1 U3953 ( .A1(n4003), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4004)
         );
  NOR2_X1 U3954 ( .A1(n3989), .A2(n5517), .ZN(n4003) );
  NOR2_X1 U3955 ( .A1(n3959), .A2(n5532), .ZN(n3986) );
  CLKBUF_X1 U3956 ( .A(n4906), .Z(n4907) );
  NAND2_X1 U3957 ( .A1(n3912), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3926)
         );
  CLKBUF_X1 U3958 ( .A(n4847), .Z(n4848) );
  NOR2_X1 U3959 ( .A1(n3909), .A2(n5574), .ZN(n3912) );
  NAND2_X1 U3960 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3909)
         );
  INV_X1 U3961 ( .A(n3884), .ZN(n3885) );
  NOR2_X1 U3962 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  INV_X1 U3963 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U3964 ( .A1(n3863), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3884)
         );
  NOR2_X1 U3965 ( .A1(n3866), .A2(n3865), .ZN(n3867) );
  INV_X1 U3966 ( .A(n3864), .ZN(n3865) );
  AOI21_X1 U3967 ( .B1(n3859), .B2(n3981), .A(n3858), .ZN(n4643) );
  NOR2_X1 U3968 ( .A1(n3819), .A2(n5617), .ZN(n3853) );
  INV_X1 U3969 ( .A(n3843), .ZN(n3820) );
  NAND2_X1 U3970 ( .A1(n3820), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3819)
         );
  NOR2_X1 U3971 ( .A1(n4477), .A2(n3152), .ZN(n4481) );
  NOR2_X1 U3972 ( .A1(n5145), .A2(n3264), .ZN(n3263) );
  INV_X1 U3973 ( .A(n3292), .ZN(n3264) );
  AND3_X1 U3974 ( .A1(n3184), .A2(STATE2_REG_0__SCAN_IN), .A3(n3719), .ZN(
        n3720) );
  NAND2_X1 U3975 ( .A1(n5059), .A2(n4382), .ZN(n5004) );
  NAND2_X1 U3976 ( .A1(n5456), .A2(n4938), .ZN(n5450) );
  AOI21_X1 U3977 ( .B1(n3270), .B2(n3268), .A(n3208), .ZN(n3267) );
  INV_X1 U3978 ( .A(n3270), .ZN(n3269) );
  OR2_X1 U3979 ( .A1(n4925), .A2(n5951), .ZN(n4891) );
  OR2_X1 U3980 ( .A1(n5944), .A2(n4315), .ZN(n4923) );
  INV_X1 U3981 ( .A(n5805), .ZN(n3259) );
  AND2_X1 U3982 ( .A1(n3235), .A2(n3233), .ZN(n3232) );
  INV_X1 U3983 ( .A(n4840), .ZN(n3233) );
  NAND2_X1 U3984 ( .A1(n4630), .A2(n4627), .ZN(n5605) );
  OR2_X1 U3985 ( .A1(n4423), .A2(n4971), .ZN(n5944) );
  NAND2_X1 U3986 ( .A1(n3256), .A2(n3255), .ZN(n3591) );
  NAND2_X1 U3987 ( .A1(n3251), .A2(n3562), .ZN(n3256) );
  XNOR2_X1 U3988 ( .A(n3254), .B(n3590), .ZN(n3592) );
  AND2_X1 U3989 ( .A1(n3534), .A2(n3291), .ZN(n3454) );
  INV_X1 U3990 ( .A(n4599), .ZN(n6485) );
  AND2_X1 U3991 ( .A1(n6033), .A2(n5970), .ZN(n5996) );
  AND2_X1 U3992 ( .A1(n6244), .A2(n6147), .ZN(n6178) );
  AND2_X1 U3993 ( .A1(n6062), .A2(n4635), .ZN(n6244) );
  NAND2_X1 U3994 ( .A1(n3491), .A2(n3501), .ZN(n3494) );
  OAI21_X1 U3995 ( .B1(n3834), .B2(STATE2_REG_0__SCAN_IN), .A(n3502), .ZN(
        n3491) );
  NOR2_X1 U3996 ( .A1(n6411), .A2(n3185), .ZN(n6330) );
  INV_X1 U3997 ( .A(n6243), .ZN(n6112) );
  NAND2_X1 U3998 ( .A1(n6585), .A2(n4659), .ZN(n4763) );
  OR2_X1 U3999 ( .A1(n4981), .A2(n4442), .ZN(n5238) );
  CLKBUF_X1 U4000 ( .A(n3496), .Z(n6597) );
  NOR2_X1 U4001 ( .A1(n6521), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6602) );
  NOR2_X1 U4002 ( .A1(n6558), .A2(n5581), .ZN(n5576) );
  NAND2_X1 U4003 ( .A1(n5630), .A2(n4451), .ZN(n5581) );
  CLKBUF_X1 U4004 ( .A(n5601), .Z(n5626) );
  INV_X1 U4005 ( .A(n5597), .ZN(n5619) );
  NOR2_X1 U4006 ( .A1(n4488), .A2(n4487), .ZN(n5601) );
  AND2_X1 U4007 ( .A1(n4942), .A2(n4494), .ZN(n5644) );
  AND2_X1 U4008 ( .A1(n5651), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5638) );
  OR2_X1 U4009 ( .A1(n5592), .A2(n4939), .ZN(n5648) );
  INV_X1 U4010 ( .A(n4496), .ZN(n4497) );
  INV_X1 U4011 ( .A(n5088), .ZN(n5671) );
  INV_X1 U4012 ( .A(n5674), .ZN(n5074) );
  AND2_X1 U4013 ( .A1(n4471), .A2(n6522), .ZN(n5674) );
  NAND2_X1 U4014 ( .A1(n5674), .A2(n5089), .ZN(n5088) );
  OAI21_X1 U4015 ( .B1(n4650), .B2(n4649), .A(n6522), .ZN(n4653) );
  INV_X1 U4016 ( .A(n5688), .ZN(n5677) );
  NAND2_X1 U4017 ( .A1(n5015), .A2(n4465), .ZN(n4257) );
  INV_X1 U4018 ( .A(n5878), .ZN(n5864) );
  NAND2_X1 U4019 ( .A1(n5050), .A2(n5040), .ZN(n5028) );
  NAND2_X1 U4020 ( .A1(n4891), .A2(n4923), .ZN(n5880) );
  NAND2_X1 U4021 ( .A1(n5812), .A2(n3726), .ZN(n5807) );
  NOR2_X1 U4022 ( .A1(n4784), .A2(n4783), .ZN(n4775) );
  OR2_X1 U4023 ( .A1(n6521), .A2(n6529), .ZN(n5937) );
  NAND2_X1 U4024 ( .A1(n4565), .A2(n4566), .ZN(n3243) );
  OR2_X1 U4025 ( .A1(n4423), .A2(n6478), .ZN(n5955) );
  NOR2_X1 U4026 ( .A1(n4954), .A2(n6251), .ZN(n4613) );
  NOR2_X1 U4027 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6405) );
  CLKBUF_X1 U4028 ( .A(n4527), .Z(n4528) );
  AND2_X1 U4029 ( .A1(n3185), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6061) );
  AND2_X1 U4030 ( .A1(n4615), .A2(n4761), .ZN(n5964) );
  INV_X1 U4031 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4954) );
  CLKBUF_X1 U4032 ( .A(n3229), .Z(n3448) );
  CLKBUF_X1 U4033 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n5224) );
  NAND2_X1 U4034 ( .A1(n4538), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6510) );
  INV_X1 U4035 ( .A(n4978), .ZN(n4538) );
  INV_X1 U4036 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6373) );
  INV_X1 U4037 ( .A(n6060), .ZN(n6035) );
  INV_X1 U4038 ( .A(n6100), .ZN(n4823) );
  AND2_X1 U4039 ( .A1(n4718), .A2(n6329), .ZN(n6108) );
  NOR2_X1 U4040 ( .A1(n6283), .A2(n6118), .ZN(n6139) );
  NOR2_X1 U4041 ( .A1(n6877), .A2(n4761), .ZN(n6269) );
  INV_X1 U4042 ( .A(n6306), .ZN(n6313) );
  INV_X1 U4043 ( .A(n6387), .ZN(n6396) );
  INV_X1 U4044 ( .A(n6269), .ZN(n6444) );
  OR2_X1 U4045 ( .A1(n6411), .A2(n6112), .ZN(n6459) );
  INV_X1 U4046 ( .A(n6476), .ZN(n6455) );
  OR2_X1 U4047 ( .A1(n6411), .A2(n6361), .ZN(n6476) );
  AND2_X1 U4048 ( .A1(n6509), .A2(n6508), .ZN(n6586) );
  NOR2_X1 U4049 ( .A1(n5869), .A2(n5337), .ZN(n5338) );
  AOI21_X1 U4050 ( .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5234), .A(n4437), 
        .ZN(n4438) );
  INV_X1 U4051 ( .A(n4436), .ZN(n4437) );
  NAND2_X1 U4052 ( .A1(n3231), .A2(n5946), .ZN(n3230) );
  NAND2_X2 U4053 ( .A1(n3532), .A2(n3531), .ZN(n4294) );
  NAND2_X1 U4054 ( .A1(n3152), .A2(n4468), .ZN(n4336) );
  NAND2_X1 U4055 ( .A1(n4933), .A2(n4935), .ZN(n4934) );
  NAND2_X1 U4056 ( .A1(n4933), .A2(n3220), .ZN(n5068) );
  NAND2_X1 U4057 ( .A1(n4496), .A2(n4495), .ZN(n4474) );
  NOR2_X1 U4058 ( .A1(n5005), .A2(n5007), .ZN(n5006) );
  AND2_X1 U4059 ( .A1(n5797), .A2(n4932), .ZN(n3208) );
  AND2_X2 U4060 ( .A1(n4534), .A2(n4604), .ZN(n3381) );
  OR2_X1 U4061 ( .A1(n3408), .A2(n6599), .ZN(n3608) );
  AND2_X1 U4062 ( .A1(n3266), .A2(n3221), .ZN(n3209) );
  OR2_X1 U4063 ( .A1(n4772), .A2(n3276), .ZN(n4838) );
  AND2_X1 U4064 ( .A1(n5040), .A2(n3245), .ZN(n3210) );
  INV_X1 U4065 ( .A(n3408), .ZN(n4467) );
  NOR2_X1 U4066 ( .A1(n5023), .A2(n5022), .ZN(n4496) );
  XOR2_X1 U4067 ( .A(n5230), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n3211) );
  AND2_X2 U4068 ( .A1(n3303), .A2(n4587), .ZN(n3386) );
  OR2_X1 U4069 ( .A1(n5005), .A2(n3282), .ZN(n3212) );
  AND2_X2 U4070 ( .A1(n3303), .A2(n4604), .ZN(n3396) );
  NAND2_X1 U4071 ( .A1(n5035), .A2(n5037), .ZN(n5030) );
  AND2_X1 U4072 ( .A1(n4333), .A2(n3240), .ZN(n3214) );
  NAND2_X2 U4073 ( .A1(n3445), .A2(n3531), .ZN(n4511) );
  NOR2_X1 U4074 ( .A1(n4996), .A2(n5020), .ZN(n4201) );
  XNOR2_X1 U4075 ( .A(n3647), .B(n3658), .ZN(n3812) );
  OR2_X1 U4076 ( .A1(n5104), .A2(n5963), .ZN(n3215) );
  NAND2_X1 U4077 ( .A1(n3177), .A2(n3551), .ZN(n3564) );
  AND2_X2 U4078 ( .A1(n3304), .A2(n3315), .ZN(n3391) );
  INV_X1 U4079 ( .A(n3438), .ZN(n3440) );
  AND2_X1 U4080 ( .A1(n4468), .A2(n4512), .ZN(n3216) );
  NAND2_X1 U4081 ( .A1(n4686), .A2(n3435), .ZN(n3523) );
  AND2_X1 U4082 ( .A1(n5050), .A2(n3210), .ZN(n3217) );
  OR2_X1 U4083 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  AND2_X1 U4084 ( .A1(n3409), .A2(n3435), .ZN(n3437) );
  NOR2_X1 U4085 ( .A1(n3252), .A2(n3563), .ZN(n3218) );
  OR2_X1 U4086 ( .A1(n4996), .A2(n3272), .ZN(n5014) );
  NAND2_X1 U4087 ( .A1(n3576), .A2(n4600), .ZN(n4576) );
  NOR2_X1 U4088 ( .A1(n5450), .A2(n5449), .ZN(n5070) );
  INV_X1 U4089 ( .A(n5869), .ZN(n5845) );
  AND2_X1 U4090 ( .A1(n4933), .A2(n3280), .ZN(n5084) );
  NOR2_X1 U4091 ( .A1(n4772), .A2(n3275), .ZN(n3219) );
  INV_X1 U4092 ( .A(n4888), .ZN(n3268) );
  AND2_X1 U4093 ( .A1(n3280), .A2(n5085), .ZN(n3220) );
  INV_X1 U4094 ( .A(n3495), .ZN(n3749) );
  OR2_X1 U4095 ( .A1(n3727), .A2(n3744), .ZN(n3221) );
  INV_X1 U4096 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3228) );
  OR2_X1 U4097 ( .A1(n3272), .A2(n5016), .ZN(n3222) );
  OR2_X1 U4098 ( .A1(n3282), .A2(n5045), .ZN(n3223) );
  OR2_X1 U4099 ( .A1(n3544), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3224)
         );
  AND2_X1 U4100 ( .A1(n3220), .A2(n3279), .ZN(n3225) );
  OR2_X1 U4101 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4232) );
  NAND2_X1 U4102 ( .A1(n3234), .A2(n3235), .ZN(n4774) );
  OR2_X1 U4103 ( .A1(n4423), .A2(n4422), .ZN(n5963) );
  NAND3_X1 U4104 ( .A1(n3575), .A2(n3572), .A3(n3574), .ZN(n4600) );
  INV_X1 U4105 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6599) );
  AND2_X1 U4106 ( .A1(n3243), .A2(n4631), .ZN(n3226) );
  OR2_X1 U4107 ( .A1(n4287), .A2(n4511), .ZN(n4651) );
  INV_X1 U4108 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5517) );
  AND2_X1 U4109 ( .A1(n3533), .A2(n3450), .ZN(n3227) );
  AND2_X2 U4110 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4604) );
  AND2_X4 U4111 ( .A1(n3229), .A2(n3228), .ZN(n4534) );
  NAND3_X1 U4112 ( .A1(n5235), .A2(n5236), .A3(n3230), .ZN(U2988) );
  INV_X2 U4113 ( .A(n3531), .ZN(n4660) );
  NAND2_X1 U4114 ( .A1(n3531), .A2(n3438), .ZN(n3495) );
  NAND2_X1 U4115 ( .A1(n3239), .A2(n3238), .ZN(n5054) );
  NOR2_X1 U4116 ( .A1(n4630), .A2(n3226), .ZN(n5927) );
  INV_X1 U4117 ( .A(n4474), .ZN(n3248) );
  NAND3_X1 U4118 ( .A1(n3576), .A2(n4600), .A3(n6599), .ZN(n3250) );
  NAND2_X1 U4119 ( .A1(n3552), .A2(n3218), .ZN(n3251) );
  NAND2_X1 U4120 ( .A1(n3250), .A2(n3253), .ZN(n3254) );
  NAND2_X1 U4121 ( .A1(n5814), .A2(n3260), .ZN(n3257) );
  NAND2_X1 U4122 ( .A1(n3257), .A2(n3258), .ZN(n4860) );
  OAI21_X1 U4123 ( .B1(n4887), .B2(n4889), .A(n4888), .ZN(n4917) );
  OR2_X2 U4124 ( .A1(n4772), .A2(n3274), .ZN(n4847) );
  NOR2_X1 U4125 ( .A1(n4772), .A2(n4773), .ZN(n4837) );
  INV_X1 U4126 ( .A(n4773), .ZN(n3277) );
  NOR2_X2 U4127 ( .A1(n5005), .A2(n3223), .ZN(n5035) );
  NAND2_X1 U4128 ( .A1(n4527), .A2(n6599), .ZN(n3552) );
  AND2_X1 U4129 ( .A1(n3524), .A2(n4660), .ZN(n3412) );
  AND4_X1 U4130 ( .A1(n3525), .A2(n3524), .A3(n3534), .A4(n3523), .ZN(n3527)
         );
  NAND2_X1 U4131 ( .A1(n3833), .A2(n3408), .ZN(n3452) );
  NAND2_X1 U4132 ( .A1(n5138), .A2(n5864), .ZN(n4212) );
  AOI21_X1 U4133 ( .B1(n5339), .B2(n5876), .A(n5338), .ZN(n5340) );
  NAND2_X1 U4135 ( .A1(n5092), .A2(n5091), .ZN(n5094) );
  NOR2_X1 U4136 ( .A1(n5408), .A2(n4326), .ZN(n3284) );
  OR2_X1 U4137 ( .A1(n4341), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4138 ( .A1(n5112), .A2(n3738), .ZN(n3286) );
  AND2_X1 U4139 ( .A1(n5797), .A2(n5435), .ZN(n3287) );
  AND2_X1 U4140 ( .A1(n5845), .A2(n4488), .ZN(n3288) );
  INV_X1 U4141 ( .A(n3501), .ZN(n3492) );
  INV_X1 U4142 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5466) );
  INV_X1 U4143 ( .A(n6573), .ZN(n6997) );
  AND2_X1 U4144 ( .A1(n4468), .A2(n5251), .ZN(n3289) );
  AND4_X1 U4145 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3290)
         );
  AND2_X1 U4146 ( .A1(n4671), .A2(n3450), .ZN(n3291) );
  OR2_X1 U4147 ( .A1(n5194), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3292)
         );
  AND2_X1 U4148 ( .A1(n5112), .A2(n3295), .ZN(n3293) );
  NAND2_X1 U4149 ( .A1(n5112), .A2(n5183), .ZN(n3294) );
  AND2_X2 U4150 ( .A1(n5878), .A2(n4204), .ZN(n5859) );
  AND2_X1 U4151 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3295) );
  INV_X1 U4152 ( .A(n3452), .ZN(n3453) );
  OR2_X1 U4153 ( .A1(n5674), .A2(n4482), .ZN(n3296) );
  INV_X1 U4154 ( .A(n5086), .ZN(n4472) );
  AND2_X1 U4155 ( .A1(n3804), .A2(n4276), .ZN(n3779) );
  INV_X1 U4156 ( .A(n3658), .ZN(n3659) );
  AND2_X1 U4157 ( .A1(n3784), .A2(n3770), .ZN(n3782) );
  INV_X1 U4158 ( .A(n3523), .ZN(n3833) );
  OR2_X1 U4159 ( .A1(n3644), .A2(n3643), .ZN(n3674) );
  INV_X1 U4160 ( .A(n3588), .ZN(n3626) );
  AND2_X1 U4161 ( .A1(n6283), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3772)
         );
  NOR2_X1 U4162 ( .A1(n4297), .A2(n3408), .ZN(n3529) );
  NAND2_X1 U4163 ( .A1(n3285), .A2(n4332), .ZN(n4333) );
  NAND2_X1 U4164 ( .A1(n3607), .A2(n3606), .ZN(n4601) );
  NAND2_X1 U4165 ( .A1(n3398), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3338)
         );
  AOI22_X1 U4166 ( .A1(n3187), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3323) );
  INV_X1 U4167 ( .A(n4403), .ZN(n4341) );
  OR2_X1 U4168 ( .A1(n6479), .A2(n6599), .ZN(n4230) );
  AND2_X1 U4169 ( .A1(n3827), .A2(EAX_REG_5__SCAN_IN), .ZN(n3851) );
  INV_X1 U4170 ( .A(n4476), .ZN(n4479) );
  INV_X1 U4171 ( .A(n3608), .ZN(n3550) );
  NAND2_X1 U4172 ( .A1(n4586), .A2(n6599), .ZN(n3625) );
  NOR2_X1 U4173 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3793), .ZN(n4282)
         );
  INV_X1 U4174 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3925) );
  INV_X1 U4175 ( .A(n4230), .ZN(n4249) );
  NOR2_X1 U4176 ( .A1(n5186), .A2(n5119), .ZN(n5165) );
  OR3_X1 U4177 ( .A1(n4526), .A2(n4525), .A3(n4650), .ZN(n4599) );
  INV_X1 U4178 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6487) );
  INV_X1 U4179 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U4180 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3989)
         );
  INV_X1 U4181 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5574) );
  AOI21_X1 U4182 ( .B1(n5845), .B2(n4489), .A(n4208), .ZN(n4209) );
  NAND2_X1 U4183 ( .A1(n4059), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4089)
         );
  NAND2_X1 U4184 ( .A1(n4004), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4031)
         );
  INV_X1 U4185 ( .A(n5194), .ZN(n5797) );
  INV_X1 U4186 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U4187 ( .A1(n5361), .A2(n3293), .ZN(n5113) );
  NOR2_X1 U4188 ( .A1(n5366), .A2(n3287), .ZN(n5361) );
  INV_X1 U4189 ( .A(n5880), .ZN(n5209) );
  INV_X1 U4190 ( .A(n5958), .ZN(n5938) );
  OR3_X1 U4191 ( .A1(n4652), .A2(n4291), .A3(n4295), .ZN(n4292) );
  INV_X1 U4192 ( .A(n4635), .ZN(n6033) );
  AND2_X1 U4193 ( .A1(n4796), .A2(n4795), .ZN(n6097) );
  INV_X1 U4194 ( .A(n4761), .ZN(n6151) );
  INV_X1 U4195 ( .A(n3657), .ZN(n4636) );
  INV_X1 U4196 ( .A(n3155), .ZN(n6147) );
  NAND2_X1 U4197 ( .A1(n3492), .A2(n3502), .ZN(n3493) );
  INV_X1 U4198 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6283) );
  AND2_X1 U4199 ( .A1(n4954), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3807) );
  INV_X1 U4200 ( .A(n6597), .ZN(n4987) );
  INV_X1 U4201 ( .A(n5641), .ZN(n5652) );
  AND2_X1 U4202 ( .A1(n5090), .A2(n5089), .ZN(n5091) );
  INV_X1 U4203 ( .A(n5090), .ZN(n5687) );
  NOR2_X1 U4204 ( .A1(n4833), .A2(n5692), .ZN(n5709) );
  OAI21_X1 U4205 ( .B1(n6597), .B2(n6896), .A(n5712), .ZN(n5740) );
  INV_X1 U4206 ( .A(n5713), .ZN(n5790) );
  OAI21_X1 U4207 ( .B1(n5097), .B2(n6412), .A(n4209), .ZN(n4210) );
  NAND2_X1 U4208 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3862)
         );
  NAND2_X1 U4209 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3843) );
  OR2_X2 U4210 ( .A1(n4978), .A2(n6519), .ZN(n4652) );
  NOR2_X1 U4211 ( .A1(n5209), .A2(n4314), .ZN(n5448) );
  NAND2_X1 U4212 ( .A1(n4313), .A2(n5955), .ZN(n5910) );
  INV_X1 U4213 ( .A(n5963), .ZN(n5946) );
  NAND2_X1 U4214 ( .A1(n4954), .A2(n6373), .ZN(n6521) );
  INV_X1 U4215 ( .A(n5982), .ZN(n5991) );
  INV_X1 U4216 ( .A(n6022), .ZN(n6024) );
  AND2_X1 U4217 ( .A1(n6033), .A2(n6032), .ZN(n6086) );
  AND2_X1 U4218 ( .A1(n4718), .A2(n6282), .ZN(n6100) );
  OAI21_X1 U4219 ( .B1(n6096), .B2(n6373), .A(n4793), .ZN(n6101) );
  OAI21_X1 U4220 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6373), .A(n6151), 
        .ZN(n6416) );
  INV_X1 U4221 ( .A(n6135), .ZN(n6138) );
  INV_X1 U4222 ( .A(n6208), .ZN(n6199) );
  OAI21_X1 U4223 ( .B1(n6217), .B2(n6247), .A(n6216), .ZN(n6237) );
  INV_X1 U4224 ( .A(n6281), .ZN(n6263) );
  AND2_X1 U4225 ( .A1(n3185), .A2(n6329), .ZN(n6243) );
  INV_X1 U4226 ( .A(n6282), .ZN(n6329) );
  AND2_X1 U4227 ( .A1(n3807), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6522) );
  INV_X1 U4228 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U4229 ( .A1(n5237), .A2(n5238), .ZN(n6604) );
  INV_X1 U4230 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6596) );
  AOI22_X1 U4231 ( .A1(n5244), .A2(n5652), .B1(REIP_REG_30__SCAN_IN), .B2(
        n5243), .ZN(n5245) );
  OR2_X1 U4232 ( .A1(n4511), .A2(n4446), .ZN(n5641) );
  INV_X1 U4233 ( .A(n5638), .ZN(n5654) );
  INV_X1 U4234 ( .A(n5592), .ZN(n5599) );
  INV_X1 U4235 ( .A(n5601), .ZN(n5655) );
  NAND2_X1 U4236 ( .A1(n4653), .A2(n5713), .ZN(n5090) );
  INV_X1 U4237 ( .A(n5692), .ZN(n5711) );
  OR2_X2 U4238 ( .A1(n4652), .A2(n6505), .ZN(n5793) );
  INV_X1 U4239 ( .A(n4210), .ZN(n4211) );
  OR2_X1 U4240 ( .A1(n5859), .A2(n5873), .ZN(n5869) );
  AND2_X1 U4241 ( .A1(n5169), .A2(n4323), .ZN(n5420) );
  NAND2_X1 U4242 ( .A1(n4703), .A2(n4546), .ZN(n5951) );
  INV_X1 U4243 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6493) );
  NOR2_X1 U4244 ( .A1(n6585), .A2(n5463), .ZN(n5223) );
  NAND2_X1 U4245 ( .A1(n5996), .A2(n6329), .ZN(n6060) );
  OR2_X1 U4246 ( .A1(n4787), .A2(n4635), .ZN(n6104) );
  NAND2_X1 U4247 ( .A1(n4710), .A2(n6210), .ZN(n6135) );
  OR2_X1 U4248 ( .A1(n6113), .A2(n6112), .ZN(n6176) );
  NAND2_X1 U4249 ( .A1(n6178), .A2(n6329), .ZN(n6241) );
  NAND2_X1 U4250 ( .A1(n6244), .A2(n6210), .ZN(n6281) );
  NAND2_X1 U4251 ( .A1(n6330), .A2(n6282), .ZN(n6351) );
  INV_X1 U4252 ( .A(n6224), .ZN(n6443) );
  INV_X1 U4253 ( .A(n6522), .ZN(n6519) );
  INV_X1 U4254 ( .A(n6583), .ZN(n6580) );
  NOR2_X1 U4255 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6915), .ZN(n6573) );
  NAND2_X1 U4256 ( .A1(n4485), .A2(n4484), .ZN(U2829) );
  NAND2_X1 U4257 ( .A1(n4212), .A2(n4211), .ZN(U2958) );
  INV_X1 U4258 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4259 ( .A1(n3188), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3302) );
  AND2_X4 U4260 ( .A1(n3298), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4587)
         );
  NOR2_X4 U4261 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3315) );
  AND2_X2 U4262 ( .A1(n4535), .A2(n4604), .ZN(n3398) );
  AOI22_X1 U4263 ( .A1(n3204), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4264 ( .A1(n3386), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3417), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3308) );
  AND2_X4 U4265 ( .A1(n4534), .A2(n3315), .ZN(n3380) );
  AOI22_X1 U4266 ( .A1(n3617), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3305) );
  NAND2_X2 U4267 ( .A1(n3310), .A2(n3309), .ZN(n3409) );
  AOI22_X1 U4268 ( .A1(n3197), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4269 ( .A1(n3617), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4270 ( .A1(n3417), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3611), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3311) );
  AND4_X2 U4271 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3321)
         );
  AOI22_X1 U4272 ( .A1(n3610), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4273 ( .A1(n3396), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4274 ( .A1(n3187), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4275 ( .A1(n3315), .A2(n4535), .ZN(n3513) );
  INV_X2 U4276 ( .A(n3513), .ZN(n3476) );
  AOI22_X1 U4277 ( .A1(n3205), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4278 ( .A1(n3617), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4279 ( .A1(n3610), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3611), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4280 ( .A1(n3205), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4281 ( .A1(n3612), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4282 ( .A1(n3512), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4283 ( .A1(n3386), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3417), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4284 ( .A1(n3157), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3326) );
  NAND2_X2 U4285 ( .A1(n3330), .A2(n3290), .ZN(n3532) );
  NAND2_X1 U4286 ( .A1(n4654), .A2(n3532), .ZN(n3524) );
  NAND2_X1 U4287 ( .A1(n3386), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4288 ( .A1(n3417), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4289 ( .A1(n3187), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4290 ( .A1(n3611), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3331)
         );
  NAND2_X1 U4291 ( .A1(n3617), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3337)
         );
  NAND2_X1 U4292 ( .A1(n3196), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3336)
         );
  NAND2_X1 U4293 ( .A1(n3381), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4294 ( .A1(n3188), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4295 ( .A1(n3512), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U4296 ( .A1(n3396), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3340)
         );
  NAND2_X1 U4297 ( .A1(n3391), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4298 ( .A1(n3198), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4299 ( .A1(n3380), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4300 ( .A1(n3610), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4301 ( .A1(n3204), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4302 ( .A1(n3612), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4303 ( .A1(n3512), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4304 ( .A1(n3396), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4305 ( .A1(n3391), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4306 ( .A1(n3197), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4307 ( .A1(n3386), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4308 ( .A1(n3417), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4309 ( .A1(n3380), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4310 ( .A1(n3617), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3362)
         );
  NAND2_X1 U4311 ( .A1(n3196), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3361)
         );
  NAND2_X1 U4312 ( .A1(n3187), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3360) );
  NAND2_X1 U4313 ( .A1(n3381), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3359)
         );
  NAND2_X1 U4314 ( .A1(n3610), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4315 ( .A1(n3611), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3365)
         );
  NAND2_X1 U4316 ( .A1(n3398), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4317 ( .A1(n3204), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4318 ( .A1(n3194), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3417), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4319 ( .A1(n3611), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4320 ( .A1(n3187), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4321 ( .A1(n3525), .A2(n3523), .ZN(n3407) );
  NAND2_X1 U4322 ( .A1(n3610), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4323 ( .A1(n3617), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3384)
         );
  NAND2_X1 U4324 ( .A1(n3380), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4325 ( .A1(n3381), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3382)
         );
  NAND2_X1 U4326 ( .A1(n3386), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4327 ( .A1(n3157), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4328 ( .A1(n3611), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4329 ( .A1(n3204), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4330 ( .A1(n3512), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4331 ( .A1(n3188), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4332 ( .A1(n3391), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4333 ( .A1(n3417), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3392) );
  NAND2_X1 U4334 ( .A1(n3195), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3402)
         );
  NAND2_X1 U4335 ( .A1(n3396), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3401)
         );
  NAND2_X1 U4336 ( .A1(n3187), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3400) );
  NAND2_X1 U4337 ( .A1(n3398), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3399)
         );
  NAND2_X1 U4338 ( .A1(n3407), .A2(n4295), .ZN(n3411) );
  NAND3_X1 U4339 ( .A1(n3412), .A2(n3411), .A3(n3526), .ZN(n3434) );
  NAND2_X1 U4340 ( .A1(n3612), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3416) );
  NAND2_X1 U4341 ( .A1(n3512), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4342 ( .A1(n3396), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3414)
         );
  NAND2_X1 U4343 ( .A1(n3391), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4344 ( .A1(n3197), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3421) );
  NAND2_X1 U4345 ( .A1(n3386), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4346 ( .A1(n3417), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3419) );
  NAND2_X1 U4347 ( .A1(n3380), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4348 ( .A1(n3617), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3425)
         );
  NAND2_X1 U4349 ( .A1(n3194), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3424)
         );
  NAND2_X1 U4350 ( .A1(n3187), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4351 ( .A1(n3381), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3422)
         );
  NAND2_X1 U4352 ( .A1(n3610), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3429) );
  NAND2_X1 U4353 ( .A1(n3611), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3428)
         );
  NAND2_X1 U4354 ( .A1(n3398), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3427)
         );
  NAND2_X1 U4355 ( .A1(n3204), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3426) );
  NAND4_X4 U4356 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), .ZN(n3445)
         );
  NAND2_X1 U4357 ( .A1(n3434), .A2(n3534), .ZN(n3451) );
  NAND2_X1 U4358 ( .A1(n3525), .A2(n3435), .ZN(n4271) );
  NAND2_X1 U4359 ( .A1(n4271), .A2(n3496), .ZN(n3436) );
  NAND2_X1 U4360 ( .A1(n3184), .A2(n3532), .ZN(n4529) );
  NAND2_X1 U4361 ( .A1(n4467), .A2(n3438), .ZN(n3752) );
  NAND2_X1 U4362 ( .A1(n3833), .A2(n3752), .ZN(n3528) );
  NAND2_X1 U4363 ( .A1(n3437), .A2(n3438), .ZN(n3439) );
  NAND2_X1 U4364 ( .A1(n3528), .A2(n3439), .ZN(n3808) );
  NAND2_X1 U4365 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6548) );
  OAI21_X1 U4366 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6548), .ZN(n4283) );
  INV_X1 U4367 ( .A(n4283), .ZN(n3536) );
  OAI21_X1 U4368 ( .B1(n3536), .B2(n3531), .A(n3440), .ZN(n3441) );
  NAND3_X1 U4369 ( .A1(n3451), .A2(n3459), .A3(n3443), .ZN(n3444) );
  NAND2_X1 U4370 ( .A1(n3444), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4371 ( .A1(n3776), .A2(n4654), .ZN(n3446) );
  INV_X1 U4372 ( .A(n3807), .ZN(n3539) );
  MUX2_X1 U4373 ( .A(n3539), .B(n6602), .S(n6283), .Z(n3449) );
  OAI22_X1 U4374 ( .A1(n3160), .A2(n3184), .B1(n3534), .B2(n3450), .ZN(n4302)
         );
  NAND2_X1 U4375 ( .A1(n3453), .A2(n3454), .ZN(n4594) );
  OR2_X1 U4376 ( .A1(n6521), .A2(n6599), .ZN(n3455) );
  AOI21_X1 U4377 ( .B1(n3524), .B2(n3496), .A(n3455), .ZN(n3460) );
  AOI21_X1 U4378 ( .B1(n4654), .B2(n3408), .A(n4671), .ZN(n3456) );
  NAND2_X1 U4379 ( .A1(n3808), .A2(n3456), .ZN(n3457) );
  NAND2_X1 U4380 ( .A1(n3457), .A2(n3531), .ZN(n3458) );
  NAND4_X1 U4381 ( .A1(n4594), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(n3461)
         );
  OR2_X2 U4382 ( .A1(n3462), .A2(n3463), .ZN(n3566) );
  NAND2_X1 U4383 ( .A1(n3462), .A2(n3463), .ZN(n3464) );
  AOI22_X1 U4384 ( .A1(n3154), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3167), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4385 ( .A1(n3203), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4386 ( .A1(n3194), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4387 ( .A1(n3994), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3465) );
  NAND4_X1 U4388 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3474)
         );
  AOI22_X1 U4389 ( .A1(n3507), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4390 ( .A1(n3157), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4391 ( .A1(n3476), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4392 ( .A1(n3190), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3469) );
  NAND4_X1 U4393 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), .ZN(n3473)
         );
  INV_X1 U4394 ( .A(n3554), .ZN(n3487) );
  AOI22_X1 U4395 ( .A1(n3154), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4396 ( .A1(n3197), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3167), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4397 ( .A1(n3869), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4398 ( .A1(n3203), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4399 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3486)
         );
  AOI22_X1 U4400 ( .A1(n3190), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4401 ( .A1(n3507), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4402 ( .A1(n3397), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4403 ( .A1(n3994), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4404 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485)
         );
  XNOR2_X1 U4405 ( .A(n3487), .B(n3719), .ZN(n3488) );
  NAND2_X1 U4406 ( .A1(n3488), .A2(n3550), .ZN(n3502) );
  NAND2_X1 U4407 ( .A1(n3776), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3490) );
  AOI21_X1 U4408 ( .B1(n3534), .B2(n3554), .A(n6599), .ZN(n3489) );
  OAI211_X1 U4409 ( .C1(n3722), .C2(n3408), .A(n3490), .B(n3489), .ZN(n3501)
         );
  NAND2_X1 U4410 ( .A1(n3534), .A2(n3532), .ZN(n3594) );
  OAI21_X1 U4411 ( .B1(n4987), .B2(n3554), .A(n3594), .ZN(n3497) );
  INV_X1 U4412 ( .A(n3497), .ZN(n3498) );
  NAND2_X1 U4413 ( .A1(n5871), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5870)
         );
  INV_X1 U4414 ( .A(n5870), .ZN(n3499) );
  INV_X1 U4415 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U4416 ( .A1(n3499), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3560)
         );
  NAND2_X1 U4417 ( .A1(n5870), .A2(n4549), .ZN(n3500) );
  AND2_X1 U4418 ( .A1(n3560), .A2(n3500), .ZN(n4545) );
  NAND2_X1 U4419 ( .A1(n3159), .A2(n6599), .ZN(n3506) );
  OR2_X1 U4420 ( .A1(n3492), .A2(n3502), .ZN(n3504) );
  NAND2_X1 U4421 ( .A1(n3550), .A2(n3719), .ZN(n3503) );
  AOI22_X1 U4422 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3154), .B1(n3507), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4423 ( .A1(n3198), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4424 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3475), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4425 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n3397), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3508) );
  NAND4_X1 U4426 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3519)
         );
  AOI22_X1 U4427 ( .A1(n3203), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4428 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3190), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4429 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n3199), .B1(n3380), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4430 ( .A1(n3476), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U4431 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3518)
         );
  INV_X1 U4432 ( .A(n3555), .ZN(n3522) );
  NAND2_X1 U4433 ( .A1(n3776), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3521) );
  NAND2_X1 U4434 ( .A1(n3550), .A2(n3722), .ZN(n3520) );
  OAI211_X1 U4435 ( .C1(n3522), .C2(n3609), .A(n3521), .B(n3520), .ZN(n3563)
         );
  INV_X1 U4436 ( .A(n3528), .ZN(n3530) );
  INV_X1 U4437 ( .A(n4651), .ZN(n4516) );
  NOR2_X1 U4438 ( .A1(n4287), .A2(n3534), .ZN(n4441) );
  NOR2_X1 U4439 ( .A1(n3438), .A2(n3532), .ZN(n3533) );
  INV_X1 U4440 ( .A(n4977), .ZN(n3535) );
  INV_X1 U4441 ( .A(n4656), .ZN(n4288) );
  NAND2_X1 U4442 ( .A1(n4421), .A2(n3537), .ZN(n3538) );
  INV_X1 U4443 ( .A(n3545), .ZN(n3542) );
  XNOR2_X1 U4444 ( .A(n6487), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6364)
         );
  NAND2_X1 U4445 ( .A1(n6602), .A2(n6364), .ZN(n3541) );
  NAND2_X1 U4446 ( .A1(n3539), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U4447 ( .A1(n3541), .A2(n3540), .ZN(n3544) );
  NAND2_X1 U4448 ( .A1(n3542), .A2(n3224), .ZN(n3565) );
  INV_X1 U4449 ( .A(n3567), .ZN(n3547) );
  INV_X1 U4450 ( .A(n3544), .ZN(n3546) );
  OAI211_X2 U4451 ( .C1(n3547), .C2(n3543), .A(n3546), .B(n3545), .ZN(n3572)
         );
  NAND2_X1 U4452 ( .A1(n3565), .A2(n3572), .ZN(n3549) );
  INV_X1 U4453 ( .A(n3172), .ZN(n3548) );
  NAND2_X1 U4454 ( .A1(n3550), .A2(n3555), .ZN(n3551) );
  NAND2_X1 U4455 ( .A1(n3155), .A2(n3749), .ZN(n3559) );
  NAND2_X1 U4456 ( .A1(n3554), .A2(n3555), .ZN(n3627) );
  OAI21_X1 U4457 ( .B1(n3555), .B2(n3554), .A(n3627), .ZN(n3556) );
  OAI211_X1 U4458 ( .C1(n3556), .C2(n4987), .A(n3809), .B(n3438), .ZN(n3557)
         );
  INV_X1 U4459 ( .A(n3557), .ZN(n3558) );
  NAND2_X1 U4460 ( .A1(n3559), .A2(n3558), .ZN(n4544) );
  NAND2_X1 U4461 ( .A1(n4545), .A2(n4544), .ZN(n3561) );
  AND2_X1 U4462 ( .A1(n3561), .A2(n3560), .ZN(n5863) );
  NAND2_X1 U4463 ( .A1(n3575), .A2(n3572), .ZN(n3571) );
  BUF_X1 U4464 ( .A(n3567), .Z(n3602) );
  INV_X1 U4465 ( .A(n6602), .ZN(n3604) );
  OR2_X1 U4466 ( .A1(n6487), .A2(n6283), .ZN(n3569) );
  NAND3_X1 U4467 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6209), .ZN(n6242) );
  INV_X1 U4468 ( .A(n6242), .ZN(n3568) );
  AOI21_X1 U4469 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3569), .A(n3568), 
        .ZN(n4666) );
  OAI22_X1 U4470 ( .A1(n3604), .A2(n4666), .B1(n3807), .B2(n6209), .ZN(n3570)
         );
  NAND2_X1 U4471 ( .A1(n3571), .A2(n3573), .ZN(n3576) );
  INV_X1 U4472 ( .A(n3573), .ZN(n3574) );
  AOI22_X1 U4473 ( .A1(n3154), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4474 ( .A1(n3199), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4475 ( .A1(n3994), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4476 ( .A1(n3157), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4477 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3587)
         );
  AOI22_X1 U4478 ( .A1(n3203), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4479 ( .A1(n3190), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4480 ( .A1(n3476), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4481 ( .A1(n3397), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4482 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  INV_X1 U4483 ( .A(n3609), .ZN(n3589) );
  AOI22_X1 U4484 ( .A1(n3776), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3589), 
        .B2(n3588), .ZN(n3590) );
  NAND2_X1 U4485 ( .A1(n4634), .A2(n3749), .ZN(n3597) );
  XNOR2_X1 U4486 ( .A(n3627), .B(n3626), .ZN(n3595) );
  INV_X1 U4487 ( .A(n3594), .ZN(n4303) );
  AOI21_X1 U4488 ( .B1(n3595), .B2(n6597), .A(n4303), .ZN(n3596) );
  NAND2_X1 U4489 ( .A1(n3597), .A2(n3596), .ZN(n5861) );
  NAND2_X1 U4490 ( .A1(n5861), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3598)
         );
  NAND2_X1 U4491 ( .A1(n5863), .A2(n3598), .ZN(n3601) );
  INV_X1 U4492 ( .A(n5861), .ZN(n3599) );
  INV_X1 U4493 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U4494 ( .A1(n3599), .A2(n5936), .ZN(n3600) );
  AND2_X2 U4495 ( .A1(n3601), .A2(n3600), .ZN(n5851) );
  NAND2_X1 U4496 ( .A1(n3602), .A2(n5224), .ZN(n3607) );
  NAND3_X1 U4497 ( .A1(n6493), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6118) );
  NAND3_X1 U4498 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6418) );
  NOR2_X1 U4499 ( .A1(n6283), .A2(n6418), .ZN(n6469) );
  INV_X1 U4500 ( .A(n6469), .ZN(n6446) );
  NAND2_X1 U4501 ( .A1(n3603), .A2(n6446), .ZN(n6144) );
  OAI22_X1 U4502 ( .A1(n6144), .A2(n3604), .B1(n3807), .B2(n6493), .ZN(n3605)
         );
  INV_X1 U4503 ( .A(n3605), .ZN(n3606) );
  XNOR2_X1 U4504 ( .A(n4600), .B(n4601), .ZN(n4586) );
  AOI22_X1 U4505 ( .A1(n4216), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4506 ( .A1(n3203), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4507 ( .A1(n3661), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4508 ( .A1(n3154), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4509 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3623)
         );
  AOI22_X1 U4510 ( .A1(n3199), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4511 ( .A1(n3190), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4512 ( .A1(n3195), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4513 ( .A1(n3157), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3618) );
  NAND4_X1 U4514 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3622)
         );
  AOI22_X1 U4515 ( .A1(n3804), .A2(n3648), .B1(n3776), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3624) );
  NAND2_X2 U4516 ( .A1(n3625), .A2(n3624), .ZN(n3657) );
  XNOR2_X2 U4517 ( .A(n3656), .B(n3657), .ZN(n4635) );
  NAND2_X1 U4518 ( .A1(n4635), .A2(n3749), .ZN(n3631) );
  NAND2_X1 U4519 ( .A1(n3627), .A2(n3626), .ZN(n3649) );
  INV_X1 U4520 ( .A(n3648), .ZN(n3628) );
  XNOR2_X1 U4521 ( .A(n3649), .B(n3628), .ZN(n3629) );
  NAND2_X1 U4522 ( .A1(n3629), .A2(n6597), .ZN(n3630) );
  NAND2_X1 U4523 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  INV_X1 U4524 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U4525 ( .A(n3632), .B(n5934), .ZN(n5852) );
  NAND2_X1 U4526 ( .A1(n5851), .A2(n5852), .ZN(n5850) );
  NAND2_X1 U4527 ( .A1(n3632), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3633)
         );
  NAND2_X1 U4528 ( .A1(n5850), .A2(n3633), .ZN(n4701) );
  INV_X1 U4529 ( .A(n3656), .ZN(n3634) );
  NAND2_X1 U4530 ( .A1(n3634), .A2(n3657), .ZN(n3647) );
  AOI22_X1 U4531 ( .A1(n3507), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3638) );
  INV_X1 U4532 ( .A(n3964), .ZN(n3661) );
  AOI22_X1 U4533 ( .A1(n3661), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4534 ( .A1(n3192), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4535 ( .A1(n3190), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3635) );
  NAND4_X1 U4536 ( .A1(n3638), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3644)
         );
  AOI22_X1 U4537 ( .A1(n3154), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4538 ( .A1(n3197), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4539 ( .A1(n3203), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4540 ( .A1(n3186), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4541 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3643)
         );
  NAND2_X1 U4542 ( .A1(n3804), .A2(n3674), .ZN(n3646) );
  NAND2_X1 U4543 ( .A1(n3776), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4544 ( .A1(n3812), .A2(n3749), .ZN(n3653) );
  AND2_X1 U4545 ( .A1(n3649), .A2(n3648), .ZN(n3675) );
  INV_X1 U4546 ( .A(n3674), .ZN(n3650) );
  XNOR2_X1 U4547 ( .A(n3675), .B(n3650), .ZN(n3651) );
  NAND2_X1 U4548 ( .A1(n3651), .A2(n6597), .ZN(n3652) );
  NAND2_X1 U4549 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  INV_X1 U4550 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4704) );
  XNOR2_X1 U4551 ( .A(n3654), .B(n4704), .ZN(n4700) );
  NAND2_X1 U4552 ( .A1(n3654), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3655)
         );
  NAND2_X1 U4553 ( .A1(n4699), .A2(n3655), .ZN(n5836) );
  AOI22_X1 U4554 ( .A1(n3154), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4555 ( .A1(n3199), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4556 ( .A1(n3661), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4557 ( .A1(n3157), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4558 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4559 ( .A1(n3203), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4560 ( .A1(n3190), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4561 ( .A1(n3476), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4562 ( .A1(n3397), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4563 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NAND2_X1 U4564 ( .A1(n3804), .A2(n3700), .ZN(n3673) );
  NAND2_X1 U4565 ( .A1(n3776), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4566 ( .A1(n3852), .A2(n3749), .ZN(n3678) );
  NAND2_X1 U4567 ( .A1(n3675), .A2(n3674), .ZN(n3701) );
  XNOR2_X1 U4568 ( .A(n3700), .B(n3701), .ZN(n3676) );
  NAND2_X1 U4569 ( .A1(n6597), .A2(n3676), .ZN(n3677) );
  NAND2_X1 U4570 ( .A1(n3678), .A2(n3677), .ZN(n3679) );
  INV_X1 U4571 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5912) );
  XNOR2_X1 U4572 ( .A(n3679), .B(n5912), .ZN(n5835) );
  NAND2_X1 U4573 ( .A1(n5836), .A2(n5835), .ZN(n5838) );
  NAND2_X1 U4574 ( .A1(n3679), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3680)
         );
  AOI22_X1 U4575 ( .A1(n3154), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4576 ( .A1(n3199), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4577 ( .A1(n3661), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4578 ( .A1(n3197), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4579 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4580 ( .A1(n3203), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4581 ( .A1(n3190), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4582 ( .A1(n3476), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4583 ( .A1(n3397), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4584 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  NAND2_X1 U4585 ( .A1(n3804), .A2(n3712), .ZN(n3695) );
  NAND2_X1 U4586 ( .A1(n3776), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4587 ( .A1(n3699), .A2(n3698), .ZN(n3859) );
  NAND3_X1 U4588 ( .A1(n3711), .A2(n3749), .A3(n3859), .ZN(n3705) );
  INV_X1 U4589 ( .A(n3700), .ZN(n3702) );
  NOR2_X1 U4590 ( .A1(n3702), .A2(n3701), .ZN(n3713) );
  XOR2_X1 U4591 ( .A(n3712), .B(n3713), .Z(n3703) );
  NAND2_X1 U4592 ( .A1(n3703), .A2(n6597), .ZN(n3704) );
  NAND2_X1 U4593 ( .A1(n3705), .A2(n3704), .ZN(n3706) );
  INV_X1 U4594 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U4595 ( .A(n3706), .B(n5917), .ZN(n5829) );
  NAND2_X1 U4596 ( .A1(n3164), .A2(n3180), .ZN(n5828) );
  NAND2_X1 U4597 ( .A1(n3706), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3707)
         );
  NAND2_X1 U4598 ( .A1(n5828), .A2(n3707), .ZN(n5822) );
  NAND2_X1 U4599 ( .A1(n3804), .A2(n3719), .ZN(n3709) );
  NAND2_X1 U4600 ( .A1(n3776), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4601 ( .A1(n3709), .A2(n3708), .ZN(n3710) );
  NAND2_X1 U4602 ( .A1(n3860), .A2(n3749), .ZN(n3716) );
  NAND2_X1 U4603 ( .A1(n3713), .A2(n3712), .ZN(n3721) );
  XNOR2_X1 U4604 ( .A(n3719), .B(n3721), .ZN(n3714) );
  NAND2_X1 U4605 ( .A1(n3714), .A2(n6597), .ZN(n3715) );
  NAND2_X1 U4606 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5906) );
  XNOR2_X1 U4608 ( .A(n3717), .B(n5906), .ZN(n5821) );
  NAND2_X1 U4609 ( .A1(n5822), .A2(n5821), .ZN(n5820) );
  NAND2_X1 U4610 ( .A1(n3717), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3718)
         );
  NOR2_X1 U4611 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  NAND2_X1 U4612 ( .A1(n3723), .A2(n6597), .ZN(n3724) );
  NAND2_X1 U4613 ( .A1(n3727), .A2(n3724), .ZN(n3725) );
  INV_X1 U4614 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U4615 ( .A(n3725), .B(n5900), .ZN(n5813) );
  NAND2_X1 U4616 ( .A1(n3725), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3726)
         );
  INV_X2 U4617 ( .A(n5194), .ZN(n5112) );
  INV_X1 U4618 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U4619 ( .A1(n5112), .A2(n5892), .ZN(n5804) );
  OR2_X1 U4620 ( .A1(n5112), .A2(n5892), .ZN(n5805) );
  INV_X1 U4621 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4622 ( .A1(n5112), .A2(n3728), .ZN(n4859) );
  NAND2_X1 U4623 ( .A1(n4860), .A2(n4859), .ZN(n5796) );
  AND2_X1 U4624 ( .A1(n5112), .A2(n5884), .ZN(n3731) );
  OR2_X1 U4625 ( .A1(n5112), .A2(n3728), .ZN(n5795) );
  OAI21_X1 U4626 ( .B1(n5884), .B2(n3727), .A(n5795), .ZN(n3729) );
  INV_X1 U4627 ( .A(n3729), .ZN(n3730) );
  INV_X1 U4628 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3732) );
  NOR2_X1 U4629 ( .A1(n5112), .A2(n3732), .ZN(n4889) );
  NAND2_X1 U4630 ( .A1(n5797), .A2(n3732), .ZN(n4888) );
  XNOR2_X1 U4631 ( .A(n5797), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4918)
         );
  INV_X1 U4632 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4932) );
  INV_X1 U4633 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3733) );
  AND2_X1 U4634 ( .A1(n5112), .A2(n3733), .ZN(n3735) );
  OR2_X1 U4635 ( .A1(n5112), .A2(n3733), .ZN(n3734) );
  INV_X1 U4636 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5201) );
  NOR2_X1 U4637 ( .A1(n3727), .A2(n5201), .ZN(n3737) );
  NAND2_X1 U4638 ( .A1(n5797), .A2(n5201), .ZN(n3736) );
  INV_X1 U4639 ( .A(n5195), .ZN(n3739) );
  NAND3_X1 U4640 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3738) );
  NAND2_X1 U4641 ( .A1(n3739), .A2(n3286), .ZN(n5123) );
  INV_X1 U4642 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5200) );
  INV_X1 U4643 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5442) );
  INV_X1 U4644 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5447) );
  AND3_X1 U4645 ( .A1(n5200), .A2(n5442), .A3(n5447), .ZN(n3740) );
  OR2_X1 U4646 ( .A1(n5112), .A2(n3740), .ZN(n3741) );
  AND2_X1 U4647 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5178) );
  AND2_X1 U4648 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U4649 ( .A1(n5178), .A2(n3742), .ZN(n5119) );
  NAND2_X1 U4650 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4321) );
  OAI21_X1 U4651 ( .B1(n5119), .B2(n4321), .A(n3727), .ZN(n3745) );
  NOR2_X1 U4652 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5177) );
  NOR2_X1 U4653 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3743) );
  INV_X1 U4654 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5435) );
  INV_X1 U4655 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5168) );
  AND4_X1 U4656 ( .A1(n5177), .A2(n3743), .A3(n5435), .A4(n5168), .ZN(n3744)
         );
  OR2_X1 U4657 ( .A1(n5112), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5146)
         );
  NOR2_X1 U4658 ( .A1(n5146), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3746)
         );
  XNOR2_X1 U4659 ( .A(n5797), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5354)
         );
  INV_X1 U4660 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5409) );
  OAI22_X1 U4661 ( .A1(n5342), .A2(n3747), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5409), .ZN(n3748) );
  XNOR2_X1 U4662 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(n3748), .ZN(n5138)
         );
  AND2_X1 U4663 ( .A1(n3448), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3750)
         );
  NOR2_X1 U4664 ( .A1(n3772), .A2(n3750), .ZN(n3755) );
  NAND2_X1 U4665 ( .A1(n3804), .A2(n3755), .ZN(n3751) );
  NAND2_X1 U4666 ( .A1(n3797), .A2(n3751), .ZN(n3759) );
  INV_X1 U4667 ( .A(n3753), .ZN(n3754) );
  AOI21_X1 U4668 ( .B1(n3752), .B2(n3755), .A(n3754), .ZN(n3757) );
  NAND2_X1 U4669 ( .A1(n4660), .A2(n3438), .ZN(n3756) );
  NAND2_X1 U4670 ( .A1(n4977), .A2(n3756), .ZN(n3778) );
  OR2_X1 U4671 ( .A1(n3757), .A2(n3778), .ZN(n3758) );
  NAND2_X1 U4672 ( .A1(n3759), .A2(n3758), .ZN(n3765) );
  NAND2_X1 U4673 ( .A1(n3804), .A2(n3531), .ZN(n3764) );
  XNOR2_X1 U4674 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3771) );
  INV_X1 U4675 ( .A(n3771), .ZN(n3760) );
  XNOR2_X1 U4676 ( .A(n3760), .B(n3772), .ZN(n4277) );
  NAND4_X1 U4677 ( .A1(n3765), .A2(n3438), .A3(n3764), .A4(n4277), .ZN(n3763)
         );
  NAND2_X1 U4678 ( .A1(n4277), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4679 ( .A1(n3797), .A2(n3761), .ZN(n3762) );
  NAND2_X1 U4680 ( .A1(n3763), .A2(n3762), .ZN(n3769) );
  INV_X1 U4681 ( .A(n3764), .ZN(n3767) );
  INV_X1 U4682 ( .A(n3765), .ZN(n3766) );
  OAI21_X1 U4683 ( .B1(n3440), .B2(n3767), .A(n3766), .ZN(n3768) );
  NAND2_X1 U4684 ( .A1(n3769), .A2(n3768), .ZN(n3781) );
  NAND2_X1 U4685 ( .A1(n6209), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4686 ( .A1(n3166), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3770) );
  INV_X1 U4687 ( .A(n3782), .ZN(n3775) );
  NAND2_X1 U4688 ( .A1(n3772), .A2(n3771), .ZN(n3774) );
  NAND2_X1 U4689 ( .A1(n6487), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4690 ( .A1(n3774), .A2(n3773), .ZN(n3783) );
  XNOR2_X1 U4691 ( .A(n3775), .B(n3783), .ZN(n4276) );
  NOR2_X1 U4692 ( .A1(n3794), .A2(n4276), .ZN(n3777) );
  AOI22_X1 U4693 ( .A1(n3781), .A2(n3780), .B1(n3779), .B2(n3778), .ZN(n3788)
         );
  NAND2_X1 U4694 ( .A1(n3783), .A2(n3782), .ZN(n3785) );
  NAND2_X1 U4695 ( .A1(n3785), .A2(n3784), .ZN(n3789) );
  XNOR2_X1 U4696 ( .A(n3297), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3790)
         );
  XNOR2_X1 U4697 ( .A(n3789), .B(n3790), .ZN(n4278) );
  INV_X1 U4698 ( .A(n4278), .ZN(n3786) );
  OAI22_X1 U4699 ( .A1(n3788), .A2(n3787), .B1(n4278), .B2(n3797), .ZN(n3796)
         );
  INV_X1 U4700 ( .A(n3789), .ZN(n3791) );
  NAND2_X1 U4701 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3800), .ZN(n3793) );
  NAND2_X1 U4702 ( .A1(n4282), .A2(n3794), .ZN(n3795) );
  NAND2_X1 U4703 ( .A1(n3796), .A2(n3795), .ZN(n3799) );
  AOI22_X1 U4704 ( .A1(n4282), .A2(n3801), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6599), .ZN(n3798) );
  NAND2_X1 U4705 ( .A1(n3799), .A2(n3798), .ZN(n3803) );
  AOI222_X1 U4706 ( .A1(n3800), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n3800), .B2(n5466), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n5466), 
        .ZN(n4279) );
  NAND2_X1 U4707 ( .A1(n4279), .A2(n3801), .ZN(n3802) );
  NAND2_X1 U4708 ( .A1(n4279), .A2(n3804), .ZN(n3805) );
  NAND2_X1 U4709 ( .A1(n3453), .A2(n3438), .ZN(n6479) );
  NAND2_X1 U4710 ( .A1(n6479), .A2(n3534), .ZN(n3811) );
  AND2_X1 U4711 ( .A1(n3808), .A2(n3809), .ZN(n3810) );
  NAND2_X1 U4712 ( .A1(n3811), .A2(n3810), .ZN(n4419) );
  NAND2_X1 U4713 ( .A1(n3812), .A2(n3981), .ZN(n3818) );
  NAND2_X1 U4714 ( .A1(n4656), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3846) );
  OAI21_X1 U4715 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6596), .A(n6251), 
        .ZN(n3814) );
  NOR2_X2 U4716 ( .A1(n3435), .A2(n6251), .ZN(n3827) );
  NAND2_X1 U4717 ( .A1(n4181), .A2(EAX_REG_4__SCAN_IN), .ZN(n3813) );
  OAI211_X1 U4718 ( .C1(n3846), .C2(n5466), .A(n3814), .B(n3813), .ZN(n3816)
         );
  AOI21_X1 U4719 ( .B1(n3819), .B2(n5617), .A(n3853), .ZN(n5844) );
  NAND2_X1 U4720 ( .A1(n5844), .A2(n4253), .ZN(n3815) );
  NAND2_X1 U4721 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  NAND2_X1 U4722 ( .A1(n3818), .A2(n3817), .ZN(n4623) );
  NAND2_X1 U4723 ( .A1(n4635), .A2(n3981), .ZN(n3825) );
  INV_X2 U4724 ( .A(n4232), .ZN(n4253) );
  OAI21_X1 U4725 ( .B1(n3820), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3819), 
        .ZN(n5858) );
  AOI22_X1 U4726 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4254), .B1(n4253), 
        .B2(n5858), .ZN(n3822) );
  NAND2_X1 U4727 ( .A1(n4181), .A2(EAX_REG_3__SCAN_IN), .ZN(n3821) );
  OAI211_X1 U4728 ( .C1(n3846), .C2(n3297), .A(n3822), .B(n3821), .ZN(n3823)
         );
  INV_X1 U4729 ( .A(n3823), .ZN(n3824) );
  NAND2_X1 U4730 ( .A1(n3825), .A2(n3824), .ZN(n4632) );
  NAND2_X1 U4731 ( .A1(n4634), .A2(n3981), .ZN(n3826) );
  INV_X1 U4732 ( .A(n4254), .ZN(n3985) );
  NAND2_X1 U4733 ( .A1(n3826), .A2(n3985), .ZN(n3848) );
  NAND2_X1 U4734 ( .A1(n3185), .A2(n3981), .ZN(n3832) );
  NAND2_X1 U4735 ( .A1(n4181), .A2(EAX_REG_1__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4736 ( .A1(n6251), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3828)
         );
  OAI211_X1 U4737 ( .C1(n3846), .C2(n3228), .A(n3829), .B(n3828), .ZN(n3830)
         );
  INV_X1 U4738 ( .A(n3830), .ZN(n3831) );
  AOI21_X1 U4739 ( .B1(n6282), .B2(n3833), .A(n6251), .ZN(n4557) );
  INV_X1 U4740 ( .A(n3981), .ZN(n3835) );
  OR2_X1 U4741 ( .A1(n6482), .A2(n3835), .ZN(n3840) );
  AOI22_X1 U4742 ( .A1(n4181), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6251), .ZN(n3838) );
  INV_X1 U4743 ( .A(n3846), .ZN(n3836) );
  NAND2_X1 U4744 ( .A1(n3836), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3837) );
  AND2_X1 U4745 ( .A1(n3838), .A2(n3837), .ZN(n3839) );
  NAND2_X1 U4746 ( .A1(n3840), .A2(n3839), .ZN(n4556) );
  NAND2_X1 U4747 ( .A1(n4557), .A2(n4556), .ZN(n4558) );
  INV_X1 U4748 ( .A(n4556), .ZN(n3841) );
  NAND2_X1 U4749 ( .A1(n3841), .A2(n4253), .ZN(n3842) );
  NAND2_X1 U4750 ( .A1(n4558), .A2(n3842), .ZN(n4507) );
  AND2_X2 U4751 ( .A1(n4508), .A2(n4507), .ZN(n3847) );
  OAI21_X1 U4752 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3843), .ZN(n5868) );
  AOI22_X1 U4753 ( .A1(n5868), .A2(n4253), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3845) );
  NAND2_X1 U4754 ( .A1(n4181), .A2(EAX_REG_2__SCAN_IN), .ZN(n3844) );
  OAI211_X1 U4755 ( .C1(n3846), .C2(n3166), .A(n3845), .B(n3844), .ZN(n4562)
         );
  NAND2_X1 U4756 ( .A1(n4563), .A2(n4562), .ZN(n3850) );
  NAND2_X1 U4757 ( .A1(n3847), .A2(n3848), .ZN(n3849) );
  AOI21_X1 U4758 ( .B1(n3852), .B2(n3981), .A(n3851), .ZN(n3855) );
  OAI21_X1 U4759 ( .B1(n3853), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3862), 
        .ZN(n5842) );
  AOI22_X1 U4760 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4254), .B1(n4253), 
        .B2(n5842), .ZN(n3854) );
  NAND2_X1 U4761 ( .A1(n3855), .A2(n3854), .ZN(n4696) );
  NAND2_X1 U4762 ( .A1(n4181), .A2(EAX_REG_6__SCAN_IN), .ZN(n3857) );
  OAI21_X1 U4763 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6596), .A(n6251), 
        .ZN(n3856) );
  XNOR2_X1 U4764 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3862), .ZN(n5831) );
  AOI22_X1 U4765 ( .A1(n3857), .A2(n3856), .B1(n4253), .B2(n5831), .ZN(n3858)
         );
  NAND2_X1 U4766 ( .A1(n3860), .A2(n3981), .ZN(n3868) );
  OAI21_X1 U4767 ( .B1(n3863), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3884), 
        .ZN(n5827) );
  AOI22_X1 U4768 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4254), .B1(n4253), 
        .B2(n5827), .ZN(n3864) );
  NAND2_X1 U4769 ( .A1(n4780), .A2(n4781), .ZN(n4772) );
  INV_X1 U4770 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4771 ( .A1(n3507), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4772 ( .A1(n3661), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4773 ( .A1(n3869), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4774 ( .A1(n3195), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4775 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3879)
         );
  AOI22_X1 U4776 ( .A1(n3154), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4777 ( .A1(n3198), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4778 ( .A1(n3190), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4779 ( .A1(n3203), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4780 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3878)
         );
  OAI21_X1 U4781 ( .B1(n3879), .B2(n3878), .A(n3981), .ZN(n3880) );
  OAI21_X1 U4782 ( .B1(n3881), .B2(n3985), .A(n3880), .ZN(n3883) );
  XNOR2_X1 U4783 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3884), .ZN(n5816) );
  NOR2_X1 U4784 ( .A1(n5816), .A2(n4232), .ZN(n3882) );
  AOI211_X1 U4785 ( .C1(n3827), .C2(EAX_REG_8__SCAN_IN), .A(n3883), .B(n3882), 
        .ZN(n4773) );
  XNOR2_X1 U4786 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3909), .ZN(n5808) );
  AOI22_X1 U4787 ( .A1(n4181), .A2(EAX_REG_9__SCAN_IN), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4788 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3190), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4789 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3199), .B1(n3189), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4790 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3869), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4791 ( .A1(n3194), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4792 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3895)
         );
  AOI22_X1 U4793 ( .A1(n3154), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4794 ( .A1(n3157), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4795 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3661), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4796 ( .A1(n3203), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4797 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  OAI21_X1 U4798 ( .B1(n3895), .B2(n3894), .A(n3981), .ZN(n3896) );
  OAI211_X1 U4799 ( .C1(n5808), .C2(n4232), .A(n3897), .B(n3896), .ZN(n4839)
         );
  INV_X1 U4800 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4873) );
  AOI22_X1 U4801 ( .A1(n3199), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4802 ( .A1(n3661), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4803 ( .A1(n3397), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4804 ( .A1(n3196), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4805 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3907)
         );
  AOI22_X1 U4806 ( .A1(n3154), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4807 ( .A1(n3157), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4808 ( .A1(n3203), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4809 ( .A1(n3190), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4810 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  OAI21_X1 U4811 ( .B1(n3907), .B2(n3906), .A(n3981), .ZN(n3908) );
  OAI21_X1 U4812 ( .B1(n4873), .B2(n3985), .A(n3908), .ZN(n3911) );
  XNOR2_X1 U4813 ( .A(n4873), .B(n3912), .ZN(n5565) );
  NOR2_X1 U4814 ( .A1(n5565), .A2(n4232), .ZN(n3910) );
  AOI211_X1 U4815 ( .C1(n3827), .C2(EAX_REG_10__SCAN_IN), .A(n3911), .B(n3910), 
        .ZN(n4843) );
  XNOR2_X1 U4816 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3926), .ZN(n5800)
         );
  AOI22_X1 U4817 ( .A1(n4181), .A2(EAX_REG_11__SCAN_IN), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4818 ( .A1(n3154), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4819 ( .A1(n3203), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4820 ( .A1(n3476), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4821 ( .A1(n3397), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4822 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3922)
         );
  AOI22_X1 U4823 ( .A1(n3507), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4824 ( .A1(n3157), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4825 ( .A1(n3190), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4826 ( .A1(n3869), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4827 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3921)
         );
  OAI21_X1 U4828 ( .B1(n3922), .B2(n3921), .A(n3981), .ZN(n3923) );
  OAI211_X1 U4829 ( .C1(n5800), .C2(n4232), .A(n3924), .B(n3923), .ZN(n4849)
         );
  XOR2_X1 U4830 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3940), .Z(n5550) );
  INV_X1 U4831 ( .A(n5550), .ZN(n4900) );
  AOI22_X1 U4832 ( .A1(n4181), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6251), .ZN(n3938) );
  AOI22_X1 U4833 ( .A1(n3154), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4834 ( .A1(n3199), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4835 ( .A1(n3203), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4836 ( .A1(n3186), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4837 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3936)
         );
  AOI22_X1 U4838 ( .A1(n3994), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4839 ( .A1(n3157), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4840 ( .A1(n3475), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4841 ( .A1(n3190), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4842 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3935)
         );
  OAI21_X1 U4843 ( .B1(n3936), .B2(n3935), .A(n3981), .ZN(n3937) );
  OAI21_X1 U4844 ( .B1(n3938), .B2(n4253), .A(n3937), .ZN(n3939) );
  AOI21_X1 U4845 ( .B1(n4900), .B2(n4253), .A(n3939), .ZN(n4854) );
  XOR2_X1 U4846 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3959), .Z(n5401) );
  NAND2_X1 U4847 ( .A1(n4181), .A2(EAX_REG_13__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4848 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n4254), .ZN(n3941)
         );
  NAND2_X1 U4849 ( .A1(n3942), .A2(n3941), .ZN(n3943) );
  AOI21_X1 U4850 ( .B1(n5401), .B2(n4253), .A(n3943), .ZN(n3956) );
  XNOR2_X1 U4851 ( .A(n3955), .B(n3956), .ZN(n4878) );
  AOI22_X1 U4852 ( .A1(n3154), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4853 ( .A1(n3199), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4854 ( .A1(n3994), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4855 ( .A1(n3157), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4856 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3953)
         );
  AOI22_X1 U4857 ( .A1(n3203), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4858 ( .A1(n3190), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4859 ( .A1(n3476), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4860 ( .A1(n3186), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3948) );
  NAND4_X1 U4861 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3952)
         );
  OR2_X1 U4862 ( .A1(n3953), .A2(n3952), .ZN(n3954) );
  AND2_X1 U4863 ( .A1(n3981), .A2(n3954), .ZN(n4879) );
  NAND2_X1 U4864 ( .A1(n4878), .A2(n4879), .ZN(n4880) );
  INV_X1 U4865 ( .A(n3956), .ZN(n3957) );
  NAND2_X1 U4866 ( .A1(n3955), .A2(n3957), .ZN(n3958) );
  NAND2_X1 U4867 ( .A1(n4880), .A2(n3958), .ZN(n4905) );
  XOR2_X1 U4868 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3986), .Z(n5527) );
  AOI22_X1 U4869 ( .A1(n4181), .A2(EAX_REG_14__SCAN_IN), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4870 ( .A1(n3197), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4871 ( .A1(n3869), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4872 ( .A1(n3476), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4873 ( .A1(n3196), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4874 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3970)
         );
  AOI22_X1 U4875 ( .A1(n3154), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3968) );
  INV_X1 U4876 ( .A(n3386), .ZN(n3964) );
  INV_X1 U4877 ( .A(n3964), .ZN(n3994) );
  AOI22_X1 U4878 ( .A1(n3203), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4879 ( .A1(n3190), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4880 ( .A1(n3199), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4881 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3969)
         );
  OAI21_X1 U4882 ( .B1(n3970), .B2(n3969), .A(n3981), .ZN(n3971) );
  OAI211_X1 U4883 ( .C1(n5527), .C2(n4232), .A(n3972), .B(n3971), .ZN(n4908)
         );
  NAND2_X1 U4884 ( .A1(n4905), .A2(n4908), .ZN(n4906) );
  AOI22_X1 U4885 ( .A1(n3869), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4886 ( .A1(n3507), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4887 ( .A1(n3397), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4888 ( .A1(n3196), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3973) );
  NAND4_X1 U4889 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3983)
         );
  AOI22_X1 U4890 ( .A1(n3157), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4891 ( .A1(n3203), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4892 ( .A1(n3154), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4893 ( .A1(n3190), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3977) );
  NAND4_X1 U4894 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3982)
         );
  OAI21_X1 U4895 ( .B1(n3983), .B2(n3982), .A(n3981), .ZN(n3984) );
  OAI21_X1 U4896 ( .B1(n5517), .B2(n3985), .A(n3984), .ZN(n3988) );
  XNOR2_X1 U4897 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3989), .ZN(n5515)
         );
  NOR2_X1 U4898 ( .A1(n5515), .A2(n4232), .ZN(n3987) );
  AOI211_X1 U4899 ( .C1(n3827), .C2(EAX_REG_15__SCAN_IN), .A(n3988), .B(n3987), 
        .ZN(n5131) );
  INV_X1 U4900 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5510) );
  XNOR2_X1 U4901 ( .A(n5510), .B(n4003), .ZN(n5508) );
  AOI22_X1 U4902 ( .A1(n4181), .A2(EAX_REG_16__SCAN_IN), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4903 ( .A1(n3197), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4904 ( .A1(n3869), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4905 ( .A1(n3203), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4906 ( .A1(n3397), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U4907 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n4000)
         );
  AOI22_X1 U4908 ( .A1(n3507), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4909 ( .A1(n3190), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4910 ( .A1(n3199), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4911 ( .A1(n3994), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4912 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  OAI21_X1 U4913 ( .B1(n4000), .B2(n3999), .A(n4249), .ZN(n4001) );
  OAI211_X1 U4914 ( .C1(n5508), .C2(n4232), .A(n4002), .B(n4001), .ZN(n4935)
         );
  OAI21_X1 U4915 ( .B1(n4004), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n4031), 
        .ZN(n5496) );
  AOI22_X1 U4916 ( .A1(n3827), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6251), .ZN(n4016) );
  AOI22_X1 U4917 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3167), .B1(n3154), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4918 ( .A1(n3203), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4919 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n3397), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4920 ( .A1(n3190), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4921 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4014)
         );
  AOI22_X1 U4922 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n3507), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4923 ( .A1(n3157), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4924 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3869), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4925 ( .A1(n3195), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4926 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  OAI21_X1 U4927 ( .B1(n4014), .B2(n4013), .A(n4249), .ZN(n4015) );
  NAND3_X1 U4928 ( .A1(n4232), .A2(n4016), .A3(n4015), .ZN(n4017) );
  OAI21_X1 U4929 ( .B1(n4232), .B2(n5496), .A(n4017), .ZN(n5389) );
  XNOR2_X1 U4930 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4031), .ZN(n5488)
         );
  AOI22_X1 U4931 ( .A1(n3827), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6251), .ZN(n4029) );
  AOI22_X1 U4932 ( .A1(n3661), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4933 ( .A1(n3203), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4934 ( .A1(n3190), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4935 ( .A1(n3476), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4936 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4027)
         );
  AOI22_X1 U4937 ( .A1(n3198), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3167), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4938 ( .A1(n3154), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4939 ( .A1(n3869), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4940 ( .A1(n3397), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U4941 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4026)
         );
  AOI221_X1 U4942 ( .B1(n4027), .B2(n4249), .C1(n4026), .C2(n4249), .A(n4253), 
        .ZN(n4028) );
  AOI22_X1 U4943 ( .A1(n4253), .A2(n5488), .B1(n4029), .B2(n4028), .ZN(n5085)
         );
  INV_X1 U4944 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4030) );
  OAI21_X1 U4945 ( .B1(n4032), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n4058), 
        .ZN(n5383) );
  AOI22_X1 U4946 ( .A1(n3827), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6251), .ZN(n4044) );
  AOI22_X1 U4947 ( .A1(n3167), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4948 ( .A1(n3203), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4949 ( .A1(n3661), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4950 ( .A1(n3617), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4033) );
  NAND4_X1 U4951 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(n4042)
         );
  AOI22_X1 U4952 ( .A1(n3154), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4953 ( .A1(n3198), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4954 ( .A1(n3192), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4955 ( .A1(n3476), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U4956 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4041)
         );
  OAI21_X1 U4957 ( .B1(n4042), .B2(n4041), .A(n4249), .ZN(n4043) );
  NAND3_X1 U4958 ( .A1(n4232), .A2(n4044), .A3(n4043), .ZN(n4045) );
  OAI21_X1 U4959 ( .B1(n4232), .B2(n5383), .A(n4045), .ZN(n5069) );
  XNOR2_X1 U4960 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4058), .ZN(n5374)
         );
  AOI22_X1 U4961 ( .A1(n3827), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6251), .ZN(n4057) );
  AOI22_X1 U4962 ( .A1(n3154), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4963 ( .A1(n3167), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4964 ( .A1(n3203), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4965 ( .A1(n3196), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U4966 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4055)
         );
  AOI22_X1 U4967 ( .A1(n3157), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4968 ( .A1(n3190), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4969 ( .A1(n3661), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4970 ( .A1(n3397), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4050) );
  NAND4_X1 U4971 ( .A1(n4053), .A2(n4052), .A3(n4051), .A4(n4050), .ZN(n4054)
         );
  AOI221_X1 U4972 ( .B1(n4055), .B2(n4249), .C1(n4054), .C2(n4249), .A(n4253), 
        .ZN(n4056) );
  AOI22_X1 U4973 ( .A1(n4253), .A2(n5374), .B1(n4057), .B2(n4056), .ZN(n5066)
         );
  INV_X1 U4974 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5303) );
  OAI21_X1 U4975 ( .B1(n4059), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4089), 
        .ZN(n5369) );
  AOI22_X1 U4976 ( .A1(n3827), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6251), .ZN(n4071) );
  AOI22_X1 U4977 ( .A1(n3199), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U4978 ( .A1(n3157), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4979 ( .A1(n3617), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4980 ( .A1(n3397), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4060) );
  NAND4_X1 U4981 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(n4069)
         );
  AOI22_X1 U4982 ( .A1(n3154), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4983 ( .A1(n3203), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4984 ( .A1(n3661), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4985 ( .A1(n3195), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4064) );
  NAND4_X1 U4986 ( .A1(n4067), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(n4068)
         );
  OAI21_X1 U4987 ( .B1(n4069), .B2(n4068), .A(n4249), .ZN(n4070) );
  NAND3_X1 U4988 ( .A1(n4232), .A2(n4071), .A3(n4070), .ZN(n4072) );
  OAI21_X1 U4989 ( .B1(n4232), .B2(n5369), .A(n4072), .ZN(n5007) );
  NAND2_X1 U4990 ( .A1(n4181), .A2(EAX_REG_22__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4991 ( .A1(n3507), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4992 ( .A1(n3197), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U4993 ( .A1(n3869), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U4994 ( .A1(n4187), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3617), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U4995 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4082)
         );
  AOI22_X1 U4996 ( .A1(n3380), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U4997 ( .A1(n3203), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U4998 ( .A1(n3476), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U4999 ( .A1(n3194), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5000 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4081)
         );
  AOI221_X1 U5001 ( .B1(n4082), .B2(n4249), .C1(n4081), .C2(n4249), .A(n4253), 
        .ZN(n4083) );
  INV_X1 U5002 ( .A(n4083), .ZN(n4084) );
  AOI21_X1 U5003 ( .B1(n6251), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4084), 
        .ZN(n4086) );
  XNOR2_X1 U5004 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .B(n4089), .ZN(n5362)
         );
  AOI21_X1 U5005 ( .B1(n4087), .B2(n4086), .A(n4085), .ZN(n5052) );
  INV_X1 U5006 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4088) );
  OR2_X1 U5007 ( .A1(n4090), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4091)
         );
  NAND2_X1 U5008 ( .A1(n4135), .A2(n4091), .ZN(n5281) );
  AOI22_X1 U5009 ( .A1(n3154), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5010 ( .A1(n3661), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5011 ( .A1(n3190), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5012 ( .A1(n3203), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4092) );
  NAND4_X1 U5013 ( .A1(n4095), .A2(n4094), .A3(n4093), .A4(n4092), .ZN(n4101)
         );
  AOI22_X1 U5014 ( .A1(n3199), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5015 ( .A1(n3197), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5016 ( .A1(n3869), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5017 ( .A1(n3397), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4096) );
  NAND4_X1 U5018 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(n4100)
         );
  NOR2_X1 U5019 ( .A1(n4101), .A2(n4100), .ZN(n4117) );
  AOI22_X1 U5020 ( .A1(n3154), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5021 ( .A1(n3661), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5022 ( .A1(n3203), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5023 ( .A1(n3190), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4102) );
  NAND4_X1 U5024 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4111)
         );
  AOI22_X1 U5025 ( .A1(n3198), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5026 ( .A1(n3195), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5027 ( .A1(n3869), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5028 ( .A1(n3475), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5029 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4110)
         );
  NOR2_X1 U5030 ( .A1(n4111), .A2(n4110), .ZN(n4118) );
  XNOR2_X1 U5031 ( .A(n4117), .B(n4118), .ZN(n4115) );
  INV_X1 U5032 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4112) );
  OAI21_X1 U5033 ( .B1(n4112), .B2(STATE2_REG_2__SCAN_IN), .A(n4232), .ZN(
        n4113) );
  AOI21_X1 U5034 ( .B1(n3827), .B2(EAX_REG_23__SCAN_IN), .A(n4113), .ZN(n4114)
         );
  OAI21_X1 U5035 ( .B1(n4230), .B2(n4115), .A(n4114), .ZN(n4116) );
  OAI21_X1 U5036 ( .B1(n5281), .B2(n4232), .A(n4116), .ZN(n5045) );
  XNOR2_X1 U5037 ( .A(n4135), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5274)
         );
  OR2_X1 U5038 ( .A1(n4118), .A2(n4117), .ZN(n4138) );
  AOI22_X1 U5039 ( .A1(n3198), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5040 ( .A1(n3203), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5041 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n3475), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5042 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3869), .B1(n3476), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U5043 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4128)
         );
  AOI22_X1 U5044 ( .A1(n3190), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5045 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3154), .B1(n3397), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5046 ( .A1(n3199), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5047 ( .A1(n4216), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5048 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4127)
         );
  NOR2_X1 U5049 ( .A1(n4128), .A2(n4127), .ZN(n4137) );
  AOI21_X1 U5050 ( .B1(n4137), .B2(n4138), .A(n4230), .ZN(n4129) );
  OAI21_X1 U5051 ( .B1(n4138), .B2(n4137), .A(n4129), .ZN(n4131) );
  AOI22_X1 U5052 ( .A1(n4181), .A2(EAX_REG_24__SCAN_IN), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4130) );
  AND2_X1 U5053 ( .A1(n4131), .A2(n4130), .ZN(n4132) );
  NAND2_X1 U5054 ( .A1(n4133), .A2(n4132), .ZN(n5037) );
  INV_X1 U5055 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4134) );
  OAI21_X1 U5056 ( .B1(n4136), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n4167), 
        .ZN(n5358) );
  AOI22_X1 U5057 ( .A1(n3507), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5058 ( .A1(n3869), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5059 ( .A1(n3195), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5060 ( .A1(n3157), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U5061 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4148)
         );
  AOI22_X1 U5062 ( .A1(n3154), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5063 ( .A1(n3203), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5064 ( .A1(n3476), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5065 ( .A1(n3617), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U5066 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4147)
         );
  NOR2_X1 U5067 ( .A1(n4148), .A2(n4147), .ZN(n4153) );
  XNOR2_X1 U5068 ( .A(n4152), .B(n4153), .ZN(n4150) );
  AOI22_X1 U5069 ( .A1(n3827), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6251), .ZN(n4149) );
  OAI21_X1 U5070 ( .B1(n4150), .B2(n4230), .A(n4149), .ZN(n4151) );
  AOI22_X1 U5071 ( .A1(n4253), .A2(n5358), .B1(n4151), .B2(n4232), .ZN(n5031)
         );
  XNOR2_X1 U5072 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4167), .ZN(n5349)
         );
  AOI22_X1 U5073 ( .A1(n3827), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6251), .ZN(n4166) );
  NOR2_X1 U5074 ( .A1(n4153), .A2(n4152), .ZN(n4180) );
  AOI22_X1 U5075 ( .A1(n3203), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3611), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5076 ( .A1(n3190), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5077 ( .A1(n3476), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5078 ( .A1(n3186), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4154) );
  NAND4_X1 U5079 ( .A1(n4157), .A2(n4156), .A3(n4155), .A4(n4154), .ZN(n4163)
         );
  AOI22_X1 U5080 ( .A1(n3154), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5081 ( .A1(n3167), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5082 ( .A1(n3661), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5083 ( .A1(n3198), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U5084 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4162)
         );
  OR2_X1 U5085 ( .A1(n4163), .A2(n4162), .ZN(n4179) );
  XOR2_X1 U5086 ( .A(n4180), .B(n4179), .Z(n4164) );
  AOI21_X1 U5087 ( .B1(n4164), .B2(n4249), .A(n4253), .ZN(n4165) );
  INV_X1 U5088 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4993) );
  OAI21_X1 U5089 ( .B1(n4168), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4214), 
        .ZN(n5348) );
  AOI22_X1 U5090 ( .A1(n3154), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5091 ( .A1(n3197), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5092 ( .A1(n3199), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5093 ( .A1(n3869), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4169) );
  NAND4_X1 U5094 ( .A1(n4172), .A2(n4171), .A3(n4170), .A4(n4169), .ZN(n4178)
         );
  AOI22_X1 U5095 ( .A1(n3190), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5096 ( .A1(n3611), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5097 ( .A1(n3203), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5098 ( .A1(n3397), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4173) );
  NAND4_X1 U5099 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4177)
         );
  NOR2_X1 U5100 ( .A1(n4178), .A2(n4177), .ZN(n4186) );
  NAND2_X1 U5101 ( .A1(n4180), .A2(n4179), .ZN(n4185) );
  XNOR2_X1 U5102 ( .A(n4186), .B(n4185), .ZN(n4183) );
  AOI22_X1 U5103 ( .A1(n4181), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6251), .ZN(n4182) );
  OAI21_X1 U5104 ( .B1(n4183), .B2(n4230), .A(n4182), .ZN(n4184) );
  AOI22_X1 U5105 ( .A1(n4253), .A2(n5348), .B1(n4184), .B2(n4232), .ZN(n5020)
         );
  XNOR2_X1 U5106 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n4214), .ZN(n4489)
         );
  AOI22_X1 U5107 ( .A1(n3827), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6251), .ZN(n4200) );
  NOR2_X1 U5108 ( .A1(n4186), .A2(n4185), .ZN(n4228) );
  AOI22_X1 U5109 ( .A1(n3203), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3611), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5110 ( .A1(n3617), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3192), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5111 ( .A1(n3476), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5112 ( .A1(n3186), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4188) );
  NAND4_X1 U5113 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4197)
         );
  AOI22_X1 U5114 ( .A1(n3154), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5115 ( .A1(n3167), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5116 ( .A1(n3661), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5117 ( .A1(n3157), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4192) );
  NAND4_X1 U5118 ( .A1(n4195), .A2(n4194), .A3(n4193), .A4(n4192), .ZN(n4196)
         );
  OR2_X1 U5119 ( .A1(n4197), .A2(n4196), .ZN(n4227) );
  XOR2_X1 U5120 ( .A(n4228), .B(n4227), .Z(n4198) );
  AOI21_X1 U5121 ( .B1(n4249), .B2(n4198), .A(n4253), .ZN(n4199) );
  NAND3_X1 U5122 ( .A1(n6599), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6530) );
  INV_X1 U5123 ( .A(n6530), .ZN(n4203) );
  AND2_X2 U5124 ( .A1(n4203), .A2(n6603), .ZN(n5876) );
  INV_X1 U5125 ( .A(n5876), .ZN(n6412) );
  OAI21_X1 U5126 ( .B1(n6602), .B2(n6603), .A(n6599), .ZN(n4204) );
  NAND2_X1 U5127 ( .A1(n6599), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5128 ( .A1(n6596), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4205) );
  AND2_X1 U5129 ( .A1(n4206), .A2(n4205), .ZN(n5873) );
  NAND2_X1 U5130 ( .A1(n6599), .A2(n6251), .ZN(n6529) );
  INV_X2 U5131 ( .A(n5937), .ZN(n5860) );
  AOI22_X1 U5132 ( .A1(n5860), .A2(REIP_REG_28__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4207) );
  INV_X1 U5133 ( .A(n4207), .ZN(n4208) );
  INV_X1 U5134 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4213) );
  NAND2_X1 U5135 ( .A1(n4215), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4258)
         );
  OAI21_X1 U5136 ( .B1(n4215), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4258), 
        .ZN(n5248) );
  AOI22_X1 U5137 ( .A1(n3203), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5138 ( .A1(n3154), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5139 ( .A1(n3869), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5140 ( .A1(n3186), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U5141 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4226)
         );
  AOI22_X1 U5142 ( .A1(n3197), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3661), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5143 ( .A1(n3199), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U5144 ( .A1(n3611), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5145 ( .A1(n3196), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4221) );
  NAND4_X1 U5146 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4225)
         );
  NOR2_X1 U5147 ( .A1(n4226), .A2(n4225), .ZN(n4235) );
  NAND2_X1 U5148 ( .A1(n4228), .A2(n4227), .ZN(n4234) );
  XNOR2_X1 U5149 ( .A(n4235), .B(n4234), .ZN(n4231) );
  AOI22_X1 U5150 ( .A1(n3827), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6251), .ZN(n4229) );
  OAI21_X1 U5151 ( .B1(n4231), .B2(n4230), .A(n4229), .ZN(n4233) );
  AOI22_X1 U5152 ( .A1(n4253), .A2(n5248), .B1(n4233), .B2(n4232), .ZN(n5016)
         );
  XNOR2_X1 U5153 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4258), .ZN(n5336)
         );
  AOI22_X1 U5154 ( .A1(n3827), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6251), .ZN(n4252) );
  NOR2_X1 U5155 ( .A1(n4235), .A2(n4234), .ZN(n4248) );
  AOI22_X1 U5156 ( .A1(n3154), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3507), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U5157 ( .A1(n3190), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5158 ( .A1(n3661), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5159 ( .A1(n3194), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4237) );
  NAND4_X1 U5160 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), .ZN(n4246)
         );
  AOI22_X1 U5161 ( .A1(n3167), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U5162 ( .A1(n3198), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3869), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5163 ( .A1(n3203), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3611), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5164 ( .A1(n3476), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4241) );
  NAND4_X1 U5165 ( .A1(n4244), .A2(n4243), .A3(n4242), .A4(n4241), .ZN(n4245)
         );
  NOR2_X1 U5166 ( .A1(n4246), .A2(n4245), .ZN(n4247) );
  XNOR2_X1 U5167 ( .A(n4248), .B(n4247), .ZN(n4250) );
  AOI21_X1 U5168 ( .B1(n4250), .B2(n4249), .A(n4253), .ZN(n4251) );
  AOI22_X1 U5169 ( .A1(n3827), .A2(EAX_REG_31__SCAN_IN), .B1(n4254), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4255) );
  INV_X1 U5170 ( .A(n4255), .ZN(n4256) );
  NAND2_X1 U5171 ( .A1(n5092), .A2(n5876), .ZN(n4269) );
  INV_X1 U5172 ( .A(n4258), .ZN(n4259) );
  NAND2_X1 U5173 ( .A1(n4259), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4260)
         );
  AOI22_X1 U5174 ( .A1(n5860), .A2(REIP_REG_31__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4261) );
  INV_X1 U5175 ( .A(n4261), .ZN(n4262) );
  NOR2_X1 U5176 ( .A1(n3288), .A2(n4262), .ZN(n4268) );
  NAND2_X1 U5177 ( .A1(n5797), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5145) );
  AND2_X1 U5178 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5139) );
  INV_X1 U5179 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4264) );
  INV_X1 U5180 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4408) );
  NOR2_X1 U5181 ( .A1(n4264), .A2(n4408), .ZN(n4433) );
  INV_X1 U5182 ( .A(n4433), .ZN(n4434) );
  NOR3_X1 U5183 ( .A1(n5146), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4417) );
  NAND3_X1 U5184 ( .A1(n4417), .A2(n4264), .A3(n4408), .ZN(n4265) );
  OAI22_X1 U5185 ( .A1(n5227), .A2(n4434), .B1(n4263), .B2(n4265), .ZN(n4266)
         );
  XNOR2_X1 U5186 ( .A(n4266), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4440)
         );
  NAND3_X1 U5187 ( .A1(n4269), .A2(n4268), .A3(n4267), .ZN(U2955) );
  INV_X1 U5188 ( .A(n5178), .ZN(n4311) );
  NAND2_X1 U5189 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U5190 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4868) );
  NOR2_X1 U5191 ( .A1(n4867), .A2(n4868), .ZN(n4310) );
  NAND2_X1 U5192 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4309) );
  NAND4_X1 U5193 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5918) );
  NOR2_X1 U5194 ( .A1(n4309), .A2(n5918), .ZN(n4862) );
  NAND2_X1 U5195 ( .A1(n4310), .A2(n4862), .ZN(n4925) );
  OR2_X1 U5196 ( .A1(n6479), .A2(n4660), .ZN(n4308) );
  INV_X1 U5197 ( .A(n4308), .ZN(n4270) );
  NAND2_X1 U5198 ( .A1(n4978), .A2(n4270), .ZN(n4285) );
  INV_X1 U5199 ( .A(n4419), .ZN(n4273) );
  NAND2_X1 U5200 ( .A1(n4271), .A2(n3445), .ZN(n4272) );
  MUX2_X1 U5201 ( .A(n4987), .B(n4272), .S(n4654), .Z(n4300) );
  NAND2_X1 U5202 ( .A1(n4273), .A2(n4300), .ZN(n4275) );
  INV_X1 U5203 ( .A(n4274), .ZN(n4980) );
  NAND2_X1 U5204 ( .A1(n4275), .A2(n4980), .ZN(n4519) );
  NAND3_X1 U5205 ( .A1(n4278), .A2(n4277), .A3(n4276), .ZN(n4281) );
  INV_X1 U5206 ( .A(n4279), .ZN(n4280) );
  OAI21_X1 U5207 ( .B1(n4282), .B2(n4281), .A(n4280), .ZN(n4981) );
  NOR2_X1 U5208 ( .A1(READY_N), .A2(n4981), .ZN(n4522) );
  OR2_X1 U5209 ( .A1(n4283), .A2(STATE_REG_0__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U5210 ( .A1(n3531), .A2(n6538), .ZN(n4984) );
  NAND3_X1 U5211 ( .A1(n4295), .A2(n4522), .A3(n4984), .ZN(n4284) );
  NAND3_X1 U5212 ( .A1(n4285), .A2(n4519), .A3(n4284), .ZN(n4286) );
  NAND2_X1 U5213 ( .A1(n4286), .A2(n6522), .ZN(n4293) );
  NAND2_X1 U5214 ( .A1(n4660), .A2(n6538), .ZN(n4448) );
  INV_X1 U5215 ( .A(READY_N), .ZN(n6896) );
  NAND2_X1 U5216 ( .A1(n4448), .A2(n6896), .ZN(n4289) );
  OAI211_X1 U5217 ( .C1(n4287), .C2(n4289), .A(n3445), .B(n4288), .ZN(n4290)
         );
  INV_X1 U5218 ( .A(n4290), .ZN(n4291) );
  NAND2_X1 U5219 ( .A1(n3534), .A2(n3531), .ZN(n4940) );
  OR2_X1 U5220 ( .A1(n4940), .A2(n4295), .ZN(n4518) );
  NAND2_X1 U5221 ( .A1(n4555), .A2(n4518), .ZN(n4298) );
  NOR2_X1 U5222 ( .A1(n4656), .A2(n3450), .ZN(n4296) );
  AOI21_X1 U5223 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n4299) );
  OAI211_X1 U5224 ( .C1(n3808), .C2(n4294), .A(n4300), .B(n4299), .ZN(n4301)
         );
  OR2_X1 U5225 ( .A1(n4302), .A2(n4301), .ZN(n4533) );
  NAND2_X1 U5226 ( .A1(n3184), .A2(n4303), .ZN(n4305) );
  NAND2_X1 U5227 ( .A1(n4594), .A2(n4305), .ZN(n4306) );
  NOR2_X1 U5228 ( .A1(n4533), .A2(n4306), .ZN(n4307) );
  NAND2_X1 U5229 ( .A1(n4274), .A2(n3531), .ZN(n6478) );
  NAND2_X1 U5230 ( .A1(n4919), .A2(n5955), .ZN(n4703) );
  INV_X1 U5231 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U5232 ( .A1(n5953), .A2(n5955), .ZN(n4546) );
  INV_X1 U5233 ( .A(n4579), .ZN(n4971) );
  NAND2_X1 U5234 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U5235 ( .A1(n5936), .A2(n5943), .ZN(n5928) );
  NAND3_X1 U5236 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n5928), .ZN(n5919) );
  NOR2_X1 U5237 ( .A1(n5919), .A2(n4309), .ZN(n4866) );
  NAND2_X1 U5238 ( .A1(n4866), .A2(n4310), .ZN(n4315) );
  NAND3_X1 U5239 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5208) );
  NOR2_X1 U5240 ( .A1(n3733), .A2(n5208), .ZN(n5199) );
  NAND3_X1 U5241 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5199), .ZN(n4314) );
  NAND3_X1 U5242 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5448), .ZN(n5186) );
  NOR2_X1 U5243 ( .A1(n4311), .A2(n5186), .ZN(n5432) );
  NAND2_X1 U5244 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4312) );
  NAND2_X1 U5245 ( .A1(n5432), .A2(n4312), .ZN(n5423) );
  NAND2_X1 U5246 ( .A1(n5944), .A2(n4919), .ZN(n4914) );
  INV_X1 U5247 ( .A(n4914), .ZN(n4313) );
  INV_X1 U5248 ( .A(n4314), .ZN(n4318) );
  NAND2_X1 U5249 ( .A1(n4423), .A2(n5937), .ZN(n5954) );
  OAI21_X1 U5250 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4919), .A(n5954), 
        .ZN(n4865) );
  INV_X1 U5251 ( .A(n4315), .ZN(n4316) );
  INV_X1 U5252 ( .A(n4703), .ZN(n4863) );
  INV_X1 U5253 ( .A(n4925), .ZN(n4920) );
  OAI22_X1 U5254 ( .A1(n4316), .A2(n5944), .B1(n4863), .B2(n4920), .ZN(n4317)
         );
  NOR2_X1 U5255 ( .A1(n4865), .A2(n4317), .ZN(n5885) );
  OAI21_X1 U5256 ( .B1(n5197), .B2(n4318), .A(n5885), .ZN(n5446) );
  NAND3_X1 U5257 ( .A1(n5178), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4319) );
  AND2_X1 U5258 ( .A1(n5910), .A2(n4319), .ZN(n4320) );
  NOR2_X1 U5259 ( .A1(n5446), .A2(n4320), .ZN(n5436) );
  AND2_X1 U5260 ( .A1(n5423), .A2(n5436), .ZN(n5169) );
  NAND2_X1 U5261 ( .A1(n5951), .A2(n5944), .ZN(n4322) );
  NAND2_X1 U5262 ( .A1(n4322), .A2(n4321), .ZN(n4323) );
  NAND2_X1 U5263 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U5264 ( .A1(n5910), .A2(n5150), .ZN(n4324) );
  NAND2_X1 U5265 ( .A1(n5420), .A2(n4324), .ZN(n5408) );
  INV_X1 U5266 ( .A(n5139), .ZN(n4325) );
  AND2_X1 U5267 ( .A1(n5910), .A2(n4325), .ZN(n4326) );
  NAND3_X1 U5268 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5165), .ZN(n5413) );
  NOR2_X1 U5269 ( .A1(n5150), .A2(n5413), .ZN(n5410) );
  NAND2_X1 U5270 ( .A1(n5410), .A2(n5139), .ZN(n5231) );
  OR2_X1 U5271 ( .A1(n4287), .A2(n4987), .ZN(n6505) );
  NAND2_X1 U5272 ( .A1(n4327), .A2(n4467), .ZN(n4328) );
  AND2_X1 U5273 ( .A1(n6505), .A2(n4328), .ZN(n4329) );
  NOR2_X2 U5274 ( .A1(n4423), .A2(n4329), .ZN(n5958) );
  INV_X1 U5275 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5884) );
  INV_X1 U5276 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U5277 ( .A1(n4468), .A2(n5558), .ZN(n4330) );
  OAI211_X1 U5278 ( .C1(n3152), .C2(n5884), .A(n4330), .B(n4403), .ZN(n4331)
         );
  OAI21_X1 U5279 ( .B1(n4402), .B2(EBX_REG_11__SCAN_IN), .A(n4331), .ZN(n4851)
         );
  INV_X1 U5280 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5281 ( .A1(n4403), .A2(EBX_REG_0__SCAN_IN), .ZN(n4335) );
  INV_X1 U5282 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U5283 ( .A1(n4294), .A2(n5657), .ZN(n4334) );
  NAND2_X1 U5284 ( .A1(n4335), .A2(n4334), .ZN(n4553) );
  NOR2_X1 U5285 ( .A1(n5642), .A2(n4511), .ZN(n4510) );
  INV_X1 U5286 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5287 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4511), .ZN(n4337)
         );
  OAI21_X1 U5288 ( .B1(n4336), .B2(EBX_REG_2__SCAN_IN), .A(n4337), .ZN(n4338)
         );
  INV_X1 U5289 ( .A(n4338), .ZN(n4339) );
  OAI211_X1 U5290 ( .C1(n4403), .C2(n4567), .A(n4339), .B(n4394), .ZN(n4566)
         );
  INV_X1 U5291 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5292 ( .A1(n4407), .A2(n4633), .B1(n4555), .B2(n5934), .ZN(n4340)
         );
  OAI21_X1 U5293 ( .B1(n4294), .B2(n4633), .A(n4340), .ZN(n4631) );
  INV_X1 U5294 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5623) );
  AOI21_X1 U5295 ( .B1(n4468), .B2(n5623), .A(n3152), .ZN(n4342) );
  OAI21_X1 U5296 ( .B1(n4341), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4342), 
        .ZN(n4343) );
  OAI21_X1 U5297 ( .B1(EBX_REG_4__SCAN_IN), .B2(n4336), .A(n4343), .ZN(n4627)
         );
  OR2_X1 U5298 ( .A1(n4402), .A2(EBX_REG_5__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U5299 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4344)
         );
  OAI211_X1 U5300 ( .C1(n4511), .C2(EBX_REG_5__SCAN_IN), .A(n4403), .B(n4344), 
        .ZN(n4345) );
  NAND2_X1 U5301 ( .A1(n4346), .A2(n4345), .ZN(n5606) );
  INV_X1 U5302 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5604) );
  AOI21_X1 U5303 ( .B1(n4468), .B2(n5604), .A(n3152), .ZN(n4347) );
  OAI21_X1 U5304 ( .B1(n4341), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4347), 
        .ZN(n4348) );
  OAI21_X1 U5305 ( .B1(EBX_REG_6__SCAN_IN), .B2(n4336), .A(n4348), .ZN(n4645)
         );
  INV_X1 U5306 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5307 ( .A1(n4407), .A2(n4785), .B1(n4555), .B2(n5906), .ZN(n4349)
         );
  OAI21_X1 U5308 ( .B1(n4294), .B2(n4785), .A(n4349), .ZN(n4783) );
  INV_X1 U5309 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5579) );
  AOI21_X1 U5310 ( .B1(n4468), .B2(n5579), .A(n3152), .ZN(n4350) );
  OAI21_X1 U5311 ( .B1(n4341), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4350), 
        .ZN(n4351) );
  OAI21_X1 U5312 ( .B1(EBX_REG_8__SCAN_IN), .B2(n4336), .A(n4351), .ZN(n4776)
         );
  INV_X1 U5313 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U5314 ( .A1(n4407), .A2(n4353), .B1(n4555), .B2(n5892), .ZN(n4352)
         );
  OAI21_X1 U5315 ( .B1(n4294), .B2(n4353), .A(n4352), .ZN(n4840) );
  INV_X1 U5316 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U5317 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4511), .ZN(n4354) );
  OAI21_X1 U5318 ( .B1(n4336), .B2(EBX_REG_10__SCAN_IN), .A(n4354), .ZN(n4355)
         );
  INV_X1 U5319 ( .A(n4355), .ZN(n4356) );
  OAI211_X1 U5320 ( .C1(n4403), .C2(n4846), .A(n4356), .B(n4394), .ZN(n4844)
         );
  INV_X1 U5321 ( .A(n4394), .ZN(n4357) );
  AOI21_X1 U5322 ( .B1(n4341), .B2(EBX_REG_12__SCAN_IN), .A(n4357), .ZN(n4359)
         );
  NAND2_X1 U5323 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4511), .ZN(n4358) );
  OAI211_X1 U5324 ( .C1(EBX_REG_12__SCAN_IN), .C2(n4336), .A(n4359), .B(n4358), 
        .ZN(n4855) );
  INV_X1 U5325 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5534) );
  AOI21_X1 U5326 ( .B1(n4468), .B2(n5534), .A(n4341), .ZN(n4360) );
  OAI21_X1 U5327 ( .B1(n3152), .B2(n4932), .A(n4360), .ZN(n4361) );
  OAI21_X1 U5328 ( .B1(EBX_REG_13__SCAN_IN), .B2(n4402), .A(n4361), .ZN(n4882)
         );
  NOR2_X2 U5329 ( .A1(n4883), .A2(n4882), .ZN(n4911) );
  INV_X1 U5330 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5331 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4511), .ZN(n4362) );
  OAI21_X1 U5332 ( .B1(n4336), .B2(EBX_REG_14__SCAN_IN), .A(n4362), .ZN(n4363)
         );
  INV_X1 U5333 ( .A(n4363), .ZN(n4364) );
  OAI211_X1 U5334 ( .C1(n4403), .C2(n4365), .A(n4364), .B(n4394), .ZN(n4912)
         );
  NAND2_X1 U5335 ( .A1(n4911), .A2(n4912), .ZN(n4910) );
  INV_X1 U5336 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U5337 ( .A1(n4468), .A2(n5670), .ZN(n4366) );
  OAI211_X1 U5338 ( .C1(n3152), .C2(n5201), .A(n4366), .B(n4403), .ZN(n4367)
         );
  OAI21_X1 U5339 ( .B1(n4402), .B2(EBX_REG_15__SCAN_IN), .A(n4367), .ZN(n5457)
         );
  NOR2_X2 U5340 ( .A1(n4910), .A2(n5457), .ZN(n5456) );
  INV_X1 U5341 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4371) );
  NAND2_X1 U5342 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4511), .ZN(n4368) );
  OAI21_X1 U5343 ( .B1(n4336), .B2(EBX_REG_16__SCAN_IN), .A(n4368), .ZN(n4369)
         );
  INV_X1 U5344 ( .A(n4369), .ZN(n4370) );
  OAI211_X1 U5345 ( .C1(n4403), .C2(n4371), .A(n4370), .B(n4394), .ZN(n4938)
         );
  OR2_X1 U5346 ( .A1(n4402), .A2(EBX_REG_17__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U5347 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4372) );
  OAI211_X1 U5348 ( .C1(n4511), .C2(EBX_REG_17__SCAN_IN), .A(n4403), .B(n4372), 
        .ZN(n4373) );
  NAND2_X1 U5349 ( .A1(n4374), .A2(n4373), .ZN(n5449) );
  INV_X1 U5350 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U5351 ( .A1(n4403), .A2(n5190), .ZN(n4376) );
  INV_X1 U5352 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U5353 ( .A1(n4468), .A2(n5314), .ZN(n4375) );
  NAND3_X1 U5354 ( .A1(n4376), .A2(n4375), .A3(n4294), .ZN(n4377) );
  OAI21_X1 U5355 ( .B1(EBX_REG_19__SCAN_IN), .B2(n4336), .A(n4377), .ZN(n5073)
         );
  INV_X1 U5356 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5183) );
  NOR2_X1 U5357 ( .A1(n4511), .A2(EBX_REG_20__SCAN_IN), .ZN(n4378) );
  AOI21_X1 U5358 ( .B1(n4555), .B2(n5183), .A(n4378), .ZN(n5062) );
  NAND2_X1 U5359 ( .A1(n4555), .A2(n5442), .ZN(n4379) );
  OR2_X1 U5360 ( .A1(n4511), .A2(EBX_REG_18__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U5361 ( .A1(n4379), .A2(n5077), .ZN(n5080) );
  NAND2_X1 U5362 ( .A1(n3152), .A2(EBX_REG_20__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5363 ( .A1(n5080), .A2(n4294), .ZN(n5072) );
  OAI211_X1 U5364 ( .C1(n5062), .C2(n5080), .A(n4380), .B(n5072), .ZN(n4381)
         );
  INV_X1 U5365 ( .A(n4381), .ZN(n4382) );
  NAND2_X1 U5366 ( .A1(n4555), .A2(n5435), .ZN(n4384) );
  NAND2_X1 U5367 ( .A1(n3152), .A2(EBX_REG_21__SCAN_IN), .ZN(n4383) );
  OAI211_X1 U5368 ( .C1(n4402), .C2(EBX_REG_21__SCAN_IN), .A(n4384), .B(n4383), 
        .ZN(n5003) );
  INV_X1 U5369 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U5370 ( .A1(n4511), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4385) );
  OAI211_X1 U5371 ( .C1(n4386), .C2(n4403), .A(n4394), .B(n4385), .ZN(n4388)
         );
  NOR2_X1 U5372 ( .A1(n4336), .A2(EBX_REG_22__SCAN_IN), .ZN(n4387) );
  NOR2_X1 U5373 ( .A1(n4388), .A2(n4387), .ZN(n5053) );
  OR2_X2 U5374 ( .A1(n5054), .A2(n5053), .ZN(n5056) );
  OR2_X1 U5375 ( .A1(n4402), .A2(EBX_REG_23__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U5376 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4389) );
  OAI211_X1 U5377 ( .C1(n4511), .C2(EBX_REG_23__SCAN_IN), .A(n4403), .B(n4389), 
        .ZN(n4390) );
  NAND2_X1 U5378 ( .A1(n4391), .A2(n4390), .ZN(n5048) );
  NOR2_X4 U5379 ( .A1(n5056), .A2(n5048), .ZN(n5050) );
  INV_X1 U5380 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U5381 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4511), .ZN(n4392) );
  OAI21_X1 U5382 ( .B1(n4336), .B2(EBX_REG_24__SCAN_IN), .A(n4392), .ZN(n4393)
         );
  INV_X1 U5383 ( .A(n4393), .ZN(n4395) );
  OAI211_X1 U5384 ( .C1(n4403), .C2(n5043), .A(n4395), .B(n4394), .ZN(n5040)
         );
  INV_X1 U5385 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5033) );
  INV_X1 U5386 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5419) );
  AOI22_X1 U5387 ( .A1(n4407), .A2(n5033), .B1(n4555), .B2(n5419), .ZN(n4396)
         );
  OAI21_X1 U5388 ( .B1(n5033), .B2(n4294), .A(n4396), .ZN(n5029) );
  INV_X1 U5389 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U5390 ( .A1(n4403), .A2(n5152), .ZN(n4398) );
  INV_X1 U5391 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U5392 ( .A1(n4468), .A2(n4994), .ZN(n4397) );
  NAND3_X1 U5393 ( .A1(n4398), .A2(n4397), .A3(n4294), .ZN(n4399) );
  OAI21_X1 U5394 ( .B1(EBX_REG_26__SCAN_IN), .B2(n4336), .A(n4399), .ZN(n4991)
         );
  NAND2_X1 U5395 ( .A1(n4555), .A2(n5409), .ZN(n4401) );
  NAND2_X1 U5396 ( .A1(n3152), .A2(EBX_REG_27__SCAN_IN), .ZN(n4400) );
  OAI211_X1 U5397 ( .C1(n4402), .C2(EBX_REG_27__SCAN_IN), .A(n4401), .B(n4400), 
        .ZN(n5022) );
  INV_X1 U5398 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U5399 ( .A1(n4403), .A2(n5143), .ZN(n4405) );
  NAND2_X1 U5400 ( .A1(n4468), .A2(n4499), .ZN(n4404) );
  NAND3_X1 U5401 ( .A1(n4405), .A2(n4404), .A3(n4294), .ZN(n4406) );
  OAI21_X1 U5402 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4336), .A(n4406), .ZN(n4495)
         );
  INV_X1 U5403 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5251) );
  AOI22_X1 U5404 ( .A1(n4407), .A2(n5251), .B1(n3152), .B2(EBX_REG_29__SCAN_IN), .ZN(n4410) );
  AND2_X1 U5405 ( .A1(n4555), .A2(n4408), .ZN(n4427) );
  INV_X1 U5406 ( .A(n4427), .ZN(n4409) );
  NAND2_X1 U5407 ( .A1(n4410), .A2(n4409), .ZN(n4411) );
  NOR2_X1 U5408 ( .A1(n4474), .A2(n4411), .ZN(n4429) );
  AND2_X1 U5409 ( .A1(n4474), .A2(n4411), .ZN(n4412) );
  NOR2_X1 U5410 ( .A1(n4429), .A2(n4412), .ZN(n5249) );
  INV_X1 U5411 ( .A(REIP_REG_29__SCAN_IN), .ZN(n4413) );
  NOR2_X1 U5412 ( .A1(n5937), .A2(n4413), .ZN(n5106) );
  AOI21_X1 U5413 ( .B1(n5958), .B2(n5249), .A(n5106), .ZN(n4414) );
  OAI21_X1 U5414 ( .B1(n5231), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4414), 
        .ZN(n4415) );
  INV_X1 U5415 ( .A(n4415), .ZN(n4424) );
  NAND2_X1 U5416 ( .A1(n4416), .A2(n4417), .ZN(n5226) );
  NAND2_X1 U5417 ( .A1(n5227), .A2(n5226), .ZN(n4418) );
  XNOR2_X1 U5418 ( .A(n4418), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5104)
         );
  OR2_X1 U5419 ( .A1(n4419), .A2(n4977), .ZN(n4577) );
  AND2_X1 U5420 ( .A1(n4577), .A2(n6495), .ZN(n4972) );
  NAND2_X1 U5421 ( .A1(n4327), .A2(n3408), .ZN(n4420) );
  AND3_X1 U5422 ( .A1(n4421), .A2(n4972), .A3(n4420), .ZN(n4422) );
  OAI211_X1 U5423 ( .C1(n4408), .C2(n3284), .A(n4424), .B(n3215), .ZN(U2989)
         );
  INV_X1 U5424 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4482) );
  OR2_X1 U5425 ( .A1(n4555), .A2(n4482), .ZN(n4426) );
  NAND2_X1 U5426 ( .A1(n4511), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4425) );
  NAND2_X1 U5427 ( .A1(n4426), .A2(n4425), .ZN(n4473) );
  INV_X1 U5428 ( .A(n4473), .ZN(n4475) );
  INV_X1 U5429 ( .A(n4555), .ZN(n4430) );
  OAI22_X1 U5430 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4511), .ZN(n4431) );
  XNOR2_X1 U5431 ( .A(n4432), .B(n4431), .ZN(n5011) );
  NAND2_X1 U5432 ( .A1(n5011), .A2(n5958), .ZN(n4439) );
  OAI21_X1 U5433 ( .B1(n5197), .B2(n4433), .A(n3284), .ZN(n5234) );
  NOR3_X1 U5434 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n5231), .A3(n4434), 
        .ZN(n4435) );
  AOI21_X1 U5435 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5860), .A(n4435), .ZN(n4436) );
  OAI211_X1 U5436 ( .C1(n5963), .C2(n4440), .A(n4439), .B(n4438), .ZN(U2987)
         );
  INV_X1 U5437 ( .A(n4441), .ZN(n4979) );
  NAND2_X1 U5438 ( .A1(n4274), .A2(n6522), .ZN(n4442) );
  NAND2_X1 U5439 ( .A1(n4954), .A2(n6251), .ZN(n6598) );
  NOR3_X1 U5440 ( .A1(n6599), .A2(n6373), .A3(n6598), .ZN(n6512) );
  NOR3_X1 U5441 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6529), .A3(n4954), .ZN(
        n6524) );
  NOR2_X1 U5442 ( .A1(n6512), .A2(n6524), .ZN(n4443) );
  NAND2_X1 U5443 ( .A1(n5937), .A2(n4443), .ZN(n4444) );
  OR2_X4 U5444 ( .A1(n6604), .A2(n4444), .ZN(n5651) );
  NAND2_X1 U5445 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5651), .ZN(n4487) );
  NAND2_X1 U5446 ( .A1(n5092), .A2(n5592), .ZN(n4464) );
  NOR2_X1 U5447 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4447) );
  INV_X1 U5448 ( .A(n4447), .ZN(n4491) );
  AND2_X2 U5449 ( .A1(n5651), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4942) );
  AND2_X1 U5450 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4942), .ZN(n4457) );
  NAND2_X1 U5451 ( .A1(n4491), .A2(n4457), .ZN(n4446) );
  INV_X1 U5452 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6576) );
  INV_X1 U5453 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6952) );
  INV_X1 U5454 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6565) );
  INV_X1 U5455 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6562) );
  INV_X1 U5456 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6558) );
  AND3_X1 U5457 ( .A1(n4448), .A2(n4447), .A3(n3445), .ZN(n4449) );
  NAND2_X2 U5458 ( .A1(n4942), .A2(n4449), .ZN(n5611) );
  INV_X1 U5459 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6557) );
  INV_X1 U5460 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6555) );
  INV_X1 U5461 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6588) );
  INV_X1 U5462 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6553) );
  INV_X1 U5463 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6551) );
  NOR3_X1 U5464 ( .A1(n6588), .A2(n6553), .A3(n6551), .ZN(n5621) );
  NAND2_X1 U5465 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5621), .ZN(n5610) );
  NOR2_X1 U5466 ( .A1(n6555), .A2(n5610), .ZN(n5593) );
  NAND2_X1 U5467 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5593), .ZN(n5586) );
  NOR2_X1 U5468 ( .A1(n6557), .A2(n5586), .ZN(n4451) );
  NAND4_X1 U5469 ( .A1(n5576), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n5552) );
  NAND3_X1 U5470 ( .A1(n5537), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n5507) );
  NOR2_X2 U5471 ( .A1(n6565), .A2(n5507), .ZN(n5505) );
  NAND3_X1 U5472 ( .A1(n5505), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n5495) );
  NAND3_X1 U5473 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4453) );
  NOR2_X2 U5474 ( .A1(n5495), .A2(n4453), .ZN(n5284) );
  NAND4_X1 U5475 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5284), .ZN(n5269) );
  NAND3_X1 U5476 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U5477 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5263), .ZN(n4486) );
  NOR2_X2 U5478 ( .A1(n6952), .A2(n4486), .ZN(n4456) );
  NAND2_X1 U5479 ( .A1(REIP_REG_29__SCAN_IN), .A2(n4456), .ZN(n4450) );
  OR3_X2 U5480 ( .A1(n6576), .A2(n4450), .A3(REIP_REG_31__SCAN_IN), .ZN(n4461)
         );
  NOR2_X1 U5481 ( .A1(REIP_REG_30__SCAN_IN), .A2(n4450), .ZN(n5242) );
  INV_X1 U5482 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6569) );
  INV_X1 U5483 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6906) );
  INV_X1 U5484 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6568) );
  NOR3_X1 U5485 ( .A1(n6569), .A2(n6906), .A3(n6568), .ZN(n4454) );
  NAND2_X1 U5486 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n4452) );
  AND3_X1 U5487 ( .A1(n5651), .A2(REIP_REG_8__SCAN_IN), .A3(n4451), .ZN(n5566)
         );
  NAND4_X1 U5488 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n5566), .ZN(n5538) );
  NOR3_X1 U5489 ( .A1(n6562), .A2(n4452), .A3(n5538), .ZN(n5506) );
  NAND4_X1 U5490 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5506), .ZN(n5305) );
  NAND2_X1 U5491 ( .A1(n5611), .A2(n5651), .ZN(n5653) );
  OAI21_X1 U5492 ( .B1(n5305), .B2(n4453), .A(n5653), .ZN(n5296) );
  OAI21_X1 U5493 ( .B1(n4454), .B2(n5611), .A(n5296), .ZN(n5286) );
  AOI21_X1 U5494 ( .B1(n5630), .B2(n4455), .A(n5286), .ZN(n4999) );
  NAND2_X1 U5495 ( .A1(REIP_REG_27__SCAN_IN), .A2(n4999), .ZN(n5262) );
  OAI21_X1 U5496 ( .B1(n6952), .B2(n5262), .A(n5653), .ZN(n5252) );
  NAND2_X1 U5497 ( .A1(n4456), .A2(n4413), .ZN(n5257) );
  NAND2_X1 U5498 ( .A1(n5252), .A2(n5257), .ZN(n5243) );
  OAI21_X1 U5499 ( .B1(n5242), .B2(n5243), .A(REIP_REG_31__SCAN_IN), .ZN(n4460) );
  NOR2_X1 U5500 ( .A1(n6538), .A2(n4491), .ZN(n6506) );
  OR2_X1 U5501 ( .A1(n4987), .A2(n6506), .ZN(n4493) );
  INV_X1 U5502 ( .A(n4493), .ZN(n4458) );
  AOI22_X1 U5503 ( .A1(n5638), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n4458), 
        .B2(n4457), .ZN(n4459) );
  NAND3_X1 U5504 ( .A1(n4461), .A2(n4460), .A3(n4459), .ZN(n4462) );
  AOI21_X1 U5505 ( .B1(n5011), .B2(n5652), .A(n4462), .ZN(n4463) );
  NAND2_X1 U5506 ( .A1(n4464), .A2(n4463), .ZN(U2796) );
  NAND2_X1 U5507 ( .A1(n4978), .A2(n4579), .ZN(n4515) );
  INV_X1 U5508 ( .A(n3435), .ZN(n5089) );
  NAND3_X1 U5509 ( .A1(n5089), .A2(n4467), .A3(n3409), .ZN(n4647) );
  INV_X1 U5510 ( .A(n4647), .ZN(n4469) );
  NAND3_X1 U5511 ( .A1(n4469), .A2(n3227), .A3(n4468), .ZN(n4470) );
  NAND2_X1 U5512 ( .A1(n4515), .A2(n4470), .ZN(n4471) );
  NAND2_X1 U5513 ( .A1(n5339), .A2(n4472), .ZN(n4485) );
  OAI21_X1 U5514 ( .B1(n3248), .B2(n4294), .A(n4475), .ZN(n4476) );
  INV_X1 U5515 ( .A(n4477), .ZN(n4478) );
  OAI22_X1 U5516 ( .A1(REIP_REG_28__SCAN_IN), .A2(n4486), .B1(n5097), .B2(
        n5599), .ZN(n4502) );
  AOI22_X1 U5517 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5638), .B1(n4489), 
        .B2(n5626), .ZN(n4490) );
  OAI21_X1 U5518 ( .B1(n6952), .B2(n5252), .A(n4490), .ZN(n4501) );
  INV_X1 U5519 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5012) );
  NAND3_X1 U5520 ( .A1(n3445), .A2(n5012), .A3(n4491), .ZN(n4492) );
  NAND2_X1 U5521 ( .A1(n4493), .A2(n4492), .ZN(n4494) );
  INV_X1 U5522 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4499) );
  INV_X1 U5523 ( .A(n4495), .ZN(n4498) );
  AOI21_X1 U5524 ( .B1(n4498), .B2(n4497), .A(n3248), .ZN(n5018) );
  INV_X1 U5525 ( .A(n5018), .ZN(n5136) );
  OAI22_X1 U5526 ( .A1(n5658), .A2(n4499), .B1(n5641), .B2(n5136), .ZN(n4500)
         );
  OR3_X1 U5527 ( .A1(n4502), .A2(n4501), .A3(n4500), .ZN(U2799) );
  INV_X1 U5528 ( .A(n6538), .ZN(n4986) );
  AND2_X1 U5529 ( .A1(n5704), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NAND2_X1 U5530 ( .A1(n6603), .A2(n4954), .ZN(n5470) );
  INV_X1 U5531 ( .A(n5470), .ZN(n5304) );
  NOR2_X1 U5532 ( .A1(n5304), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4506) );
  NAND3_X1 U5533 ( .A1(n6604), .A2(n4987), .A3(n4940), .ZN(n4505) );
  OAI21_X1 U5534 ( .B1(n6604), .B2(n4506), .A(n4505), .ZN(U3474) );
  NOR2_X1 U5535 ( .A1(n4508), .A2(n4507), .ZN(n4509) );
  OR2_X1 U5536 ( .A1(n3847), .A2(n4509), .ZN(n4756) );
  INV_X1 U5537 ( .A(n4756), .ZN(n5647) );
  AOI21_X1 U5538 ( .B1(n5642), .B2(n4511), .A(n4510), .ZN(n4548) );
  OAI22_X1 U5539 ( .A1(n4548), .A2(n5088), .B1(n5674), .B2(n4512), .ZN(n4513)
         );
  AOI21_X1 U5540 ( .B1(n5647), .B2(n4472), .A(n4513), .ZN(n4514) );
  INV_X1 U5541 ( .A(n4514), .ZN(U2858) );
  NOR2_X1 U5542 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6373), .ZN(n6585) );
  INV_X1 U5543 ( .A(n4515), .ZN(n4526) );
  AOI21_X1 U5544 ( .B1(n6478), .B2(n4287), .A(n6538), .ZN(n4517) );
  OAI21_X1 U5545 ( .B1(n4517), .B2(n4516), .A(n6896), .ZN(n4520) );
  OAI211_X1 U5546 ( .C1(n4978), .C2(n4520), .A(n4519), .B(n4518), .ZN(n4525)
         );
  OR2_X1 U5547 ( .A1(n4978), .A2(n4577), .ZN(n4524) );
  NAND2_X1 U5548 ( .A1(n4521), .A2(n4522), .ZN(n4523) );
  NAND2_X1 U5549 ( .A1(n4524), .A2(n4523), .ZN(n4650) );
  NAND2_X1 U5550 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4613), .ZN(n6528) );
  INV_X1 U5551 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6843) );
  OAI22_X1 U5552 ( .A1(n6485), .A2(n6519), .B1(n6528), .B2(n6843), .ZN(n5463)
         );
  INV_X1 U5553 ( .A(n5223), .ZN(n5467) );
  INV_X1 U5554 ( .A(n4521), .ZN(n4531) );
  AND3_X1 U5555 ( .A1(n4287), .A2(n4648), .A3(n3168), .ZN(n4530) );
  NAND2_X1 U5556 ( .A1(n4531), .A2(n4530), .ZN(n4532) );
  NOR2_X1 U5557 ( .A1(n4533), .A2(n4532), .ZN(n6481) );
  INV_X1 U5558 ( .A(n6481), .ZN(n4953) );
  INV_X1 U5559 ( .A(n4534), .ZN(n4536) );
  INV_X1 U5560 ( .A(n4535), .ZN(n4964) );
  NAND2_X1 U5561 ( .A1(n4536), .A2(n4964), .ZN(n4540) );
  OAI22_X1 U5562 ( .A1(n6478), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n4540), .B2(n6479), .ZN(n4537) );
  AOI21_X1 U5563 ( .B1(n4528), .B2(n4953), .A(n4537), .ZN(n6484) );
  NOR2_X1 U5564 ( .A1(n6484), .A2(n6521), .ZN(n4542) );
  NOR2_X1 U5565 ( .A1(n4954), .A2(n5953), .ZN(n4962) );
  INV_X1 U5566 ( .A(n4962), .ZN(n4957) );
  INV_X1 U5567 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5568 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4539), .B2(n4549), .ZN(n4963)
         );
  OAI22_X1 U5569 ( .A1(n6510), .A2(n4540), .B1(n4957), .B2(n4963), .ZN(n4541)
         );
  OAI21_X1 U5570 ( .B1(n4542), .B2(n4541), .A(n5467), .ZN(n4543) );
  OAI21_X1 U5571 ( .B1(n5467), .B2(n3228), .A(n4543), .ZN(U3460) );
  XOR2_X1 U5572 ( .A(n4545), .B(n4544), .Z(n4754) );
  NAND3_X1 U5573 ( .A1(n5910), .A2(n4546), .A3(n4549), .ZN(n4547) );
  NAND2_X1 U5574 ( .A1(n5860), .A2(REIP_REG_1__SCAN_IN), .ZN(n4755) );
  OAI211_X1 U5575 ( .C1(n4548), .C2(n5938), .A(n4547), .B(n4755), .ZN(n4551)
         );
  NAND2_X1 U5576 ( .A1(n5953), .A2(n4914), .ZN(n5960) );
  AOI21_X1 U5577 ( .B1(n5954), .B2(n5960), .A(n4549), .ZN(n4550) );
  AOI211_X1 U5578 ( .C1(n5946), .C2(n4754), .A(n4551), .B(n4550), .ZN(n4552)
         );
  INV_X1 U5579 ( .A(n4552), .ZN(U3017) );
  INV_X1 U5580 ( .A(n4553), .ZN(n4554) );
  AOI21_X1 U5581 ( .B1(n4555), .B2(n5953), .A(n4554), .ZN(n5959) );
  INV_X1 U5582 ( .A(n5959), .ZN(n4560) );
  OR2_X1 U5583 ( .A1(n4557), .A2(n4556), .ZN(n4559) );
  AND2_X1 U5584 ( .A1(n4559), .A2(n4558), .ZN(n5875) );
  INV_X1 U5585 ( .A(n5875), .ZN(n5663) );
  OAI222_X1 U5586 ( .A1(n4560), .A2(n5088), .B1(n5674), .B2(n5657), .C1(n5663), 
        .C2(n5086), .ZN(U2859) );
  NOR2_X1 U5587 ( .A1(n4563), .A2(n4562), .ZN(n4564) );
  NOR2_X1 U5588 ( .A1(n4561), .A2(n4564), .ZN(n5865) );
  INV_X1 U5589 ( .A(n5865), .ZN(n4658) );
  XNOR2_X1 U5590 ( .A(n4565), .B(n4566), .ZN(n5939) );
  OAI222_X1 U5591 ( .A1(n5086), .A2(n4658), .B1(n4567), .B2(n5674), .C1(n5088), 
        .C2(n5939), .ZN(U2857) );
  INV_X1 U5592 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U5593 ( .A1(n5692), .A2(n3445), .ZN(n4836) );
  AOI22_X1 U5594 ( .A1(n4833), .A2(UWORD_REG_14__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4568) );
  OAI21_X1 U5595 ( .B1(n5744), .B2(n4836), .A(n4568), .ZN(U2893) );
  INV_X1 U5596 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5731) );
  AOI22_X1 U5597 ( .A1(n4833), .A2(UWORD_REG_8__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5598 ( .B1(n5731), .B2(n4836), .A(n4569), .ZN(U2899) );
  INV_X1 U5599 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5733) );
  AOI22_X1 U5600 ( .A1(n4833), .A2(UWORD_REG_9__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4570) );
  OAI21_X1 U5601 ( .B1(n5733), .B2(n4836), .A(n4570), .ZN(U2898) );
  INV_X1 U5602 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5735) );
  AOI22_X1 U5603 ( .A1(n4833), .A2(UWORD_REG_10__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5604 ( .B1(n5735), .B2(n4836), .A(n4571), .ZN(U2897) );
  INV_X1 U5605 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5737) );
  AOI22_X1 U5606 ( .A1(n4833), .A2(UWORD_REG_11__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4572) );
  OAI21_X1 U5607 ( .B1(n5737), .B2(n4836), .A(n4572), .ZN(U2896) );
  INV_X1 U5608 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5739) );
  AOI22_X1 U5609 ( .A1(n4833), .A2(UWORD_REG_12__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4573) );
  OAI21_X1 U5610 ( .B1(n5739), .B2(n4836), .A(n4573), .ZN(U2895) );
  INV_X1 U5611 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5742) );
  AOI22_X1 U5612 ( .A1(n4833), .A2(UWORD_REG_13__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U5613 ( .B1(n5742), .B2(n4836), .A(n4574), .ZN(U2894) );
  MUX2_X1 U5614 ( .A(n4599), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4575) );
  NOR2_X1 U5615 ( .A1(n4575), .A2(n5466), .ZN(n4609) );
  INV_X1 U5616 ( .A(n4577), .ZN(n4578) );
  OR2_X1 U5617 ( .A1(n4579), .A2(n4578), .ZN(n4597) );
  XNOR2_X1 U5618 ( .A(n4535), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4582)
         );
  XNOR2_X1 U5619 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4580) );
  OAI22_X1 U5620 ( .A1(n6478), .A2(n4580), .B1(n4594), .B2(n4582), .ZN(n4581)
         );
  AOI21_X1 U5621 ( .B1(n4597), .B2(n4582), .A(n4581), .ZN(n4583) );
  OAI21_X1 U5622 ( .B1(n4576), .B2(n6481), .A(n4583), .ZN(n4967) );
  NAND2_X1 U5623 ( .A1(n4967), .A2(n4599), .ZN(n4585) );
  NAND2_X1 U5624 ( .A1(n6485), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4584) );
  INV_X1 U5625 ( .A(n6362), .ZN(n6029) );
  INV_X1 U5626 ( .A(n4587), .ZN(n4590) );
  INV_X1 U5627 ( .A(n4588), .ZN(n4589) );
  OAI211_X1 U5628 ( .C1(n4535), .C2(n4590), .A(n3206), .B(n4589), .ZN(n4596)
         );
  AOI21_X1 U5629 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3297), .ZN(n4591) );
  NOR3_X1 U5630 ( .A1(n3157), .A2(n3611), .A3(n4591), .ZN(n5221) );
  MUX2_X1 U5631 ( .A(n5224), .B(n4588), .S(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .Z(n4592) );
  INV_X1 U5632 ( .A(n6478), .ZN(n4952) );
  OAI21_X1 U5633 ( .B1(n4587), .B2(n4592), .A(n4952), .ZN(n4593) );
  OAI21_X1 U5634 ( .B1(n5221), .B2(n4594), .A(n4593), .ZN(n4595) );
  AOI21_X1 U5635 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(n4598) );
  OAI21_X1 U5636 ( .B1(n6029), .B2(n6481), .A(n4598), .ZN(n5220) );
  MUX2_X1 U5637 ( .A(n5224), .B(n5220), .S(n4599), .Z(n6492) );
  NAND2_X1 U5638 ( .A1(n4954), .A2(n6492), .ZN(n4607) );
  INV_X1 U5639 ( .A(n4601), .ZN(n4712) );
  NOR2_X1 U5640 ( .A1(n4600), .A2(n4712), .ZN(n4602) );
  XNOR2_X1 U5641 ( .A(n4602), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5616)
         );
  NAND2_X1 U5642 ( .A1(n4521), .A2(n4954), .ZN(n4603) );
  OR2_X1 U5643 ( .A1(n5616), .A2(n4603), .ZN(n5462) );
  AND2_X1 U5644 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6843), .ZN(n4605) );
  NAND2_X1 U5645 ( .A1(n4604), .A2(n4605), .ZN(n4606) );
  OAI211_X1 U5646 ( .C1(n6489), .C2(n4607), .A(n5462), .B(n4606), .ZN(n4608)
         );
  OR2_X1 U5647 ( .A1(n4609), .A2(n4608), .ZN(n6500) );
  INV_X1 U5648 ( .A(n4609), .ZN(n4610) );
  NAND2_X1 U5649 ( .A1(n4534), .A2(n4610), .ZN(n4611) );
  NAND2_X1 U5650 ( .A1(n6500), .A2(n4611), .ZN(n6513) );
  NOR2_X1 U5651 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4954), .ZN(n5217) );
  INV_X1 U5652 ( .A(n5217), .ZN(n4620) );
  AOI222_X1 U5653 ( .A1(n6513), .A2(n4613), .B1(n3159), .B2(n4620), .C1(n6405), 
        .C2(n6329), .ZN(n4617) );
  NAND2_X1 U5654 ( .A1(n6513), .A2(n6843), .ZN(n4612) );
  INV_X1 U5655 ( .A(n6528), .ZN(n6584) );
  NAND2_X1 U5656 ( .A1(n4612), .A2(n6584), .ZN(n4615) );
  INV_X1 U5657 ( .A(n6598), .ZN(n4614) );
  NAND2_X1 U5658 ( .A1(n5964), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4616) );
  OAI21_X1 U5659 ( .B1(n4617), .B2(n5964), .A(n4616), .ZN(U3465) );
  INV_X1 U5660 ( .A(n6405), .ZN(n6417) );
  AOI211_X1 U5661 ( .C1(n6147), .C2(n6596), .A(n6417), .B(n6061), .ZN(n4619)
         );
  AOI21_X1 U5662 ( .B1(n4528), .B2(n4620), .A(n4619), .ZN(n4622) );
  NAND2_X1 U5663 ( .A1(n5964), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4621) );
  OAI21_X1 U5664 ( .B1(n4622), .B2(n5964), .A(n4621), .ZN(U3464) );
  AND2_X1 U5665 ( .A1(n4561), .A2(n4632), .ZN(n4626) );
  AND2_X1 U5666 ( .A1(n4624), .A2(n4561), .ZN(n4695) );
  INV_X1 U5667 ( .A(n4695), .ZN(n4625) );
  OAI21_X1 U5668 ( .B1(n4626), .B2(n4623), .A(n4625), .ZN(n5849) );
  OAI21_X1 U5669 ( .B1(n4627), .B2(n4630), .A(n5605), .ZN(n5622) );
  INV_X1 U5670 ( .A(n5622), .ZN(n4628) );
  AOI22_X1 U5671 ( .A1(n5671), .A2(n4628), .B1(n5074), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4629) );
  OAI21_X1 U5672 ( .B1(n5849), .B2(n5086), .A(n4629), .ZN(U2855) );
  INV_X1 U5673 ( .A(n5927), .ZN(n4944) );
  XNOR2_X1 U5674 ( .A(n4561), .B(n4632), .ZN(n5854) );
  OAI222_X1 U5675 ( .A1(n4944), .A2(n5088), .B1(n4633), .B2(n5674), .C1(n5854), 
        .C2(n5086), .ZN(U2856) );
  INV_X1 U5676 ( .A(n5964), .ZN(n4641) );
  NAND2_X1 U5677 ( .A1(n4634), .A2(n3657), .ZN(n6411) );
  NAND2_X1 U5678 ( .A1(n6330), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6324) );
  INV_X1 U5679 ( .A(n4634), .ZN(n6062) );
  INV_X1 U5680 ( .A(n6244), .ZN(n6246) );
  NAND2_X1 U5681 ( .A1(n6324), .A2(n6246), .ZN(n6064) );
  INV_X1 U5682 ( .A(n6064), .ZN(n4637) );
  NAND2_X1 U5683 ( .A1(n4634), .A2(n4636), .ZN(n6113) );
  INV_X1 U5684 ( .A(n6061), .ZN(n6245) );
  OR2_X1 U5685 ( .A1(n6113), .A2(n6245), .ZN(n6115) );
  AOI21_X1 U5686 ( .B1(n4637), .B2(n6115), .A(n6417), .ZN(n4639) );
  AND2_X1 U5687 ( .A1(n6603), .A2(n6596), .ZN(n6414) );
  INV_X1 U5688 ( .A(n6414), .ZN(n6034) );
  OAI22_X1 U5689 ( .A1(n6033), .A2(n6034), .B1(n6029), .B2(n5217), .ZN(n4638)
         );
  OAI21_X1 U5690 ( .B1(n4639), .B2(n4638), .A(n4641), .ZN(n4640) );
  OAI21_X1 U5691 ( .B1(n4641), .B2(n6493), .A(n4640), .ZN(U3462) );
  XNOR2_X1 U5692 ( .A(n4642), .B(n4643), .ZN(n5834) );
  XOR2_X1 U5693 ( .A(n4644), .B(n4645), .Z(n5911) );
  AOI22_X1 U5694 ( .A1(n5671), .A2(n5911), .B1(n5074), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4646) );
  OAI21_X1 U5695 ( .B1(n5834), .B2(n5086), .A(n4646), .ZN(U2853) );
  NOR2_X1 U5696 ( .A1(n4648), .A2(n4647), .ZN(n4649) );
  NAND2_X1 U5697 ( .A1(n4654), .A2(n3435), .ZN(n4655) );
  AND2_X1 U5698 ( .A1(n5090), .A2(n4656), .ZN(n5682) );
  AND2_X1 U5699 ( .A1(n3440), .A2(n3435), .ZN(n4657) );
  NOR2_X2 U5700 ( .A1(n5682), .A2(n5684), .ZN(n5691) );
  INV_X1 U5701 ( .A(DATAI_4_), .ZN(n6877) );
  INV_X1 U5702 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5759) );
  OAI222_X1 U5703 ( .A1(n5849), .A2(n5677), .B1(n5691), .B2(n6877), .C1(n5090), 
        .C2(n5759), .ZN(U2887) );
  INV_X1 U5704 ( .A(DATAI_3_), .ZN(n4672) );
  INV_X1 U5705 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5756) );
  OAI222_X1 U5706 ( .A1(n5854), .A2(n5677), .B1(n5691), .B2(n4672), .C1(n5090), 
        .C2(n5756), .ZN(U2888) );
  INV_X1 U5707 ( .A(DATAI_1_), .ZN(n6981) );
  INV_X1 U5708 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5750) );
  OAI222_X1 U5709 ( .A1(n4756), .A2(n5677), .B1(n5691), .B2(n6981), .C1(n5090), 
        .C2(n5750), .ZN(U2890) );
  INV_X1 U5710 ( .A(DATAI_2_), .ZN(n4676) );
  INV_X1 U5711 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5753) );
  OAI222_X1 U5712 ( .A1(n4658), .A2(n5677), .B1(n5691), .B2(n4676), .C1(n5090), 
        .C2(n5753), .ZN(U2889) );
  INV_X1 U5713 ( .A(DATAI_6_), .ZN(n6909) );
  INV_X1 U5714 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5765) );
  OAI222_X1 U5715 ( .A1(n5834), .A2(n5677), .B1(n5691), .B2(n6909), .C1(n5090), 
        .C2(n5765), .ZN(U2885) );
  INV_X1 U5716 ( .A(DATAI_0_), .ZN(n4762) );
  INV_X1 U5717 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5747) );
  OAI222_X1 U5718 ( .A1(n5663), .A2(n5677), .B1(n5691), .B2(n4762), .C1(n5090), 
        .C2(n5747), .ZN(U2891) );
  NOR2_X2 U5719 ( .A1(n4763), .A2(n4660), .ZN(n6427) );
  INV_X1 U5720 ( .A(n6427), .ZN(n4730) );
  NOR2_X1 U5721 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6118), .ZN(n6107)
         );
  INV_X1 U5722 ( .A(n6107), .ZN(n4694) );
  NOR2_X1 U5723 ( .A1(n6113), .A2(n3185), .ZN(n4718) );
  INV_X1 U5724 ( .A(n6113), .ZN(n4710) );
  OAI21_X1 U5725 ( .B1(n6108), .B2(n6138), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4662) );
  INV_X1 U5726 ( .A(n4576), .ZN(n4661) );
  NAND2_X1 U5727 ( .A1(n4661), .A2(n4528), .ZN(n6402) );
  OR2_X1 U5728 ( .A1(n6362), .A2(n6402), .ZN(n4665) );
  NAND3_X1 U5729 ( .A1(n4662), .A2(n6603), .A3(n4665), .ZN(n4664) );
  AND2_X1 U5730 ( .A1(n4666), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6368) );
  OAI21_X1 U5731 ( .B1(n6364), .B2(n6251), .A(n6151), .ZN(n6369) );
  AOI211_X1 U5732 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4694), .A(n6368), .B(
        n6369), .ZN(n4663) );
  NAND3_X1 U5733 ( .A1(n6493), .A2(n4664), .A3(n4663), .ZN(n6109) );
  NAND2_X1 U5734 ( .A1(n6109), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4670) );
  AND2_X1 U5735 ( .A1(n5876), .A2(DATAI_25_), .ZN(n6428) );
  AND2_X1 U5736 ( .A1(n5876), .A2(DATAI_17_), .ZN(n6335) );
  INV_X1 U5737 ( .A(n6335), .ZN(n6431) );
  INV_X1 U5738 ( .A(n4665), .ZN(n6114) );
  INV_X1 U5739 ( .A(n6364), .ZN(n4790) );
  OR2_X1 U5740 ( .A1(n4666), .A2(n6251), .ZN(n4794) );
  NOR3_X1 U5741 ( .A1(n4790), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4794), 
        .ZN(n4667) );
  AOI21_X1 U5742 ( .B1(n6114), .B2(n6603), .A(n4667), .ZN(n6105) );
  NOR2_X2 U5743 ( .A1(n6981), .A2(n4761), .ZN(n6426) );
  INV_X1 U5744 ( .A(n6426), .ZN(n4818) );
  OAI22_X1 U5745 ( .A1(n6135), .A2(n6431), .B1(n6105), .B2(n4818), .ZN(n4668)
         );
  AOI21_X1 U5746 ( .B1(n6428), .B2(n6108), .A(n4668), .ZN(n4669) );
  OAI211_X1 U5747 ( .C1(n4730), .C2(n4694), .A(n4670), .B(n4669), .ZN(U3069)
         );
  NOR2_X2 U5748 ( .A1(n4763), .A2(n4671), .ZN(n6439) );
  INV_X1 U5749 ( .A(n6439), .ZN(n4720) );
  NAND2_X1 U5750 ( .A1(n6109), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4675) );
  AND2_X1 U5751 ( .A1(n5876), .A2(DATAI_27_), .ZN(n6440) );
  AND2_X1 U5752 ( .A1(n5876), .A2(DATAI_19_), .ZN(n6224) );
  NOR2_X2 U5753 ( .A1(n4672), .A2(n4761), .ZN(n6438) );
  INV_X1 U5754 ( .A(n6438), .ZN(n4797) );
  OAI22_X1 U5755 ( .A1(n6135), .A2(n6443), .B1(n6105), .B2(n4797), .ZN(n4673)
         );
  AOI21_X1 U5756 ( .B1(n6440), .B2(n6108), .A(n4673), .ZN(n4674) );
  OAI211_X1 U5757 ( .C1(n4694), .C2(n4720), .A(n4675), .B(n4674), .ZN(U3071)
         );
  NOR2_X2 U5758 ( .A1(n4763), .A2(n3450), .ZN(n6433) );
  INV_X1 U5759 ( .A(n6433), .ZN(n4725) );
  NAND2_X1 U5760 ( .A1(n6109), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4679) );
  AND2_X1 U5761 ( .A1(n5876), .A2(DATAI_26_), .ZN(n6434) );
  AND2_X1 U5762 ( .A1(n5876), .A2(DATAI_18_), .ZN(n6259) );
  INV_X1 U5763 ( .A(n6259), .ZN(n6437) );
  NOR2_X2 U5764 ( .A1(n4676), .A2(n4761), .ZN(n6432) );
  INV_X1 U5765 ( .A(n6432), .ZN(n4806) );
  OAI22_X1 U5766 ( .A1(n6135), .A2(n6437), .B1(n6105), .B2(n4806), .ZN(n4677)
         );
  AOI21_X1 U5767 ( .B1(n6434), .B2(n6108), .A(n4677), .ZN(n4678) );
  OAI211_X1 U5768 ( .C1(n4694), .C2(n4725), .A(n4679), .B(n4678), .ZN(U3070)
         );
  NOR2_X2 U5769 ( .A1(n4763), .A2(n5089), .ZN(n6470) );
  INV_X1 U5770 ( .A(n6470), .ZN(n4735) );
  NAND2_X1 U5771 ( .A1(n6109), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4682) );
  AND2_X1 U5772 ( .A1(n5876), .A2(DATAI_31_), .ZN(n6397) );
  AND2_X1 U5773 ( .A1(n5876), .A2(DATAI_23_), .ZN(n6472) );
  INV_X1 U5774 ( .A(n6472), .ZN(n6401) );
  INV_X1 U5775 ( .A(DATAI_7_), .ZN(n4782) );
  NOR2_X2 U5776 ( .A1(n4782), .A2(n4761), .ZN(n6468) );
  INV_X1 U5777 ( .A(n6468), .ZN(n4814) );
  OAI22_X1 U5778 ( .A1(n6135), .A2(n6401), .B1(n6105), .B2(n4814), .ZN(n4680)
         );
  AOI21_X1 U5779 ( .B1(n6397), .B2(n6108), .A(n4680), .ZN(n4681) );
  OAI211_X1 U5780 ( .C1(n4694), .C2(n4735), .A(n4682), .B(n4681), .ZN(U3075)
         );
  NOR2_X2 U5781 ( .A1(n4763), .A2(n3440), .ZN(n6454) );
  INV_X1 U5782 ( .A(n6454), .ZN(n4745) );
  NAND2_X1 U5783 ( .A1(n6109), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4685) );
  AND2_X1 U5784 ( .A1(n5876), .A2(DATAI_29_), .ZN(n6456) );
  AND2_X1 U5785 ( .A1(n5876), .A2(DATAI_21_), .ZN(n6348) );
  INV_X1 U5786 ( .A(n6348), .ZN(n6460) );
  INV_X1 U5787 ( .A(DATAI_5_), .ZN(n4697) );
  NOR2_X2 U5788 ( .A1(n4697), .A2(n4761), .ZN(n6453) );
  INV_X1 U5789 ( .A(n6453), .ZN(n4810) );
  OAI22_X1 U5790 ( .A1(n6135), .A2(n6460), .B1(n6105), .B2(n4810), .ZN(n4683)
         );
  AOI21_X1 U5791 ( .B1(n6456), .B2(n6108), .A(n4683), .ZN(n4684) );
  OAI211_X1 U5792 ( .C1(n4694), .C2(n4745), .A(n4685), .B(n4684), .ZN(U3073)
         );
  NOR2_X2 U5793 ( .A1(n4763), .A2(n4686), .ZN(n6462) );
  INV_X1 U5794 ( .A(n6462), .ZN(n4740) );
  NAND2_X1 U5795 ( .A1(n6109), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4689) );
  AND2_X1 U5796 ( .A1(n5876), .A2(DATAI_30_), .ZN(n6390) );
  AND2_X1 U5797 ( .A1(n5876), .A2(DATAI_22_), .ZN(n6463) );
  INV_X1 U5798 ( .A(n6463), .ZN(n6393) );
  NOR2_X2 U5799 ( .A1(n6909), .A2(n4761), .ZN(n6461) );
  INV_X1 U5800 ( .A(n6461), .ZN(n4822) );
  OAI22_X1 U5801 ( .A1(n6135), .A2(n6393), .B1(n6105), .B2(n4822), .ZN(n4687)
         );
  AOI21_X1 U5802 ( .B1(n6390), .B2(n6108), .A(n4687), .ZN(n4688) );
  OAI211_X1 U5803 ( .C1(n4694), .C2(n4740), .A(n4689), .B(n4688), .ZN(U3074)
         );
  INV_X1 U5804 ( .A(n4763), .ZN(n4690) );
  NAND2_X1 U5805 ( .A1(n4690), .A2(n3408), .ZN(n6447) );
  NAND2_X1 U5806 ( .A1(n6109), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U5807 ( .A1(n5876), .A2(DATAI_28_), .ZN(n6452) );
  INV_X1 U5808 ( .A(n6452), .ZN(n4749) );
  AND2_X1 U5809 ( .A1(n5876), .A2(DATAI_20_), .ZN(n6449) );
  INV_X1 U5810 ( .A(n6449), .ZN(n6266) );
  OAI22_X1 U5811 ( .A1(n6135), .A2(n6266), .B1(n6105), .B2(n6444), .ZN(n4691)
         );
  AOI21_X1 U5812 ( .B1(n6108), .B2(n4749), .A(n4691), .ZN(n4692) );
  OAI211_X1 U5813 ( .C1(n4694), .C2(n6447), .A(n4693), .B(n4692), .ZN(U3072)
         );
  XOR2_X1 U5814 ( .A(n4696), .B(n4695), .Z(n5839) );
  INV_X1 U5815 ( .A(n5839), .ZN(n4698) );
  INV_X1 U5816 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5762) );
  OAI222_X1 U5817 ( .A1(n4698), .A2(n5677), .B1(n5691), .B2(n4697), .C1(n5090), 
        .C2(n5762), .ZN(U2886) );
  OAI21_X1 U5818 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n5843) );
  NOR2_X1 U5819 ( .A1(n5938), .A2(n5622), .ZN(n4708) );
  NOR2_X1 U5820 ( .A1(n5934), .A2(n4704), .ZN(n4706) );
  NAND2_X1 U5821 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4702) );
  OAI21_X1 U5822 ( .B1(n4702), .B2(n5951), .A(n5944), .ZN(n5929) );
  OAI211_X1 U5823 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5929), .B(n5928), .ZN(n4705) );
  NOR2_X1 U5824 ( .A1(n5944), .A2(n5928), .ZN(n5941) );
  AOI21_X1 U5825 ( .B1(n4703), .B2(n4702), .A(n4865), .ZN(n5942) );
  INV_X1 U5826 ( .A(n5942), .ZN(n5908) );
  NOR2_X1 U5827 ( .A1(n5941), .A2(n5908), .ZN(n5935) );
  OAI22_X1 U5828 ( .A1(n4706), .A2(n4705), .B1(n5935), .B2(n4704), .ZN(n4707)
         );
  AOI211_X1 U5829 ( .C1(n5860), .C2(REIP_REG_4__SCAN_IN), .A(n4708), .B(n4707), 
        .ZN(n4709) );
  OAI21_X1 U5830 ( .B1(n5963), .B2(n5843), .A(n4709), .ZN(U3014) );
  NAND2_X1 U5831 ( .A1(n6487), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6319) );
  OR2_X1 U5832 ( .A1(n6319), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4788)
         );
  NAND3_X1 U5833 ( .A1(n4710), .A2(STATEBS16_REG_SCAN_IN), .A3(n6147), .ZN(
        n4711) );
  NAND2_X1 U5834 ( .A1(n4711), .A2(n6603), .ZN(n4717) );
  NOR2_X1 U5835 ( .A1(n4576), .A2(n4528), .ZN(n6317) );
  NAND2_X1 U5836 ( .A1(n6317), .A2(n4712), .ZN(n4791) );
  OR2_X1 U5837 ( .A1(n4791), .A2(n6482), .ZN(n4713) );
  OR2_X1 U5838 ( .A1(n6283), .A2(n4788), .ZN(n4765) );
  NAND2_X1 U5839 ( .A1(n4713), .A2(n4765), .ZN(n4715) );
  NOR2_X1 U5840 ( .A1(n4717), .A2(n4715), .ZN(n4714) );
  INV_X1 U5841 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4723) );
  INV_X1 U5842 ( .A(n4715), .ZN(n4716) );
  OAI22_X1 U5843 ( .A1(n4717), .A2(n4716), .B1(n4788), .B2(n6251), .ZN(n4768)
         );
  AOI22_X1 U5844 ( .A1(n6100), .A2(n6440), .B1(n6108), .B2(n6224), .ZN(n4719)
         );
  OAI21_X1 U5845 ( .B1(n4720), .B2(n4765), .A(n4719), .ZN(n4721) );
  AOI21_X1 U5846 ( .B1(n6438), .B2(n4768), .A(n4721), .ZN(n4722) );
  OAI21_X1 U5847 ( .B1(n4771), .B2(n4723), .A(n4722), .ZN(U3063) );
  INV_X1 U5848 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5849 ( .A1(n6100), .A2(n6434), .B1(n6108), .B2(n6259), .ZN(n4724)
         );
  OAI21_X1 U5850 ( .B1(n4725), .B2(n4765), .A(n4724), .ZN(n4726) );
  AOI21_X1 U5851 ( .B1(n6432), .B2(n4768), .A(n4726), .ZN(n4727) );
  OAI21_X1 U5852 ( .B1(n4771), .B2(n4728), .A(n4727), .ZN(U3062) );
  INV_X1 U5853 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5854 ( .A1(n6100), .A2(n6428), .B1(n6108), .B2(n6335), .ZN(n4729)
         );
  OAI21_X1 U5855 ( .B1(n4730), .B2(n4765), .A(n4729), .ZN(n4731) );
  AOI21_X1 U5856 ( .B1(n6426), .B2(n4768), .A(n4731), .ZN(n4732) );
  OAI21_X1 U5857 ( .B1(n4771), .B2(n4733), .A(n4732), .ZN(U3061) );
  INV_X1 U5858 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5859 ( .A1(n6100), .A2(n6397), .B1(n6108), .B2(n6472), .ZN(n4734)
         );
  OAI21_X1 U5860 ( .B1(n4735), .B2(n4765), .A(n4734), .ZN(n4736) );
  AOI21_X1 U5861 ( .B1(n6468), .B2(n4768), .A(n4736), .ZN(n4737) );
  OAI21_X1 U5862 ( .B1(n4771), .B2(n4738), .A(n4737), .ZN(U3067) );
  INV_X1 U5863 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U5864 ( .A1(n6100), .A2(n6390), .B1(n6108), .B2(n6463), .ZN(n4739)
         );
  OAI21_X1 U5865 ( .B1(n4740), .B2(n4765), .A(n4739), .ZN(n4741) );
  AOI21_X1 U5866 ( .B1(n6461), .B2(n4768), .A(n4741), .ZN(n4742) );
  OAI21_X1 U5867 ( .B1(n4771), .B2(n4743), .A(n4742), .ZN(U3066) );
  INV_X1 U5868 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4748) );
  AOI22_X1 U5869 ( .A1(n6100), .A2(n6456), .B1(n6108), .B2(n6348), .ZN(n4744)
         );
  OAI21_X1 U5870 ( .B1(n4745), .B2(n4765), .A(n4744), .ZN(n4746) );
  AOI21_X1 U5871 ( .B1(n6453), .B2(n4768), .A(n4746), .ZN(n4747) );
  OAI21_X1 U5872 ( .B1(n4771), .B2(n4748), .A(n4747), .ZN(U3065) );
  INV_X1 U5873 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U5874 ( .A1(n6449), .A2(n6108), .B1(n6100), .B2(n4749), .ZN(n4750)
         );
  OAI21_X1 U5875 ( .B1(n6447), .B2(n4765), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5876 ( .B1(n6269), .B2(n4768), .A(n4751), .ZN(n4752) );
  OAI21_X1 U5877 ( .B1(n4771), .B2(n4753), .A(n4752), .ZN(U3064) );
  INV_X1 U5878 ( .A(n4754), .ZN(n4760) );
  INV_X1 U5879 ( .A(n4755), .ZN(n4758) );
  OAI22_X1 U5880 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n5869), .B1(n6412), 
        .B2(n4756), .ZN(n4757) );
  AOI211_X1 U5881 ( .C1(n5859), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4758), 
        .B(n4757), .ZN(n4759) );
  OAI21_X1 U5882 ( .B1(n4760), .B2(n5878), .A(n4759), .ZN(U2985) );
  INV_X1 U5883 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4770) );
  NOR2_X2 U5884 ( .A1(n4762), .A2(n4761), .ZN(n6409) );
  NOR2_X2 U5885 ( .A1(n4763), .A2(n3534), .ZN(n6410) );
  INV_X1 U5886 ( .A(n6410), .ZN(n4766) );
  AND2_X1 U5887 ( .A1(n5876), .A2(DATAI_24_), .ZN(n6422) );
  AND2_X1 U5888 ( .A1(n5876), .A2(DATAI_16_), .ZN(n6331) );
  AOI22_X1 U5889 ( .A1(n6100), .A2(n6422), .B1(n6108), .B2(n6331), .ZN(n4764)
         );
  OAI21_X1 U5890 ( .B1(n4766), .B2(n4765), .A(n4764), .ZN(n4767) );
  AOI21_X1 U5891 ( .B1(n6409), .B2(n4768), .A(n4767), .ZN(n4769) );
  OAI21_X1 U5892 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(U3060) );
  XNOR2_X1 U5893 ( .A(n4772), .B(n4773), .ZN(n5819) );
  OAI21_X1 U5894 ( .B1(n4776), .B2(n4775), .A(n4774), .ZN(n5895) );
  INV_X1 U5895 ( .A(n5895), .ZN(n4777) );
  AOI22_X1 U5896 ( .A1(n5671), .A2(n4777), .B1(n5074), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4778) );
  OAI21_X1 U5897 ( .B1(n5819), .B2(n5086), .A(n4778), .ZN(U2851) );
  INV_X1 U5898 ( .A(DATAI_8_), .ZN(n4779) );
  INV_X1 U5899 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5771) );
  OAI222_X1 U5900 ( .A1(n5819), .A2(n5677), .B1(n5691), .B2(n4779), .C1(n5090), 
        .C2(n5771), .ZN(U2883) );
  XOR2_X1 U5901 ( .A(n4781), .B(n4780), .Z(n5824) );
  INV_X1 U5902 ( .A(n5824), .ZN(n4786) );
  INV_X1 U5903 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5768) );
  OAI222_X1 U5904 ( .A1(n4786), .A2(n5677), .B1(n5691), .B2(n4782), .C1(n5090), 
        .C2(n5768), .ZN(U2884) );
  XNOR2_X1 U5905 ( .A(n4784), .B(n4783), .ZN(n5901) );
  OAI222_X1 U5906 ( .A1(n5086), .A2(n4786), .B1(n4785), .B2(n5674), .C1(n5088), 
        .C2(n5901), .ZN(U2852) );
  NAND2_X1 U5907 ( .A1(n6062), .A2(n6243), .ZN(n4787) );
  INV_X1 U5908 ( .A(n6440), .ZN(n6227) );
  NOR2_X1 U5909 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4788), .ZN(n6096)
         );
  NAND3_X1 U5910 ( .A1(n4823), .A2(n6405), .A3(n6104), .ZN(n4789) );
  NAND2_X1 U5911 ( .A1(n4789), .A2(n6034), .ZN(n4792) );
  AND2_X1 U5912 ( .A1(n6144), .A2(n4790), .ZN(n5966) );
  OAI21_X1 U5913 ( .B1(n5966), .B2(n6251), .A(n6151), .ZN(n5969) );
  AOI211_X1 U5914 ( .C1(n4792), .C2(n4791), .A(n6368), .B(n5969), .ZN(n4793)
         );
  NAND2_X1 U5915 ( .A1(n6101), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4800) );
  NAND3_X1 U5916 ( .A1(n6029), .A2(n6405), .A3(n6317), .ZN(n4796) );
  INV_X1 U5917 ( .A(n4794), .ZN(n6365) );
  NAND2_X1 U5918 ( .A1(n5966), .A2(n6365), .ZN(n4795) );
  OAI22_X1 U5919 ( .A1(n4823), .A2(n6443), .B1(n6097), .B2(n4797), .ZN(n4798)
         );
  AOI21_X1 U5920 ( .B1(n6096), .B2(n6439), .A(n4798), .ZN(n4799) );
  OAI211_X1 U5921 ( .C1(n6104), .C2(n6227), .A(n4800), .B(n4799), .ZN(U3055)
         );
  INV_X1 U5922 ( .A(n6422), .ZN(n6334) );
  NAND2_X1 U5923 ( .A1(n6101), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4805) );
  INV_X1 U5924 ( .A(n6409), .ZN(n4802) );
  NAND2_X1 U5925 ( .A1(n6100), .A2(n6331), .ZN(n4801) );
  OAI21_X1 U5926 ( .B1(n6097), .B2(n4802), .A(n4801), .ZN(n4803) );
  AOI21_X1 U5927 ( .B1(n6410), .B2(n6096), .A(n4803), .ZN(n4804) );
  OAI211_X1 U5928 ( .C1(n6334), .C2(n6104), .A(n4805), .B(n4804), .ZN(U3052)
         );
  INV_X1 U5929 ( .A(n6434), .ZN(n6262) );
  NAND2_X1 U5930 ( .A1(n6101), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4809) );
  OAI22_X1 U5931 ( .A1(n4823), .A2(n6437), .B1(n6097), .B2(n4806), .ZN(n4807)
         );
  AOI21_X1 U5932 ( .B1(n6096), .B2(n6433), .A(n4807), .ZN(n4808) );
  OAI211_X1 U5933 ( .C1(n6104), .C2(n6262), .A(n4809), .B(n4808), .ZN(U3054)
         );
  INV_X1 U5934 ( .A(n6456), .ZN(n6352) );
  NAND2_X1 U5935 ( .A1(n6101), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4813) );
  OAI22_X1 U5936 ( .A1(n4823), .A2(n6460), .B1(n6097), .B2(n4810), .ZN(n4811)
         );
  AOI21_X1 U5937 ( .B1(n6096), .B2(n6454), .A(n4811), .ZN(n4812) );
  OAI211_X1 U5938 ( .C1(n6104), .C2(n6352), .A(n4813), .B(n4812), .ZN(U3057)
         );
  INV_X1 U5939 ( .A(n6397), .ZN(n6477) );
  NAND2_X1 U5940 ( .A1(n6101), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4817) );
  OAI22_X1 U5941 ( .A1(n4823), .A2(n6401), .B1(n6097), .B2(n4814), .ZN(n4815)
         );
  AOI21_X1 U5942 ( .B1(n6096), .B2(n6470), .A(n4815), .ZN(n4816) );
  OAI211_X1 U5943 ( .C1(n6104), .C2(n6477), .A(n4817), .B(n4816), .ZN(U3059)
         );
  INV_X1 U5944 ( .A(n6428), .ZN(n6338) );
  NAND2_X1 U5945 ( .A1(n6101), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4821) );
  OAI22_X1 U5946 ( .A1(n4823), .A2(n6431), .B1(n6097), .B2(n4818), .ZN(n4819)
         );
  AOI21_X1 U5947 ( .B1(n6096), .B2(n6427), .A(n4819), .ZN(n4820) );
  OAI211_X1 U5948 ( .C1(n6104), .C2(n6338), .A(n4821), .B(n4820), .ZN(U3053)
         );
  INV_X1 U5949 ( .A(n6390), .ZN(n6466) );
  NAND2_X1 U5950 ( .A1(n6101), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4826) );
  OAI22_X1 U5951 ( .A1(n4823), .A2(n6393), .B1(n6097), .B2(n4822), .ZN(n4824)
         );
  AOI21_X1 U5952 ( .B1(n6096), .B2(n6462), .A(n4824), .ZN(n4825) );
  OAI211_X1 U5953 ( .C1(n6104), .C2(n6466), .A(n4826), .B(n4825), .ZN(U3058)
         );
  INV_X1 U5954 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5721) );
  AOI22_X1 U5955 ( .A1(n4833), .A2(UWORD_REG_3__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4827) );
  OAI21_X1 U5956 ( .B1(n5721), .B2(n4836), .A(n4827), .ZN(U2904) );
  INV_X1 U5957 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5725) );
  AOI22_X1 U5958 ( .A1(n4833), .A2(UWORD_REG_5__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4828) );
  OAI21_X1 U5959 ( .B1(n5725), .B2(n4836), .A(n4828), .ZN(U2902) );
  INV_X1 U5960 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5729) );
  AOI22_X1 U5961 ( .A1(n4833), .A2(UWORD_REG_7__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4829) );
  OAI21_X1 U5962 ( .B1(n5729), .B2(n4836), .A(n4829), .ZN(U2900) );
  INV_X1 U5963 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5717) );
  AOI22_X1 U5964 ( .A1(n4833), .A2(UWORD_REG_1__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4830) );
  OAI21_X1 U5965 ( .B1(n5717), .B2(n4836), .A(n4830), .ZN(U2906) );
  INV_X1 U5966 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5727) );
  AOI22_X1 U5967 ( .A1(n4833), .A2(UWORD_REG_6__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4831) );
  OAI21_X1 U5968 ( .B1(n5727), .B2(n4836), .A(n4831), .ZN(U2901) );
  INV_X1 U5969 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5719) );
  AOI22_X1 U5970 ( .A1(n4833), .A2(UWORD_REG_2__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4832) );
  OAI21_X1 U5971 ( .B1(n5719), .B2(n4836), .A(n4832), .ZN(U2905) );
  INV_X1 U5972 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5723) );
  AOI22_X1 U5973 ( .A1(n4833), .A2(UWORD_REG_4__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4834) );
  OAI21_X1 U5974 ( .B1(n5723), .B2(n4836), .A(n4834), .ZN(U2903) );
  INV_X1 U5975 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5715) );
  AOI22_X1 U5976 ( .A1(n4833), .A2(UWORD_REG_0__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4835) );
  OAI21_X1 U5977 ( .B1(n5715), .B2(n4836), .A(n4835), .ZN(U2907) );
  OAI21_X1 U5978 ( .B1(n4837), .B2(n4839), .A(n4838), .ZN(n5811) );
  AOI21_X1 U5979 ( .B1(n4840), .B2(n4774), .A(n3207), .ZN(n5887) );
  AOI22_X1 U5980 ( .A1(n5671), .A2(n5887), .B1(EBX_REG_9__SCAN_IN), .B2(n5074), 
        .ZN(n4841) );
  OAI21_X1 U5981 ( .B1(n5811), .B2(n5086), .A(n4841), .ZN(U2850) );
  INV_X1 U5982 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5774) );
  INV_X1 U5983 ( .A(DATAI_9_), .ZN(n4842) );
  OAI222_X1 U5984 ( .A1(n5677), .A2(n5811), .B1(n5090), .B2(n5774), .C1(n4842), 
        .C2(n5691), .ZN(U2882) );
  AOI21_X1 U5985 ( .B1(n4838), .B2(n4843), .A(n3219), .ZN(n5564) );
  INV_X1 U5986 ( .A(n5564), .ZN(n4845) );
  INV_X1 U5987 ( .A(DATAI_10_), .ZN(n6865) );
  INV_X1 U5988 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5777) );
  OAI222_X1 U5989 ( .A1(n4845), .A2(n5677), .B1(n5691), .B2(n6865), .C1(n5090), 
        .C2(n5777), .ZN(U2881) );
  OAI21_X1 U5990 ( .B1(n4844), .B2(n3207), .A(n4850), .ZN(n5562) );
  OAI222_X1 U5991 ( .A1(n5562), .A2(n5088), .B1(n4846), .B2(n5674), .C1(n4845), 
        .C2(n5086), .ZN(U2849) );
  OAI21_X1 U5992 ( .B1(n3219), .B2(n4849), .A(n4848), .ZN(n5803) );
  AOI21_X1 U5993 ( .B1(n4851), .B2(n4850), .A(n4856), .ZN(n5879) );
  AOI22_X1 U5994 ( .A1(n5671), .A2(n5879), .B1(n5074), .B2(EBX_REG_11__SCAN_IN), .ZN(n4852) );
  OAI21_X1 U5995 ( .B1(n5803), .B2(n5086), .A(n4852), .ZN(U2848) );
  INV_X1 U5996 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5780) );
  INV_X1 U5997 ( .A(DATAI_11_), .ZN(n4853) );
  OAI222_X1 U5998 ( .A1(n5677), .A2(n5803), .B1(n5090), .B2(n5780), .C1(n4853), 
        .C2(n5691), .ZN(U2880) );
  AOI21_X1 U5999 ( .B1(n4848), .B2(n4854), .A(n3955), .ZN(n4902) );
  INV_X1 U6000 ( .A(n4902), .ZN(n5548) );
  INV_X1 U6001 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4857) );
  XNOR2_X1 U6002 ( .A(n4856), .B(n4855), .ZN(n5544) );
  OAI222_X1 U6003 ( .A1(n5548), .A2(n5086), .B1(n4857), .B2(n5674), .C1(n5088), 
        .C2(n5544), .ZN(U2847) );
  INV_X1 U6004 ( .A(DATAI_12_), .ZN(n4858) );
  INV_X1 U6005 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5783) );
  OAI222_X1 U6006 ( .A1(n5548), .A2(n5677), .B1(n5691), .B2(n4858), .C1(n5090), 
        .C2(n5783), .ZN(U2879) );
  NAND2_X1 U6007 ( .A1(n5795), .A2(n4859), .ZN(n4861) );
  XOR2_X1 U6008 ( .A(n4861), .B(n4860), .Z(n4877) );
  INV_X1 U6009 ( .A(n4867), .ZN(n5894) );
  OAI22_X1 U6010 ( .A1(n4866), .A2(n5944), .B1(n4863), .B2(n4862), .ZN(n4864)
         );
  NOR2_X1 U6011 ( .A1(n4865), .A2(n4864), .ZN(n5905) );
  OAI21_X1 U6012 ( .B1(n5894), .B2(n5197), .A(n5905), .ZN(n5886) );
  INV_X1 U6013 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6560) );
  OAI22_X1 U6014 ( .A1(n5938), .A2(n5562), .B1(n6560), .B2(n5937), .ZN(n4871)
         );
  NAND2_X1 U6015 ( .A1(n4866), .A2(n5929), .ZN(n5907) );
  NOR2_X1 U6016 ( .A1(n4867), .A2(n5907), .ZN(n5888) );
  OAI211_X1 U6017 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5888), .B(n4868), .ZN(n4869) );
  INV_X1 U6018 ( .A(n4869), .ZN(n4870) );
  AOI211_X1 U6019 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n5886), .A(n4871), .B(n4870), .ZN(n4872) );
  OAI21_X1 U6020 ( .B1(n4877), .B2(n5963), .A(n4872), .ZN(U3008) );
  NAND2_X1 U6021 ( .A1(n5564), .A2(n5876), .ZN(n4876) );
  INV_X1 U6022 ( .A(n5859), .ZN(n5872) );
  OAI22_X1 U6023 ( .A1(n5872), .A2(n4873), .B1(n5937), .B2(n6560), .ZN(n4874)
         );
  AOI21_X1 U6024 ( .B1(n5845), .B2(n5565), .A(n4874), .ZN(n4875) );
  OAI211_X1 U6025 ( .C1(n4877), .C2(n5878), .A(n4876), .B(n4875), .ZN(U2976)
         );
  OR2_X1 U6026 ( .A1(n4879), .A2(n4878), .ZN(n4881) );
  NAND2_X1 U6027 ( .A1(n4881), .A2(n4880), .ZN(n5543) );
  XNOR2_X1 U6028 ( .A(n4883), .B(n4882), .ZN(n5533) );
  INV_X1 U6029 ( .A(n5533), .ZN(n4884) );
  AOI22_X1 U6030 ( .A1(n5671), .A2(n4884), .B1(n5074), .B2(EBX_REG_13__SCAN_IN), .ZN(n4885) );
  OAI21_X1 U6031 ( .B1(n5086), .B2(n5543), .A(n4885), .ZN(U2846) );
  INV_X1 U6032 ( .A(DATAI_13_), .ZN(n4886) );
  INV_X1 U6033 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5786) );
  OAI222_X1 U6034 ( .A1(n5543), .A2(n5677), .B1(n5691), .B2(n4886), .C1(n5090), 
        .C2(n5786), .ZN(U2878) );
  NOR2_X1 U6035 ( .A1(n4889), .A2(n3268), .ZN(n4890) );
  XNOR2_X1 U6036 ( .A(n4887), .B(n4890), .ZN(n4904) );
  NOR2_X1 U6037 ( .A1(n5209), .A2(n5884), .ZN(n4895) );
  NAND2_X1 U6038 ( .A1(n5944), .A2(n4891), .ZN(n5173) );
  INV_X1 U6039 ( .A(n5885), .ZN(n4892) );
  AOI21_X1 U6040 ( .B1(n5884), .B2(n5173), .A(n4892), .ZN(n4893) );
  INV_X1 U6041 ( .A(n4893), .ZN(n4894) );
  MUX2_X1 U6042 ( .A(n4895), .B(n4894), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n4897) );
  OAI22_X1 U6043 ( .A1(n5938), .A2(n5544), .B1(n6562), .B2(n5937), .ZN(n4896)
         );
  NOR2_X1 U6044 ( .A1(n4897), .A2(n4896), .ZN(n4898) );
  OAI21_X1 U6045 ( .B1(n4904), .B2(n5963), .A(n4898), .ZN(U3006) );
  AOI22_X1 U6046 ( .A1(n5859), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n5860), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n4899) );
  OAI21_X1 U6047 ( .B1(n5869), .B2(n4900), .A(n4899), .ZN(n4901) );
  AOI21_X1 U6048 ( .B1(n4902), .B2(n5876), .A(n4901), .ZN(n4903) );
  OAI21_X1 U6049 ( .B1(n4904), .B2(n5878), .A(n4903), .ZN(U2974) );
  OAI21_X1 U6050 ( .B1(n4905), .B2(n4908), .A(n4907), .ZN(n5531) );
  INV_X1 U6051 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5789) );
  INV_X1 U6052 ( .A(DATAI_14_), .ZN(n4909) );
  OAI222_X1 U6053 ( .A1(n5677), .A2(n5531), .B1(n5090), .B2(n5789), .C1(n4909), 
        .C2(n5691), .ZN(U2877) );
  OAI21_X1 U6054 ( .B1(n4912), .B2(n4911), .A(n4910), .ZN(n5523) );
  OAI222_X1 U6055 ( .A1(n5088), .A2(n5523), .B1(n5674), .B2(n4365), .C1(n5086), 
        .C2(n5531), .ZN(U2845) );
  INV_X1 U6056 ( .A(n5955), .ZN(n4915) );
  NAND2_X1 U6057 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4913) );
  AOI22_X1 U6058 ( .A1(n4915), .A2(n5208), .B1(n4914), .B2(n4913), .ZN(n4916)
         );
  NAND2_X1 U6059 ( .A1(n5885), .A2(n4916), .ZN(n5210) );
  INV_X1 U6060 ( .A(n5210), .ZN(n4931) );
  XNOR2_X1 U6061 ( .A(n4917), .B(n4918), .ZN(n5402) );
  NAND2_X1 U6062 ( .A1(n5402), .A2(n5946), .ZN(n4930) );
  INV_X1 U6063 ( .A(n4919), .ZN(n4921) );
  NAND3_X1 U6064 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4921), .A3(n4920), 
        .ZN(n4922) );
  NAND3_X1 U6065 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n4932), .ZN(n4924) );
  AOI21_X1 U6066 ( .B1(n4923), .B2(n4922), .A(n4924), .ZN(n5211) );
  NOR3_X1 U6067 ( .A1(n5955), .A2(n4925), .A3(n4924), .ZN(n4928) );
  INV_X1 U6068 ( .A(REIP_REG_13__SCAN_IN), .ZN(n4926) );
  OAI22_X1 U6069 ( .A1(n5938), .A2(n5533), .B1(n5937), .B2(n4926), .ZN(n4927)
         );
  NOR3_X1 U6070 ( .A1(n5211), .A2(n4928), .A3(n4927), .ZN(n4929) );
  OAI211_X1 U6071 ( .C1(n4932), .C2(n4931), .A(n4930), .B(n4929), .ZN(U3005)
         );
  OAI21_X1 U6072 ( .B1(n4933), .B2(n4935), .A(n4934), .ZN(n5514) );
  AOI22_X1 U6073 ( .A1(n5684), .A2(DATAI_0_), .B1(n5687), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6074 ( .A1(n5682), .A2(DATAI_16_), .ZN(n4936) );
  OAI211_X1 U6075 ( .C1(n5514), .C2(n5677), .A(n4937), .B(n4936), .ZN(U2875)
         );
  OAI21_X1 U6076 ( .B1(n4938), .B2(n5456), .A(n5450), .ZN(n5503) );
  OAI222_X1 U6077 ( .A1(n5088), .A2(n5503), .B1(n5674), .B2(n4371), .C1(n5086), 
        .C2(n5514), .ZN(U2843) );
  AND2_X1 U6078 ( .A1(n4942), .A2(n3535), .ZN(n4939) );
  INV_X1 U6079 ( .A(n5648), .ZN(n5664) );
  INV_X1 U6080 ( .A(n5858), .ZN(n4950) );
  INV_X1 U6081 ( .A(n4940), .ZN(n4941) );
  NAND2_X1 U6082 ( .A1(n4942), .A2(n4941), .ZN(n5656) );
  NOR2_X1 U6083 ( .A1(n5611), .A2(REIP_REG_1__SCAN_IN), .ZN(n5640) );
  INV_X1 U6084 ( .A(n5651), .ZN(n4943) );
  NOR3_X1 U6085 ( .A1(n5640), .A2(n4943), .A3(n6551), .ZN(n5631) );
  OAI21_X1 U6086 ( .B1(n5611), .B2(n5621), .A(n5651), .ZN(n5620) );
  OAI21_X1 U6087 ( .B1(n5631), .B2(REIP_REG_3__SCAN_IN), .A(n5620), .ZN(n4948)
         );
  INV_X1 U6088 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4945) );
  OAI22_X1 U6089 ( .A1(n5654), .A2(n4945), .B1(n5641), .B2(n4944), .ZN(n4946)
         );
  AOI21_X1 U6090 ( .B1(n5644), .B2(EBX_REG_3__SCAN_IN), .A(n4946), .ZN(n4947)
         );
  OAI211_X1 U6091 ( .C1(n6029), .C2(n5656), .A(n4948), .B(n4947), .ZN(n4949)
         );
  AOI21_X1 U6092 ( .B1(n5601), .B2(n4950), .A(n4949), .ZN(n4951) );
  OAI21_X1 U6093 ( .B1(n5664), .B2(n5854), .A(n4951), .ZN(U2824) );
  INV_X1 U6094 ( .A(n6521), .ZN(n4968) );
  AOI21_X1 U6095 ( .B1(n4952), .B2(n4968), .A(n5223), .ZN(n4960) );
  OAI21_X1 U6096 ( .B1(n6521), .B2(n6479), .A(n6510), .ZN(n4958) );
  NAND2_X1 U6097 ( .A1(n4953), .A2(n6373), .ZN(n4955) );
  OAI21_X1 U6098 ( .B1(n4955), .B2(n6482), .A(n4954), .ZN(n4956) );
  AOI22_X1 U6099 ( .A1(n4958), .A2(n3448), .B1(n4957), .B2(n4956), .ZN(n4959)
         );
  OAI22_X1 U6100 ( .A1(n4960), .A2(n3448), .B1(n5223), .B2(n4959), .ZN(U3461)
         );
  INV_X1 U6101 ( .A(n6510), .ZN(n4961) );
  AOI21_X1 U6102 ( .B1(n4961), .B2(n4964), .A(n5223), .ZN(n4970) );
  AND2_X1 U6103 ( .A1(n4963), .A2(n4962), .ZN(n4966) );
  NOR3_X1 U6104 ( .A1(n6510), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4964), 
        .ZN(n4965) );
  AOI211_X1 U6105 ( .C1(n4968), .C2(n4967), .A(n4966), .B(n4965), .ZN(n4969)
         );
  OAI22_X1 U6106 ( .A1(n4970), .A2(n3166), .B1(n5223), .B2(n4969), .ZN(U3459)
         );
  OR2_X1 U6107 ( .A1(n4978), .A2(n4971), .ZN(n4976) );
  NAND2_X1 U6108 ( .A1(n4981), .A2(n4274), .ZN(n4975) );
  NAND2_X1 U6109 ( .A1(n4972), .A2(n4979), .ZN(n4973) );
  NAND2_X1 U6110 ( .A1(n4978), .A2(n4973), .ZN(n4974) );
  AND3_X1 U6111 ( .A1(n4976), .A2(n4975), .A3(n4974), .ZN(n6496) );
  INV_X1 U6112 ( .A(n6496), .ZN(n4990) );
  NAND2_X1 U6113 ( .A1(n4978), .A2(n4977), .ZN(n4983) );
  OAI21_X1 U6114 ( .B1(n4981), .B2(n4980), .A(n4979), .ZN(n4982) );
  NAND2_X1 U6115 ( .A1(n4983), .A2(n4982), .ZN(n5468) );
  OAI21_X1 U6116 ( .B1(n4984), .B2(n3445), .A(n6896), .ZN(n4985) );
  INV_X1 U6117 ( .A(n4985), .ZN(n4989) );
  OR2_X1 U6118 ( .A1(n4987), .A2(n4986), .ZN(n4988) );
  AND2_X1 U6119 ( .A1(n4989), .A2(n4988), .ZN(n6594) );
  OR2_X1 U6120 ( .A1(n5468), .A2(n6594), .ZN(n6498) );
  AND2_X1 U6121 ( .A1(n6498), .A2(n6522), .ZN(n5474) );
  MUX2_X1 U6122 ( .A(MORE_REG_SCAN_IN), .B(n4990), .S(n5474), .Z(U3471) );
  OR2_X1 U6123 ( .A1(n4991), .A2(n3217), .ZN(n4992) );
  NAND2_X1 U6124 ( .A1(n4992), .A2(n5023), .ZN(n5149) );
  OAI22_X1 U6125 ( .A1(n4994), .A2(n5658), .B1(n4993), .B2(n5654), .ZN(n5001)
         );
  INV_X1 U6126 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6880) );
  NOR2_X1 U6127 ( .A1(n6880), .A2(n5269), .ZN(n5267) );
  AOI21_X1 U6128 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5267), .A(
        REIP_REG_26__SCAN_IN), .ZN(n4998) );
  OAI22_X1 U6129 ( .A1(n4999), .A2(n4998), .B1(n5353), .B2(n5599), .ZN(n5000)
         );
  OAI21_X1 U6130 ( .B1(n5641), .B2(n5149), .A(n5002), .ZN(U2801) );
  XNOR2_X1 U6131 ( .A(n5004), .B(n5003), .ZN(n5429) );
  AOI21_X1 U6132 ( .B1(n5005), .B2(n5007), .A(n5006), .ZN(n5371) );
  INV_X1 U6133 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5058) );
  OAI22_X1 U6134 ( .A1(n5058), .A2(n5658), .B1(n5369), .B2(n5655), .ZN(n5009)
         );
  INV_X1 U6135 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5373) );
  OAI22_X1 U6136 ( .A1(n5373), .A2(n5654), .B1(n6568), .B2(n5296), .ZN(n5008)
         );
  AOI211_X1 U6137 ( .C1(n5371), .C2(n5592), .A(n5009), .B(n5008), .ZN(n5010)
         );
  NAND2_X1 U6138 ( .A1(n5284), .A2(n6568), .ZN(n5295) );
  OAI211_X1 U6139 ( .C1(n5641), .C2(n5429), .A(n5010), .B(n5295), .ZN(U2806)
         );
  INV_X1 U6140 ( .A(n5011), .ZN(n5013) );
  OAI22_X1 U6141 ( .A1(n5013), .A2(n5088), .B1(n5674), .B2(n5012), .ZN(U2828)
         );
  AOI21_X1 U6142 ( .B1(n5014), .B2(n5016), .A(n5015), .ZN(n5317) );
  INV_X1 U6143 ( .A(n5317), .ZN(n5259) );
  AOI22_X1 U6144 ( .A1(n5671), .A2(n5249), .B1(EBX_REG_29__SCAN_IN), .B2(n5074), .ZN(n5017) );
  OAI21_X1 U6145 ( .B1(n5259), .B2(n5086), .A(n5017), .ZN(U2830) );
  AOI22_X1 U6146 ( .A1(n5671), .A2(n5018), .B1(EBX_REG_28__SCAN_IN), .B2(n5074), .ZN(n5019) );
  OAI21_X1 U6147 ( .B1(n5097), .B2(n5086), .A(n5019), .ZN(U2831) );
  AOI21_X1 U6148 ( .B1(n4996), .B2(n5020), .A(n4201), .ZN(n5345) );
  INV_X1 U6149 ( .A(n5345), .ZN(n5025) );
  AOI21_X1 U6150 ( .B1(n5023), .B2(n5022), .A(n4496), .ZN(n5405) );
  AOI22_X1 U6151 ( .A1(n5671), .A2(n5405), .B1(EBX_REG_27__SCAN_IN), .B2(n5074), .ZN(n5024) );
  OAI21_X1 U6152 ( .B1(n5025), .B2(n5086), .A(n5024), .ZN(U2832) );
  INV_X1 U6153 ( .A(n5149), .ZN(n5026) );
  AOI22_X1 U6154 ( .A1(n5671), .A2(n5026), .B1(n5074), .B2(EBX_REG_26__SCAN_IN), .ZN(n5027) );
  OAI21_X1 U6155 ( .B1(n5353), .B2(n5086), .A(n5027), .ZN(U2833) );
  AOI21_X1 U6156 ( .B1(n5029), .B2(n5028), .A(n3217), .ZN(n5415) );
  INV_X1 U6157 ( .A(n5415), .ZN(n5034) );
  AOI21_X1 U6158 ( .B1(n5030), .B2(n5031), .A(n4995), .ZN(n5355) );
  INV_X1 U6159 ( .A(n5355), .ZN(n5032) );
  OAI222_X1 U6160 ( .A1(n5034), .A2(n5088), .B1(n5033), .B2(n5674), .C1(n5032), 
        .C2(n5086), .ZN(U2834) );
  BUF_X1 U6161 ( .A(n5035), .Z(n5036) );
  INV_X1 U6162 ( .A(n5036), .ZN(n5047) );
  INV_X1 U6163 ( .A(n5037), .ZN(n5038) );
  NAND2_X1 U6164 ( .A1(n5047), .A2(n5038), .ZN(n5039) );
  AND2_X1 U6165 ( .A1(n5039), .A2(n5030), .ZN(n5324) );
  INV_X1 U6166 ( .A(n5324), .ZN(n5044) );
  INV_X1 U6167 ( .A(n5040), .ZN(n5041) );
  XNOR2_X1 U6168 ( .A(n5050), .B(n5041), .ZN(n5275) );
  INV_X1 U6169 ( .A(n5275), .ZN(n5042) );
  OAI222_X1 U6170 ( .A1(n5044), .A2(n5086), .B1(n5043), .B2(n5674), .C1(n5088), 
        .C2(n5042), .ZN(U2835) );
  NAND2_X1 U6171 ( .A1(n3212), .A2(n5045), .ZN(n5046) );
  NAND2_X1 U6172 ( .A1(n5047), .A2(n5046), .ZN(n5327) );
  AND2_X1 U6173 ( .A1(n5056), .A2(n5048), .ZN(n5049) );
  NOR2_X1 U6174 ( .A1(n5050), .A2(n5049), .ZN(n5285) );
  AOI22_X1 U6175 ( .A1(n5671), .A2(n5285), .B1(n5074), .B2(EBX_REG_23__SCAN_IN), .ZN(n5051) );
  OAI21_X1 U6176 ( .B1(n5327), .B2(n5086), .A(n5051), .ZN(U2836) );
  OAI21_X1 U6177 ( .B1(n5052), .B2(n5006), .A(n3212), .ZN(n5365) );
  NAND2_X1 U6178 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  NAND2_X1 U6179 ( .A1(n5056), .A2(n5055), .ZN(n5421) );
  OAI222_X1 U6180 ( .A1(n5365), .A2(n5086), .B1(n5674), .B2(n4386), .C1(n5421), 
        .C2(n5088), .ZN(U2837) );
  INV_X1 U6181 ( .A(n5371), .ZN(n5057) );
  OAI222_X1 U6182 ( .A1(n5088), .A2(n5429), .B1(n5674), .B2(n5058), .C1(n5086), 
        .C2(n5057), .ZN(U2838) );
  INV_X1 U6183 ( .A(n5080), .ZN(n5060) );
  NAND2_X1 U6184 ( .A1(n5059), .A2(n5060), .ZN(n5061) );
  OAI21_X1 U6185 ( .B1(n5059), .B2(n4294), .A(n5061), .ZN(n5063) );
  XNOR2_X1 U6186 ( .A(n5063), .B(n5062), .ZN(n5297) );
  BUF_X1 U6187 ( .A(n5064), .Z(n5065) );
  OAI21_X1 U6188 ( .B1(n5065), .B2(n5066), .A(n5005), .ZN(n5378) );
  INV_X1 U6189 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5067) );
  OAI222_X1 U6190 ( .A1(n5088), .A2(n5297), .B1(n5086), .B2(n5378), .C1(n5067), 
        .C2(n5674), .ZN(U2839) );
  AOI21_X1 U6191 ( .B1(n5068), .B2(n5069), .A(n5065), .ZN(n5380) );
  INV_X1 U6192 ( .A(n5380), .ZN(n5076) );
  NAND2_X1 U6193 ( .A1(n5077), .A2(n3152), .ZN(n5071) );
  NAND3_X1 U6194 ( .A1(n5070), .A2(n5072), .A3(n5071), .ZN(n5083) );
  XNOR2_X1 U6195 ( .A(n5083), .B(n5073), .ZN(n5308) );
  AOI22_X1 U6196 ( .A1(n5671), .A2(n5308), .B1(n5074), .B2(EBX_REG_19__SCAN_IN), .ZN(n5075) );
  OAI21_X1 U6197 ( .B1(n5076), .B2(n5086), .A(n5075), .ZN(U2840) );
  INV_X1 U6198 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6199 ( .A1(n5078), .A2(n3152), .ZN(n5079) );
  OAI21_X1 U6200 ( .B1(n5080), .B2(n3152), .A(n5079), .ZN(n5081) );
  OR2_X1 U6201 ( .A1(n5070), .A2(n5081), .ZN(n5082) );
  NAND2_X1 U6202 ( .A1(n5083), .A2(n5082), .ZN(n5491) );
  INV_X1 U6203 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5087) );
  OAI21_X1 U6204 ( .B1(n5084), .B2(n5085), .A(n5068), .ZN(n5678) );
  OAI222_X1 U6205 ( .A1(n5088), .A2(n5491), .B1(n5087), .B2(n5674), .C1(n5086), 
        .C2(n5678), .ZN(U2841) );
  AOI22_X1 U6206 ( .A1(n5682), .A2(DATAI_31_), .B1(n5687), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6207 ( .A1(n5094), .A2(n5093), .ZN(U2860) );
  AOI22_X1 U6208 ( .A1(n5684), .A2(DATAI_12_), .B1(n5687), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6209 ( .A1(n5682), .A2(DATAI_28_), .ZN(n5095) );
  OAI211_X1 U6210 ( .C1(n5097), .C2(n5677), .A(n5096), .B(n5095), .ZN(U2863)
         );
  AOI22_X1 U6211 ( .A1(n5684), .A2(DATAI_10_), .B1(n5687), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6212 ( .A1(n5682), .A2(DATAI_26_), .ZN(n5098) );
  OAI211_X1 U6213 ( .C1(n5353), .C2(n5677), .A(n5099), .B(n5098), .ZN(U2865)
         );
  AOI22_X1 U6214 ( .A1(n5684), .A2(DATAI_6_), .B1(n5687), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6215 ( .A1(n5682), .A2(DATAI_22_), .ZN(n5100) );
  OAI211_X1 U6216 ( .C1(n5365), .C2(n5677), .A(n5101), .B(n5100), .ZN(U2869)
         );
  AOI22_X1 U6217 ( .A1(n5684), .A2(DATAI_4_), .B1(n5687), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6218 ( .A1(n5682), .A2(DATAI_20_), .ZN(n5102) );
  OAI211_X1 U6219 ( .C1(n5378), .C2(n5677), .A(n5103), .B(n5102), .ZN(U2871)
         );
  NAND2_X1 U6220 ( .A1(n5317), .A2(n5876), .ZN(n5108) );
  NOR2_X1 U6221 ( .A1(n5248), .A2(n5869), .ZN(n5105) );
  AOI211_X1 U6222 ( .C1(n5859), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5106), 
        .B(n5105), .ZN(n5107) );
  OAI211_X1 U6223 ( .C1(n5104), .C2(n5878), .A(n5108), .B(n5107), .ZN(U2957)
         );
  XNOR2_X1 U6224 ( .A(n3727), .B(n5190), .ZN(n5184) );
  INV_X1 U6225 ( .A(n5176), .ZN(n5109) );
  NAND2_X1 U6226 ( .A1(n5109), .A2(n3294), .ZN(n5111) );
  OR2_X1 U6227 ( .A1(n5112), .A2(n5183), .ZN(n5110) );
  XNOR2_X1 U6228 ( .A(n5797), .B(n5435), .ZN(n5368) );
  NOR2_X1 U6229 ( .A1(n3727), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5359)
         );
  NAND2_X1 U6230 ( .A1(n5366), .A2(n5359), .ZN(n5121) );
  OAI21_X1 U6231 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5121), .A(n5113), 
        .ZN(n5114) );
  XNOR2_X1 U6232 ( .A(n5114), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5163)
         );
  INV_X1 U6233 ( .A(n5274), .ZN(n5116) );
  NAND2_X1 U6234 ( .A1(n5860), .A2(REIP_REG_24__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6235 ( .A1(n5859), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5115)
         );
  OAI211_X1 U6236 ( .C1(n5116), .C2(n5869), .A(n5158), .B(n5115), .ZN(n5117)
         );
  AOI21_X1 U6237 ( .B1(n5324), .B2(n5876), .A(n5117), .ZN(n5118) );
  OAI21_X1 U6238 ( .B1(n5163), .B2(n5878), .A(n5118), .ZN(U2962) );
  INV_X1 U6239 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6240 ( .A1(n5797), .A2(n5120), .ZN(n5122) );
  OAI21_X1 U6241 ( .B1(n5123), .B2(n5122), .A(n5121), .ZN(n5124) );
  XNOR2_X1 U6242 ( .A(n5124), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5172)
         );
  INV_X1 U6243 ( .A(n5327), .ZN(n5127) );
  NOR2_X1 U6244 ( .A1(n5937), .A2(n6569), .ZN(n5164) );
  AOI21_X1 U6245 ( .B1(n5859), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5164), 
        .ZN(n5125) );
  OAI21_X1 U6246 ( .B1(n5281), .B2(n5869), .A(n5125), .ZN(n5126) );
  AOI21_X1 U6247 ( .B1(n5127), .B2(n5876), .A(n5126), .ZN(n5128) );
  OAI21_X1 U6248 ( .B1(n5172), .B2(n5878), .A(n5128), .ZN(U2963) );
  XNOR2_X1 U6249 ( .A(n5797), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5130)
         );
  XNOR2_X1 U6250 ( .A(n5129), .B(n5130), .ZN(n5455) );
  AOI21_X1 U6251 ( .B1(n4907), .B2(n5131), .A(n4933), .ZN(n5689) );
  INV_X1 U6252 ( .A(n5515), .ZN(n5133) );
  AOI22_X1 U6253 ( .A1(n5859), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5860), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5132) );
  OAI21_X1 U6254 ( .B1(n5869), .B2(n5133), .A(n5132), .ZN(n5134) );
  AOI21_X1 U6255 ( .B1(n5689), .B2(n5876), .A(n5134), .ZN(n5135) );
  OAI21_X1 U6256 ( .B1(n5455), .B2(n5878), .A(n5135), .ZN(U2971) );
  INV_X1 U6257 ( .A(n5408), .ZN(n5144) );
  OAI22_X1 U6258 ( .A1(n5938), .A2(n5136), .B1(n5937), .B2(n6952), .ZN(n5137)
         );
  AOI21_X1 U6259 ( .B1(n5946), .B2(n5138), .A(n5137), .ZN(n5142) );
  AOI21_X1 U6260 ( .B1(n5143), .B2(n5409), .A(n5139), .ZN(n5140) );
  NAND2_X1 U6261 ( .A1(n5410), .A2(n5140), .ZN(n5141) );
  OAI211_X1 U6262 ( .C1(n5144), .C2(n5143), .A(n5142), .B(n5141), .ZN(U2990)
         );
  NAND2_X1 U6263 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  XNOR2_X1 U6264 ( .A(n4416), .B(n5147), .ZN(n5350) );
  INV_X1 U6265 ( .A(n5350), .ZN(n5157) );
  INV_X1 U6266 ( .A(n5420), .ZN(n5155) );
  INV_X1 U6267 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5148) );
  OAI22_X1 U6268 ( .A1(n5938), .A2(n5149), .B1(n5937), .B2(n5148), .ZN(n5154)
         );
  INV_X1 U6269 ( .A(n5150), .ZN(n5151) );
  AOI211_X1 U6270 ( .C1(n5152), .C2(n5419), .A(n5151), .B(n5413), .ZN(n5153)
         );
  AOI211_X1 U6271 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5155), .A(n5154), .B(n5153), .ZN(n5156) );
  OAI21_X1 U6272 ( .B1(n5157), .B2(n5963), .A(n5156), .ZN(U2992) );
  AOI21_X1 U6273 ( .B1(n5165), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6274 ( .A1(n5958), .A2(n5275), .ZN(n5159) );
  OAI211_X1 U6275 ( .C1(n5420), .C2(n5160), .A(n5159), .B(n5158), .ZN(n5161)
         );
  INV_X1 U6276 ( .A(n5161), .ZN(n5162) );
  OAI21_X1 U6277 ( .B1(n5163), .B2(n5963), .A(n5162), .ZN(U2994) );
  AOI21_X1 U6278 ( .B1(n5958), .B2(n5285), .A(n5164), .ZN(n5167) );
  NAND2_X1 U6279 ( .A1(n5165), .A2(n5168), .ZN(n5166) );
  OAI211_X1 U6280 ( .C1(n5169), .C2(n5168), .A(n5167), .B(n5166), .ZN(n5170)
         );
  INV_X1 U6281 ( .A(n5170), .ZN(n5171) );
  OAI21_X1 U6282 ( .B1(n5172), .B2(n5963), .A(n5171), .ZN(U2995) );
  AOI21_X1 U6283 ( .B1(n5447), .B2(n5173), .A(n5446), .ZN(n5443) );
  INV_X1 U6284 ( .A(n5443), .ZN(n5174) );
  AOI21_X1 U6285 ( .B1(n5442), .B2(n5910), .A(n5174), .ZN(n5191) );
  XNOR2_X1 U6286 ( .A(n5797), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5175)
         );
  XNOR2_X1 U6287 ( .A(n5176), .B(n5175), .ZN(n5375) );
  NAND2_X1 U6288 ( .A1(n5375), .A2(n5946), .ZN(n5182) );
  NOR3_X1 U6289 ( .A1(n5178), .A2(n5177), .A3(n5186), .ZN(n5180) );
  NOR2_X1 U6290 ( .A1(n5938), .A2(n5297), .ZN(n5179) );
  AOI211_X1 U6291 ( .C1(n5860), .C2(REIP_REG_20__SCAN_IN), .A(n5180), .B(n5179), .ZN(n5181) );
  OAI211_X1 U6292 ( .C1(n5191), .C2(n5183), .A(n5182), .B(n5181), .ZN(U2998)
         );
  XNOR2_X1 U6293 ( .A(n5185), .B(n5184), .ZN(n5379) );
  INV_X1 U6294 ( .A(n5186), .ZN(n5187) );
  AOI22_X1 U6295 ( .A1(n5860), .A2(REIP_REG_19__SCAN_IN), .B1(n5187), .B2(
        n5190), .ZN(n5189) );
  NAND2_X1 U6296 ( .A1(n5958), .A2(n5308), .ZN(n5188) );
  OAI211_X1 U6297 ( .C1(n5191), .C2(n5190), .A(n5189), .B(n5188), .ZN(n5192)
         );
  AOI21_X1 U6298 ( .B1(n5379), .B2(n5946), .A(n5192), .ZN(n5193) );
  INV_X1 U6299 ( .A(n5193), .ZN(U2999) );
  NOR2_X1 U6300 ( .A1(n5194), .A2(n5200), .ZN(n5391) );
  NOR2_X1 U6301 ( .A1(n3727), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5390)
         );
  NOR2_X1 U6302 ( .A1(n5391), .A2(n5390), .ZN(n5196) );
  XOR2_X1 U6303 ( .A(n5196), .B(n5195), .Z(n5395) );
  INV_X1 U6304 ( .A(n5395), .ZN(n5205) );
  OAI21_X1 U6305 ( .B1(n5197), .B2(n5199), .A(n5885), .ZN(n5454) );
  INV_X1 U6306 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5198) );
  OAI22_X1 U6307 ( .A1(n5938), .A2(n5503), .B1(n5937), .B2(n5198), .ZN(n5203)
         );
  NAND2_X1 U6308 ( .A1(n5199), .A2(n5880), .ZN(n5461) );
  AOI221_X1 U6309 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5201), .C2(n5200), .A(n5461), 
        .ZN(n5202) );
  AOI211_X1 U6310 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5454), .A(n5203), .B(n5202), .ZN(n5204) );
  OAI21_X1 U6311 ( .B1(n5205), .B2(n5963), .A(n5204), .ZN(U3002) );
  XNOR2_X1 U6312 ( .A(n5797), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5206)
         );
  XNOR2_X1 U6313 ( .A(n5207), .B(n5206), .ZN(n5398) );
  NOR3_X1 U6314 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5209), .A3(n5208), 
        .ZN(n5215) );
  OAI21_X1 U6315 ( .B1(n5211), .B2(n5210), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5213) );
  NAND2_X1 U6316 ( .A1(n5860), .A2(REIP_REG_14__SCAN_IN), .ZN(n5212) );
  OAI211_X1 U6317 ( .C1(n5938), .C2(n5523), .A(n5213), .B(n5212), .ZN(n5214)
         );
  AOI211_X1 U6318 ( .C1(n5398), .C2(n5946), .A(n5215), .B(n5214), .ZN(n5216)
         );
  INV_X1 U6319 ( .A(n5216), .ZN(U3004) );
  XNOR2_X1 U6320 ( .A(n4634), .B(n6061), .ZN(n5218) );
  OAI22_X1 U6321 ( .A1(n5218), .A2(n6417), .B1(n5217), .B2(n4576), .ZN(n5219)
         );
  MUX2_X1 U6322 ( .A(n5219), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(n5964), 
        .Z(U3463) );
  INV_X1 U6323 ( .A(n5220), .ZN(n5222) );
  OAI22_X1 U6324 ( .A1(n5222), .A2(n6521), .B1(n5221), .B2(n6510), .ZN(n5225)
         );
  MUX2_X1 U6325 ( .A(n5225), .B(n5224), .S(n5223), .Z(U3456) );
  NAND2_X1 U6326 ( .A1(n5226), .A2(n4408), .ZN(n5229) );
  NOR2_X1 U6327 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n5231), .ZN(n5232)
         );
  AOI22_X1 U6328 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n5232), .B1(n5860), .B2(REIP_REG_30__SCAN_IN), .ZN(n5236) );
  AOI22_X1 U6329 ( .A1(n5234), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n5244), .B2(n5958), .ZN(n5235) );
  INV_X1 U6330 ( .A(n5237), .ZN(n5712) );
  AOI21_X1 U6331 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5238), .A(n5712), .ZN(
        n5239) );
  NAND2_X1 U6332 ( .A1(n5470), .A2(n5239), .ZN(U2788) );
  INV_X1 U6333 ( .A(n5339), .ZN(n5247) );
  AOI22_X1 U6334 ( .A1(EBX_REG_30__SCAN_IN), .A2(n5644), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5638), .ZN(n5240) );
  INV_X1 U6335 ( .A(n5240), .ZN(n5241) );
  AOI211_X1 U6336 ( .C1(n5336), .C2(n5626), .A(n5242), .B(n5241), .ZN(n5246)
         );
  OAI211_X1 U6337 ( .C1(n5247), .C2(n5599), .A(n5246), .B(n5245), .ZN(U2797)
         );
  INV_X1 U6338 ( .A(n5248), .ZN(n5256) );
  INV_X1 U6339 ( .A(n5249), .ZN(n5250) );
  OAI22_X1 U6340 ( .A1(n5658), .A2(n5251), .B1(n5250), .B2(n5641), .ZN(n5255)
         );
  INV_X1 U6341 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5253) );
  OAI22_X1 U6342 ( .A1(n5253), .A2(n5654), .B1(n4413), .B2(n5252), .ZN(n5254)
         );
  OAI211_X1 U6343 ( .C1(n5259), .C2(n5599), .A(n5258), .B(n5257), .ZN(U2798)
         );
  INV_X1 U6344 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5260) );
  OAI22_X1 U6345 ( .A1(n5260), .A2(n5654), .B1(n5348), .B2(n5655), .ZN(n5261)
         );
  AOI21_X1 U6346 ( .B1(EBX_REG_27__SCAN_IN), .B2(n5644), .A(n5261), .ZN(n5266)
         );
  AOI22_X1 U6347 ( .A1(n5592), .A2(n5345), .B1(n5652), .B2(n5405), .ZN(n5265)
         );
  OAI21_X1 U6348 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5263), .A(n5262), .ZN(n5264) );
  NAND3_X1 U6349 ( .A1(n5266), .A2(n5265), .A3(n5264), .ZN(U2800) );
  AOI22_X1 U6350 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5644), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5638), .ZN(n5273) );
  INV_X1 U6351 ( .A(n5358), .ZN(n5268) );
  INV_X1 U6352 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6571) );
  AOI22_X1 U6353 ( .A1(n5268), .A2(n5601), .B1(n5267), .B2(n6571), .ZN(n5272)
         );
  AOI22_X1 U6354 ( .A1(n5355), .A2(n5592), .B1(n5652), .B2(n5415), .ZN(n5271)
         );
  NOR2_X1 U6355 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5269), .ZN(n5276) );
  OAI21_X1 U6356 ( .B1(n5276), .B2(n5286), .A(REIP_REG_25__SCAN_IN), .ZN(n5270) );
  NAND4_X1 U6357 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(U2802)
         );
  AOI22_X1 U6358 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5644), .B1(n5274), .B2(n5601), .ZN(n5280) );
  AOI22_X1 U6359 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5286), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5638), .ZN(n5279) );
  AOI22_X1 U6360 ( .A1(n5324), .A2(n5592), .B1(n5652), .B2(n5275), .ZN(n5278)
         );
  INV_X1 U6361 ( .A(n5276), .ZN(n5277) );
  NAND4_X1 U6362 ( .A1(n5280), .A2(n5279), .A3(n5278), .A4(n5277), .ZN(U2803)
         );
  INV_X1 U6363 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5282) );
  OAI22_X1 U6364 ( .A1(n5282), .A2(n5658), .B1(n5281), .B2(n5655), .ZN(n5283)
         );
  AOI21_X1 U6365 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5638), .A(n5283), 
        .ZN(n5289) );
  NAND2_X1 U6366 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5284), .ZN(n5291) );
  OAI21_X1 U6367 ( .B1(n6906), .B2(n5291), .A(n6569), .ZN(n5287) );
  AOI22_X1 U6368 ( .A1(n5287), .A2(n5286), .B1(n5652), .B2(n5285), .ZN(n5288)
         );
  OAI211_X1 U6369 ( .C1(n5327), .C2(n5599), .A(n5289), .B(n5288), .ZN(U2804)
         );
  AOI22_X1 U6370 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5638), .B1(n5362), 
        .B2(n5626), .ZN(n5290) );
  OAI21_X1 U6371 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5291), .A(n5290), .ZN(n5293) );
  OAI22_X1 U6372 ( .A1(n5365), .A2(n5599), .B1(n5641), .B2(n5421), .ZN(n5292)
         );
  AOI211_X1 U6373 ( .C1(EBX_REG_22__SCAN_IN), .C2(n5644), .A(n5293), .B(n5292), 
        .ZN(n5294) );
  OAI221_X1 U6374 ( .B1(n6906), .B2(n5296), .C1(n6906), .C2(n5295), .A(n5294), 
        .ZN(U2805) );
  AOI22_X1 U6375 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5644), .B1(n5374), .B2(n5626), .ZN(n5302) );
  INV_X1 U6376 ( .A(n5296), .ZN(n5300) );
  NAND2_X1 U6377 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5307) );
  INV_X1 U6378 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6961) );
  OAI21_X1 U6379 ( .B1(n5495), .B2(n5307), .A(n6961), .ZN(n5299) );
  OAI22_X1 U6380 ( .A1(n5378), .A2(n5599), .B1(n5297), .B2(n5641), .ZN(n5298)
         );
  AOI21_X1 U6381 ( .B1(n5300), .B2(n5299), .A(n5298), .ZN(n5301) );
  OAI211_X1 U6382 ( .C1(n5303), .C2(n5654), .A(n5302), .B(n5301), .ZN(U2807)
         );
  NAND2_X1 U6383 ( .A1(n5651), .A2(n5304), .ZN(n5597) );
  INV_X1 U6384 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6746) );
  NAND2_X1 U6385 ( .A1(n5653), .A2(n5305), .ZN(n5501) );
  OAI22_X1 U6386 ( .A1(n5383), .A2(n5655), .B1(n6746), .B2(n5501), .ZN(n5306)
         );
  AOI211_X1 U6387 ( .C1(n5638), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5619), 
        .B(n5306), .ZN(n5313) );
  OAI21_X1 U6388 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5307), .ZN(n5310) );
  INV_X1 U6389 ( .A(n5308), .ZN(n5309) );
  OAI22_X1 U6390 ( .A1(n5495), .A2(n5310), .B1(n5309), .B2(n5641), .ZN(n5311)
         );
  AOI21_X1 U6391 ( .B1(n5592), .B2(n5380), .A(n5311), .ZN(n5312) );
  OAI211_X1 U6392 ( .C1(n5314), .C2(n5658), .A(n5313), .B(n5312), .ZN(U2808)
         );
  AOI22_X1 U6393 ( .A1(n5339), .A2(n5688), .B1(n5682), .B2(DATAI_30_), .ZN(
        n5316) );
  AOI22_X1 U6394 ( .A1(n5684), .A2(DATAI_14_), .B1(n5687), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6395 ( .A1(n5316), .A2(n5315), .ZN(U2861) );
  AOI22_X1 U6396 ( .A1(n5317), .A2(n5688), .B1(n5682), .B2(DATAI_29_), .ZN(
        n5319) );
  AOI22_X1 U6397 ( .A1(n5684), .A2(DATAI_13_), .B1(n5687), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6398 ( .A1(n5319), .A2(n5318), .ZN(U2862) );
  AOI22_X1 U6399 ( .A1(n5345), .A2(n5688), .B1(n5682), .B2(DATAI_27_), .ZN(
        n5321) );
  AOI22_X1 U6400 ( .A1(n5684), .A2(DATAI_11_), .B1(n5687), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6401 ( .A1(n5321), .A2(n5320), .ZN(U2864) );
  AOI22_X1 U6402 ( .A1(n5355), .A2(n5688), .B1(n5682), .B2(DATAI_25_), .ZN(
        n5323) );
  AOI22_X1 U6403 ( .A1(n5684), .A2(DATAI_9_), .B1(n5687), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6404 ( .A1(n5323), .A2(n5322), .ZN(U2866) );
  AOI22_X1 U6405 ( .A1(n5324), .A2(n5688), .B1(n5682), .B2(DATAI_24_), .ZN(
        n5326) );
  AOI22_X1 U6406 ( .A1(n5684), .A2(DATAI_8_), .B1(n5687), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6407 ( .A1(n5326), .A2(n5325), .ZN(U2867) );
  OR2_X1 U6408 ( .A1(n5327), .A2(n5677), .ZN(n5329) );
  NAND2_X1 U6409 ( .A1(n5682), .A2(DATAI_23_), .ZN(n5328) );
  AND2_X1 U6410 ( .A1(n5329), .A2(n5328), .ZN(n5331) );
  AOI22_X1 U6411 ( .A1(n5684), .A2(DATAI_7_), .B1(n5687), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6412 ( .A1(n5331), .A2(n5330), .ZN(U2868) );
  AOI22_X1 U6413 ( .A1(n5371), .A2(n5688), .B1(n5682), .B2(DATAI_21_), .ZN(
        n5333) );
  AOI22_X1 U6414 ( .A1(n5684), .A2(DATAI_5_), .B1(n5687), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6415 ( .A1(n5333), .A2(n5332), .ZN(U2870) );
  AOI22_X1 U6416 ( .A1(n5380), .A2(n5688), .B1(n5682), .B2(DATAI_19_), .ZN(
        n5335) );
  AOI22_X1 U6417 ( .A1(n5684), .A2(DATAI_3_), .B1(n5687), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6418 ( .A1(n5335), .A2(n5334), .ZN(U2872) );
  AOI22_X1 U6419 ( .A1(n5860), .A2(REIP_REG_30__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5341) );
  INV_X1 U6420 ( .A(n5336), .ZN(n5337) );
  OAI211_X1 U6421 ( .C1(n3211), .C2(n5878), .A(n5341), .B(n5340), .ZN(U2956)
         );
  AOI22_X1 U6422 ( .A1(n5860), .A2(REIP_REG_27__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5347) );
  NOR2_X1 U6423 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  XNOR2_X1 U6424 ( .A(n5344), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5406)
         );
  AOI22_X1 U6425 ( .A1(n5864), .A2(n5406), .B1(n5876), .B2(n5345), .ZN(n5346)
         );
  OAI211_X1 U6426 ( .C1(n5869), .C2(n5348), .A(n5347), .B(n5346), .ZN(U2959)
         );
  AOI22_X1 U6427 ( .A1(n5860), .A2(REIP_REG_26__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5352) );
  AOI22_X1 U6428 ( .A1(n5350), .A2(n5864), .B1(n5845), .B2(n5349), .ZN(n5351)
         );
  OAI211_X1 U6429 ( .C1(n6412), .C2(n5353), .A(n5352), .B(n5351), .ZN(U2960)
         );
  AOI22_X1 U6430 ( .A1(n5860), .A2(REIP_REG_25__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5357) );
  OAI21_X1 U6431 ( .B1(n3209), .B2(n5354), .A(n4263), .ZN(n5416) );
  AOI22_X1 U6432 ( .A1(n5355), .A2(n5876), .B1(n5864), .B2(n5416), .ZN(n5356)
         );
  OAI211_X1 U6433 ( .C1(n5869), .C2(n5358), .A(n5357), .B(n5356), .ZN(U2961)
         );
  AOI22_X1 U6434 ( .A1(n5860), .A2(REIP_REG_22__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5364) );
  AOI21_X1 U6435 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3727), .A(n5359), 
        .ZN(n5360) );
  XNOR2_X1 U6436 ( .A(n5361), .B(n5360), .ZN(n5425) );
  AOI22_X1 U6437 ( .A1(n5425), .A2(n5864), .B1(n5845), .B2(n5362), .ZN(n5363)
         );
  OAI211_X1 U6438 ( .C1(n6412), .C2(n5365), .A(n5364), .B(n5363), .ZN(U2964)
         );
  OAI22_X1 U6439 ( .A1(n5430), .A2(n5878), .B1(n5369), .B2(n5869), .ZN(n5370)
         );
  AOI21_X1 U6440 ( .B1(n5876), .B2(n5371), .A(n5370), .ZN(n5372) );
  NAND2_X1 U6441 ( .A1(n5860), .A2(REIP_REG_21__SCAN_IN), .ZN(n5433) );
  OAI211_X1 U6442 ( .C1(n5373), .C2(n5872), .A(n5372), .B(n5433), .ZN(U2965)
         );
  AOI22_X1 U6443 ( .A1(n5860), .A2(REIP_REG_20__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5377) );
  AOI22_X1 U6444 ( .A1(n5375), .A2(n5864), .B1(n5845), .B2(n5374), .ZN(n5376)
         );
  OAI211_X1 U6445 ( .C1(n6412), .C2(n5378), .A(n5377), .B(n5376), .ZN(U2966)
         );
  AOI22_X1 U6446 ( .A1(n5860), .A2(REIP_REG_19__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5382) );
  AOI22_X1 U6447 ( .A1(n5380), .A2(n5876), .B1(n5864), .B2(n5379), .ZN(n5381)
         );
  OAI211_X1 U6448 ( .C1(n5869), .C2(n5383), .A(n5382), .B(n5381), .ZN(U2967)
         );
  AOI22_X1 U6449 ( .A1(n5860), .A2(REIP_REG_18__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6450 ( .A1(n5391), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5385) );
  NAND3_X1 U6451 ( .A1(n5195), .A2(n5390), .A3(n5447), .ZN(n5384) );
  OAI21_X1 U6452 ( .B1(n5195), .B2(n5385), .A(n5384), .ZN(n5386) );
  XNOR2_X1 U6453 ( .A(n5386), .B(n5442), .ZN(n5439) );
  AOI22_X1 U6454 ( .A1(n5864), .A2(n5439), .B1(n5845), .B2(n5488), .ZN(n5387)
         );
  OAI211_X1 U6455 ( .C1(n6412), .C2(n5678), .A(n5388), .B(n5387), .ZN(U2968)
         );
  INV_X1 U6456 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5497) );
  AOI21_X1 U6457 ( .B1(n4934), .B2(n5389), .A(n5084), .ZN(n5683) );
  MUX2_X1 U6458 ( .A(n5391), .B(n5390), .S(n5195), .Z(n5392) );
  XNOR2_X1 U6459 ( .A(n5392), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5453)
         );
  OAI22_X1 U6460 ( .A1(n5453), .A2(n5878), .B1(n5869), .B2(n5496), .ZN(n5393)
         );
  AOI21_X1 U6461 ( .B1(n5876), .B2(n5683), .A(n5393), .ZN(n5394) );
  NAND2_X1 U6462 ( .A1(n5860), .A2(REIP_REG_17__SCAN_IN), .ZN(n5444) );
  OAI211_X1 U6463 ( .C1(n5497), .C2(n5872), .A(n5394), .B(n5444), .ZN(U2969)
         );
  AOI22_X1 U6464 ( .A1(n5860), .A2(REIP_REG_16__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5397) );
  AOI22_X1 U6465 ( .A1(n5395), .A2(n5864), .B1(n5845), .B2(n5508), .ZN(n5396)
         );
  OAI211_X1 U6466 ( .C1(n6412), .C2(n5514), .A(n5397), .B(n5396), .ZN(U2970)
         );
  AOI22_X1 U6467 ( .A1(n5860), .A2(REIP_REG_14__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5400) );
  AOI22_X1 U6468 ( .A1(n5398), .A2(n5864), .B1(n5845), .B2(n5527), .ZN(n5399)
         );
  OAI211_X1 U6469 ( .C1(n6412), .C2(n5531), .A(n5400), .B(n5399), .ZN(U2972)
         );
  AOI22_X1 U6470 ( .A1(n5860), .A2(REIP_REG_13__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5404) );
  INV_X1 U6471 ( .A(n5401), .ZN(n5540) );
  AOI22_X1 U6472 ( .A1(n5402), .A2(n5864), .B1(n5845), .B2(n5540), .ZN(n5403)
         );
  OAI211_X1 U6473 ( .C1(n6412), .C2(n5543), .A(n5404), .B(n5403), .ZN(U2973)
         );
  AOI22_X1 U6474 ( .A1(n5406), .A2(n5946), .B1(n5405), .B2(n5958), .ZN(n5412)
         );
  INV_X1 U6475 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6846) );
  NOR2_X1 U6476 ( .A1(n5937), .A2(n6846), .ZN(n5407) );
  AOI221_X1 U6477 ( .B1(n5410), .B2(n5409), .C1(n5408), .C2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5407), .ZN(n5411) );
  NAND2_X1 U6478 ( .A1(n5412), .A2(n5411), .ZN(U2991) );
  INV_X1 U6479 ( .A(n5413), .ZN(n5414) );
  AOI22_X1 U6480 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5860), .B1(n5414), .B2(
        n5419), .ZN(n5418) );
  AOI22_X1 U6481 ( .A1(n5416), .A2(n5946), .B1(n5958), .B2(n5415), .ZN(n5417)
         );
  OAI211_X1 U6482 ( .C1(n5420), .C2(n5419), .A(n5418), .B(n5417), .ZN(U2993)
         );
  INV_X1 U6483 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5428) );
  NOR2_X1 U6484 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5422) );
  OAI22_X1 U6485 ( .A1(n5423), .A2(n5422), .B1(n5421), .B2(n5938), .ZN(n5424)
         );
  AOI21_X1 U6486 ( .B1(n5425), .B2(n5946), .A(n5424), .ZN(n5427) );
  NAND2_X1 U6487 ( .A1(n5860), .A2(REIP_REG_22__SCAN_IN), .ZN(n5426) );
  OAI211_X1 U6488 ( .C1(n5436), .C2(n5428), .A(n5427), .B(n5426), .ZN(U2996)
         );
  OAI22_X1 U6489 ( .A1(n5430), .A2(n5963), .B1(n5938), .B2(n5429), .ZN(n5431)
         );
  AOI21_X1 U6490 ( .B1(n5432), .B2(n5435), .A(n5431), .ZN(n5434) );
  OAI211_X1 U6491 ( .C1(n5436), .C2(n5435), .A(n5434), .B(n5433), .ZN(U2997)
         );
  NOR2_X1 U6492 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5447), .ZN(n5437)
         );
  AOI22_X1 U6493 ( .A1(n5860), .A2(REIP_REG_18__SCAN_IN), .B1(n5448), .B2(
        n5437), .ZN(n5441) );
  INV_X1 U6494 ( .A(n5491), .ZN(n5438) );
  AOI22_X1 U6495 ( .A1(n5439), .A2(n5946), .B1(n5958), .B2(n5438), .ZN(n5440)
         );
  OAI211_X1 U6496 ( .C1(n5443), .C2(n5442), .A(n5441), .B(n5440), .ZN(U3000)
         );
  INV_X1 U6497 ( .A(n5444), .ZN(n5445) );
  AOI221_X1 U6498 ( .B1(n5448), .B2(n5447), .C1(n5446), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5445), .ZN(n5452) );
  AOI21_X1 U6499 ( .B1(n5450), .B2(n5449), .A(n5070), .ZN(n5665) );
  NAND2_X1 U6500 ( .A1(n5958), .A2(n5665), .ZN(n5451) );
  OAI211_X1 U6501 ( .C1(n5453), .C2(n5963), .A(n5452), .B(n5451), .ZN(U3001)
         );
  AOI22_X1 U6502 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5454), .B1(n5860), .B2(REIP_REG_15__SCAN_IN), .ZN(n5460) );
  INV_X1 U6503 ( .A(n5455), .ZN(n5458) );
  AOI21_X1 U6504 ( .B1(n5457), .B2(n4910), .A(n5456), .ZN(n5668) );
  AOI22_X1 U6505 ( .A1(n5458), .A2(n5946), .B1(n5958), .B2(n5668), .ZN(n5459)
         );
  OAI211_X1 U6506 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5461), .A(n5460), .B(n5459), .ZN(U3003) );
  INV_X1 U6507 ( .A(n5462), .ZN(n5464) );
  NAND3_X1 U6508 ( .A1(n5464), .A2(n6373), .A3(n5463), .ZN(n5465) );
  OAI21_X1 U6509 ( .B1(n5467), .B2(n5466), .A(n5465), .ZN(U3455) );
  INV_X1 U6510 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6550) );
  INV_X1 U6511 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6844) );
  AOI21_X1 U6512 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6550), .A(n6844), .ZN(n5472) );
  INV_X1 U6513 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6847) );
  AOI21_X1 U6514 ( .B1(n5472), .B2(n6847), .A(n6998), .ZN(U2789) );
  OAI21_X1 U6515 ( .B1(n5468), .B2(n6519), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5469) );
  OAI21_X1 U6516 ( .B1(n5470), .B2(n6599), .A(n5469), .ZN(U2790) );
  INV_X1 U6517 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6875) );
  NOR2_X1 U6518 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5473) );
  NOR2_X1 U6519 ( .A1(n6998), .A2(n5473), .ZN(n5471) );
  AOI22_X1 U6520 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6998), .B1(n6875), .B2(
        n5471), .ZN(U2791) );
  NOR2_X2 U6521 ( .A1(n6998), .A2(n5472), .ZN(n6583) );
  OAI21_X1 U6522 ( .B1(BS16_N), .B2(n5473), .A(n6583), .ZN(n6582) );
  OAI21_X1 U6523 ( .B1(n6583), .B2(n6596), .A(n6582), .ZN(U2792) );
  OAI21_X1 U6524 ( .B1(n5474), .B2(n6843), .A(n5878), .ZN(U2793) );
  NOR4_X1 U6525 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(n5478) );
  NOR4_X1 U6526 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5477) );
  NOR4_X1 U6527 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5476) );
  NOR4_X1 U6528 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5475) );
  NAND4_X1 U6529 ( .A1(n5478), .A2(n5477), .A3(n5476), .A4(n5475), .ZN(n5484)
         );
  NOR4_X1 U6530 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(DATAWIDTH_REG_18__SCAN_IN), .ZN(n5482)
         );
  AOI211_X1 U6531 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_23__SCAN_IN), .B(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n5481) );
  NOR4_X1 U6532 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n5480) );
  NOR4_X1 U6533 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_22__SCAN_IN), .ZN(n5479) );
  NAND4_X1 U6534 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n5483)
         );
  NOR2_X1 U6535 ( .A1(n5484), .A2(n5483), .ZN(n6593) );
  INV_X1 U6536 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6963) );
  NOR3_X1 U6537 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U6538 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5486), .A(n6593), .ZN(n5485)
         );
  OAI21_X1 U6539 ( .B1(n6593), .B2(n6963), .A(n5485), .ZN(U2794) );
  INV_X1 U6540 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6927) );
  AOI21_X1 U6541 ( .B1(n6588), .B2(n6927), .A(n5486), .ZN(n5487) );
  INV_X1 U6542 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6694) );
  INV_X1 U6543 ( .A(n6593), .ZN(n6590) );
  AOI22_X1 U6544 ( .A1(n6593), .A2(n5487), .B1(n6694), .B2(n6590), .ZN(U2795)
         );
  INV_X1 U6545 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U6546 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5644), .B1(n5488), .B2(n5626), .ZN(n5489) );
  OAI21_X1 U6547 ( .B1(n6759), .B2(n5501), .A(n5489), .ZN(n5490) );
  AOI211_X1 U6548 ( .C1(n5638), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5619), 
        .B(n5490), .ZN(n5494) );
  OAI22_X1 U6549 ( .A1(n5678), .A2(n5599), .B1(n5641), .B2(n5491), .ZN(n5492)
         );
  INV_X1 U6550 ( .A(n5492), .ZN(n5493) );
  OAI211_X1 U6551 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5495), .A(n5494), .B(n5493), .ZN(U2809) );
  AOI21_X1 U6552 ( .B1(n5505), .B2(REIP_REG_16__SCAN_IN), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5502) );
  OAI22_X1 U6553 ( .A1(n5497), .A2(n5654), .B1(n5496), .B2(n5655), .ZN(n5498)
         );
  AOI211_X1 U6554 ( .C1(n5644), .C2(EBX_REG_17__SCAN_IN), .A(n5619), .B(n5498), 
        .ZN(n5500) );
  AOI22_X1 U6555 ( .A1(n5683), .A2(n5592), .B1(n5652), .B2(n5665), .ZN(n5499)
         );
  OAI211_X1 U6556 ( .C1(n5502), .C2(n5501), .A(n5500), .B(n5499), .ZN(U2810)
         );
  NOR2_X1 U6557 ( .A1(n5503), .A2(n5641), .ZN(n5504) );
  AOI21_X1 U6558 ( .B1(n5505), .B2(n5198), .A(n5504), .ZN(n5513) );
  INV_X1 U6559 ( .A(n5653), .ZN(n5567) );
  NOR2_X1 U6560 ( .A1(n5506), .A2(n5567), .ZN(n5528) );
  NOR2_X1 U6561 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5507), .ZN(n5519) );
  AOI22_X1 U6562 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5644), .B1(n5508), .B2(n5626), .ZN(n5509) );
  OAI211_X1 U6563 ( .C1(n5654), .C2(n5510), .A(n5509), .B(n5597), .ZN(n5511)
         );
  AOI221_X1 U6564 ( .B1(n5528), .B2(REIP_REG_16__SCAN_IN), .C1(n5519), .C2(
        REIP_REG_16__SCAN_IN), .A(n5511), .ZN(n5512) );
  OAI211_X1 U6565 ( .C1(n5599), .C2(n5514), .A(n5513), .B(n5512), .ZN(U2811)
         );
  AOI22_X1 U6566 ( .A1(n5515), .A2(n5626), .B1(n5592), .B2(n5689), .ZN(n5521)
         );
  AOI22_X1 U6567 ( .A1(n5528), .A2(REIP_REG_15__SCAN_IN), .B1(n5652), .B2(
        n5668), .ZN(n5516) );
  OAI211_X1 U6568 ( .C1(n5654), .C2(n5517), .A(n5516), .B(n5597), .ZN(n5518)
         );
  AOI211_X1 U6569 ( .C1(n5644), .C2(EBX_REG_15__SCAN_IN), .A(n5519), .B(n5518), 
        .ZN(n5520) );
  NAND2_X1 U6570 ( .A1(n5521), .A2(n5520), .ZN(U2812) );
  NAND2_X1 U6571 ( .A1(n5638), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5522)
         );
  OAI211_X1 U6572 ( .C1(n5523), .C2(n5641), .A(n5522), .B(n5597), .ZN(n5524)
         );
  AOI21_X1 U6573 ( .B1(n5644), .B2(EBX_REG_14__SCAN_IN), .A(n5524), .ZN(n5525)
         );
  INV_X1 U6574 ( .A(n5525), .ZN(n5526) );
  AOI21_X1 U6575 ( .B1(n5527), .B2(n5626), .A(n5526), .ZN(n5530) );
  OAI221_X1 U6576 ( .B1(REIP_REG_14__SCAN_IN), .B2(n5537), .C1(
        REIP_REG_14__SCAN_IN), .C2(REIP_REG_13__SCAN_IN), .A(n5528), .ZN(n5529) );
  OAI211_X1 U6577 ( .C1(n5531), .C2(n5599), .A(n5530), .B(n5529), .ZN(U2813)
         );
  OAI21_X1 U6578 ( .B1(n5654), .B2(n5532), .A(n5597), .ZN(n5536) );
  OAI22_X1 U6579 ( .A1(n5658), .A2(n5534), .B1(n5533), .B2(n5641), .ZN(n5535)
         );
  AOI211_X1 U6580 ( .C1(n5537), .C2(n4926), .A(n5536), .B(n5535), .ZN(n5542)
         );
  NAND2_X1 U6581 ( .A1(n5653), .A2(n5538), .ZN(n5554) );
  OAI21_X1 U6582 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5552), .A(n5554), .ZN(n5539) );
  AOI22_X1 U6583 ( .A1(n5540), .A2(n5601), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5539), .ZN(n5541) );
  OAI211_X1 U6584 ( .C1(n5599), .C2(n5543), .A(n5542), .B(n5541), .ZN(U2814)
         );
  AOI22_X1 U6585 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5644), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5638), .ZN(n5547) );
  INV_X1 U6586 ( .A(n5544), .ZN(n5545) );
  AOI21_X1 U6587 ( .B1(n5652), .B2(n5545), .A(n5619), .ZN(n5546) );
  OAI211_X1 U6588 ( .C1(n5599), .C2(n5548), .A(n5547), .B(n5546), .ZN(n5549)
         );
  AOI21_X1 U6589 ( .B1(n5550), .B2(n5601), .A(n5549), .ZN(n5551) );
  OAI221_X1 U6590 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5552), .C1(n6562), .C2(
        n5554), .A(n5551), .ZN(U2815) );
  INV_X1 U6591 ( .A(n5576), .ZN(n5553) );
  NAND2_X1 U6592 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5568) );
  NOR2_X1 U6593 ( .A1(n5553), .A2(n5568), .ZN(n5556) );
  INV_X1 U6594 ( .A(n5554), .ZN(n5555) );
  MUX2_X1 U6595 ( .A(n5556), .B(n5555), .S(REIP_REG_11__SCAN_IN), .Z(n5560) );
  AOI22_X1 U6596 ( .A1(n5638), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5652), 
        .B2(n5879), .ZN(n5557) );
  OAI211_X1 U6597 ( .C1(n5658), .C2(n5558), .A(n5557), .B(n5597), .ZN(n5559)
         );
  AOI211_X1 U6598 ( .C1(n5800), .C2(n5626), .A(n5560), .B(n5559), .ZN(n5561)
         );
  OAI21_X1 U6599 ( .B1(n5599), .B2(n5803), .A(n5561), .ZN(U2816) );
  OAI22_X1 U6600 ( .A1(n5654), .A2(n4873), .B1(n5641), .B2(n5562), .ZN(n5563)
         );
  AOI211_X1 U6601 ( .C1(n5644), .C2(EBX_REG_10__SCAN_IN), .A(n5619), .B(n5563), 
        .ZN(n5572) );
  AOI22_X1 U6602 ( .A1(n5565), .A2(n5626), .B1(n5592), .B2(n5564), .ZN(n5571)
         );
  NOR2_X1 U6603 ( .A1(n5567), .A2(n5566), .ZN(n5583) );
  NAND2_X1 U6604 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5583), .ZN(n5570) );
  OAI211_X1 U6605 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n5576), .B(n5568), .ZN(n5569) );
  NAND4_X1 U6606 ( .A1(n5572), .A2(n5571), .A3(n5570), .A4(n5569), .ZN(U2817)
         );
  INV_X1 U6607 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6559) );
  AOI22_X1 U6608 ( .A1(n5644), .A2(EBX_REG_9__SCAN_IN), .B1(n5652), .B2(n5887), 
        .ZN(n5573) );
  OAI211_X1 U6609 ( .C1(n5654), .C2(n5574), .A(n5573), .B(n5597), .ZN(n5575)
         );
  AOI221_X1 U6610 ( .B1(n5576), .B2(n6559), .C1(n5583), .C2(
        REIP_REG_9__SCAN_IN), .A(n5575), .ZN(n5578) );
  NAND2_X1 U6611 ( .A1(n5808), .A2(n5626), .ZN(n5577) );
  OAI211_X1 U6612 ( .C1(n5811), .C2(n5599), .A(n5578), .B(n5577), .ZN(U2818)
         );
  OAI22_X1 U6613 ( .A1(n5658), .A2(n5579), .B1(n5641), .B2(n5895), .ZN(n5580)
         );
  AOI211_X1 U6614 ( .C1(n5638), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5619), 
        .B(n5580), .ZN(n5585) );
  NAND2_X1 U6615 ( .A1(n6558), .A2(n5581), .ZN(n5582) );
  AOI22_X1 U6616 ( .A1(n5816), .A2(n5601), .B1(n5583), .B2(n5582), .ZN(n5584)
         );
  OAI211_X1 U6617 ( .C1(n5599), .C2(n5819), .A(n5585), .B(n5584), .ZN(U2819)
         );
  NOR3_X1 U6618 ( .A1(n5611), .A2(REIP_REG_7__SCAN_IN), .A3(n5586), .ZN(n5591)
         );
  INV_X1 U6619 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5589) );
  INV_X1 U6620 ( .A(n5901), .ZN(n5587) );
  AOI22_X1 U6621 ( .A1(n5644), .A2(EBX_REG_7__SCAN_IN), .B1(n5652), .B2(n5587), 
        .ZN(n5588) );
  OAI211_X1 U6622 ( .C1(n5654), .C2(n5589), .A(n5588), .B(n5597), .ZN(n5590)
         );
  AOI211_X1 U6623 ( .C1(n5824), .C2(n5592), .A(n5591), .B(n5590), .ZN(n5595)
         );
  OAI21_X1 U6624 ( .B1(n5611), .B2(n5593), .A(n5651), .ZN(n5613) );
  INV_X1 U6625 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6556) );
  AND3_X1 U6626 ( .A1(n5630), .A2(n5593), .A3(n6556), .ZN(n5596) );
  OAI21_X1 U6627 ( .B1(n5613), .B2(n5596), .A(REIP_REG_7__SCAN_IN), .ZN(n5594)
         );
  OAI211_X1 U6628 ( .C1(n5655), .C2(n5827), .A(n5595), .B(n5594), .ZN(U2820)
         );
  AOI21_X1 U6629 ( .B1(n5613), .B2(REIP_REG_6__SCAN_IN), .A(n5596), .ZN(n5603)
         );
  AOI22_X1 U6630 ( .A1(n5638), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n5652), 
        .B2(n5911), .ZN(n5598) );
  OAI211_X1 U6631 ( .C1(n5599), .C2(n5834), .A(n5598), .B(n5597), .ZN(n5600)
         );
  AOI21_X1 U6632 ( .B1(n5831), .B2(n5601), .A(n5600), .ZN(n5602) );
  OAI211_X1 U6633 ( .C1(n5604), .C2(n5658), .A(n5603), .B(n5602), .ZN(U2821)
         );
  INV_X1 U6634 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5608) );
  AOI21_X1 U6635 ( .B1(n5606), .B2(n5605), .A(n4644), .ZN(n5921) );
  AOI21_X1 U6636 ( .B1(n5921), .B2(n5652), .A(n5619), .ZN(n5607) );
  OAI21_X1 U6637 ( .B1(n5608), .B2(n5654), .A(n5607), .ZN(n5609) );
  AOI21_X1 U6638 ( .B1(n5644), .B2(EBX_REG_5__SCAN_IN), .A(n5609), .ZN(n5615)
         );
  OAI21_X1 U6639 ( .B1(n5611), .B2(n5610), .A(n6555), .ZN(n5612) );
  AOI22_X1 U6640 ( .A1(n5613), .A2(n5612), .B1(n5839), .B2(n5648), .ZN(n5614)
         );
  OAI211_X1 U6641 ( .C1(n5842), .C2(n5655), .A(n5615), .B(n5614), .ZN(U2822)
         );
  OAI22_X1 U6642 ( .A1(n5617), .A2(n5654), .B1(n5616), .B2(n5656), .ZN(n5618)
         );
  AOI211_X1 U6643 ( .C1(REIP_REG_4__SCAN_IN), .C2(n5620), .A(n5619), .B(n5618), 
        .ZN(n5628) );
  INV_X1 U6644 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6554) );
  AND3_X1 U6645 ( .A1(n5630), .A2(n5621), .A3(n6554), .ZN(n5625) );
  OAI22_X1 U6646 ( .A1(n5658), .A2(n5623), .B1(n5641), .B2(n5622), .ZN(n5624)
         );
  AOI211_X1 U6647 ( .C1(n5626), .C2(n5844), .A(n5625), .B(n5624), .ZN(n5627)
         );
  OAI211_X1 U6648 ( .C1(n5664), .C2(n5849), .A(n5628), .B(n5627), .ZN(U2823)
         );
  INV_X1 U6649 ( .A(n5939), .ZN(n5629) );
  AOI22_X1 U6650 ( .A1(n5652), .A2(n5629), .B1(n5644), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5637) );
  NAND2_X1 U6651 ( .A1(n5630), .A2(REIP_REG_1__SCAN_IN), .ZN(n5632) );
  AOI21_X1 U6652 ( .B1(n6551), .B2(n5632), .A(n5631), .ZN(n5635) );
  INV_X1 U6653 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5633) );
  OAI22_X1 U6654 ( .A1(n4576), .A2(n5656), .B1(n5654), .B2(n5633), .ZN(n5634)
         );
  AOI211_X1 U6655 ( .C1(n5648), .C2(n5865), .A(n5635), .B(n5634), .ZN(n5636)
         );
  OAI211_X1 U6656 ( .C1(n5868), .C2(n5655), .A(n5637), .B(n5636), .ZN(U2825)
         );
  AND2_X1 U6657 ( .A1(n5638), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5639)
         );
  NOR2_X1 U6658 ( .A1(n5640), .A2(n5639), .ZN(n5650) );
  INV_X1 U6659 ( .A(n4528), .ZN(n5965) );
  OAI22_X1 U6660 ( .A1(n5642), .A2(n5641), .B1(n5655), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5643) );
  AOI21_X1 U6661 ( .B1(n5644), .B2(EBX_REG_1__SCAN_IN), .A(n5643), .ZN(n5645)
         );
  OAI21_X1 U6662 ( .B1(n5965), .B2(n5656), .A(n5645), .ZN(n5646) );
  AOI21_X1 U6663 ( .B1(n5648), .B2(n5647), .A(n5646), .ZN(n5649) );
  OAI211_X1 U6664 ( .C1(n5651), .C2(n6588), .A(n5650), .B(n5649), .ZN(U2826)
         );
  AOI22_X1 U6665 ( .A1(n5653), .A2(REIP_REG_0__SCAN_IN), .B1(n5652), .B2(n5959), .ZN(n5662) );
  NAND2_X1 U6666 ( .A1(n5655), .A2(n5654), .ZN(n5660) );
  OAI22_X1 U6667 ( .A1(n5658), .A2(n5657), .B1(n6482), .B2(n5656), .ZN(n5659)
         );
  AOI21_X1 U6668 ( .B1(n5660), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5659), 
        .ZN(n5661) );
  OAI211_X1 U6669 ( .C1(n5664), .C2(n5663), .A(n5662), .B(n5661), .ZN(U2827)
         );
  INV_X1 U6670 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5667) );
  AOI22_X1 U6671 ( .A1(n5683), .A2(n4472), .B1(n5671), .B2(n5665), .ZN(n5666)
         );
  OAI21_X1 U6672 ( .B1(n5674), .B2(n5667), .A(n5666), .ZN(U2842) );
  AOI22_X1 U6673 ( .A1(n5689), .A2(n4472), .B1(n5671), .B2(n5668), .ZN(n5669)
         );
  OAI21_X1 U6674 ( .B1(n5674), .B2(n5670), .A(n5669), .ZN(U2844) );
  INV_X1 U6675 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5673) );
  AOI22_X1 U6676 ( .A1(n5839), .A2(n4472), .B1(n5671), .B2(n5921), .ZN(n5672)
         );
  OAI21_X1 U6677 ( .B1(n5674), .B2(n5673), .A(n5672), .ZN(U2854) );
  INV_X1 U6678 ( .A(n5682), .ZN(n5676) );
  INV_X1 U6679 ( .A(DATAI_18_), .ZN(n5675) );
  OAI22_X1 U6680 ( .A1(n5678), .A2(n5677), .B1(n5676), .B2(n5675), .ZN(n5679)
         );
  INV_X1 U6681 ( .A(n5679), .ZN(n5681) );
  AOI22_X1 U6682 ( .A1(n5684), .A2(DATAI_2_), .B1(n5687), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U6683 ( .A1(n5681), .A2(n5680), .ZN(U2873) );
  AOI22_X1 U6684 ( .A1(n5683), .A2(n5688), .B1(n5682), .B2(DATAI_17_), .ZN(
        n5686) );
  AOI22_X1 U6685 ( .A1(n5684), .A2(DATAI_1_), .B1(n5687), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U6686 ( .A1(n5686), .A2(n5685), .ZN(U2874) );
  INV_X1 U6687 ( .A(DATAI_15_), .ZN(n6698) );
  AOI22_X1 U6688 ( .A1(n5689), .A2(n5688), .B1(n5687), .B2(EAX_REG_15__SCAN_IN), .ZN(n5690) );
  OAI21_X1 U6689 ( .B1(n5691), .B2(n6698), .A(n5690), .ZN(U2876) );
  INV_X1 U6690 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5794) );
  AOI22_X1 U6691 ( .A1(n4833), .A2(LWORD_REG_15__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5693) );
  OAI21_X1 U6692 ( .B1(n5794), .B2(n5711), .A(n5693), .ZN(U2908) );
  AOI22_X1 U6693 ( .A1(n4833), .A2(LWORD_REG_14__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5694) );
  OAI21_X1 U6694 ( .B1(n5789), .B2(n5711), .A(n5694), .ZN(U2909) );
  AOI22_X1 U6695 ( .A1(n4833), .A2(LWORD_REG_13__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5695) );
  OAI21_X1 U6696 ( .B1(n5786), .B2(n5711), .A(n5695), .ZN(U2910) );
  AOI22_X1 U6697 ( .A1(n4833), .A2(LWORD_REG_12__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5696) );
  OAI21_X1 U6698 ( .B1(n5783), .B2(n5711), .A(n5696), .ZN(U2911) );
  AOI22_X1 U6699 ( .A1(n4833), .A2(LWORD_REG_11__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5697) );
  OAI21_X1 U6700 ( .B1(n5780), .B2(n5711), .A(n5697), .ZN(U2912) );
  AOI22_X1 U6701 ( .A1(n4833), .A2(LWORD_REG_10__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5698) );
  OAI21_X1 U6702 ( .B1(n5777), .B2(n5711), .A(n5698), .ZN(U2913) );
  AOI22_X1 U6703 ( .A1(n4833), .A2(LWORD_REG_9__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5699) );
  OAI21_X1 U6704 ( .B1(n5774), .B2(n5711), .A(n5699), .ZN(U2914) );
  AOI22_X1 U6705 ( .A1(n4833), .A2(LWORD_REG_8__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5700) );
  OAI21_X1 U6706 ( .B1(n5771), .B2(n5711), .A(n5700), .ZN(U2915) );
  AOI22_X1 U6707 ( .A1(n4833), .A2(LWORD_REG_7__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5701) );
  OAI21_X1 U6708 ( .B1(n5768), .B2(n5711), .A(n5701), .ZN(U2916) );
  AOI22_X1 U6709 ( .A1(n4833), .A2(LWORD_REG_6__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5702) );
  OAI21_X1 U6710 ( .B1(n5765), .B2(n5711), .A(n5702), .ZN(U2917) );
  AOI22_X1 U6711 ( .A1(n4833), .A2(LWORD_REG_5__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5703) );
  OAI21_X1 U6712 ( .B1(n5762), .B2(n5711), .A(n5703), .ZN(U2918) );
  AOI22_X1 U6713 ( .A1(n4833), .A2(LWORD_REG_4__SCAN_IN), .B1(n5704), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5705) );
  OAI21_X1 U6714 ( .B1(n5759), .B2(n5711), .A(n5705), .ZN(U2919) );
  AOI22_X1 U6715 ( .A1(n4833), .A2(LWORD_REG_3__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5706) );
  OAI21_X1 U6716 ( .B1(n5756), .B2(n5711), .A(n5706), .ZN(U2920) );
  AOI22_X1 U6717 ( .A1(n4833), .A2(LWORD_REG_2__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5707) );
  OAI21_X1 U6718 ( .B1(n5753), .B2(n5711), .A(n5707), .ZN(U2921) );
  AOI22_X1 U6719 ( .A1(n4833), .A2(LWORD_REG_1__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5708) );
  OAI21_X1 U6720 ( .B1(n5750), .B2(n5711), .A(n5708), .ZN(U2922) );
  AOI22_X1 U6721 ( .A1(n4833), .A2(LWORD_REG_0__SCAN_IN), .B1(n5709), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5710) );
  OAI21_X1 U6722 ( .B1(n5747), .B2(n5711), .A(n5710), .ZN(U2923) );
  AND2_X1 U6723 ( .A1(n5790), .A2(DATAI_0_), .ZN(n5745) );
  AOI21_X1 U6724 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n5791), .A(n5745), .ZN(n5714) );
  OAI21_X1 U6725 ( .B1(n5715), .B2(n5793), .A(n5714), .ZN(U2924) );
  AND2_X1 U6726 ( .A1(n5790), .A2(DATAI_1_), .ZN(n5748) );
  AOI21_X1 U6727 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n5791), .A(n5748), .ZN(n5716) );
  OAI21_X1 U6728 ( .B1(n5717), .B2(n5793), .A(n5716), .ZN(U2925) );
  AND2_X1 U6729 ( .A1(n5790), .A2(DATAI_2_), .ZN(n5751) );
  AOI21_X1 U6730 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n5791), .A(n5751), .ZN(n5718) );
  OAI21_X1 U6731 ( .B1(n5719), .B2(n5793), .A(n5718), .ZN(U2926) );
  AND2_X1 U6732 ( .A1(n5790), .A2(DATAI_3_), .ZN(n5754) );
  AOI21_X1 U6733 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n5791), .A(n5754), .ZN(n5720) );
  OAI21_X1 U6734 ( .B1(n5721), .B2(n5793), .A(n5720), .ZN(U2927) );
  AND2_X1 U6735 ( .A1(n5790), .A2(DATAI_4_), .ZN(n5757) );
  AOI21_X1 U6736 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n5791), .A(n5757), .ZN(n5722) );
  OAI21_X1 U6737 ( .B1(n5723), .B2(n5793), .A(n5722), .ZN(U2928) );
  AND2_X1 U6738 ( .A1(n5790), .A2(DATAI_5_), .ZN(n5760) );
  AOI21_X1 U6739 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n5791), .A(n5760), .ZN(n5724) );
  OAI21_X1 U6740 ( .B1(n5725), .B2(n5793), .A(n5724), .ZN(U2929) );
  AND2_X1 U6741 ( .A1(n5790), .A2(DATAI_6_), .ZN(n5763) );
  AOI21_X1 U6742 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n5791), .A(n5763), .ZN(n5726) );
  OAI21_X1 U6743 ( .B1(n5727), .B2(n5793), .A(n5726), .ZN(U2930) );
  AND2_X1 U6744 ( .A1(n5790), .A2(DATAI_7_), .ZN(n5766) );
  AOI21_X1 U6745 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n5791), .A(n5766), .ZN(n5728) );
  OAI21_X1 U6746 ( .B1(n5729), .B2(n5793), .A(n5728), .ZN(U2931) );
  AND2_X1 U6747 ( .A1(n5790), .A2(DATAI_8_), .ZN(n5769) );
  AOI21_X1 U6748 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n5791), .A(n5769), .ZN(n5730) );
  OAI21_X1 U6749 ( .B1(n5731), .B2(n5793), .A(n5730), .ZN(U2932) );
  AND2_X1 U6750 ( .A1(n5790), .A2(DATAI_9_), .ZN(n5772) );
  AOI21_X1 U6751 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n5740), .A(n5772), .ZN(n5732) );
  OAI21_X1 U6752 ( .B1(n5733), .B2(n5793), .A(n5732), .ZN(U2933) );
  AND2_X1 U6753 ( .A1(n5790), .A2(DATAI_10_), .ZN(n5775) );
  AOI21_X1 U6754 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n5740), .A(n5775), .ZN(
        n5734) );
  OAI21_X1 U6755 ( .B1(n5735), .B2(n5793), .A(n5734), .ZN(U2934) );
  AND2_X1 U6756 ( .A1(n5790), .A2(DATAI_11_), .ZN(n5778) );
  AOI21_X1 U6757 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n5740), .A(n5778), .ZN(
        n5736) );
  OAI21_X1 U6758 ( .B1(n5737), .B2(n5793), .A(n5736), .ZN(U2935) );
  AND2_X1 U6759 ( .A1(n5790), .A2(DATAI_12_), .ZN(n5781) );
  AOI21_X1 U6760 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n5740), .A(n5781), .ZN(
        n5738) );
  OAI21_X1 U6761 ( .B1(n5739), .B2(n5793), .A(n5738), .ZN(U2936) );
  AND2_X1 U6762 ( .A1(n5790), .A2(DATAI_13_), .ZN(n5784) );
  AOI21_X1 U6763 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n5740), .A(n5784), .ZN(
        n5741) );
  OAI21_X1 U6764 ( .B1(n5742), .B2(n5793), .A(n5741), .ZN(U2937) );
  AND2_X1 U6765 ( .A1(n5790), .A2(DATAI_14_), .ZN(n5787) );
  AOI21_X1 U6766 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n5791), .A(n5787), .ZN(
        n5743) );
  OAI21_X1 U6767 ( .B1(n5744), .B2(n5793), .A(n5743), .ZN(U2938) );
  AOI21_X1 U6768 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n5791), .A(n5745), .ZN(n5746) );
  OAI21_X1 U6769 ( .B1(n5747), .B2(n5793), .A(n5746), .ZN(U2939) );
  AOI21_X1 U6770 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n5791), .A(n5748), .ZN(n5749) );
  OAI21_X1 U6771 ( .B1(n5750), .B2(n5793), .A(n5749), .ZN(U2940) );
  AOI21_X1 U6772 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n5791), .A(n5751), .ZN(n5752) );
  OAI21_X1 U6773 ( .B1(n5753), .B2(n5793), .A(n5752), .ZN(U2941) );
  AOI21_X1 U6774 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n5791), .A(n5754), .ZN(n5755) );
  OAI21_X1 U6775 ( .B1(n5756), .B2(n5793), .A(n5755), .ZN(U2942) );
  AOI21_X1 U6776 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n5791), .A(n5757), .ZN(n5758) );
  OAI21_X1 U6777 ( .B1(n5759), .B2(n5793), .A(n5758), .ZN(U2943) );
  AOI21_X1 U6778 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n5791), .A(n5760), .ZN(n5761) );
  OAI21_X1 U6779 ( .B1(n5762), .B2(n5793), .A(n5761), .ZN(U2944) );
  AOI21_X1 U6780 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n5791), .A(n5763), .ZN(n5764) );
  OAI21_X1 U6781 ( .B1(n5765), .B2(n5793), .A(n5764), .ZN(U2945) );
  AOI21_X1 U6782 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n5791), .A(n5766), .ZN(n5767) );
  OAI21_X1 U6783 ( .B1(n5768), .B2(n5793), .A(n5767), .ZN(U2946) );
  AOI21_X1 U6784 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n5791), .A(n5769), .ZN(n5770) );
  OAI21_X1 U6785 ( .B1(n5771), .B2(n5793), .A(n5770), .ZN(U2947) );
  AOI21_X1 U6786 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n5791), .A(n5772), .ZN(n5773) );
  OAI21_X1 U6787 ( .B1(n5774), .B2(n5793), .A(n5773), .ZN(U2948) );
  AOI21_X1 U6788 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n5791), .A(n5775), .ZN(
        n5776) );
  OAI21_X1 U6789 ( .B1(n5777), .B2(n5793), .A(n5776), .ZN(U2949) );
  AOI21_X1 U6790 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n5791), .A(n5778), .ZN(
        n5779) );
  OAI21_X1 U6791 ( .B1(n5780), .B2(n5793), .A(n5779), .ZN(U2950) );
  AOI21_X1 U6792 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n5791), .A(n5781), .ZN(
        n5782) );
  OAI21_X1 U6793 ( .B1(n5783), .B2(n5793), .A(n5782), .ZN(U2951) );
  AOI21_X1 U6794 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n5791), .A(n5784), .ZN(
        n5785) );
  OAI21_X1 U6795 ( .B1(n5786), .B2(n5793), .A(n5785), .ZN(U2952) );
  AOI21_X1 U6796 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n5791), .A(n5787), .ZN(
        n5788) );
  OAI21_X1 U6797 ( .B1(n5789), .B2(n5793), .A(n5788), .ZN(U2953) );
  AOI22_X1 U6798 ( .A1(n5791), .A2(LWORD_REG_15__SCAN_IN), .B1(n5790), .B2(
        DATAI_15_), .ZN(n5792) );
  OAI21_X1 U6799 ( .B1(n5794), .B2(n5793), .A(n5792), .ZN(U2954) );
  AOI22_X1 U6800 ( .A1(n5860), .A2(REIP_REG_11__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U6801 ( .A1(n5796), .A2(n5795), .ZN(n5799) );
  XNOR2_X1 U6802 ( .A(n5797), .B(n5884), .ZN(n5798) );
  XNOR2_X1 U6803 ( .A(n5799), .B(n5798), .ZN(n5881) );
  AOI22_X1 U6804 ( .A1(n5864), .A2(n5881), .B1(n5845), .B2(n5800), .ZN(n5801)
         );
  OAI211_X1 U6805 ( .C1(n6412), .C2(n5803), .A(n5802), .B(n5801), .ZN(U2975)
         );
  AOI22_X1 U6806 ( .A1(n5860), .A2(REIP_REG_9__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6807 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  XNOR2_X1 U6808 ( .A(n5807), .B(n5806), .ZN(n5889) );
  AOI22_X1 U6809 ( .A1(n5889), .A2(n5864), .B1(n5845), .B2(n5808), .ZN(n5809)
         );
  OAI211_X1 U6810 ( .C1(n6412), .C2(n5811), .A(n5810), .B(n5809), .ZN(U2977)
         );
  AOI22_X1 U6811 ( .A1(n5860), .A2(REIP_REG_8__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U6812 ( .B1(n3179), .B2(n5813), .A(n5812), .ZN(n5815) );
  INV_X1 U6813 ( .A(n5815), .ZN(n5898) );
  AOI22_X1 U6814 ( .A1(n5898), .A2(n5864), .B1(n5845), .B2(n5816), .ZN(n5817)
         );
  OAI211_X1 U6815 ( .C1(n6412), .C2(n5819), .A(n5818), .B(n5817), .ZN(U2978)
         );
  AOI22_X1 U6816 ( .A1(n5860), .A2(REIP_REG_7__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5826) );
  OAI21_X1 U6817 ( .B1(n5822), .B2(n5821), .A(n5820), .ZN(n5823) );
  INV_X1 U6818 ( .A(n5823), .ZN(n5903) );
  AOI22_X1 U6819 ( .A1(n5824), .A2(n5876), .B1(n5864), .B2(n5903), .ZN(n5825)
         );
  OAI211_X1 U6820 ( .C1(n5869), .C2(n5827), .A(n5826), .B(n5825), .ZN(U2979)
         );
  AOI22_X1 U6821 ( .A1(n5860), .A2(REIP_REG_6__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5833) );
  OAI21_X1 U6822 ( .B1(n3165), .B2(n5829), .A(n5828), .ZN(n5830) );
  INV_X1 U6823 ( .A(n5830), .ZN(n5914) );
  AOI22_X1 U6824 ( .A1(n5914), .A2(n5864), .B1(n5845), .B2(n5831), .ZN(n5832)
         );
  OAI211_X1 U6825 ( .C1(n6412), .C2(n5834), .A(n5833), .B(n5832), .ZN(U2980)
         );
  AOI22_X1 U6826 ( .A1(n5860), .A2(REIP_REG_5__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5841) );
  OR2_X1 U6827 ( .A1(n5836), .A2(n5835), .ZN(n5837) );
  AND2_X1 U6828 ( .A1(n5838), .A2(n5837), .ZN(n5922) );
  AOI22_X1 U6829 ( .A1(n5839), .A2(n5876), .B1(n5864), .B2(n5922), .ZN(n5840)
         );
  OAI211_X1 U6830 ( .C1(n5869), .C2(n5842), .A(n5841), .B(n5840), .ZN(U2981)
         );
  AOI22_X1 U6831 ( .A1(n5860), .A2(REIP_REG_4__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5848) );
  INV_X1 U6832 ( .A(n5843), .ZN(n5846) );
  AOI22_X1 U6833 ( .A1(n5846), .A2(n5864), .B1(n5845), .B2(n5844), .ZN(n5847)
         );
  OAI211_X1 U6834 ( .C1(n6412), .C2(n5849), .A(n5848), .B(n5847), .ZN(U2982)
         );
  AOI22_X1 U6835 ( .A1(n5860), .A2(REIP_REG_3__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5857) );
  OAI21_X1 U6836 ( .B1(n5852), .B2(n5851), .A(n5850), .ZN(n5853) );
  INV_X1 U6837 ( .A(n5853), .ZN(n5930) );
  INV_X1 U6838 ( .A(n5854), .ZN(n5855) );
  AOI22_X1 U6839 ( .A1(n5864), .A2(n5930), .B1(n5855), .B2(n5876), .ZN(n5856)
         );
  OAI211_X1 U6840 ( .C1(n5869), .C2(n5858), .A(n5857), .B(n5856), .ZN(U2983)
         );
  AOI22_X1 U6841 ( .A1(n5860), .A2(REIP_REG_2__SCAN_IN), .B1(n5859), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5867) );
  XNOR2_X1 U6842 ( .A(n5861), .B(n5936), .ZN(n5862) );
  XNOR2_X1 U6843 ( .A(n5863), .B(n5862), .ZN(n5945) );
  AOI22_X1 U6844 ( .A1(n5865), .A2(n5876), .B1(n5945), .B2(n5864), .ZN(n5866)
         );
  OAI211_X1 U6845 ( .C1(n5869), .C2(n5868), .A(n5867), .B(n5866), .ZN(U2984)
         );
  OAI21_X1 U6846 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5871), .A(n5870), 
        .ZN(n5962) );
  NAND2_X1 U6847 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AOI22_X1 U6848 ( .A1(n5876), .A2(n5875), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5874), .ZN(n5877) );
  NAND2_X1 U6849 ( .A1(n5860), .A2(REIP_REG_0__SCAN_IN), .ZN(n5952) );
  OAI211_X1 U6850 ( .C1(n5878), .C2(n5962), .A(n5877), .B(n5952), .ZN(U2986)
         );
  AOI22_X1 U6851 ( .A1(n5958), .A2(n5879), .B1(n5860), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5883) );
  AOI22_X1 U6852 ( .A1(n5946), .A2(n5881), .B1(n5884), .B2(n5880), .ZN(n5882)
         );
  OAI211_X1 U6853 ( .C1(n5885), .C2(n5884), .A(n5883), .B(n5882), .ZN(U3007)
         );
  INV_X1 U6854 ( .A(n5886), .ZN(n5893) );
  AOI22_X1 U6855 ( .A1(n5958), .A2(n5887), .B1(n5860), .B2(REIP_REG_9__SCAN_IN), .ZN(n5891) );
  AOI22_X1 U6856 ( .A1(n5889), .A2(n5946), .B1(n5888), .B2(n5892), .ZN(n5890)
         );
  OAI211_X1 U6857 ( .C1(n5893), .C2(n5892), .A(n5891), .B(n5890), .ZN(U3009)
         );
  AOI211_X1 U6858 ( .C1(n5906), .C2(n5900), .A(n5894), .B(n5907), .ZN(n5897)
         );
  OAI22_X1 U6859 ( .A1(n5938), .A2(n5895), .B1(n6558), .B2(n5937), .ZN(n5896)
         );
  AOI211_X1 U6860 ( .C1(n5898), .C2(n5946), .A(n5897), .B(n5896), .ZN(n5899)
         );
  OAI21_X1 U6861 ( .B1(n5905), .B2(n5900), .A(n5899), .ZN(U3010) );
  OAI22_X1 U6862 ( .A1(n5938), .A2(n5901), .B1(n6557), .B2(n5937), .ZN(n5902)
         );
  AOI21_X1 U6863 ( .B1(n5903), .B2(n5946), .A(n5902), .ZN(n5904) );
  OAI221_X1 U6864 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5907), .C1(n5906), .C2(n5905), .A(n5904), .ZN(U3011) );
  OR2_X1 U6865 ( .A1(n5912), .A2(n5919), .ZN(n5909) );
  AOI21_X1 U6866 ( .B1(n5910), .B2(n5909), .A(n5908), .ZN(n5926) );
  AOI22_X1 U6867 ( .A1(n5958), .A2(n5911), .B1(n5860), .B2(REIP_REG_6__SCAN_IN), .ZN(n5916) );
  NOR3_X1 U6868 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5912), .A3(n5919), 
        .ZN(n5913) );
  AOI22_X1 U6869 ( .A1(n5914), .A2(n5946), .B1(n5913), .B2(n5929), .ZN(n5915)
         );
  OAI211_X1 U6870 ( .C1(n5926), .C2(n5917), .A(n5916), .B(n5915), .ZN(U3012)
         );
  OAI22_X1 U6871 ( .A1(n5944), .A2(n5919), .B1(n5918), .B2(n5951), .ZN(n5920)
         );
  NOR2_X1 U6872 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5920), .ZN(n5925)
         );
  AOI22_X1 U6873 ( .A1(n5922), .A2(n5946), .B1(n5958), .B2(n5921), .ZN(n5924)
         );
  NAND2_X1 U6874 ( .A1(n5860), .A2(REIP_REG_5__SCAN_IN), .ZN(n5923) );
  OAI211_X1 U6875 ( .C1(n5926), .C2(n5925), .A(n5924), .B(n5923), .ZN(U3013)
         );
  AOI22_X1 U6876 ( .A1(n5958), .A2(n5927), .B1(n5860), .B2(REIP_REG_3__SCAN_IN), .ZN(n5933) );
  AND2_X1 U6877 ( .A1(n5929), .A2(n5928), .ZN(n5931) );
  AOI22_X1 U6878 ( .A1(n5931), .A2(n5934), .B1(n5930), .B2(n5946), .ZN(n5932)
         );
  OAI211_X1 U6879 ( .C1(n5935), .C2(n5934), .A(n5933), .B(n5932), .ZN(U3015)
         );
  NAND2_X1 U6880 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5936), .ZN(n5950)
         );
  OAI22_X1 U6881 ( .A1(n5939), .A2(n5938), .B1(n6551), .B2(n5937), .ZN(n5940)
         );
  NOR2_X1 U6882 ( .A1(n5941), .A2(n5940), .ZN(n5949) );
  OAI21_X1 U6883 ( .B1(n5944), .B2(n5943), .A(n5942), .ZN(n5947) );
  AOI22_X1 U6884 ( .A1(n5947), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n5946), 
        .B2(n5945), .ZN(n5948) );
  OAI211_X1 U6885 ( .C1(n5951), .C2(n5950), .A(n5949), .B(n5948), .ZN(U3016)
         );
  INV_X1 U6886 ( .A(n5952), .ZN(n5957) );
  AOI21_X1 U6887 ( .B1(n5955), .B2(n5954), .A(n5953), .ZN(n5956) );
  AOI211_X1 U6888 ( .C1(n5959), .C2(n5958), .A(n5957), .B(n5956), .ZN(n5961)
         );
  OAI211_X1 U6889 ( .C1(n5963), .C2(n5962), .A(n5961), .B(n5960), .ZN(U3018)
         );
  AND2_X1 U6890 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5964), .ZN(U3019)
         );
  NAND3_X1 U6891 ( .A1(n6493), .A2(n6209), .A3(n6487), .ZN(n6002) );
  NOR2_X1 U6892 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6002), .ZN(n5992)
         );
  AND2_X1 U6893 ( .A1(n5965), .A2(n4576), .ZN(n6177) );
  NAND2_X1 U6894 ( .A1(n6029), .A2(n6177), .ZN(n5998) );
  OR2_X1 U6895 ( .A1(n5998), .A2(n6417), .ZN(n5968) );
  NAND2_X1 U6896 ( .A1(n5966), .A2(n6368), .ZN(n5967) );
  AND2_X1 U6897 ( .A1(n5968), .A2(n5967), .ZN(n5982) );
  AOI22_X1 U6898 ( .A1(n6410), .A2(n5992), .B1(n6409), .B2(n5991), .ZN(n5975)
         );
  INV_X1 U6899 ( .A(n5992), .ZN(n5983) );
  AOI211_X1 U6900 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5983), .A(n6365), .B(
        n5969), .ZN(n5973) );
  NOR2_X1 U6901 ( .A1(n4634), .A2(n3155), .ZN(n5970) );
  NAND2_X1 U6902 ( .A1(n5996), .A2(n6282), .ZN(n6022) );
  INV_X1 U6903 ( .A(n6459), .ZN(n6471) );
  NOR3_X1 U6904 ( .A1(n6024), .A2(n6471), .A3(n6417), .ZN(n5971) );
  OAI21_X1 U6905 ( .B1(n5971), .B2(n6414), .A(n5998), .ZN(n5972) );
  NAND2_X1 U6906 ( .A1(n5973), .A2(n5972), .ZN(n5993) );
  AOI22_X1 U6907 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5993), .B1(n6331), 
        .B2(n6024), .ZN(n5974) );
  OAI211_X1 U6908 ( .C1(n6334), .C2(n6459), .A(n5975), .B(n5974), .ZN(U3020)
         );
  AOI22_X1 U6909 ( .A1(n6427), .A2(n5992), .B1(n6426), .B2(n5991), .ZN(n5977)
         );
  AOI22_X1 U6910 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5993), .B1(n6335), 
        .B2(n6024), .ZN(n5976) );
  OAI211_X1 U6911 ( .C1(n6338), .C2(n6459), .A(n5977), .B(n5976), .ZN(U3021)
         );
  AOI22_X1 U6912 ( .A1(n6433), .A2(n5992), .B1(n6432), .B2(n5991), .ZN(n5979)
         );
  AOI22_X1 U6913 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5993), .B1(n6259), 
        .B2(n6024), .ZN(n5978) );
  OAI211_X1 U6914 ( .C1(n6262), .C2(n6459), .A(n5979), .B(n5978), .ZN(U3022)
         );
  AOI22_X1 U6915 ( .A1(n6439), .A2(n5992), .B1(n6438), .B2(n5991), .ZN(n5981)
         );
  AOI22_X1 U6916 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5993), .B1(n6224), 
        .B2(n6024), .ZN(n5980) );
  OAI211_X1 U6917 ( .C1(n6227), .C2(n6459), .A(n5981), .B(n5980), .ZN(U3023)
         );
  OAI22_X1 U6918 ( .A1(n6447), .A2(n5983), .B1(n5982), .B2(n6444), .ZN(n5984)
         );
  INV_X1 U6919 ( .A(n5984), .ZN(n5986) );
  AOI22_X1 U6920 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5993), .B1(n6449), 
        .B2(n6024), .ZN(n5985) );
  OAI211_X1 U6921 ( .C1(n6452), .C2(n6459), .A(n5986), .B(n5985), .ZN(U3024)
         );
  AOI22_X1 U6922 ( .A1(n6454), .A2(n5992), .B1(n6453), .B2(n5991), .ZN(n5988)
         );
  AOI22_X1 U6923 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5993), .B1(n6348), 
        .B2(n6024), .ZN(n5987) );
  OAI211_X1 U6924 ( .C1(n6352), .C2(n6459), .A(n5988), .B(n5987), .ZN(U3025)
         );
  AOI22_X1 U6925 ( .A1(n6462), .A2(n5992), .B1(n6461), .B2(n5991), .ZN(n5990)
         );
  AOI22_X1 U6926 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5993), .B1(n6463), 
        .B2(n6024), .ZN(n5989) );
  OAI211_X1 U6927 ( .C1(n6466), .C2(n6459), .A(n5990), .B(n5989), .ZN(U3026)
         );
  AOI22_X1 U6928 ( .A1(n6470), .A2(n5992), .B1(n6468), .B2(n5991), .ZN(n5995)
         );
  AOI22_X1 U6929 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5993), .B1(n6472), 
        .B2(n6024), .ZN(n5994) );
  OAI211_X1 U6930 ( .C1(n6477), .C2(n6459), .A(n5995), .B(n5994), .ZN(U3027)
         );
  NOR2_X1 U6931 ( .A1(n6283), .A2(n6002), .ZN(n6023) );
  AOI22_X1 U6932 ( .A1(n6035), .A2(n6331), .B1(n6410), .B2(n6023), .ZN(n6006)
         );
  INV_X1 U6933 ( .A(n5996), .ZN(n5997) );
  OAI21_X1 U6934 ( .B1(n5997), .B2(n6596), .A(n6603), .ZN(n6004) );
  OR2_X1 U6935 ( .A1(n5998), .A2(n6482), .ZN(n5999) );
  INV_X1 U6936 ( .A(n6023), .ZN(n6013) );
  AND2_X1 U6937 ( .A1(n5999), .A2(n6013), .ZN(n6003) );
  INV_X1 U6938 ( .A(n6003), .ZN(n6001) );
  AOI21_X1 U6939 ( .B1(n6417), .B2(n6002), .A(n6416), .ZN(n6000) );
  OAI21_X1 U6940 ( .B1(n6004), .B2(n6001), .A(n6000), .ZN(n6026) );
  OAI22_X1 U6941 ( .A1(n6004), .A2(n6003), .B1(n6251), .B2(n6002), .ZN(n6025)
         );
  AOI22_X1 U6942 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6026), .B1(n6409), 
        .B2(n6025), .ZN(n6005) );
  OAI211_X1 U6943 ( .C1(n6334), .C2(n6022), .A(n6006), .B(n6005), .ZN(U3028)
         );
  AOI22_X1 U6944 ( .A1(n6035), .A2(n6335), .B1(n6427), .B2(n6023), .ZN(n6008)
         );
  AOI22_X1 U6945 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6026), .B1(n6426), 
        .B2(n6025), .ZN(n6007) );
  OAI211_X1 U6946 ( .C1(n6338), .C2(n6022), .A(n6008), .B(n6007), .ZN(U3029)
         );
  AOI22_X1 U6947 ( .A1(n6024), .A2(n6434), .B1(n6433), .B2(n6023), .ZN(n6010)
         );
  AOI22_X1 U6948 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6026), .B1(n6432), 
        .B2(n6025), .ZN(n6009) );
  OAI211_X1 U6949 ( .C1(n6060), .C2(n6437), .A(n6010), .B(n6009), .ZN(U3030)
         );
  AOI22_X1 U6950 ( .A1(n6024), .A2(n6440), .B1(n6439), .B2(n6023), .ZN(n6012)
         );
  AOI22_X1 U6951 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6026), .B1(n6438), 
        .B2(n6025), .ZN(n6011) );
  OAI211_X1 U6952 ( .C1(n6060), .C2(n6443), .A(n6012), .B(n6011), .ZN(U3031)
         );
  OR2_X1 U6953 ( .A1(n6447), .A2(n6013), .ZN(n6014) );
  OAI21_X1 U6954 ( .B1(n6060), .B2(n6266), .A(n6014), .ZN(n6015) );
  INV_X1 U6955 ( .A(n6015), .ZN(n6017) );
  AOI22_X1 U6956 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6026), .B1(n6269), 
        .B2(n6025), .ZN(n6016) );
  OAI211_X1 U6957 ( .C1(n6452), .C2(n6022), .A(n6017), .B(n6016), .ZN(U3032)
         );
  AOI22_X1 U6958 ( .A1(n6035), .A2(n6348), .B1(n6454), .B2(n6023), .ZN(n6019)
         );
  AOI22_X1 U6959 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6026), .B1(n6453), 
        .B2(n6025), .ZN(n6018) );
  OAI211_X1 U6960 ( .C1(n6352), .C2(n6022), .A(n6019), .B(n6018), .ZN(U3033)
         );
  AOI22_X1 U6961 ( .A1(n6035), .A2(n6463), .B1(n6462), .B2(n6023), .ZN(n6021)
         );
  AOI22_X1 U6962 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6026), .B1(n6461), 
        .B2(n6025), .ZN(n6020) );
  OAI211_X1 U6963 ( .C1(n6466), .C2(n6022), .A(n6021), .B(n6020), .ZN(U3034)
         );
  AOI22_X1 U6964 ( .A1(n6024), .A2(n6397), .B1(n6470), .B2(n6023), .ZN(n6028)
         );
  AOI22_X1 U6965 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6026), .B1(n6468), 
        .B2(n6025), .ZN(n6027) );
  OAI211_X1 U6966 ( .C1(n6060), .C2(n6401), .A(n6028), .B(n6027), .ZN(U3035)
         );
  NAND3_X1 U6967 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6493), .A3(n6209), .ZN(n6069) );
  NOR2_X1 U6968 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6069), .ZN(n6056)
         );
  AND2_X1 U6969 ( .A1(n4576), .A2(n4528), .ZN(n6212) );
  NAND2_X1 U6970 ( .A1(n6029), .A2(n6212), .ZN(n6065) );
  OR2_X1 U6971 ( .A1(n6065), .A2(n6417), .ZN(n6031) );
  NAND3_X1 U6972 ( .A1(n6368), .A2(n6364), .A3(n6493), .ZN(n6030) );
  AND2_X1 U6973 ( .A1(n6031), .A2(n6030), .ZN(n6046) );
  INV_X1 U6974 ( .A(n6046), .ZN(n6055) );
  AOI22_X1 U6975 ( .A1(n6410), .A2(n6056), .B1(n6409), .B2(n6055), .ZN(n6039)
         );
  INV_X1 U6976 ( .A(n6210), .ZN(n6361) );
  NOR2_X1 U6977 ( .A1(n6361), .A2(n4634), .ZN(n6032) );
  OAI21_X1 U6978 ( .B1(n6035), .B2(n6086), .A(n6034), .ZN(n6036) );
  NAND2_X1 U6979 ( .A1(n6036), .A2(n6065), .ZN(n6037) );
  NOR2_X1 U6980 ( .A1(n6365), .A2(n6369), .ZN(n6214) );
  OAI221_X1 U6981 ( .B1(n6056), .B2(n6373), .C1(n6056), .C2(n6037), .A(n6214), 
        .ZN(n6057) );
  AOI22_X1 U6982 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n6057), .B1(n6331), 
        .B2(n6086), .ZN(n6038) );
  OAI211_X1 U6983 ( .C1(n6334), .C2(n6060), .A(n6039), .B(n6038), .ZN(U3036)
         );
  AOI22_X1 U6984 ( .A1(n6427), .A2(n6056), .B1(n6426), .B2(n6055), .ZN(n6041)
         );
  AOI22_X1 U6985 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6335), .ZN(n6040) );
  OAI211_X1 U6986 ( .C1(n6060), .C2(n6338), .A(n6041), .B(n6040), .ZN(U3037)
         );
  AOI22_X1 U6987 ( .A1(n6433), .A2(n6056), .B1(n6432), .B2(n6055), .ZN(n6043)
         );
  AOI22_X1 U6988 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6259), .ZN(n6042) );
  OAI211_X1 U6989 ( .C1(n6060), .C2(n6262), .A(n6043), .B(n6042), .ZN(U3038)
         );
  AOI22_X1 U6990 ( .A1(n6439), .A2(n6056), .B1(n6438), .B2(n6055), .ZN(n6045)
         );
  AOI22_X1 U6991 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6224), .ZN(n6044) );
  OAI211_X1 U6992 ( .C1(n6060), .C2(n6227), .A(n6045), .B(n6044), .ZN(U3039)
         );
  INV_X1 U6993 ( .A(n6056), .ZN(n6047) );
  OAI22_X1 U6994 ( .A1(n6447), .A2(n6047), .B1(n6046), .B2(n6444), .ZN(n6048)
         );
  INV_X1 U6995 ( .A(n6048), .ZN(n6050) );
  AOI22_X1 U6996 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6449), .ZN(n6049) );
  OAI211_X1 U6997 ( .C1(n6060), .C2(n6452), .A(n6050), .B(n6049), .ZN(U3040)
         );
  AOI22_X1 U6998 ( .A1(n6454), .A2(n6056), .B1(n6453), .B2(n6055), .ZN(n6052)
         );
  AOI22_X1 U6999 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6348), .ZN(n6051) );
  OAI211_X1 U7000 ( .C1(n6060), .C2(n6352), .A(n6052), .B(n6051), .ZN(U3041)
         );
  AOI22_X1 U7001 ( .A1(n6462), .A2(n6056), .B1(n6461), .B2(n6055), .ZN(n6054)
         );
  AOI22_X1 U7002 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6463), .ZN(n6053) );
  OAI211_X1 U7003 ( .C1(n6060), .C2(n6466), .A(n6054), .B(n6053), .ZN(U3042)
         );
  AOI22_X1 U7004 ( .A1(n6470), .A2(n6056), .B1(n6468), .B2(n6055), .ZN(n6059)
         );
  AOI22_X1 U7005 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n6057), .B1(n6086), 
        .B2(n6472), .ZN(n6058) );
  OAI211_X1 U7006 ( .C1(n6060), .C2(n6477), .A(n6059), .B(n6058), .ZN(U3043)
         );
  INV_X1 U7007 ( .A(n6086), .ZN(n6095) );
  NOR2_X1 U7008 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6242), .ZN(n6090)
         );
  INV_X1 U7009 ( .A(n6104), .ZN(n6089) );
  AOI22_X1 U7010 ( .A1(n6410), .A2(n6090), .B1(n6089), .B2(n6331), .ZN(n6073)
         );
  NAND2_X1 U7011 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  OAI21_X1 U7012 ( .B1(n6064), .B2(n6063), .A(n6405), .ZN(n6071) );
  OR2_X1 U7013 ( .A1(n6065), .A2(n6482), .ZN(n6066) );
  INV_X1 U7014 ( .A(n6090), .ZN(n6080) );
  NAND2_X1 U7015 ( .A1(n6066), .A2(n6080), .ZN(n6068) );
  AOI21_X1 U7016 ( .B1(n6069), .B2(n6417), .A(n6416), .ZN(n6067) );
  OAI21_X1 U7017 ( .B1(n6071), .B2(n6068), .A(n6067), .ZN(n6092) );
  INV_X1 U7018 ( .A(n6068), .ZN(n6070) );
  OAI22_X1 U7019 ( .A1(n6071), .A2(n6070), .B1(n6069), .B2(n6251), .ZN(n6091)
         );
  AOI22_X1 U7020 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6092), .B1(n6409), 
        .B2(n6091), .ZN(n6072) );
  OAI211_X1 U7021 ( .C1(n6334), .C2(n6095), .A(n6073), .B(n6072), .ZN(U3044)
         );
  AOI22_X1 U7022 ( .A1(n6427), .A2(n6090), .B1(n6089), .B2(n6335), .ZN(n6075)
         );
  AOI22_X1 U7023 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6092), .B1(n6426), 
        .B2(n6091), .ZN(n6074) );
  OAI211_X1 U7024 ( .C1(n6095), .C2(n6338), .A(n6075), .B(n6074), .ZN(U3045)
         );
  AOI22_X1 U7025 ( .A1(n6433), .A2(n6090), .B1(n6434), .B2(n6086), .ZN(n6077)
         );
  AOI22_X1 U7026 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6092), .B1(n6432), 
        .B2(n6091), .ZN(n6076) );
  OAI211_X1 U7027 ( .C1(n6437), .C2(n6104), .A(n6077), .B(n6076), .ZN(U3046)
         );
  AOI22_X1 U7028 ( .A1(n6439), .A2(n6090), .B1(n6440), .B2(n6086), .ZN(n6079)
         );
  AOI22_X1 U7029 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6092), .B1(n6438), 
        .B2(n6091), .ZN(n6078) );
  OAI211_X1 U7030 ( .C1(n6443), .C2(n6104), .A(n6079), .B(n6078), .ZN(U3047)
         );
  OAI22_X1 U7031 ( .A1(n6447), .A2(n6080), .B1(n6266), .B2(n6104), .ZN(n6081)
         );
  INV_X1 U7032 ( .A(n6081), .ZN(n6083) );
  AOI22_X1 U7033 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6092), .B1(n6269), 
        .B2(n6091), .ZN(n6082) );
  OAI211_X1 U7034 ( .C1(n6095), .C2(n6452), .A(n6083), .B(n6082), .ZN(U3048)
         );
  AOI22_X1 U7035 ( .A1(n6454), .A2(n6090), .B1(n6456), .B2(n6086), .ZN(n6085)
         );
  AOI22_X1 U7036 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6092), .B1(n6453), 
        .B2(n6091), .ZN(n6084) );
  OAI211_X1 U7037 ( .C1(n6460), .C2(n6104), .A(n6085), .B(n6084), .ZN(U3049)
         );
  AOI22_X1 U7038 ( .A1(n6462), .A2(n6090), .B1(n6390), .B2(n6086), .ZN(n6088)
         );
  AOI22_X1 U7039 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6092), .B1(n6461), 
        .B2(n6091), .ZN(n6087) );
  OAI211_X1 U7040 ( .C1(n6393), .C2(n6104), .A(n6088), .B(n6087), .ZN(U3050)
         );
  AOI22_X1 U7041 ( .A1(n6470), .A2(n6090), .B1(n6089), .B2(n6472), .ZN(n6094)
         );
  AOI22_X1 U7042 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6092), .B1(n6468), 
        .B2(n6091), .ZN(n6093) );
  OAI211_X1 U7043 ( .C1(n6095), .C2(n6477), .A(n6094), .B(n6093), .ZN(U3051)
         );
  INV_X1 U7044 ( .A(n6096), .ZN(n6098) );
  OAI22_X1 U7045 ( .A1(n6447), .A2(n6098), .B1(n6097), .B2(n6444), .ZN(n6099)
         );
  INV_X1 U7046 ( .A(n6099), .ZN(n6103) );
  AOI22_X1 U7047 ( .A1(n6101), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6449), 
        .B2(n6100), .ZN(n6102) );
  OAI211_X1 U7048 ( .C1(n6452), .C2(n6104), .A(n6103), .B(n6102), .ZN(U3056)
         );
  INV_X1 U7049 ( .A(n6331), .ZN(n6425) );
  INV_X1 U7050 ( .A(n6105), .ZN(n6106) );
  AOI22_X1 U7051 ( .A1(n6410), .A2(n6107), .B1(n6409), .B2(n6106), .ZN(n6111)
         );
  AOI22_X1 U7052 ( .A1(n6109), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6422), 
        .B2(n6108), .ZN(n6110) );
  OAI211_X1 U7053 ( .C1(n6425), .C2(n6135), .A(n6111), .B(n6110), .ZN(U3068)
         );
  AOI22_X1 U7054 ( .A1(n6410), .A2(n6139), .B1(n6138), .B2(n6422), .ZN(n6122)
         );
  AOI21_X1 U7055 ( .B1(n6114), .B2(n3159), .A(n6139), .ZN(n6120) );
  INV_X1 U7056 ( .A(n6120), .ZN(n6117) );
  NAND2_X1 U7057 ( .A1(n6603), .A2(n6115), .ZN(n6119) );
  AOI21_X1 U7058 ( .B1(n6118), .B2(n6417), .A(n6416), .ZN(n6116) );
  OAI21_X1 U7059 ( .B1(n6117), .B2(n6119), .A(n6116), .ZN(n6141) );
  OAI22_X1 U7060 ( .A1(n6120), .A2(n6119), .B1(n6251), .B2(n6118), .ZN(n6140)
         );
  AOI22_X1 U7061 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6141), .B1(n6409), 
        .B2(n6140), .ZN(n6121) );
  OAI211_X1 U7062 ( .C1(n6425), .C2(n6176), .A(n6122), .B(n6121), .ZN(U3076)
         );
  INV_X1 U7063 ( .A(n6176), .ZN(n6148) );
  AOI22_X1 U7064 ( .A1(n6427), .A2(n6139), .B1(n6335), .B2(n6148), .ZN(n6124)
         );
  AOI22_X1 U7065 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6141), .B1(n6426), 
        .B2(n6140), .ZN(n6123) );
  OAI211_X1 U7066 ( .C1(n6338), .C2(n6135), .A(n6124), .B(n6123), .ZN(U3077)
         );
  AOI22_X1 U7067 ( .A1(n6433), .A2(n6139), .B1(n6259), .B2(n6148), .ZN(n6126)
         );
  AOI22_X1 U7068 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6141), .B1(n6432), 
        .B2(n6140), .ZN(n6125) );
  OAI211_X1 U7069 ( .C1(n6262), .C2(n6135), .A(n6126), .B(n6125), .ZN(U3078)
         );
  AOI22_X1 U7070 ( .A1(n6439), .A2(n6139), .B1(n6138), .B2(n6440), .ZN(n6128)
         );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6141), .B1(n6438), 
        .B2(n6140), .ZN(n6127) );
  OAI211_X1 U7072 ( .C1(n6443), .C2(n6176), .A(n6128), .B(n6127), .ZN(U3079)
         );
  INV_X1 U7073 ( .A(n6139), .ZN(n6129) );
  OAI22_X1 U7074 ( .A1(n6447), .A2(n6129), .B1(n6266), .B2(n6176), .ZN(n6130)
         );
  INV_X1 U7075 ( .A(n6130), .ZN(n6132) );
  AOI22_X1 U7076 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6141), .B1(n6269), 
        .B2(n6140), .ZN(n6131) );
  OAI211_X1 U7077 ( .C1(n6452), .C2(n6135), .A(n6132), .B(n6131), .ZN(U3080)
         );
  AOI22_X1 U7078 ( .A1(n6454), .A2(n6139), .B1(n6348), .B2(n6148), .ZN(n6134)
         );
  AOI22_X1 U7079 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6141), .B1(n6453), 
        .B2(n6140), .ZN(n6133) );
  OAI211_X1 U7080 ( .C1(n6352), .C2(n6135), .A(n6134), .B(n6133), .ZN(U3081)
         );
  AOI22_X1 U7081 ( .A1(n6462), .A2(n6139), .B1(n6138), .B2(n6390), .ZN(n6137)
         );
  AOI22_X1 U7082 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6141), .B1(n6461), 
        .B2(n6140), .ZN(n6136) );
  OAI211_X1 U7083 ( .C1(n6393), .C2(n6176), .A(n6137), .B(n6136), .ZN(U3082)
         );
  AOI22_X1 U7084 ( .A1(n6470), .A2(n6139), .B1(n6138), .B2(n6397), .ZN(n6143)
         );
  AOI22_X1 U7085 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6141), .B1(n6468), 
        .B2(n6140), .ZN(n6142) );
  OAI211_X1 U7086 ( .C1(n6401), .C2(n6176), .A(n6143), .B(n6142), .ZN(U3083)
         );
  NAND3_X1 U7087 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6209), .A3(n6487), .ZN(n6182) );
  NOR2_X1 U7088 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6182), .ZN(n6172)
         );
  NAND2_X1 U7089 ( .A1(n6177), .A2(n6362), .ZN(n6149) );
  OR2_X1 U7090 ( .A1(n6149), .A2(n6417), .ZN(n6146) );
  NOR2_X1 U7091 ( .A1(n6144), .A2(n6364), .ZN(n6284) );
  NAND2_X1 U7092 ( .A1(n6284), .A2(n6368), .ZN(n6145) );
  AND2_X1 U7093 ( .A1(n6146), .A2(n6145), .ZN(n6162) );
  INV_X1 U7094 ( .A(n6162), .ZN(n6171) );
  AOI22_X1 U7095 ( .A1(n6410), .A2(n6172), .B1(n6409), .B2(n6171), .ZN(n6155)
         );
  NAND2_X1 U7096 ( .A1(n6178), .A2(n6282), .ZN(n6208) );
  NOR3_X1 U7097 ( .A1(n6199), .A2(n6148), .A3(n6417), .ZN(n6150) );
  OAI21_X1 U7098 ( .B1(n6150), .B2(n6414), .A(n6149), .ZN(n6153) );
  INV_X1 U7099 ( .A(n6172), .ZN(n6163) );
  OAI21_X1 U7100 ( .B1(n6284), .B2(n6251), .A(n6151), .ZN(n6290) );
  AOI211_X1 U7101 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6163), .A(n6365), .B(
        n6290), .ZN(n6152) );
  NAND2_X1 U7102 ( .A1(n6153), .A2(n6152), .ZN(n6173) );
  AOI22_X1 U7103 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n6173), .B1(n6331), 
        .B2(n6199), .ZN(n6154) );
  OAI211_X1 U7104 ( .C1(n6334), .C2(n6176), .A(n6155), .B(n6154), .ZN(U3084)
         );
  AOI22_X1 U7105 ( .A1(n6427), .A2(n6172), .B1(n6426), .B2(n6171), .ZN(n6157)
         );
  AOI22_X1 U7106 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n6173), .B1(n6335), 
        .B2(n6199), .ZN(n6156) );
  OAI211_X1 U7107 ( .C1(n6338), .C2(n6176), .A(n6157), .B(n6156), .ZN(U3085)
         );
  AOI22_X1 U7108 ( .A1(n6433), .A2(n6172), .B1(n6432), .B2(n6171), .ZN(n6159)
         );
  AOI22_X1 U7109 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n6173), .B1(n6259), 
        .B2(n6199), .ZN(n6158) );
  OAI211_X1 U7110 ( .C1(n6262), .C2(n6176), .A(n6159), .B(n6158), .ZN(U3086)
         );
  AOI22_X1 U7111 ( .A1(n6439), .A2(n6172), .B1(n6438), .B2(n6171), .ZN(n6161)
         );
  AOI22_X1 U7112 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n6173), .B1(n6224), 
        .B2(n6199), .ZN(n6160) );
  OAI211_X1 U7113 ( .C1(n6227), .C2(n6176), .A(n6161), .B(n6160), .ZN(U3087)
         );
  OAI22_X1 U7114 ( .A1(n6447), .A2(n6163), .B1(n6162), .B2(n6444), .ZN(n6164)
         );
  INV_X1 U7115 ( .A(n6164), .ZN(n6166) );
  AOI22_X1 U7116 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n6173), .B1(n6449), 
        .B2(n6199), .ZN(n6165) );
  OAI211_X1 U7117 ( .C1(n6452), .C2(n6176), .A(n6166), .B(n6165), .ZN(U3088)
         );
  AOI22_X1 U7118 ( .A1(n6454), .A2(n6172), .B1(n6453), .B2(n6171), .ZN(n6168)
         );
  AOI22_X1 U7119 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n6173), .B1(n6348), 
        .B2(n6199), .ZN(n6167) );
  OAI211_X1 U7120 ( .C1(n6352), .C2(n6176), .A(n6168), .B(n6167), .ZN(U3089)
         );
  AOI22_X1 U7121 ( .A1(n6462), .A2(n6172), .B1(n6461), .B2(n6171), .ZN(n6170)
         );
  AOI22_X1 U7122 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n6173), .B1(n6463), 
        .B2(n6199), .ZN(n6169) );
  OAI211_X1 U7123 ( .C1(n6466), .C2(n6176), .A(n6170), .B(n6169), .ZN(U3090)
         );
  AOI22_X1 U7124 ( .A1(n6470), .A2(n6172), .B1(n6468), .B2(n6171), .ZN(n6175)
         );
  AOI22_X1 U7125 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n6173), .B1(n6472), 
        .B2(n6199), .ZN(n6174) );
  OAI211_X1 U7126 ( .C1(n6477), .C2(n6176), .A(n6175), .B(n6174), .ZN(U3091)
         );
  NOR2_X1 U7127 ( .A1(n6283), .A2(n6182), .ZN(n6202) );
  AOI22_X1 U7128 ( .A1(n6199), .A2(n6422), .B1(n6410), .B2(n6202), .ZN(n6186)
         );
  NAND2_X1 U7129 ( .A1(n6362), .A2(n3159), .ZN(n6403) );
  INV_X1 U7130 ( .A(n6403), .ZN(n6318) );
  AOI21_X1 U7131 ( .B1(n6318), .B2(n6177), .A(n6202), .ZN(n6184) );
  INV_X1 U7132 ( .A(n6184), .ZN(n6181) );
  INV_X1 U7133 ( .A(n6178), .ZN(n6179) );
  OAI21_X1 U7134 ( .B1(n6179), .B2(n6596), .A(n6603), .ZN(n6183) );
  AOI21_X1 U7135 ( .B1(n6417), .B2(n6182), .A(n6416), .ZN(n6180) );
  OAI21_X1 U7136 ( .B1(n6181), .B2(n6183), .A(n6180), .ZN(n6205) );
  OAI22_X1 U7137 ( .A1(n6184), .A2(n6183), .B1(n6251), .B2(n6182), .ZN(n6204)
         );
  AOI22_X1 U7138 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6205), .B1(n6409), 
        .B2(n6204), .ZN(n6185) );
  OAI211_X1 U7139 ( .C1(n6425), .C2(n6241), .A(n6186), .B(n6185), .ZN(U3092)
         );
  AOI22_X1 U7140 ( .A1(n6199), .A2(n6428), .B1(n6427), .B2(n6202), .ZN(n6188)
         );
  AOI22_X1 U7141 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6205), .B1(n6426), 
        .B2(n6204), .ZN(n6187) );
  OAI211_X1 U7142 ( .C1(n6431), .C2(n6241), .A(n6188), .B(n6187), .ZN(U3093)
         );
  AOI22_X1 U7143 ( .A1(n6199), .A2(n6434), .B1(n6433), .B2(n6202), .ZN(n6190)
         );
  AOI22_X1 U7144 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6205), .B1(n6432), 
        .B2(n6204), .ZN(n6189) );
  OAI211_X1 U7145 ( .C1(n6437), .C2(n6241), .A(n6190), .B(n6189), .ZN(U3094)
         );
  AOI22_X1 U7146 ( .A1(n6199), .A2(n6440), .B1(n6439), .B2(n6202), .ZN(n6192)
         );
  AOI22_X1 U7147 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6205), .B1(n6438), 
        .B2(n6204), .ZN(n6191) );
  OAI211_X1 U7148 ( .C1(n6443), .C2(n6241), .A(n6192), .B(n6191), .ZN(U3095)
         );
  INV_X1 U7149 ( .A(n6202), .ZN(n6193) );
  OAI22_X1 U7150 ( .A1(n6241), .A2(n6266), .B1(n6447), .B2(n6193), .ZN(n6194)
         );
  INV_X1 U7151 ( .A(n6194), .ZN(n6196) );
  AOI22_X1 U7152 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6205), .B1(n6269), 
        .B2(n6204), .ZN(n6195) );
  OAI211_X1 U7153 ( .C1(n6452), .C2(n6208), .A(n6196), .B(n6195), .ZN(U3096)
         );
  AOI22_X1 U7154 ( .A1(n6199), .A2(n6456), .B1(n6454), .B2(n6202), .ZN(n6198)
         );
  AOI22_X1 U7155 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6205), .B1(n6453), 
        .B2(n6204), .ZN(n6197) );
  OAI211_X1 U7156 ( .C1(n6460), .C2(n6241), .A(n6198), .B(n6197), .ZN(U3097)
         );
  AOI22_X1 U7157 ( .A1(n6199), .A2(n6390), .B1(n6462), .B2(n6202), .ZN(n6201)
         );
  AOI22_X1 U7158 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6205), .B1(n6461), 
        .B2(n6204), .ZN(n6200) );
  OAI211_X1 U7159 ( .C1(n6393), .C2(n6241), .A(n6201), .B(n6200), .ZN(U3098)
         );
  INV_X1 U7160 ( .A(n6241), .ZN(n6203) );
  AOI22_X1 U7161 ( .A1(n6203), .A2(n6472), .B1(n6470), .B2(n6202), .ZN(n6207)
         );
  AOI22_X1 U7162 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6205), .B1(n6468), 
        .B2(n6204), .ZN(n6206) );
  OAI211_X1 U7163 ( .C1(n6477), .C2(n6208), .A(n6207), .B(n6206), .ZN(U3099)
         );
  NAND3_X1 U7164 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6209), .ZN(n6252) );
  NOR2_X1 U7165 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6252), .ZN(n6236)
         );
  AOI22_X1 U7166 ( .A1(n6410), .A2(n6236), .B1(n6263), .B2(n6331), .ZN(n6219)
         );
  NAND2_X1 U7167 ( .A1(n6241), .A2(n6281), .ZN(n6211) );
  AOI21_X1 U7168 ( .B1(n6211), .B2(STATEBS16_REG_SCAN_IN), .A(n6417), .ZN(
        n6215) );
  NAND2_X1 U7169 ( .A1(n6212), .A2(n6362), .ZN(n6247) );
  INV_X1 U7170 ( .A(n6236), .ZN(n6228) );
  AOI22_X1 U7171 ( .A1(n6215), .A2(n6247), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6228), .ZN(n6213) );
  OAI211_X1 U7172 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6251), .A(n6214), .B(n6213), .ZN(n6238) );
  INV_X1 U7173 ( .A(n6215), .ZN(n6217) );
  NAND3_X1 U7174 ( .A1(n6368), .A2(n6364), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6238), .B1(n6409), 
        .B2(n6237), .ZN(n6218) );
  OAI211_X1 U7176 ( .C1(n6334), .C2(n6241), .A(n6219), .B(n6218), .ZN(U3100)
         );
  AOI22_X1 U7177 ( .A1(n6427), .A2(n6236), .B1(n6263), .B2(n6335), .ZN(n6221)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6238), .B1(n6426), 
        .B2(n6237), .ZN(n6220) );
  OAI211_X1 U7179 ( .C1(n6338), .C2(n6241), .A(n6221), .B(n6220), .ZN(U3101)
         );
  AOI22_X1 U7180 ( .A1(n6433), .A2(n6236), .B1(n6263), .B2(n6259), .ZN(n6223)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6238), .B1(n6432), 
        .B2(n6237), .ZN(n6222) );
  OAI211_X1 U7182 ( .C1(n6262), .C2(n6241), .A(n6223), .B(n6222), .ZN(U3102)
         );
  AOI22_X1 U7183 ( .A1(n6439), .A2(n6236), .B1(n6263), .B2(n6224), .ZN(n6226)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6238), .B1(n6438), 
        .B2(n6237), .ZN(n6225) );
  OAI211_X1 U7185 ( .C1(n6227), .C2(n6241), .A(n6226), .B(n6225), .ZN(U3103)
         );
  OAI22_X1 U7186 ( .A1(n6447), .A2(n6228), .B1(n6266), .B2(n6281), .ZN(n6229)
         );
  INV_X1 U7187 ( .A(n6229), .ZN(n6231) );
  AOI22_X1 U7188 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6238), .B1(n6269), 
        .B2(n6237), .ZN(n6230) );
  OAI211_X1 U7189 ( .C1(n6452), .C2(n6241), .A(n6231), .B(n6230), .ZN(U3104)
         );
  AOI22_X1 U7190 ( .A1(n6454), .A2(n6236), .B1(n6263), .B2(n6348), .ZN(n6233)
         );
  AOI22_X1 U7191 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6238), .B1(n6453), 
        .B2(n6237), .ZN(n6232) );
  OAI211_X1 U7192 ( .C1(n6352), .C2(n6241), .A(n6233), .B(n6232), .ZN(U3105)
         );
  AOI22_X1 U7193 ( .A1(n6462), .A2(n6236), .B1(n6263), .B2(n6463), .ZN(n6235)
         );
  AOI22_X1 U7194 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6238), .B1(n6461), 
        .B2(n6237), .ZN(n6234) );
  OAI211_X1 U7195 ( .C1(n6466), .C2(n6241), .A(n6235), .B(n6234), .ZN(U3106)
         );
  AOI22_X1 U7196 ( .A1(n6470), .A2(n6236), .B1(n6263), .B2(n6472), .ZN(n6240)
         );
  AOI22_X1 U7197 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6238), .B1(n6468), 
        .B2(n6237), .ZN(n6239) );
  OAI211_X1 U7198 ( .C1(n6477), .C2(n6241), .A(n6240), .B(n6239), .ZN(U3107)
         );
  NOR2_X1 U7199 ( .A1(n6493), .A2(n6242), .ZN(n6276) );
  NAND2_X1 U7200 ( .A1(n6244), .A2(n6243), .ZN(n6306) );
  AOI22_X1 U7201 ( .A1(n6410), .A2(n6276), .B1(n6313), .B2(n6331), .ZN(n6256)
         );
  OAI21_X1 U7202 ( .B1(n6246), .B2(n6245), .A(n6405), .ZN(n6254) );
  OR2_X1 U7203 ( .A1(n6247), .A2(n6482), .ZN(n6248) );
  INV_X1 U7204 ( .A(n6276), .ZN(n6267) );
  NAND2_X1 U7205 ( .A1(n6248), .A2(n6267), .ZN(n6250) );
  INV_X1 U7206 ( .A(n6416), .ZN(n6326) );
  NAND2_X1 U7207 ( .A1(n6417), .A2(n6252), .ZN(n6249) );
  OAI211_X1 U7208 ( .C1(n6254), .C2(n6250), .A(n6326), .B(n6249), .ZN(n6278)
         );
  INV_X1 U7209 ( .A(n6250), .ZN(n6253) );
  OAI22_X1 U7210 ( .A1(n6254), .A2(n6253), .B1(n6252), .B2(n6251), .ZN(n6277)
         );
  AOI22_X1 U7211 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6278), .B1(n6409), 
        .B2(n6277), .ZN(n6255) );
  OAI211_X1 U7212 ( .C1(n6334), .C2(n6281), .A(n6256), .B(n6255), .ZN(U3108)
         );
  AOI22_X1 U7213 ( .A1(n6427), .A2(n6276), .B1(n6263), .B2(n6428), .ZN(n6258)
         );
  AOI22_X1 U7214 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6278), .B1(n6426), 
        .B2(n6277), .ZN(n6257) );
  OAI211_X1 U7215 ( .C1(n6431), .C2(n6306), .A(n6258), .B(n6257), .ZN(U3109)
         );
  AOI22_X1 U7216 ( .A1(n6433), .A2(n6276), .B1(n6313), .B2(n6259), .ZN(n6261)
         );
  AOI22_X1 U7217 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6278), .B1(n6432), 
        .B2(n6277), .ZN(n6260) );
  OAI211_X1 U7218 ( .C1(n6262), .C2(n6281), .A(n6261), .B(n6260), .ZN(U3110)
         );
  AOI22_X1 U7219 ( .A1(n6439), .A2(n6276), .B1(n6263), .B2(n6440), .ZN(n6265)
         );
  AOI22_X1 U7220 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6278), .B1(n6438), 
        .B2(n6277), .ZN(n6264) );
  OAI211_X1 U7221 ( .C1(n6443), .C2(n6306), .A(n6265), .B(n6264), .ZN(U3111)
         );
  OAI22_X1 U7222 ( .A1(n6447), .A2(n6267), .B1(n6266), .B2(n6306), .ZN(n6268)
         );
  INV_X1 U7223 ( .A(n6268), .ZN(n6271) );
  AOI22_X1 U7224 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6278), .B1(n6269), 
        .B2(n6277), .ZN(n6270) );
  OAI211_X1 U7225 ( .C1(n6452), .C2(n6281), .A(n6271), .B(n6270), .ZN(U3112)
         );
  AOI22_X1 U7226 ( .A1(n6454), .A2(n6276), .B1(n6313), .B2(n6348), .ZN(n6273)
         );
  AOI22_X1 U7227 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6278), .B1(n6453), 
        .B2(n6277), .ZN(n6272) );
  OAI211_X1 U7228 ( .C1(n6352), .C2(n6281), .A(n6273), .B(n6272), .ZN(U3113)
         );
  AOI22_X1 U7229 ( .A1(n6462), .A2(n6276), .B1(n6313), .B2(n6463), .ZN(n6275)
         );
  AOI22_X1 U7230 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6278), .B1(n6461), 
        .B2(n6277), .ZN(n6274) );
  OAI211_X1 U7231 ( .C1(n6466), .C2(n6281), .A(n6275), .B(n6274), .ZN(U3114)
         );
  AOI22_X1 U7232 ( .A1(n6470), .A2(n6276), .B1(n6313), .B2(n6472), .ZN(n6280)
         );
  AOI22_X1 U7233 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6278), .B1(n6468), 
        .B2(n6277), .ZN(n6279) );
  OAI211_X1 U7234 ( .C1(n6477), .C2(n6281), .A(n6280), .B(n6279), .ZN(U3115)
         );
  NOR2_X1 U7235 ( .A1(n6493), .A2(n6319), .ZN(n6328) );
  NAND2_X1 U7236 ( .A1(n6283), .A2(n6328), .ZN(n6302) );
  INV_X1 U7237 ( .A(n6302), .ZN(n6312) );
  AND2_X1 U7238 ( .A1(n6317), .A2(n6362), .ZN(n6287) );
  NAND2_X1 U7239 ( .A1(n6287), .A2(n6603), .ZN(n6286) );
  NAND2_X1 U7240 ( .A1(n6284), .A2(n6365), .ZN(n6285) );
  AND2_X1 U7241 ( .A1(n6286), .A2(n6285), .ZN(n6301) );
  INV_X1 U7242 ( .A(n6301), .ZN(n6311) );
  AOI22_X1 U7243 ( .A1(n6410), .A2(n6312), .B1(n6409), .B2(n6311), .ZN(n6294)
         );
  AOI21_X1 U7244 ( .B1(n6351), .B2(n6306), .A(n6596), .ZN(n6288) );
  NOR3_X1 U7245 ( .A1(n6288), .A2(n6287), .A3(n6417), .ZN(n6289) );
  AOI211_X1 U7246 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6302), .A(n6290), .B(
        n6289), .ZN(n6292) );
  INV_X1 U7247 ( .A(n6368), .ZN(n6291) );
  NAND2_X1 U7248 ( .A1(n6292), .A2(n6291), .ZN(n6314) );
  AOI22_X1 U7249 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6314), .B1(n6422), 
        .B2(n6313), .ZN(n6293) );
  OAI211_X1 U7250 ( .C1(n6425), .C2(n6351), .A(n6294), .B(n6293), .ZN(U3116)
         );
  AOI22_X1 U7251 ( .A1(n6427), .A2(n6312), .B1(n6426), .B2(n6311), .ZN(n6296)
         );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6314), .B1(n6428), 
        .B2(n6313), .ZN(n6295) );
  OAI211_X1 U7253 ( .C1(n6431), .C2(n6351), .A(n6296), .B(n6295), .ZN(U3117)
         );
  AOI22_X1 U7254 ( .A1(n6433), .A2(n6312), .B1(n6432), .B2(n6311), .ZN(n6298)
         );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6314), .B1(n6434), 
        .B2(n6313), .ZN(n6297) );
  OAI211_X1 U7256 ( .C1(n6437), .C2(n6351), .A(n6298), .B(n6297), .ZN(U3118)
         );
  AOI22_X1 U7257 ( .A1(n6439), .A2(n6312), .B1(n6438), .B2(n6311), .ZN(n6300)
         );
  AOI22_X1 U7258 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6314), .B1(n6440), 
        .B2(n6313), .ZN(n6299) );
  OAI211_X1 U7259 ( .C1(n6443), .C2(n6351), .A(n6300), .B(n6299), .ZN(U3119)
         );
  OAI22_X1 U7260 ( .A1(n6447), .A2(n6302), .B1(n6301), .B2(n6444), .ZN(n6303)
         );
  INV_X1 U7261 ( .A(n6303), .ZN(n6305) );
  INV_X1 U7262 ( .A(n6351), .ZN(n6357) );
  AOI22_X1 U7263 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6314), .B1(n6449), 
        .B2(n6357), .ZN(n6304) );
  OAI211_X1 U7264 ( .C1(n6452), .C2(n6306), .A(n6305), .B(n6304), .ZN(U3120)
         );
  AOI22_X1 U7265 ( .A1(n6454), .A2(n6312), .B1(n6453), .B2(n6311), .ZN(n6308)
         );
  AOI22_X1 U7266 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6314), .B1(n6456), 
        .B2(n6313), .ZN(n6307) );
  OAI211_X1 U7267 ( .C1(n6460), .C2(n6351), .A(n6308), .B(n6307), .ZN(U3121)
         );
  AOI22_X1 U7268 ( .A1(n6462), .A2(n6312), .B1(n6461), .B2(n6311), .ZN(n6310)
         );
  AOI22_X1 U7269 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6314), .B1(n6390), 
        .B2(n6313), .ZN(n6309) );
  OAI211_X1 U7270 ( .C1(n6393), .C2(n6351), .A(n6310), .B(n6309), .ZN(U3122)
         );
  AOI22_X1 U7271 ( .A1(n6470), .A2(n6312), .B1(n6468), .B2(n6311), .ZN(n6316)
         );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6314), .B1(n6397), 
        .B2(n6313), .ZN(n6315) );
  OAI211_X1 U7273 ( .C1(n6401), .C2(n6351), .A(n6316), .B(n6315), .ZN(U3123)
         );
  AND2_X1 U7274 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6328), .ZN(n6356)
         );
  AOI21_X1 U7275 ( .B1(n6318), .B2(n6317), .A(n6356), .ZN(n6325) );
  OR2_X1 U7276 ( .A1(n6325), .A2(n6417), .ZN(n6323) );
  INV_X1 U7277 ( .A(n6319), .ZN(n6321) );
  AND2_X1 U7278 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7279 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  AND2_X1 U7280 ( .A1(n6323), .A2(n6322), .ZN(n6343) );
  INV_X1 U7281 ( .A(n6343), .ZN(n6355) );
  AOI22_X1 U7282 ( .A1(n6410), .A2(n6356), .B1(n6409), .B2(n6355), .ZN(n6333)
         );
  NAND2_X1 U7283 ( .A1(n6325), .A2(n6324), .ZN(n6327) );
  OAI221_X1 U7284 ( .B1(n6405), .B2(n6328), .C1(n6417), .C2(n6327), .A(n6326), 
        .ZN(n6358) );
  NAND2_X1 U7285 ( .A1(n6330), .A2(n6329), .ZN(n6387) );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6358), .B1(n6331), 
        .B2(n6396), .ZN(n6332) );
  OAI211_X1 U7287 ( .C1(n6334), .C2(n6351), .A(n6333), .B(n6332), .ZN(U3124)
         );
  AOI22_X1 U7288 ( .A1(n6427), .A2(n6356), .B1(n6426), .B2(n6355), .ZN(n6337)
         );
  AOI22_X1 U7289 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6358), .B1(n6335), 
        .B2(n6396), .ZN(n6336) );
  OAI211_X1 U7290 ( .C1(n6338), .C2(n6351), .A(n6337), .B(n6336), .ZN(U3125)
         );
  AOI22_X1 U7291 ( .A1(n6433), .A2(n6356), .B1(n6432), .B2(n6355), .ZN(n6340)
         );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6358), .B1(n6434), 
        .B2(n6357), .ZN(n6339) );
  OAI211_X1 U7293 ( .C1(n6437), .C2(n6387), .A(n6340), .B(n6339), .ZN(U3126)
         );
  AOI22_X1 U7294 ( .A1(n6439), .A2(n6356), .B1(n6438), .B2(n6355), .ZN(n6342)
         );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6358), .B1(n6440), 
        .B2(n6357), .ZN(n6341) );
  OAI211_X1 U7296 ( .C1(n6443), .C2(n6387), .A(n6342), .B(n6341), .ZN(U3127)
         );
  INV_X1 U7297 ( .A(n6356), .ZN(n6344) );
  OAI22_X1 U7298 ( .A1(n6447), .A2(n6344), .B1(n6343), .B2(n6444), .ZN(n6345)
         );
  INV_X1 U7299 ( .A(n6345), .ZN(n6347) );
  AOI22_X1 U7300 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6358), .B1(n6449), 
        .B2(n6396), .ZN(n6346) );
  OAI211_X1 U7301 ( .C1(n6452), .C2(n6351), .A(n6347), .B(n6346), .ZN(U3128)
         );
  AOI22_X1 U7302 ( .A1(n6454), .A2(n6356), .B1(n6453), .B2(n6355), .ZN(n6350)
         );
  AOI22_X1 U7303 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6358), .B1(n6348), 
        .B2(n6396), .ZN(n6349) );
  OAI211_X1 U7304 ( .C1(n6352), .C2(n6351), .A(n6350), .B(n6349), .ZN(U3129)
         );
  AOI22_X1 U7305 ( .A1(n6462), .A2(n6356), .B1(n6461), .B2(n6355), .ZN(n6354)
         );
  AOI22_X1 U7306 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6358), .B1(n6390), 
        .B2(n6357), .ZN(n6353) );
  OAI211_X1 U7307 ( .C1(n6393), .C2(n6387), .A(n6354), .B(n6353), .ZN(U3130)
         );
  AOI22_X1 U7308 ( .A1(n6470), .A2(n6356), .B1(n6468), .B2(n6355), .ZN(n6360)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6358), .B1(n6397), 
        .B2(n6357), .ZN(n6359) );
  OAI211_X1 U7310 ( .C1(n6401), .C2(n6387), .A(n6360), .B(n6359), .ZN(U3131)
         );
  NOR2_X1 U7311 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6418), .ZN(n6395)
         );
  INV_X1 U7312 ( .A(n6402), .ZN(n6363) );
  NAND3_X1 U7313 ( .A1(n6363), .A2(n6405), .A3(n6362), .ZN(n6367) );
  NAND3_X1 U7314 ( .A1(n6365), .A2(n6364), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6366) );
  AND2_X1 U7315 ( .A1(n6367), .A2(n6366), .ZN(n6382) );
  INV_X1 U7316 ( .A(n6382), .ZN(n6394) );
  AOI22_X1 U7317 ( .A1(n6410), .A2(n6395), .B1(n6409), .B2(n6394), .ZN(n6375)
         );
  NOR3_X1 U7318 ( .A1(n6369), .A2(n6493), .A3(n6368), .ZN(n6372) );
  OAI21_X1 U7319 ( .B1(n6396), .B2(n6455), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6370) );
  NAND3_X1 U7320 ( .A1(n6402), .A2(n6603), .A3(n6370), .ZN(n6371) );
  OAI211_X1 U7321 ( .C1(n6395), .C2(n6373), .A(n6372), .B(n6371), .ZN(n6398)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6398), .B1(n6422), 
        .B2(n6396), .ZN(n6374) );
  OAI211_X1 U7323 ( .C1(n6425), .C2(n6476), .A(n6375), .B(n6374), .ZN(U3132)
         );
  AOI22_X1 U7324 ( .A1(n6427), .A2(n6395), .B1(n6426), .B2(n6394), .ZN(n6377)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6398), .B1(n6428), 
        .B2(n6396), .ZN(n6376) );
  OAI211_X1 U7326 ( .C1(n6431), .C2(n6476), .A(n6377), .B(n6376), .ZN(U3133)
         );
  AOI22_X1 U7327 ( .A1(n6433), .A2(n6395), .B1(n6432), .B2(n6394), .ZN(n6379)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6398), .B1(n6434), 
        .B2(n6396), .ZN(n6378) );
  OAI211_X1 U7329 ( .C1(n6437), .C2(n6476), .A(n6379), .B(n6378), .ZN(U3134)
         );
  AOI22_X1 U7330 ( .A1(n6439), .A2(n6395), .B1(n6438), .B2(n6394), .ZN(n6381)
         );
  AOI22_X1 U7331 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6398), .B1(n6440), 
        .B2(n6396), .ZN(n6380) );
  OAI211_X1 U7332 ( .C1(n6443), .C2(n6476), .A(n6381), .B(n6380), .ZN(U3135)
         );
  INV_X1 U7333 ( .A(n6395), .ZN(n6383) );
  OAI22_X1 U7334 ( .A1(n6447), .A2(n6383), .B1(n6382), .B2(n6444), .ZN(n6384)
         );
  INV_X1 U7335 ( .A(n6384), .ZN(n6386) );
  AOI22_X1 U7336 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6398), .B1(n6449), 
        .B2(n6455), .ZN(n6385) );
  OAI211_X1 U7337 ( .C1(n6452), .C2(n6387), .A(n6386), .B(n6385), .ZN(U3136)
         );
  AOI22_X1 U7338 ( .A1(n6454), .A2(n6395), .B1(n6453), .B2(n6394), .ZN(n6389)
         );
  AOI22_X1 U7339 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6398), .B1(n6456), 
        .B2(n6396), .ZN(n6388) );
  OAI211_X1 U7340 ( .C1(n6460), .C2(n6476), .A(n6389), .B(n6388), .ZN(U3137)
         );
  AOI22_X1 U7341 ( .A1(n6462), .A2(n6395), .B1(n6461), .B2(n6394), .ZN(n6392)
         );
  AOI22_X1 U7342 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6398), .B1(n6390), 
        .B2(n6396), .ZN(n6391) );
  OAI211_X1 U7343 ( .C1(n6393), .C2(n6476), .A(n6392), .B(n6391), .ZN(U3138)
         );
  AOI22_X1 U7344 ( .A1(n6470), .A2(n6395), .B1(n6468), .B2(n6394), .ZN(n6400)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6398), .B1(n6397), 
        .B2(n6396), .ZN(n6399) );
  OAI211_X1 U7346 ( .C1(n6401), .C2(n6476), .A(n6400), .B(n6399), .ZN(U3139)
         );
  OR2_X1 U7347 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  NAND2_X1 U7348 ( .A1(n6404), .A2(n6446), .ZN(n6420) );
  NAND2_X1 U7349 ( .A1(n6420), .A2(n6405), .ZN(n6408) );
  INV_X1 U7350 ( .A(n6418), .ZN(n6406) );
  NAND2_X1 U7351 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6406), .ZN(n6407) );
  AND2_X1 U7352 ( .A1(n6408), .A2(n6407), .ZN(n6445) );
  INV_X1 U7353 ( .A(n6445), .ZN(n6467) );
  AOI22_X1 U7354 ( .A1(n6410), .A2(n6469), .B1(n6409), .B2(n6467), .ZN(n6424)
         );
  INV_X1 U7355 ( .A(n6411), .ZN(n6413) );
  AOI21_X1 U7356 ( .B1(n6413), .B2(n3155), .A(n6412), .ZN(n6415) );
  NOR2_X1 U7357 ( .A1(n6415), .A2(n6414), .ZN(n6421) );
  AOI21_X1 U7358 ( .B1(n6418), .B2(n6417), .A(n6416), .ZN(n6419) );
  OAI21_X1 U7359 ( .B1(n6421), .B2(n6420), .A(n6419), .ZN(n6473) );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6473), .B1(n6422), 
        .B2(n6455), .ZN(n6423) );
  OAI211_X1 U7361 ( .C1(n6425), .C2(n6459), .A(n6424), .B(n6423), .ZN(U3140)
         );
  AOI22_X1 U7362 ( .A1(n6427), .A2(n6469), .B1(n6426), .B2(n6467), .ZN(n6430)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6473), .B1(n6428), 
        .B2(n6455), .ZN(n6429) );
  OAI211_X1 U7364 ( .C1(n6431), .C2(n6459), .A(n6430), .B(n6429), .ZN(U3141)
         );
  AOI22_X1 U7365 ( .A1(n6433), .A2(n6469), .B1(n6432), .B2(n6467), .ZN(n6436)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6473), .B1(n6434), 
        .B2(n6455), .ZN(n6435) );
  OAI211_X1 U7367 ( .C1(n6437), .C2(n6459), .A(n6436), .B(n6435), .ZN(U3142)
         );
  AOI22_X1 U7368 ( .A1(n6439), .A2(n6469), .B1(n6438), .B2(n6467), .ZN(n6442)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6473), .B1(n6440), 
        .B2(n6455), .ZN(n6441) );
  OAI211_X1 U7370 ( .C1(n6443), .C2(n6459), .A(n6442), .B(n6441), .ZN(U3143)
         );
  OAI22_X1 U7371 ( .A1(n6447), .A2(n6446), .B1(n6445), .B2(n6444), .ZN(n6448)
         );
  INV_X1 U7372 ( .A(n6448), .ZN(n6451) );
  AOI22_X1 U7373 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6473), .B1(n6449), 
        .B2(n6471), .ZN(n6450) );
  OAI211_X1 U7374 ( .C1(n6452), .C2(n6476), .A(n6451), .B(n6450), .ZN(U3144)
         );
  AOI22_X1 U7375 ( .A1(n6454), .A2(n6469), .B1(n6453), .B2(n6467), .ZN(n6458)
         );
  AOI22_X1 U7376 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6473), .B1(n6456), 
        .B2(n6455), .ZN(n6457) );
  OAI211_X1 U7377 ( .C1(n6460), .C2(n6459), .A(n6458), .B(n6457), .ZN(U3145)
         );
  AOI22_X1 U7378 ( .A1(n6462), .A2(n6469), .B1(n6461), .B2(n6467), .ZN(n6465)
         );
  AOI22_X1 U7379 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6473), .B1(n6463), 
        .B2(n6471), .ZN(n6464) );
  OAI211_X1 U7380 ( .C1(n6466), .C2(n6476), .A(n6465), .B(n6464), .ZN(U3146)
         );
  AOI22_X1 U7381 ( .A1(n6470), .A2(n6469), .B1(n6468), .B2(n6467), .ZN(n6475)
         );
  AOI22_X1 U7382 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6473), .B1(n6472), 
        .B2(n6471), .ZN(n6474) );
  OAI211_X1 U7383 ( .C1(n6477), .C2(n6476), .A(n6475), .B(n6474), .ZN(U3147)
         );
  MUX2_X1 U7384 ( .A(n6479), .B(n6478), .S(INSTQUEUERD_ADDR_REG_0__SCAN_IN), 
        .Z(n6480) );
  OAI211_X1 U7385 ( .C1(n6482), .C2(n6481), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6480), .ZN(n6488) );
  INV_X1 U7386 ( .A(n6488), .ZN(n6483) );
  OAI22_X1 U7387 ( .A1(n6485), .A2(n6484), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6483), .ZN(n6486) );
  OAI21_X1 U7388 ( .B1(n6488), .B2(n6487), .A(n6486), .ZN(n6490) );
  AOI222_X1 U7389 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6490), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6489), .C1(n6490), .C2(n6489), 
        .ZN(n6491) );
  AOI222_X1 U7390 ( .A1(n6493), .A2(n6492), .B1(n6493), .B2(n6491), .C1(n6492), 
        .C2(n6491), .ZN(n6494) );
  OR2_X1 U7391 ( .A1(n6494), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6502)
         );
  NOR2_X1 U7392 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6497) );
  OAI211_X1 U7393 ( .C1(n6498), .C2(n6497), .A(n6496), .B(n6495), .ZN(n6499)
         );
  NOR2_X1 U7394 ( .A1(n6500), .A2(n6499), .ZN(n6501) );
  NOR2_X1 U7395 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6896), .ZN(n6532) );
  NAND2_X1 U7396 ( .A1(n6520), .A2(n6522), .ZN(n6504) );
  NAND2_X1 U7397 ( .A1(READY_N), .A2(n4833), .ZN(n6503) );
  NAND2_X1 U7398 ( .A1(n6504), .A2(n6503), .ZN(n6509) );
  INV_X1 U7399 ( .A(n6505), .ZN(n6507) );
  NAND2_X1 U7400 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  NOR2_X1 U7401 ( .A1(n6532), .A2(n6586), .ZN(n6516) );
  OAI21_X1 U7402 ( .B1(n6598), .B2(n6510), .A(n6599), .ZN(n6511) );
  OR2_X1 U7403 ( .A1(n6586), .A2(n6511), .ZN(n6515) );
  AOI21_X1 U7404 ( .B1(n6513), .B2(n6584), .A(n6512), .ZN(n6514) );
  OAI211_X1 U7405 ( .C1(n6516), .C2(n6599), .A(n6515), .B(n6514), .ZN(n6517)
         );
  INV_X1 U7406 ( .A(n6517), .ZN(n6518) );
  OAI21_X1 U7407 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(U3148) );
  NOR2_X1 U7408 ( .A1(n6599), .A2(n6521), .ZN(n6523) );
  AOI21_X1 U7409 ( .B1(n6523), .B2(n6896), .A(n6522), .ZN(n6527) );
  INV_X1 U7410 ( .A(n6524), .ZN(n6526) );
  OAI211_X1 U7411 ( .C1(n6586), .C2(n6532), .A(STATE2_REG_1__SCAN_IN), .B(
        n6529), .ZN(n6525) );
  OAI211_X1 U7412 ( .C1(n6586), .C2(n6527), .A(n6526), .B(n6525), .ZN(U3149)
         );
  NAND3_X1 U7413 ( .A1(n6529), .A2(n6598), .A3(n6528), .ZN(n6531) );
  OAI21_X1 U7414 ( .B1(n6532), .B2(n6531), .A(n6530), .ZN(U3150) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6580), .ZN(U3151) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6580), .ZN(U3152) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6580), .ZN(U3153) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6580), .ZN(U3154) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6580), .ZN(U3155) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6580), .ZN(U3156) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6580), .ZN(U3157) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6580), .ZN(U3158) );
  INV_X1 U7423 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6979) );
  NOR2_X1 U7424 ( .A1(n6583), .A2(n6979), .ZN(U3159) );
  AND2_X1 U7425 ( .A1(n6580), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  AND2_X1 U7426 ( .A1(n6580), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7427 ( .A1(n6580), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7428 ( .A1(n6580), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7429 ( .A1(n6580), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  INV_X1 U7430 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U7431 ( .A1(n6583), .A2(n6932), .ZN(U3165) );
  INV_X1 U7432 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6913) );
  NOR2_X1 U7433 ( .A1(n6583), .A2(n6913), .ZN(U3166) );
  INV_X1 U7434 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6890) );
  NOR2_X1 U7435 ( .A1(n6583), .A2(n6890), .ZN(U3167) );
  INV_X1 U7436 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6974) );
  NOR2_X1 U7437 ( .A1(n6583), .A2(n6974), .ZN(U3168) );
  AND2_X1 U7438 ( .A1(n6580), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  INV_X1 U7439 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6948) );
  NOR2_X1 U7440 ( .A1(n6583), .A2(n6948), .ZN(U3170) );
  INV_X1 U7441 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6982) );
  NOR2_X1 U7442 ( .A1(n6583), .A2(n6982), .ZN(U3171) );
  INV_X1 U7443 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U7444 ( .A1(n6583), .A2(n6912), .ZN(U3172) );
  INV_X1 U7445 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U7446 ( .A1(n6583), .A2(n6754), .ZN(U3173) );
  AND2_X1 U7447 ( .A1(n6580), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  INV_X1 U7448 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6964) );
  NOR2_X1 U7449 ( .A1(n6583), .A2(n6964), .ZN(U3175) );
  AND2_X1 U7450 ( .A1(n6580), .A2(DATAWIDTH_REG_6__SCAN_IN), .ZN(U3176) );
  INV_X1 U7451 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6864) );
  NOR2_X1 U7452 ( .A1(n6583), .A2(n6864), .ZN(U3177) );
  INV_X1 U7453 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U7454 ( .A1(n6583), .A2(n6899), .ZN(U3178) );
  INV_X1 U7455 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6897) );
  NOR2_X1 U7456 ( .A1(n6583), .A2(n6897), .ZN(U3179) );
  INV_X1 U7457 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U7458 ( .A1(n6583), .A2(n6945), .ZN(U3180) );
  INV_X1 U7459 ( .A(n6548), .ZN(n6535) );
  NOR2_X1 U7460 ( .A1(n6896), .A2(n6915), .ZN(n6545) );
  AOI21_X1 U7461 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6545), .ZN(n6549)
         );
  INV_X1 U7462 ( .A(HOLD), .ZN(n6541) );
  NOR2_X1 U7463 ( .A1(n6915), .A2(n6541), .ZN(n6536) );
  INV_X1 U7464 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6533) );
  OAI21_X1 U7465 ( .B1(n6536), .B2(n6533), .A(n6997), .ZN(n6534) );
  OAI211_X1 U7466 ( .C1(NA_N), .C2(n6550), .A(n6844), .B(n6548), .ZN(n6543) );
  OAI211_X1 U7467 ( .C1(n6535), .C2(n6549), .A(n6534), .B(n6543), .ZN(U3181)
         );
  NOR2_X1 U7468 ( .A1(n6550), .A2(n6541), .ZN(n6540) );
  AOI21_X1 U7469 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6536), .ZN(n6539) );
  INV_X1 U7470 ( .A(n6545), .ZN(n6537) );
  OAI211_X1 U7471 ( .C1(n6540), .C2(n6539), .A(n6538), .B(n6537), .ZN(U3182)
         );
  INV_X1 U7472 ( .A(NA_N), .ZN(n6916) );
  AOI21_X1 U7473 ( .B1(n6916), .B2(READY_N), .A(n6915), .ZN(n6542) );
  AOI211_X1 U7474 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6550), .A(n6542), 
        .B(n6541), .ZN(n6544) );
  OAI21_X1 U7475 ( .B1(n6544), .B2(n6844), .A(n6543), .ZN(n6547) );
  NAND4_X1 U7476 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6545), .A4(n6916), .ZN(n6546) );
  OAI211_X1 U7477 ( .C1(n6549), .C2(n6548), .A(n6547), .B(n6546), .ZN(U3183)
         );
  NAND2_X1 U7478 ( .A1(n6998), .A2(n6550), .ZN(n6572) );
  INV_X1 U7479 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6930) );
  INV_X2 U7480 ( .A(n6997), .ZN(n6998) );
  OAI222_X1 U7481 ( .A1(n6572), .A2(n6551), .B1(n6930), .B2(n6998), .C1(n6588), 
        .C2(n6575), .ZN(U3184) );
  INV_X1 U7482 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6910) );
  OAI222_X1 U7483 ( .A1(n6575), .A2(n6551), .B1(n6910), .B2(n6998), .C1(n6553), 
        .C2(n6577), .ZN(U3185) );
  INV_X1 U7484 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6552) );
  OAI222_X1 U7485 ( .A1(n6575), .A2(n6553), .B1(n6552), .B2(n6998), .C1(n6554), 
        .C2(n6577), .ZN(U3186) );
  INV_X1 U7486 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6730) );
  OAI222_X1 U7487 ( .A1(n6575), .A2(n6554), .B1(n6730), .B2(n6998), .C1(n6555), 
        .C2(n6577), .ZN(U3187) );
  INV_X1 U7488 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6894) );
  OAI222_X1 U7489 ( .A1(n6575), .A2(n6555), .B1(n6894), .B2(n6998), .C1(n6556), 
        .C2(n6577), .ZN(U3188) );
  INV_X1 U7490 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6907) );
  OAI222_X1 U7491 ( .A1(n6575), .A2(n6556), .B1(n6907), .B2(n6998), .C1(n6557), 
        .C2(n6577), .ZN(U3189) );
  INV_X1 U7492 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6860) );
  OAI222_X1 U7493 ( .A1(n6575), .A2(n6557), .B1(n6860), .B2(n6998), .C1(n6558), 
        .C2(n6577), .ZN(U3190) );
  INV_X1 U7494 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6723) );
  OAI222_X1 U7495 ( .A1(n6572), .A2(n6559), .B1(n6723), .B2(n6998), .C1(n6558), 
        .C2(n6575), .ZN(U3191) );
  INV_X1 U7496 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6862) );
  OAI222_X1 U7497 ( .A1(n6575), .A2(n6559), .B1(n6862), .B2(n6998), .C1(n6560), 
        .C2(n6577), .ZN(U3192) );
  INV_X1 U7498 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6973) );
  INV_X1 U7499 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6561) );
  OAI222_X1 U7500 ( .A1(n6575), .A2(n6560), .B1(n6973), .B2(n6573), .C1(n6561), 
        .C2(n6577), .ZN(U3193) );
  INV_X1 U7501 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6881) );
  OAI222_X1 U7502 ( .A1(n6575), .A2(n6561), .B1(n6881), .B2(n6998), .C1(n6562), 
        .C2(n6577), .ZN(U3194) );
  INV_X1 U7503 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6958) );
  OAI222_X1 U7504 ( .A1(n6577), .A2(n4926), .B1(n6958), .B2(n6573), .C1(n6562), 
        .C2(n6575), .ZN(U3195) );
  INV_X1 U7505 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6967) );
  INV_X1 U7506 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6564) );
  OAI222_X1 U7507 ( .A1(n6575), .A2(n4926), .B1(n6967), .B2(n6998), .C1(n6564), 
        .C2(n6577), .ZN(U3196) );
  INV_X1 U7508 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6563) );
  OAI222_X1 U7509 ( .A1(n6575), .A2(n6564), .B1(n6563), .B2(n6998), .C1(n6565), 
        .C2(n6572), .ZN(U3197) );
  INV_X1 U7510 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6841) );
  OAI222_X1 U7511 ( .A1(n6572), .A2(n5198), .B1(n6841), .B2(n6573), .C1(n6565), 
        .C2(n6575), .ZN(U3198) );
  INV_X1 U7512 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6900) );
  INV_X1 U7513 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6949) );
  OAI222_X1 U7514 ( .A1(n6575), .A2(n5198), .B1(n6900), .B2(n6573), .C1(n6949), 
        .C2(n6572), .ZN(U3199) );
  INV_X1 U7515 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6566) );
  OAI222_X1 U7516 ( .A1(n6577), .A2(n6759), .B1(n6566), .B2(n6573), .C1(n6949), 
        .C2(n6575), .ZN(U3200) );
  INV_X1 U7517 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6883) );
  OAI222_X1 U7518 ( .A1(n6575), .A2(n6759), .B1(n6883), .B2(n6573), .C1(n6746), 
        .C2(n6572), .ZN(U3201) );
  INV_X1 U7519 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6758) );
  OAI222_X1 U7520 ( .A1(n6575), .A2(n6746), .B1(n6758), .B2(n6573), .C1(n6961), 
        .C2(n6572), .ZN(U3202) );
  INV_X1 U7521 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6567) );
  OAI222_X1 U7522 ( .A1(n6575), .A2(n6961), .B1(n6567), .B2(n6998), .C1(n6568), 
        .C2(n6572), .ZN(U3203) );
  INV_X1 U7523 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6978) );
  OAI222_X1 U7524 ( .A1(n6575), .A2(n6568), .B1(n6978), .B2(n6573), .C1(n6906), 
        .C2(n6572), .ZN(U3204) );
  INV_X1 U7525 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6733) );
  OAI222_X1 U7526 ( .A1(n6575), .A2(n6906), .B1(n6733), .B2(n6998), .C1(n6569), 
        .C2(n6577), .ZN(U3205) );
  INV_X1 U7527 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6725) );
  OAI222_X1 U7528 ( .A1(n6575), .A2(n6569), .B1(n6725), .B2(n6573), .C1(n6880), 
        .C2(n6577), .ZN(U3206) );
  INV_X1 U7529 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6743) );
  OAI222_X1 U7530 ( .A1(n6572), .A2(n6571), .B1(n6743), .B2(n6998), .C1(n6880), 
        .C2(n6575), .ZN(U3207) );
  INV_X1 U7531 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6570) );
  OAI222_X1 U7532 ( .A1(n6575), .A2(n6571), .B1(n6570), .B2(n6998), .C1(n5148), 
        .C2(n6577), .ZN(U3208) );
  INV_X1 U7533 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6849) );
  OAI222_X1 U7534 ( .A1(n6575), .A2(n5148), .B1(n6849), .B2(n6998), .C1(n6846), 
        .C2(n6572), .ZN(U3209) );
  INV_X1 U7535 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6753) );
  OAI222_X1 U7536 ( .A1(n6575), .A2(n6846), .B1(n6753), .B2(n6998), .C1(n6952), 
        .C2(n6572), .ZN(U3210) );
  INV_X1 U7537 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6867) );
  OAI222_X1 U7538 ( .A1(n6575), .A2(n6952), .B1(n6867), .B2(n6998), .C1(n4413), 
        .C2(n6577), .ZN(U3211) );
  INV_X1 U7539 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6574) );
  OAI222_X1 U7540 ( .A1(n6575), .A2(n4413), .B1(n6574), .B2(n6573), .C1(n6576), 
        .C2(n6577), .ZN(U3212) );
  INV_X1 U7541 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6929) );
  INV_X1 U7542 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6706) );
  OAI222_X1 U7543 ( .A1(n6577), .A2(n6929), .B1(n6706), .B2(n6998), .C1(n6576), 
        .C2(n6575), .ZN(U3213) );
  INV_X1 U7544 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6951) );
  INV_X1 U7545 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U7546 ( .A1(n6998), .A2(n6951), .B1(n6578), .B2(n6997), .ZN(U3446)
         );
  INV_X1 U7547 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6868) );
  AOI22_X1 U7548 ( .A1(n6998), .A2(n6963), .B1(n6868), .B2(n6997), .ZN(U3447)
         );
  INV_X1 U7549 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6976) );
  INV_X1 U7550 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6966) );
  AOI22_X1 U7551 ( .A1(n6998), .A2(n6976), .B1(n6966), .B2(n6997), .ZN(U3448)
         );
  INV_X1 U7552 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6581) );
  INV_X1 U7553 ( .A(n6582), .ZN(n6579) );
  AOI21_X1 U7554 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(U3451) );
  OAI21_X1 U7555 ( .B1(n6583), .B2(n6927), .A(n6582), .ZN(U3452) );
  AOI211_X1 U7556 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6586), .A(n6585), .B(
        n6584), .ZN(n6587) );
  INV_X1 U7557 ( .A(n6587), .ZN(U3453) );
  AOI21_X1 U7558 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6589) );
  AOI22_X1 U7559 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6589), .B2(n6588), .ZN(n6591) );
  AOI22_X1 U7560 ( .A1(n6593), .A2(n6591), .B1(n6951), .B2(n6590), .ZN(U3468)
         );
  OAI21_X1 U7561 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6593), .ZN(n6592) );
  OAI21_X1 U7562 ( .B1(n6593), .B2(n6976), .A(n6592), .ZN(U3469) );
  INV_X1 U7563 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6893) );
  AOI22_X1 U7564 ( .A1(n6998), .A2(READREQUEST_REG_SCAN_IN), .B1(n6893), .B2(
        n6997), .ZN(U3470) );
  INV_X1 U7565 ( .A(n6594), .ZN(n6595) );
  AOI211_X1 U7566 ( .C1(n6597), .C2(n6596), .A(n6251), .B(n6595), .ZN(n6600)
         );
  OAI21_X1 U7567 ( .B1(n6600), .B2(n6599), .A(n6598), .ZN(n6606) );
  AND2_X1 U7568 ( .A1(n6896), .A2(n4833), .ZN(n6601) );
  NOR4_X1 U7569 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6605)
         );
  MUX2_X1 U7570 ( .A(n6606), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6605), .Z(
        U3472) );
  INV_X1 U7571 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6780) );
  INV_X1 U7572 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6850) );
  AOI22_X1 U7573 ( .A1(n6998), .A2(n6780), .B1(n6850), .B2(n6997), .ZN(U3473)
         );
  OAI22_X1 U7574 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(keyinput_f80), .ZN(n6607) );
  AOI221_X1 U7575 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(keyinput_f80), .C2(
        ADDRESS_REG_20__SCAN_IN), .A(n6607), .ZN(n6613) );
  OAI22_X1 U7576 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(keyinput_f76), .ZN(n6608) );
  AOI221_X1 U7577 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f76), .C2(ADDRESS_REG_24__SCAN_IN), .A(n6608), .ZN(n6612) );
  OAI22_X1 U7578 ( .A1(keyinput_f87), .A2(ADDRESS_REG_13__SCAN_IN), .B1(
        keyinput_f127), .B2(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6609) );
  AOI221_X1 U7579 ( .B1(keyinput_f87), .B2(ADDRESS_REG_13__SCAN_IN), .C1(
        DATAWIDTH_REG_23__SCAN_IN), .C2(keyinput_f127), .A(n6609), .ZN(n6611)
         );
  XNOR2_X1 U7580 ( .A(ADDRESS_REG_5__SCAN_IN), .B(keyinput_f95), .ZN(n6610) );
  NAND4_X1 U7581 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .ZN(n6641)
         );
  OAI22_X1 U7582 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(BE_N_REG_1__SCAN_IN), 
        .B2(keyinput_f69), .ZN(n6614) );
  AOI221_X1 U7583 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(keyinput_f69), .C2(
        BE_N_REG_1__SCAN_IN), .A(n6614), .ZN(n6621) );
  OAI22_X1 U7584 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f42), .B1(
        M_IO_N_REG_SCAN_IN), .B2(keyinput_f40), .ZN(n6615) );
  AOI221_X1 U7585 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .C1(
        keyinput_f40), .C2(M_IO_N_REG_SCAN_IN), .A(n6615), .ZN(n6620) );
  OAI22_X1 U7586 ( .A1(DATAI_14_), .A2(keyinput_f17), .B1(keyinput_f112), .B2(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n6616) );
  AOI221_X1 U7587 ( .B1(DATAI_14_), .B2(keyinput_f17), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput_f112), .A(n6616), .ZN(n6619)
         );
  OAI22_X1 U7588 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(keyinput_f118), .B2(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6617) );
  AOI221_X1 U7589 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(
        DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput_f118), .A(n6617), .ZN(n6618)
         );
  NAND4_X1 U7590 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6640)
         );
  OAI22_X1 U7591 ( .A1(keyinput_f110), .A2(DATAWIDTH_REG_6__SCAN_IN), .B1(
        keyinput_f98), .B2(ADDRESS_REG_2__SCAN_IN), .ZN(n6622) );
  AOI221_X1 U7592 ( .B1(keyinput_f110), .B2(DATAWIDTH_REG_6__SCAN_IN), .C1(
        ADDRESS_REG_2__SCAN_IN), .C2(keyinput_f98), .A(n6622), .ZN(n6629) );
  OAI22_X1 U7593 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(keyinput_f96), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n6623) );
  AOI221_X1 U7594 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(
        ADDRESS_REG_4__SCAN_IN), .C2(keyinput_f96), .A(n6623), .ZN(n6628) );
  OAI22_X1 U7595 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_f57), .B1(
        keyinput_f84), .B2(ADDRESS_REG_16__SCAN_IN), .ZN(n6624) );
  AOI221_X1 U7596 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .C1(
        ADDRESS_REG_16__SCAN_IN), .C2(keyinput_f84), .A(n6624), .ZN(n6627) );
  OAI22_X1 U7597 ( .A1(keyinput_f119), .A2(DATAWIDTH_REG_15__SCAN_IN), .B1(
        keyinput_f122), .B2(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6625) );
  AOI221_X1 U7598 ( .B1(keyinput_f119), .B2(DATAWIDTH_REG_15__SCAN_IN), .C1(
        DATAWIDTH_REG_18__SCAN_IN), .C2(keyinput_f122), .A(n6625), .ZN(n6626)
         );
  NAND4_X1 U7599 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n6639)
         );
  OAI22_X1 U7600 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f104), .B2(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6630) );
  AOI221_X1 U7601 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput_f104), .A(n6630), .ZN(n6637)
         );
  OAI22_X1 U7602 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(keyinput_f5), .B2(
        DATAI_26_), .ZN(n6631) );
  AOI221_X1 U7603 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(DATAI_26_), .C2(
        keyinput_f5), .A(n6631), .ZN(n6636) );
  OAI22_X1 U7604 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_f52), .B1(
        keyinput_f125), .B2(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6632) );
  AOI221_X1 U7605 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput_f125), .A(n6632), .ZN(n6635)
         );
  OAI22_X1 U7606 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(keyinput_f72), .ZN(n6633) );
  AOI221_X1 U7607 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(keyinput_f72), .C2(
        ADDRESS_REG_28__SCAN_IN), .A(n6633), .ZN(n6634) );
  NAND4_X1 U7608 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6638)
         );
  NOR4_X1 U7609 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n6775)
         );
  OAI22_X1 U7610 ( .A1(READY_N), .A2(keyinput_f35), .B1(keyinput_f83), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n6642) );
  AOI221_X1 U7611 ( .B1(READY_N), .B2(keyinput_f35), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput_f83), .A(n6642), .ZN(n6649) );
  OAI22_X1 U7612 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_f61), .B1(DATAI_11_), .B2(keyinput_f20), .ZN(n6643) );
  AOI221_X1 U7613 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .C1(
        keyinput_f20), .C2(DATAI_11_), .A(n6643), .ZN(n6648) );
  OAI22_X1 U7614 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(
        DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput_f108), .ZN(n6644) );
  AOI221_X1 U7615 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(keyinput_f108), 
        .C2(DATAWIDTH_REG_4__SCAN_IN), .A(n6644), .ZN(n6647) );
  OAI22_X1 U7616 ( .A1(keyinput_f99), .A2(ADDRESS_REG_1__SCAN_IN), .B1(
        keyinput_f90), .B2(ADDRESS_REG_10__SCAN_IN), .ZN(n6645) );
  AOI221_X1 U7617 ( .B1(keyinput_f99), .B2(ADDRESS_REG_1__SCAN_IN), .C1(
        ADDRESS_REG_10__SCAN_IN), .C2(keyinput_f90), .A(n6645), .ZN(n6646) );
  NAND4_X1 U7618 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6677)
         );
  OAI22_X1 U7619 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(keyinput_f81), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n6650) );
  AOI221_X1 U7620 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(
        ADDRESS_REG_19__SCAN_IN), .C2(keyinput_f81), .A(n6650), .ZN(n6657) );
  OAI22_X1 U7621 ( .A1(keyinput_f111), .A2(DATAWIDTH_REG_7__SCAN_IN), .B1(
        keyinput_f126), .B2(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6651) );
  AOI221_X1 U7622 ( .B1(keyinput_f111), .B2(DATAWIDTH_REG_7__SCAN_IN), .C1(
        DATAWIDTH_REG_22__SCAN_IN), .C2(keyinput_f126), .A(n6651), .ZN(n6656)
         );
  OAI22_X1 U7623 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(D_C_N_REG_SCAN_IN), 
        .B2(keyinput_f41), .ZN(n6652) );
  AOI221_X1 U7624 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(keyinput_f41), .C2(
        D_C_N_REG_SCAN_IN), .A(n6652), .ZN(n6655) );
  OAI22_X1 U7625 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(DATAI_7_), .B2(keyinput_f24), .ZN(n6653) );
  AOI221_X1 U7626 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f24), .C2(DATAI_7_), .A(n6653), .ZN(n6654) );
  NAND4_X1 U7627 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6676)
         );
  OAI22_X1 U7628 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(
        READREQUEST_REG_SCAN_IN), .B2(keyinput_f37), .ZN(n6658) );
  AOI221_X1 U7629 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(keyinput_f37), .C2(
        READREQUEST_REG_SCAN_IN), .A(n6658), .ZN(n6665) );
  OAI22_X1 U7630 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(
        DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_f124), .ZN(n6659) );
  AOI221_X1 U7631 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(keyinput_f124), 
        .C2(DATAWIDTH_REG_20__SCAN_IN), .A(n6659), .ZN(n6664) );
  OAI22_X1 U7632 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_f59), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_f121), .ZN(n6660) );
  AOI221_X1 U7633 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_f59), .C1(
        keyinput_f121), .C2(DATAWIDTH_REG_17__SCAN_IN), .A(n6660), .ZN(n6663)
         );
  OAI22_X1 U7634 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(keyinput_f38), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6661) );
  AOI221_X1 U7635 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(ADS_N_REG_SCAN_IN), 
        .C2(keyinput_f38), .A(n6661), .ZN(n6662) );
  NAND4_X1 U7636 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6675)
         );
  OAI22_X1 U7637 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(keyinput_f86), .ZN(n6666) );
  AOI221_X1 U7638 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(keyinput_f86), .C2(
        ADDRESS_REG_14__SCAN_IN), .A(n6666), .ZN(n6673) );
  OAI22_X1 U7639 ( .A1(keyinput_f85), .A2(ADDRESS_REG_15__SCAN_IN), .B1(
        keyinput_f34), .B2(BS16_N), .ZN(n6667) );
  AOI221_X1 U7640 ( .B1(keyinput_f85), .B2(ADDRESS_REG_15__SCAN_IN), .C1(
        BS16_N), .C2(keyinput_f34), .A(n6667), .ZN(n6672) );
  OAI22_X1 U7641 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(BE_N_REG_2__SCAN_IN), 
        .B2(keyinput_f68), .ZN(n6668) );
  AOI221_X1 U7642 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(keyinput_f68), .C2(
        BE_N_REG_2__SCAN_IN), .A(n6668), .ZN(n6671) );
  OAI22_X1 U7643 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f89), .B2(ADDRESS_REG_11__SCAN_IN), .ZN(n6669) );
  AOI221_X1 U7644 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_f101), .C1(
        ADDRESS_REG_11__SCAN_IN), .C2(keyinput_f89), .A(n6669), .ZN(n6670) );
  NAND4_X1 U7645 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .ZN(n6674)
         );
  NOR4_X1 U7646 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6774)
         );
  OAI22_X1 U7647 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(DATAI_5_), .B2(
        keyinput_f26), .ZN(n6678) );
  AOI221_X1 U7648 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(keyinput_f26), .C2(
        DATAI_5_), .A(n6678), .ZN(n6685) );
  OAI22_X1 U7649 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(keyinput_f47), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6679) );
  AOI221_X1 U7650 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_f47), .A(n6679), .ZN(n6684)
         );
  OAI22_X1 U7651 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(keyinput_f123), .B2(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6680) );
  AOI221_X1 U7652 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput_f123), .A(n6680), .ZN(n6683)
         );
  OAI22_X1 U7653 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(keyinput_f116), .B2(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n6681) );
  AOI221_X1 U7654 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(keyinput_f116), .A(n6681), .ZN(n6682)
         );
  NAND4_X1 U7655 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6719)
         );
  AOI22_X1 U7656 ( .A1(keyinput_f115), .A2(DATAWIDTH_REG_11__SCAN_IN), .B1(
        REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .ZN(n6686) );
  OAI221_X1 U7657 ( .B1(keyinput_f115), .B2(DATAWIDTH_REG_11__SCAN_IN), .C1(
        REIP_REG_17__SCAN_IN), .C2(keyinput_f65), .A(n6686), .ZN(n6718) );
  OAI22_X1 U7658 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f30), .B2(DATAI_1_), .ZN(n6687) );
  AOI221_X1 U7659 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_f66), .C1(DATAI_1_), .C2(keyinput_f30), .A(n6687), .ZN(n6692) );
  OAI22_X1 U7660 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_f117), .ZN(n6688) );
  AOI221_X1 U7661 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f117), .C2(DATAWIDTH_REG_13__SCAN_IN), .A(n6688), .ZN(n6691)
         );
  XNOR2_X1 U7662 ( .A(keyinput_f67), .B(BE_N_REG_3__SCAN_IN), .ZN(n6690) );
  XNOR2_X1 U7663 ( .A(keyinput_f36), .B(HOLD), .ZN(n6689) );
  NAND4_X1 U7664 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6717)
         );
  OAI22_X1 U7665 ( .A1(keyinput_f50), .A2(n6694), .B1(n6867), .B2(keyinput_f73), .ZN(n6693) );
  AOI221_X1 U7666 ( .B1(n6694), .B2(keyinput_f50), .C1(n6867), .C2(
        keyinput_f73), .A(n6693), .ZN(n6715) );
  AOI22_X1 U7667 ( .A1(n6973), .A2(keyinput_f91), .B1(n6909), .B2(keyinput_f25), .ZN(n6695) );
  OAI221_X1 U7668 ( .B1(n6973), .B2(keyinput_f91), .C1(n6909), .C2(
        keyinput_f25), .A(n6695), .ZN(n6703) );
  INV_X1 U7669 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6697) );
  AOI22_X1 U7670 ( .A1(n6698), .A2(keyinput_f16), .B1(keyinput_f39), .B2(n6697), .ZN(n6696) );
  OAI221_X1 U7671 ( .B1(n6698), .B2(keyinput_f16), .C1(n6697), .C2(
        keyinput_f39), .A(n6696), .ZN(n6702) );
  INV_X1 U7672 ( .A(DATAI_27_), .ZN(n6700) );
  AOI22_X1 U7673 ( .A1(n6700), .A2(keyinput_f4), .B1(keyinput_f21), .B2(n6865), 
        .ZN(n6699) );
  OAI221_X1 U7674 ( .B1(n6700), .B2(keyinput_f4), .C1(n6865), .C2(keyinput_f21), .A(n6699), .ZN(n6701) );
  NOR3_X1 U7675 ( .A1(n6703), .A2(n6702), .A3(n6701), .ZN(n6714) );
  OAI22_X1 U7676 ( .A1(n6906), .A2(keyinput_f60), .B1(n6860), .B2(keyinput_f94), .ZN(n6704) );
  AOI221_X1 U7677 ( .B1(n6906), .B2(keyinput_f60), .C1(keyinput_f94), .C2(
        n6860), .A(n6704), .ZN(n6713) );
  XOR2_X1 U7678 ( .A(keyinput_f109), .B(DATAWIDTH_REG_5__SCAN_IN), .Z(n6711)
         );
  XOR2_X1 U7679 ( .A(keyinput_f33), .B(NA_N), .Z(n6710) );
  INV_X1 U7680 ( .A(DATAI_21_), .ZN(n6936) );
  AOI22_X1 U7681 ( .A1(n6706), .A2(keyinput_f71), .B1(n6936), .B2(keyinput_f10), .ZN(n6705) );
  OAI221_X1 U7682 ( .B1(n6706), .B2(keyinput_f71), .C1(n6936), .C2(
        keyinput_f10), .A(n6705), .ZN(n6709) );
  AOI22_X1 U7683 ( .A1(n6849), .A2(keyinput_f75), .B1(n6961), .B2(keyinput_f62), .ZN(n6707) );
  OAI221_X1 U7684 ( .B1(n6849), .B2(keyinput_f75), .C1(n6961), .C2(
        keyinput_f62), .A(n6707), .ZN(n6708) );
  NOR4_X1 U7685 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n6712)
         );
  NAND4_X1 U7686 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6716)
         );
  NOR4_X1 U7687 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6773)
         );
  INV_X1 U7688 ( .A(DATAI_20_), .ZN(n6878) );
  INV_X1 U7689 ( .A(keyinput_f107), .ZN(n6721) );
  AOI22_X1 U7690 ( .A1(n6878), .A2(keyinput_f11), .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(n6721), .ZN(n6720) );
  OAI221_X1 U7691 ( .B1(n6878), .B2(keyinput_f11), .C1(n6721), .C2(
        DATAWIDTH_REG_3__SCAN_IN), .A(n6720), .ZN(n6771) );
  INV_X1 U7692 ( .A(DATAI_23_), .ZN(n6960) );
  AOI22_X1 U7693 ( .A1(n6723), .A2(keyinput_f93), .B1(n6960), .B2(keyinput_f8), 
        .ZN(n6722) );
  OAI221_X1 U7694 ( .B1(n6723), .B2(keyinput_f93), .C1(n6960), .C2(keyinput_f8), .A(n6722), .ZN(n6770) );
  OAI22_X1 U7695 ( .A1(n6725), .A2(keyinput_f78), .B1(n6963), .B2(keyinput_f48), .ZN(n6724) );
  AOI221_X1 U7696 ( .B1(n6725), .B2(keyinput_f78), .C1(keyinput_f48), .C2(
        n6963), .A(n6724), .ZN(n6728) );
  XOR2_X1 U7697 ( .A(keyinput_f106), .B(DATAWIDTH_REG_2__SCAN_IN), .Z(n6726)
         );
  AOI21_X1 U7698 ( .B1(keyinput_f120), .B2(n6913), .A(n6726), .ZN(n6727) );
  OAI211_X1 U7699 ( .C1(keyinput_f120), .C2(n6913), .A(n6728), .B(n6727), .ZN(
        n6769) );
  AOI22_X1 U7700 ( .A1(n6967), .A2(keyinput_f88), .B1(keyinput_f97), .B2(n6730), .ZN(n6729) );
  OAI221_X1 U7701 ( .B1(n6967), .B2(keyinput_f88), .C1(n6730), .C2(
        keyinput_f97), .A(n6729), .ZN(n6740) );
  INV_X1 U7702 ( .A(keyinput_f114), .ZN(n6732) );
  AOI22_X1 U7703 ( .A1(n6733), .A2(keyinput_f79), .B1(
        DATAWIDTH_REG_10__SCAN_IN), .B2(n6732), .ZN(n6731) );
  OAI221_X1 U7704 ( .B1(n6733), .B2(keyinput_f79), .C1(n6732), .C2(
        DATAWIDTH_REG_10__SCAN_IN), .A(n6731), .ZN(n6739) );
  AOI22_X1 U7705 ( .A1(n6893), .A2(keyinput_f46), .B1(n5148), .B2(keyinput_f56), .ZN(n6734) );
  OAI221_X1 U7706 ( .B1(n6893), .B2(keyinput_f46), .C1(n5148), .C2(
        keyinput_f56), .A(n6734), .ZN(n6738) );
  INV_X1 U7707 ( .A(keyinput_f49), .ZN(n6736) );
  AOI22_X1 U7708 ( .A1(n6846), .A2(keyinput_f55), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(n6736), .ZN(n6735) );
  OAI221_X1 U7709 ( .B1(n6846), .B2(keyinput_f55), .C1(n6736), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n6735), .ZN(n6737) );
  NOR4_X1 U7710 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6767)
         );
  INV_X1 U7711 ( .A(DATAI_17_), .ZN(n6742) );
  AOI22_X1 U7712 ( .A1(n6743), .A2(keyinput_f77), .B1(n6742), .B2(keyinput_f14), .ZN(n6741) );
  OAI221_X1 U7713 ( .B1(n6743), .B2(keyinput_f77), .C1(n6742), .C2(
        keyinput_f14), .A(n6741), .ZN(n6751) );
  AOI22_X1 U7714 ( .A1(n6843), .A2(keyinput_f45), .B1(keyinput_f105), .B2(
        n6927), .ZN(n6744) );
  OAI221_X1 U7715 ( .B1(n6843), .B2(keyinput_f45), .C1(n6927), .C2(
        keyinput_f105), .A(n6744), .ZN(n6750) );
  AOI22_X1 U7716 ( .A1(n6746), .A2(keyinput_f63), .B1(keyinput_f100), .B2(
        n6930), .ZN(n6745) );
  OAI221_X1 U7717 ( .B1(n6746), .B2(keyinput_f63), .C1(n6930), .C2(
        keyinput_f100), .A(n6745), .ZN(n6749) );
  AOI22_X1 U7718 ( .A1(n6915), .A2(keyinput_f102), .B1(n6844), .B2(
        keyinput_f103), .ZN(n6747) );
  OAI221_X1 U7719 ( .B1(n6915), .B2(keyinput_f102), .C1(n6844), .C2(
        keyinput_f103), .A(n6747), .ZN(n6748) );
  NOR4_X1 U7720 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6766)
         );
  OAI22_X1 U7721 ( .A1(keyinput_f113), .A2(n6754), .B1(n6753), .B2(
        keyinput_f74), .ZN(n6752) );
  AOI221_X1 U7722 ( .B1(n6754), .B2(keyinput_f113), .C1(n6753), .C2(
        keyinput_f74), .A(n6752), .ZN(n6765) );
  INV_X1 U7723 ( .A(MORE_REG_SCAN_IN), .ZN(n6756) );
  AOI22_X1 U7724 ( .A1(n6756), .A2(keyinput_f44), .B1(n6952), .B2(keyinput_f54), .ZN(n6755) );
  OAI221_X1 U7725 ( .B1(n6756), .B2(keyinput_f44), .C1(n6952), .C2(
        keyinput_f54), .A(n6755), .ZN(n6763) );
  AOI22_X1 U7726 ( .A1(n6759), .A2(keyinput_f64), .B1(keyinput_f82), .B2(n6758), .ZN(n6757) );
  OAI221_X1 U7727 ( .B1(n6759), .B2(keyinput_f64), .C1(n6758), .C2(
        keyinput_f82), .A(n6757), .ZN(n6762) );
  AOI22_X1 U7728 ( .A1(n6966), .A2(keyinput_f70), .B1(keyinput_f92), .B2(n6862), .ZN(n6760) );
  OAI221_X1 U7729 ( .B1(n6966), .B2(keyinput_f70), .C1(n6862), .C2(
        keyinput_f92), .A(n6760), .ZN(n6761) );
  NOR3_X1 U7730 ( .A1(n6763), .A2(n6762), .A3(n6761), .ZN(n6764) );
  NAND4_X1 U7731 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6768)
         );
  NOR4_X1 U7732 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6772)
         );
  NAND4_X1 U7733 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6777)
         );
  AOI21_X1 U7734 ( .B1(keyinput_f32), .B2(n6777), .A(keyinput_g32), .ZN(n6779)
         );
  INV_X1 U7735 ( .A(keyinput_f32), .ZN(n6776) );
  AOI21_X1 U7736 ( .B1(n6777), .B2(n6776), .A(n6780), .ZN(n6778) );
  AOI22_X1 U7737 ( .A1(n6780), .A2(n6779), .B1(keyinput_g32), .B2(n6778), .ZN(
        n6996) );
  XOR2_X1 U7738 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_g74), .Z(n6787) );
  AOI22_X1 U7739 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(keyinput_g71), .B1(
        DATAI_8_), .B2(keyinput_g23), .ZN(n6781) );
  OAI221_X1 U7740 ( .B1(ADDRESS_REG_29__SCAN_IN), .B2(keyinput_g71), .C1(
        DATAI_8_), .C2(keyinput_g23), .A(n6781), .ZN(n6786) );
  AOI22_X1 U7741 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput_g124), .B1(
        DATAI_12_), .B2(keyinput_g19), .ZN(n6782) );
  OAI221_X1 U7742 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_g124), .C1(
        DATAI_12_), .C2(keyinput_g19), .A(n6782), .ZN(n6785) );
  AOI22_X1 U7743 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6783) );
  OAI221_X1 U7744 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6783), .ZN(n6784) );
  NOR4_X1 U7745 ( .A1(n6787), .A2(n6786), .A3(n6785), .A4(n6784), .ZN(n6815)
         );
  AOI22_X1 U7746 ( .A1(ADDRESS_REG_2__SCAN_IN), .A2(keyinput_g98), .B1(
        DATAI_0_), .B2(keyinput_g31), .ZN(n6788) );
  OAI221_X1 U7747 ( .B1(ADDRESS_REG_2__SCAN_IN), .B2(keyinput_g98), .C1(
        DATAI_0_), .C2(keyinput_g31), .A(n6788), .ZN(n6795) );
  AOI22_X1 U7748 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput_g77), .B1(
        DATAI_27_), .B2(keyinput_g4), .ZN(n6789) );
  OAI221_X1 U7749 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput_g77), .C1(
        DATAI_27_), .C2(keyinput_g4), .A(n6789), .ZN(n6794) );
  AOI22_X1 U7750 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(DATAI_2_), .B2(
        keyinput_g29), .ZN(n6790) );
  OAI221_X1 U7751 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n6790), .ZN(n6793) );
  AOI22_X1 U7752 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(STATE_REG_2__SCAN_IN), 
        .B2(keyinput_g101), .ZN(n6791) );
  OAI221_X1 U7753 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(STATE_REG_2__SCAN_IN), .C2(keyinput_g101), .A(n6791), .ZN(n6792) );
  NOR4_X1 U7754 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6814)
         );
  AOI22_X1 U7755 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput_g122), .B1(
        DATAI_3_), .B2(keyinput_g28), .ZN(n6796) );
  OAI221_X1 U7756 ( .B1(DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_g122), .C1(
        DATAI_3_), .C2(keyinput_g28), .A(n6796), .ZN(n6803) );
  AOI22_X1 U7757 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(keyinput_g87), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n6797) );
  OAI221_X1 U7758 ( .B1(ADDRESS_REG_13__SCAN_IN), .B2(keyinput_g87), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g42), .A(n6797), .ZN(n6802)
         );
  AOI22_X1 U7759 ( .A1(HOLD), .A2(keyinput_g36), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n6798) );
  OAI221_X1 U7760 ( .B1(HOLD), .B2(keyinput_g36), .C1(REIP_REG_19__SCAN_IN), 
        .C2(keyinput_g63), .A(n6798), .ZN(n6801) );
  AOI22_X1 U7761 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(REIP_REG_25__SCAN_IN), 
        .B2(keyinput_g57), .ZN(n6799) );
  OAI221_X1 U7762 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6799), .ZN(n6800) );
  NOR4_X1 U7763 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6813)
         );
  AOI22_X1 U7764 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput_g117), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_g112), .ZN(n6804) );
  OAI221_X1 U7765 ( .B1(DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_g117), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput_g112), .A(n6804), .ZN(n6811)
         );
  AOI22_X1 U7766 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        REIP_REG_18__SCAN_IN), .B2(keyinput_g64), .ZN(n6805) );
  OAI221_X1 U7767 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        REIP_REG_18__SCAN_IN), .C2(keyinput_g64), .A(n6805), .ZN(n6810) );
  AOI22_X1 U7768 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .ZN(n6806) );
  OAI221_X1 U7769 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6806), .ZN(n6809) );
  AOI22_X1 U7770 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(keyinput_g125), .B1(
        DATAI_16_), .B2(keyinput_g15), .ZN(n6807) );
  OAI221_X1 U7771 ( .B1(DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_g125), .C1(
        DATAI_16_), .C2(keyinput_g15), .A(n6807), .ZN(n6808) );
  NOR4_X1 U7772 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6812)
         );
  NAND4_X1 U7773 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6994)
         );
  AOI22_X1 U7774 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput_g76), .B1(
        DATAI_13_), .B2(keyinput_g18), .ZN(n6816) );
  OAI221_X1 U7775 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput_g76), .C1(
        DATAI_13_), .C2(keyinput_g18), .A(n6816), .ZN(n6823) );
  AOI22_X1 U7776 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(keyinput_g81), .ZN(n6817) );
  OAI221_X1 U7777 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        ADDRESS_REG_19__SCAN_IN), .C2(keyinput_g81), .A(n6817), .ZN(n6822) );
  AOI22_X1 U7778 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput_g84), .B1(
        DATAI_15_), .B2(keyinput_g16), .ZN(n6818) );
  OAI221_X1 U7779 ( .B1(ADDRESS_REG_16__SCAN_IN), .B2(keyinput_g84), .C1(
        DATAI_15_), .C2(keyinput_g16), .A(n6818), .ZN(n6821) );
  AOI22_X1 U7780 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_31_), .B2(
        keyinput_g0), .ZN(n6819) );
  OAI221_X1 U7781 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(DATAI_31_), .C2(
        keyinput_g0), .A(n6819), .ZN(n6820) );
  NOR4_X1 U7782 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6858)
         );
  AOI22_X1 U7783 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput_g93), .B1(
        DATAI_5_), .B2(keyinput_g26), .ZN(n6824) );
  OAI221_X1 U7784 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput_g93), .C1(
        DATAI_5_), .C2(keyinput_g26), .A(n6824), .ZN(n6831) );
  AOI22_X1 U7785 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput_g110), .B1(
        DATAI_14_), .B2(keyinput_g17), .ZN(n6825) );
  OAI221_X1 U7786 ( .B1(DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_g110), .C1(
        DATAI_14_), .C2(keyinput_g17), .A(n6825), .ZN(n6830) );
  AOI22_X1 U7787 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(keyinput_g126), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6826) );
  OAI221_X1 U7788 ( .B1(DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput_g126), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6826), .ZN(n6829) );
  AOI22_X1 U7789 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(keyinput_g113), .B1(
        DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_g123), .ZN(n6827) );
  OAI221_X1 U7790 ( .B1(DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput_g113), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput_g123), .A(n6827), .ZN(n6828)
         );
  NOR4_X1 U7791 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n6857)
         );
  AOI22_X1 U7792 ( .A1(BE_N_REG_2__SCAN_IN), .A2(keyinput_g68), .B1(
        DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .ZN(n6832) );
  OAI221_X1 U7793 ( .B1(BE_N_REG_2__SCAN_IN), .B2(keyinput_g68), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput_g104), .A(n6832), .ZN(n6839)
         );
  AOI22_X1 U7794 ( .A1(ADDRESS_REG_3__SCAN_IN), .A2(keyinput_g97), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(keyinput_g78), .ZN(n6833) );
  OAI221_X1 U7795 ( .B1(ADDRESS_REG_3__SCAN_IN), .B2(keyinput_g97), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput_g78), .A(n6833), .ZN(n6838) );
  AOI22_X1 U7796 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(keyinput_g72), .B1(
        DATAI_9_), .B2(keyinput_g22), .ZN(n6834) );
  OAI221_X1 U7797 ( .B1(ADDRESS_REG_28__SCAN_IN), .B2(keyinput_g72), .C1(
        DATAI_9_), .C2(keyinput_g22), .A(n6834), .ZN(n6837) );
  AOI22_X1 U7798 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput_g79), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_g52), .ZN(n6835) );
  OAI221_X1 U7799 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput_g79), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_g52), .A(n6835), .ZN(n6836) );
  NOR4_X1 U7800 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6856)
         );
  AOI22_X1 U7801 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput_g82), .B1(n6841), 
        .B2(keyinput_g86), .ZN(n6840) );
  OAI221_X1 U7802 ( .B1(ADDRESS_REG_18__SCAN_IN), .B2(keyinput_g82), .C1(n6841), .C2(keyinput_g86), .A(n6840), .ZN(n6854) );
  AOI22_X1 U7803 ( .A1(n6844), .A2(keyinput_g103), .B1(keyinput_g45), .B2(
        n6843), .ZN(n6842) );
  OAI221_X1 U7804 ( .B1(n6844), .B2(keyinput_g103), .C1(n6843), .C2(
        keyinput_g45), .A(n6842), .ZN(n6853) );
  AOI22_X1 U7805 ( .A1(n6847), .A2(keyinput_g38), .B1(n6846), .B2(keyinput_g55), .ZN(n6845) );
  OAI221_X1 U7806 ( .B1(n6847), .B2(keyinput_g38), .C1(n6846), .C2(
        keyinput_g55), .A(n6845), .ZN(n6852) );
  AOI22_X1 U7807 ( .A1(n6850), .A2(keyinput_g40), .B1(keyinput_g75), .B2(n6849), .ZN(n6848) );
  OAI221_X1 U7808 ( .B1(n6850), .B2(keyinput_g40), .C1(n6849), .C2(
        keyinput_g75), .A(n6848), .ZN(n6851) );
  NOR4_X1 U7809 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6855)
         );
  NAND4_X1 U7810 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6993)
         );
  AOI22_X1 U7811 ( .A1(n6860), .A2(keyinput_g94), .B1(n5198), .B2(keyinput_g66), .ZN(n6859) );
  OAI221_X1 U7812 ( .B1(n6860), .B2(keyinput_g94), .C1(n5198), .C2(
        keyinput_g66), .A(n6859), .ZN(n6872) );
  AOI22_X1 U7813 ( .A1(n6862), .A2(keyinput_g92), .B1(n5675), .B2(keyinput_g13), .ZN(n6861) );
  OAI221_X1 U7814 ( .B1(n6862), .B2(keyinput_g92), .C1(n5675), .C2(
        keyinput_g13), .A(n6861), .ZN(n6871) );
  AOI22_X1 U7815 ( .A1(n6865), .A2(keyinput_g21), .B1(keyinput_g109), .B2(
        n6864), .ZN(n6863) );
  OAI221_X1 U7816 ( .B1(n6865), .B2(keyinput_g21), .C1(n6864), .C2(
        keyinput_g109), .A(n6863), .ZN(n6870) );
  AOI22_X1 U7817 ( .A1(n6868), .A2(keyinput_g69), .B1(keyinput_g73), .B2(n6867), .ZN(n6866) );
  OAI221_X1 U7818 ( .B1(n6868), .B2(keyinput_g69), .C1(n6867), .C2(
        keyinput_g73), .A(n6866), .ZN(n6869) );
  NOR4_X1 U7819 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6924)
         );
  INV_X1 U7820 ( .A(DATAI_25_), .ZN(n6874) );
  AOI22_X1 U7821 ( .A1(n6875), .A2(keyinput_g41), .B1(n6874), .B2(keyinput_g6), 
        .ZN(n6873) );
  OAI221_X1 U7822 ( .B1(n6875), .B2(keyinput_g41), .C1(n6874), .C2(keyinput_g6), .A(n6873), .ZN(n6888) );
  AOI22_X1 U7823 ( .A1(n6878), .A2(keyinput_g11), .B1(n6877), .B2(keyinput_g27), .ZN(n6876) );
  OAI221_X1 U7824 ( .B1(n6878), .B2(keyinput_g11), .C1(n6877), .C2(
        keyinput_g27), .A(n6876), .ZN(n6887) );
  AOI22_X1 U7825 ( .A1(n6881), .A2(keyinput_g90), .B1(n6880), .B2(keyinput_g58), .ZN(n6879) );
  OAI221_X1 U7826 ( .B1(n6881), .B2(keyinput_g90), .C1(n6880), .C2(
        keyinput_g58), .A(n6879), .ZN(n6886) );
  INV_X1 U7827 ( .A(DATAI_22_), .ZN(n6884) );
  AOI22_X1 U7828 ( .A1(n6884), .A2(keyinput_g9), .B1(keyinput_g83), .B2(n6883), 
        .ZN(n6882) );
  OAI221_X1 U7829 ( .B1(n6884), .B2(keyinput_g9), .C1(n6883), .C2(keyinput_g83), .A(n6882), .ZN(n6885) );
  NOR4_X1 U7830 ( .A1(n6888), .A2(n6887), .A3(n6886), .A4(n6885), .ZN(n6923)
         );
  INV_X1 U7831 ( .A(DATAI_24_), .ZN(n6891) );
  AOI22_X1 U7832 ( .A1(n6891), .A2(keyinput_g7), .B1(keyinput_g119), .B2(n6890), .ZN(n6889) );
  OAI221_X1 U7833 ( .B1(n6891), .B2(keyinput_g7), .C1(n6890), .C2(
        keyinput_g119), .A(n6889), .ZN(n6904) );
  AOI22_X1 U7834 ( .A1(n6894), .A2(keyinput_g96), .B1(keyinput_g46), .B2(n6893), .ZN(n6892) );
  OAI221_X1 U7835 ( .B1(n6894), .B2(keyinput_g96), .C1(n6893), .C2(
        keyinput_g46), .A(n6892), .ZN(n6903) );
  AOI22_X1 U7836 ( .A1(n6897), .A2(keyinput_g107), .B1(n6896), .B2(
        keyinput_g35), .ZN(n6895) );
  OAI221_X1 U7837 ( .B1(n6897), .B2(keyinput_g107), .C1(n6896), .C2(
        keyinput_g35), .A(n6895), .ZN(n6902) );
  AOI22_X1 U7838 ( .A1(n6900), .A2(keyinput_g85), .B1(n6899), .B2(
        keyinput_g108), .ZN(n6898) );
  OAI221_X1 U7839 ( .B1(n6900), .B2(keyinput_g85), .C1(n6899), .C2(
        keyinput_g108), .A(n6898), .ZN(n6901) );
  NOR4_X1 U7840 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6922)
         );
  AOI22_X1 U7841 ( .A1(n6907), .A2(keyinput_g95), .B1(n6906), .B2(keyinput_g60), .ZN(n6905) );
  OAI221_X1 U7842 ( .B1(n6907), .B2(keyinput_g95), .C1(n6906), .C2(
        keyinput_g60), .A(n6905), .ZN(n6920) );
  AOI22_X1 U7843 ( .A1(n6910), .A2(keyinput_g99), .B1(n6909), .B2(keyinput_g25), .ZN(n6908) );
  OAI221_X1 U7844 ( .B1(n6910), .B2(keyinput_g99), .C1(n6909), .C2(
        keyinput_g25), .A(n6908), .ZN(n6919) );
  AOI22_X1 U7845 ( .A1(n6913), .A2(keyinput_g120), .B1(keyinput_g114), .B2(
        n6912), .ZN(n6911) );
  OAI221_X1 U7846 ( .B1(n6913), .B2(keyinput_g120), .C1(n6912), .C2(
        keyinput_g114), .A(n6911), .ZN(n6918) );
  AOI22_X1 U7847 ( .A1(n6916), .A2(keyinput_g33), .B1(n6915), .B2(
        keyinput_g102), .ZN(n6914) );
  OAI221_X1 U7848 ( .B1(n6916), .B2(keyinput_g33), .C1(n6915), .C2(
        keyinput_g102), .A(n6914), .ZN(n6917) );
  NOR4_X1 U7849 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6921)
         );
  NAND4_X1 U7850 ( .A1(n6924), .A2(n6923), .A3(n6922), .A4(n6921), .ZN(n6992)
         );
  INV_X1 U7851 ( .A(DATAI_19_), .ZN(n6926) );
  AOI22_X1 U7852 ( .A1(n6927), .A2(keyinput_g105), .B1(n6926), .B2(
        keyinput_g12), .ZN(n6925) );
  OAI221_X1 U7853 ( .B1(n6927), .B2(keyinput_g105), .C1(n6926), .C2(
        keyinput_g12), .A(n6925), .ZN(n6940) );
  AOI22_X1 U7854 ( .A1(n6930), .A2(keyinput_g100), .B1(n6929), .B2(
        keyinput_g51), .ZN(n6928) );
  OAI221_X1 U7855 ( .B1(n6930), .B2(keyinput_g100), .C1(n6929), .C2(
        keyinput_g51), .A(n6928), .ZN(n6939) );
  INV_X1 U7856 ( .A(DATAI_30_), .ZN(n6933) );
  AOI22_X1 U7857 ( .A1(n6933), .A2(keyinput_g1), .B1(keyinput_g121), .B2(n6932), .ZN(n6931) );
  OAI221_X1 U7858 ( .B1(n6933), .B2(keyinput_g1), .C1(n6932), .C2(
        keyinput_g121), .A(n6931), .ZN(n6938) );
  INV_X1 U7859 ( .A(BS16_N), .ZN(n6935) );
  AOI22_X1 U7860 ( .A1(n6936), .A2(keyinput_g10), .B1(keyinput_g34), .B2(n6935), .ZN(n6934) );
  OAI221_X1 U7861 ( .B1(n6936), .B2(keyinput_g10), .C1(n6935), .C2(
        keyinput_g34), .A(n6934), .ZN(n6937) );
  NOR4_X1 U7862 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6990)
         );
  INV_X1 U7863 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6943) );
  INV_X1 U7864 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7865 ( .A1(n6943), .A2(keyinput_g67), .B1(n6942), .B2(keyinput_g37), .ZN(n6941) );
  OAI221_X1 U7866 ( .B1(n6943), .B2(keyinput_g67), .C1(n6942), .C2(
        keyinput_g37), .A(n6941), .ZN(n6956) );
  INV_X1 U7867 ( .A(DATAI_29_), .ZN(n6946) );
  AOI22_X1 U7868 ( .A1(n6946), .A2(keyinput_g2), .B1(keyinput_g106), .B2(n6945), .ZN(n6944) );
  OAI221_X1 U7869 ( .B1(n6946), .B2(keyinput_g2), .C1(n6945), .C2(
        keyinput_g106), .A(n6944), .ZN(n6955) );
  AOI22_X1 U7870 ( .A1(n6949), .A2(keyinput_g65), .B1(keyinput_g116), .B2(
        n6948), .ZN(n6947) );
  OAI221_X1 U7871 ( .B1(n6949), .B2(keyinput_g65), .C1(n6948), .C2(
        keyinput_g116), .A(n6947), .ZN(n6954) );
  AOI22_X1 U7872 ( .A1(n6952), .A2(keyinput_g54), .B1(keyinput_g49), .B2(n6951), .ZN(n6950) );
  OAI221_X1 U7873 ( .B1(n6952), .B2(keyinput_g54), .C1(n6951), .C2(
        keyinput_g49), .A(n6950), .ZN(n6953) );
  NOR4_X1 U7874 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6989)
         );
  AOI22_X1 U7875 ( .A1(n4413), .A2(keyinput_g53), .B1(keyinput_g89), .B2(n6958), .ZN(n6957) );
  OAI221_X1 U7876 ( .B1(n4413), .B2(keyinput_g53), .C1(n6958), .C2(
        keyinput_g89), .A(n6957), .ZN(n6971) );
  AOI22_X1 U7877 ( .A1(n6961), .A2(keyinput_g62), .B1(keyinput_g8), .B2(n6960), 
        .ZN(n6959) );
  OAI221_X1 U7878 ( .B1(n6961), .B2(keyinput_g62), .C1(n6960), .C2(keyinput_g8), .A(n6959), .ZN(n6970) );
  AOI22_X1 U7879 ( .A1(n6964), .A2(keyinput_g111), .B1(keyinput_g48), .B2(
        n6963), .ZN(n6962) );
  OAI221_X1 U7880 ( .B1(n6964), .B2(keyinput_g111), .C1(n6963), .C2(
        keyinput_g48), .A(n6962), .ZN(n6969) );
  AOI22_X1 U7881 ( .A1(n6967), .A2(keyinput_g88), .B1(keyinput_g70), .B2(n6966), .ZN(n6965) );
  OAI221_X1 U7882 ( .B1(n6967), .B2(keyinput_g88), .C1(n6966), .C2(
        keyinput_g70), .A(n6965), .ZN(n6968) );
  NOR4_X1 U7883 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n6988)
         );
  AOI22_X1 U7884 ( .A1(n6974), .A2(keyinput_g118), .B1(keyinput_g91), .B2(
        n6973), .ZN(n6972) );
  OAI221_X1 U7885 ( .B1(n6974), .B2(keyinput_g118), .C1(n6973), .C2(
        keyinput_g91), .A(n6972), .ZN(n6986) );
  AOI22_X1 U7886 ( .A1(n6976), .A2(keyinput_g47), .B1(n5148), .B2(keyinput_g56), .ZN(n6975) );
  OAI221_X1 U7887 ( .B1(n6976), .B2(keyinput_g47), .C1(n5148), .C2(
        keyinput_g56), .A(n6975), .ZN(n6985) );
  AOI22_X1 U7888 ( .A1(n6979), .A2(keyinput_g127), .B1(n6978), .B2(
        keyinput_g80), .ZN(n6977) );
  OAI221_X1 U7889 ( .B1(n6979), .B2(keyinput_g127), .C1(n6978), .C2(
        keyinput_g80), .A(n6977), .ZN(n6984) );
  AOI22_X1 U7890 ( .A1(n6982), .A2(keyinput_g115), .B1(n6981), .B2(
        keyinput_g30), .ZN(n6980) );
  OAI221_X1 U7891 ( .B1(n6982), .B2(keyinput_g115), .C1(n6981), .C2(
        keyinput_g30), .A(n6980), .ZN(n6983) );
  NOR4_X1 U7892 ( .A1(n6986), .A2(n6985), .A3(n6984), .A4(n6983), .ZN(n6987)
         );
  NAND4_X1 U7893 ( .A1(n6990), .A2(n6989), .A3(n6988), .A4(n6987), .ZN(n6991)
         );
  NOR4_X1 U7894 ( .A1(n6994), .A2(n6993), .A3(n6992), .A4(n6991), .ZN(n6995)
         );
  NOR2_X1 U7895 ( .A1(n6996), .A2(n6995), .ZN(n7000) );
  AOI22_X1 U7896 ( .A1(n6998), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6997), .ZN(n6999) );
  XNOR2_X1 U7897 ( .A(n7000), .B(n6999), .ZN(U3445) );
  CLKBUF_X1 U3606 ( .A(n3827), .Z(n4181) );
  CLKBUF_X1 U3609 ( .A(n3437), .Z(n4656) );
  CLKBUF_X2 U3617 ( .A(n4618), .Z(n3155) );
  NAND4_X2 U3619 ( .A1(n3369), .A2(n3213), .A3(n3368), .A4(n3367), .ZN(n3408)
         );
  CLKBUF_X1 U3626 ( .A(n5709), .Z(n5704) );
  AOI211_X2 U3643 ( .C1(n4788), .C2(n6417), .A(n4714), .B(n6416), .ZN(n4771)
         );
  CLKBUF_X3 U3670 ( .A(n3581), .Z(n3194) );
endmodule

