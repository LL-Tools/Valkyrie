

module b22_C_gen_AntiSAT_k_128_8 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6471, n6472, n6474, n6475, n6476, n6477, n6478, n6479, n6481, n6482,
         n6483, n6484, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15308;

  INV_X1 U7219 ( .A(n13252), .ZN(n13424) );
  NOR2_X2 U7220 ( .A1(n14411), .A2(n14412), .ZN(n11619) );
  CLKBUF_X2 U7221 ( .A(n9533), .Z(n12586) );
  NAND2_X1 U7222 ( .A1(n8980), .A2(n8979), .ZN(n9293) );
  CLKBUF_X2 U7223 ( .A(n9160), .Z(n12338) );
  BUF_X2 U7224 ( .A(n9153), .Z(n12341) );
  OAI211_X1 U7225 ( .C1(SI_5_), .C2(n9165), .A(n9164), .B(n9163), .ZN(n10971)
         );
  INV_X2 U7226 ( .A(n9102), .ZN(n9279) );
  BUF_X2 U7227 ( .A(n7571), .Z(n7965) );
  XNOR2_X1 U7228 ( .A(n9091), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U7229 ( .A1(n7097), .A2(n6852), .ZN(n9053) );
  CLKBUF_X2 U7230 ( .A(n8844), .Z(n6655) );
  AND3_X1 U7231 ( .A1(n7748), .A2(n7462), .A3(n7405), .ZN(n7019) );
  XNOR2_X1 U7232 ( .A(n8142), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8552) );
  INV_X2 U7233 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8154) );
  NOR2_X1 U7234 ( .A1(n13233), .A2(n6835), .ZN(n6834) );
  CLKBUF_X2 U7235 ( .A(n8867), .Z(n6643) );
  AND2_X1 U7236 ( .A1(n8551), .A2(n11023), .ZN(n8666) );
  INV_X1 U7237 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8149) );
  INV_X1 U7238 ( .A(n9590), .ZN(n10737) );
  OR2_X1 U7239 ( .A1(n10033), .A2(n8553), .ZN(n9956) );
  INV_X1 U7240 ( .A(n10334), .ZN(n12152) );
  NAND2_X1 U7241 ( .A1(n11573), .A2(n9619), .ZN(n12230) );
  INV_X1 U7242 ( .A(n12341), .ZN(n9489) );
  INV_X1 U7243 ( .A(n6471), .ZN(n6482) );
  AND2_X1 U7244 ( .A1(n12607), .A2(n12606), .ZN(n14307) );
  INV_X1 U7245 ( .A(n12504), .ZN(n12514) );
  INV_X1 U7246 ( .A(n9382), .ZN(n12340) );
  NOR2_X1 U7247 ( .A1(n9329), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n9331) );
  INV_X1 U7248 ( .A(n9956), .ZN(n12001) );
  INV_X1 U7249 ( .A(n11854), .ZN(n8105) );
  NAND2_X2 U7250 ( .A1(n8098), .A2(n14157), .ZN(n9746) );
  INV_X1 U7251 ( .A(n13843), .ZN(n11688) );
  NAND2_X1 U7252 ( .A1(n9153), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9107) );
  XNOR2_X1 U7253 ( .A(n8550), .B(n8923), .ZN(n13216) );
  XNOR2_X1 U7254 ( .A(n7057), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7467) );
  XNOR2_X1 U7255 ( .A(n7615), .B(n7613), .ZN(n9764) );
  INV_X2 U7256 ( .A(n7495), .ZN(n9735) );
  NAND4_X1 U7257 ( .A1(n9129), .A2(n9128), .A3(n9127), .A4(n9126), .ZN(n12552)
         );
  INV_X1 U7258 ( .A(n12398), .ZN(n10709) );
  INV_X1 U7259 ( .A(n11714), .ZN(n13720) );
  INV_X2 U7260 ( .A(n14047), .ZN(n14041) );
  NAND2_X1 U7261 ( .A1(n9094), .A2(n12965), .ZN(n6471) );
  BUF_X2 U7262 ( .A(n8668), .Z(n13131) );
  NAND2_X1 U7263 ( .A1(n13254), .A2(n13253), .ZN(n13422) );
  INV_X2 U7264 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13201) );
  NAND2_X2 U7265 ( .A1(n6944), .A2(n7633), .ZN(n7648) );
  INV_X1 U7266 ( .A(n8004), .ZN(n6472) );
  NAND2_X2 U7267 ( .A1(n13995), .A2(n7865), .ZN(n13967) );
  NAND2_X2 U7268 ( .A1(n13992), .A2(n7864), .ZN(n13995) );
  XNOR2_X2 U7269 ( .A(n12053), .B(n12051), .ZN(n13690) );
  NAND2_X2 U7270 ( .A1(n14456), .A2(n6675), .ZN(n12053) );
  NAND2_X2 U7271 ( .A1(n7705), .A2(n7446), .ZN(n7707) );
  XNOR2_X2 U7272 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14217) );
  MUX2_X2 U7273 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12908), .S(n15076), .Z(
        n12909) );
  MUX2_X2 U7274 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12908), .S(n15085), .Z(
        n12851) );
  XNOR2_X2 U7275 ( .A(n13721), .B(n7516), .ZN(n11891) );
  OR2_X2 U7276 ( .A1(n10060), .A2(n12958), .ZN(n9123) );
  OR2_X2 U7277 ( .A1(n8844), .A2(n8158), .ZN(n8163) );
  NAND2_X2 U7278 ( .A1(n12667), .A2(n7445), .ZN(n9524) );
  NAND2_X2 U7279 ( .A1(n9668), .A2(n12265), .ZN(n12240) );
  NAND2_X2 U7284 ( .A1(n8203), .A2(n8202), .ZN(n10305) );
  OAI21_X2 U7285 ( .B1(n8964), .B2(n7244), .A(n7242), .ZN(n9213) );
  NOR2_X2 U7286 ( .A1(n8134), .A2(n8133), .ZN(n8551) );
  NAND2_X2 U7287 ( .A1(n8141), .A2(n8140), .ZN(n11023) );
  NAND2_X4 U7288 ( .A1(n8238), .A2(n8237), .ZN(n14803) );
  NAND2_X2 U7289 ( .A1(n8147), .A2(n8653), .ZN(n10023) );
  OAI21_X2 U7290 ( .B1(n7651), .B2(n6516), .A(n7192), .ZN(n7689) );
  XNOR2_X2 U7291 ( .A(n13128), .B(n10689), .ZN(n10266) );
  AND2_X1 U7292 ( .A1(n13127), .A2(n9956), .ZN(n10365) );
  AOI21_X2 U7293 ( .B1(n8495), .B2(n6545), .A(n7129), .ZN(n13254) );
  NAND2_X2 U7294 ( .A1(n13321), .A2(n8474), .ZN(n13317) );
  AOI21_X2 U7295 ( .B1(n11942), .B2(n7027), .A(n7026), .ZN(n7025) );
  NAND2_X2 U7296 ( .A1(n8297), .A2(n8296), .ZN(n11133) );
  NAND4_X1 U7297 ( .A1(n9099), .A2(n9098), .A3(n9097), .A4(n9096), .ZN(n12555)
         );
  XNOR2_X2 U7298 ( .A(n8025), .B(n8024), .ZN(n8031) );
  OAI21_X2 U7299 ( .B1(n8023), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8025) );
  AND2_X1 U7300 ( .A1(n11264), .A2(n11261), .ZN(n7347) );
  XNOR2_X2 U7301 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9111) );
  NOR2_X2 U7302 ( .A1(n14522), .A2(n14521), .ZN(n14520) );
  OAI21_X2 U7303 ( .B1(n14246), .B2(n14245), .A(n14285), .ZN(n14521) );
  AND2_X1 U7304 ( .A1(n6680), .A2(n11904), .ZN(n7221) );
  NAND2_X2 U7305 ( .A1(n7951), .A2(n7950), .ZN(n14079) );
  NAND2_X2 U7307 ( .A1(n7115), .A2(n7116), .ZN(n11244) );
  NAND2_X4 U7308 ( .A1(n8310), .A2(n8309), .ZN(n11263) );
  NAND2_X2 U7309 ( .A1(n8555), .A2(n8554), .ZN(n10249) );
  NAND2_X2 U7310 ( .A1(n7607), .A2(n7606), .ZN(n11734) );
  BUF_X2 U7311 ( .A(n8206), .Z(n6474) );
  AOI21_X2 U7312 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9972), .A(n10011), .ZN(
        n9984) );
  OAI21_X1 U7313 ( .B1(n13043), .B2(n7317), .A(n7315), .ZN(n11986) );
  INV_X1 U7314 ( .A(n12586), .ZN(n6475) );
  XNOR2_X2 U7315 ( .A(n7016), .B(n9021), .ZN(n9533) );
  AOI211_X1 U7316 ( .C1(n14069), .C2(n13999), .A(n13876), .B(n13875), .ZN(
        n13877) );
  INV_X2 U7317 ( .A(n12511), .ZN(n12378) );
  OR2_X1 U7318 ( .A1(n12647), .A2(n12655), .ZN(n12393) );
  OR2_X1 U7319 ( .A1(n9001), .A2(n13560), .ZN(n9003) );
  NAND2_X1 U7320 ( .A1(n9613), .A2(n9612), .ZN(n11364) );
  NAND2_X1 U7321 ( .A1(n11774), .A2(n11775), .ZN(n7738) );
  OAI21_X1 U7322 ( .B1(n10894), .B2(n10893), .A(n10892), .ZN(n10898) );
  NAND2_X1 U7323 ( .A1(n6854), .A2(n6855), .ZN(n7631) );
  INV_X2 U7324 ( .A(n10737), .ZN(n9675) );
  INV_X1 U7325 ( .A(n12356), .ZN(n6476) );
  NAND2_X1 U7326 ( .A1(n12416), .A2(n12422), .ZN(n12414) );
  INV_X1 U7327 ( .A(n10821), .ZN(n10833) );
  INV_X1 U7328 ( .A(n11232), .ZN(n12548) );
  INV_X1 U7329 ( .A(n9547), .ZN(n12524) );
  INV_X1 U7330 ( .A(n13722), .ZN(n14046) );
  NAND2_X2 U7331 ( .A1(n14013), .A2(n12147), .ZN(n10334) );
  INV_X1 U7332 ( .A(n12551), .ZN(n11093) );
  AND4_X1 U7333 ( .A1(n9190), .A2(n9189), .A3(n9188), .A4(n9187), .ZN(n11232)
         );
  INV_X1 U7334 ( .A(n12147), .ZN(n12161) );
  CLKBUF_X1 U7335 ( .A(n12623), .Z(n6490) );
  CLKBUF_X3 U7336 ( .A(n10024), .Z(n13129) );
  BUF_X2 U7337 ( .A(n9483), .Z(n9529) );
  INV_X1 U7339 ( .A(n11694), .ZN(n7408) );
  NAND2_X1 U7340 ( .A1(n6489), .A2(n7495), .ZN(n9381) );
  CLKBUF_X2 U7341 ( .A(n8545), .Z(n6666) );
  NAND2_X1 U7342 ( .A1(n13843), .A2(n14168), .ZN(n11689) );
  CLKBUF_X2 U7343 ( .A(n8456), .Z(n8615) );
  AND2_X1 U7344 ( .A1(n9746), .A2(n9735), .ZN(n7531) );
  BUF_X1 U7345 ( .A(n8552), .Z(n8935) );
  NAND2_X1 U7346 ( .A1(n6684), .A2(n6683), .ZN(n8035) );
  NAND2_X1 U7347 ( .A1(n7817), .A2(n7816), .ZN(n7834) );
  INV_X4 U7348 ( .A(n7495), .ZN(n7777) );
  NOR2_X1 U7349 ( .A1(n8201), .A2(n8207), .ZN(n9880) );
  INV_X1 U7350 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7816) );
  AOI22_X1 U7351 ( .A1(n11848), .A2(n11847), .B1(n11846), .B2(n11845), .ZN(
        n11863) );
  AOI21_X1 U7352 ( .B1(n7012), .B2(n15038), .A(n6621), .ZN(n7011) );
  AOI211_X1 U7353 ( .C1(n14490), .C2(n14084), .A(n13613), .B(n13612), .ZN(
        n13614) );
  AND2_X1 U7354 ( .A1(n9537), .A2(n9536), .ZN(n12652) );
  AOI21_X1 U7355 ( .B1(n6987), .B2(n6989), .A(n6565), .ZN(n6985) );
  AND2_X1 U7356 ( .A1(n7079), .A2(n7077), .ZN(n9575) );
  AND2_X1 U7357 ( .A1(n14067), .A2(n14066), .ZN(n6662) );
  NAND2_X1 U7358 ( .A1(n9661), .A2(n9660), .ZN(n7385) );
  AND2_X1 U7359 ( .A1(n12516), .A2(n12519), .ZN(n12379) );
  OR2_X1 U7360 ( .A1(n9578), .A2(n9565), .ZN(n12516) );
  NAND2_X1 U7361 ( .A1(n11993), .A2(n11992), .ZN(n13035) );
  AOI21_X1 U7362 ( .B1(n12339), .B2(n12338), .A(n6617), .ZN(n12907) );
  NAND2_X1 U7363 ( .A1(n9573), .A2(n9481), .ZN(n12658) );
  NAND2_X1 U7364 ( .A1(n12682), .A2(n12681), .ZN(n12680) );
  NAND2_X1 U7365 ( .A1(n9474), .A2(n9473), .ZN(n9676) );
  NAND2_X1 U7366 ( .A1(n9463), .A2(n9462), .ZN(n12506) );
  NAND2_X1 U7367 ( .A1(n6729), .A2(n6734), .ZN(n13885) );
  NOR3_X1 U7368 ( .A1(n14063), .A2(n6892), .A3(n14064), .ZN(n14066) );
  NOR3_X1 U7369 ( .A1(n6893), .A2(n13855), .A3(n14509), .ZN(n14063) );
  NAND2_X1 U7370 ( .A1(n7279), .A2(n7280), .ZN(n9562) );
  OR2_X1 U7371 ( .A1(n14297), .A2(n14296), .ZN(n6909) );
  AND2_X1 U7372 ( .A1(n6913), .A2(n6914), .ZN(n14297) );
  OR2_X1 U7373 ( .A1(n14341), .A2(n12566), .ZN(n7105) );
  OR2_X1 U7374 ( .A1(n6495), .A2(n12396), .ZN(n12716) );
  XNOR2_X1 U7375 ( .A(n6517), .B(n6698), .ZN(n13194) );
  NAND2_X1 U7376 ( .A1(n9426), .A2(n9425), .ZN(n12395) );
  INV_X1 U7377 ( .A(n12250), .ZN(n7390) );
  AND2_X1 U7378 ( .A1(n6917), .A2(n6916), .ZN(n14538) );
  XNOR2_X1 U7379 ( .A(n7995), .B(n7994), .ZN(n11684) );
  NAND2_X1 U7380 ( .A1(n9404), .A2(n9403), .ZN(n12731) );
  NAND2_X1 U7381 ( .A1(n8999), .A2(n8998), .ZN(n9414) );
  OAI21_X1 U7382 ( .B1(n6950), .B2(n6946), .A(n6945), .ZN(n7995) );
  OR2_X1 U7383 ( .A1(n14534), .A2(n14533), .ZN(n6916) );
  NAND2_X1 U7384 ( .A1(n11611), .A2(n7147), .ZN(n13490) );
  OR2_X1 U7385 ( .A1(n7948), .A2(n6956), .ZN(n6949) );
  NAND2_X1 U7386 ( .A1(n13647), .A2(n13646), .ZN(n13645) );
  AND2_X1 U7387 ( .A1(n6920), .A2(n6919), .ZN(n14534) );
  NAND2_X1 U7388 ( .A1(n7929), .A2(n7928), .ZN(n7948) );
  NAND2_X1 U7389 ( .A1(n11612), .A2(n8384), .ZN(n11611) );
  NAND2_X1 U7390 ( .A1(n7838), .A2(n7837), .ZN(n14119) );
  AND2_X1 U7391 ( .A1(n14729), .A2(n14730), .ZN(n14726) );
  NOR2_X1 U7392 ( .A1(n6651), .A2(n14525), .ZN(n14528) );
  NAND2_X1 U7393 ( .A1(n8994), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U7394 ( .A1(n11467), .A2(n11466), .ZN(n11471) );
  NAND2_X1 U7395 ( .A1(n7181), .A2(n7179), .ZN(n11467) );
  OAI21_X1 U7396 ( .B1(n7911), .B2(n10934), .A(n7914), .ZN(n7927) );
  NAND2_X1 U7397 ( .A1(n7820), .A2(n7819), .ZN(n14125) );
  XNOR2_X1 U7398 ( .A(n7896), .B(SI_22_), .ZN(n8465) );
  XNOR2_X1 U7399 ( .A(n7745), .B(n7744), .ZN(n10469) );
  NAND2_X2 U7400 ( .A1(n8360), .A2(n8359), .ZN(n14412) );
  OAI21_X1 U7401 ( .B1(n7810), .B2(n6970), .A(n6968), .ZN(n7896) );
  NAND2_X1 U7402 ( .A1(n7797), .A2(n7796), .ZN(n7810) );
  XNOR2_X1 U7403 ( .A(n7741), .B(n7771), .ZN(n10387) );
  INV_X1 U7404 ( .A(n11903), .ZN(n6477) );
  OAI21_X1 U7405 ( .B1(n7707), .B2(n7196), .A(n7194), .ZN(n7770) );
  XNOR2_X1 U7406 ( .A(n7705), .B(n7446), .ZN(n10020) );
  NAND2_X1 U7407 ( .A1(n6869), .A2(n7188), .ZN(n7705) );
  NAND2_X1 U7408 ( .A1(n10236), .A2(n10237), .ZN(n10339) );
  XNOR2_X1 U7409 ( .A(n7668), .B(n7652), .ZN(n9910) );
  NAND2_X1 U7410 ( .A1(n7638), .A2(n7637), .ZN(n11748) );
  NAND2_X1 U7411 ( .A1(n7651), .A2(n7650), .ZN(n7668) );
  NAND2_X2 U7412 ( .A1(n8269), .A2(n8268), .ZN(n14820) );
  INV_X2 U7413 ( .A(n15045), .ZN(n12844) );
  NAND2_X1 U7414 ( .A1(n7618), .A2(n7617), .ZN(n11739) );
  NAND2_X1 U7415 ( .A1(n7648), .A2(n7647), .ZN(n7651) );
  XNOR2_X1 U7416 ( .A(n7631), .B(n7629), .ZN(n9775) );
  AOI21_X1 U7417 ( .B1(n10622), .B2(n10621), .A(n6845), .ZN(n10757) );
  AND3_X1 U7418 ( .A1(n9200), .A2(n9199), .A3(n9198), .ZN(n14848) );
  AND2_X1 U7419 ( .A1(n12425), .A2(n12428), .ZN(n12356) );
  NAND2_X2 U7420 ( .A1(n10278), .A2(n13300), .ZN(n13336) );
  NOR2_X1 U7421 ( .A1(n14901), .A2(n14900), .ZN(n14899) );
  AND2_X1 U7423 ( .A1(n12407), .A2(n12410), .ZN(n12357) );
  AND2_X1 U7424 ( .A1(n7557), .A2(n7556), .ZN(n11713) );
  NAND2_X1 U7425 ( .A1(n8212), .A2(n8211), .ZN(n10413) );
  NAND2_X1 U7426 ( .A1(n6943), .A2(n7570), .ZN(n7584) );
  MUX2_X1 U7427 ( .A(n10265), .B(n13128), .S(n8867), .Z(n8682) );
  OAI211_X1 U7428 ( .C1(n9763), .C2(n9381), .A(n6524), .B(n9179), .ZN(n10947)
         );
  INV_X2 U7429 ( .A(n10305), .ZN(n8204) );
  INV_X1 U7430 ( .A(n10579), .ZN(n6478) );
  CLKBUF_X1 U7431 ( .A(n12129), .Z(n6648) );
  NOR2_X1 U7432 ( .A1(n10264), .A2(n10265), .ZN(n10303) );
  NAND2_X1 U7433 ( .A1(n9175), .A2(n8962), .ZN(n8964) );
  AND3_X1 U7434 ( .A1(n9105), .A2(n9104), .A3(n9103), .ZN(n11678) );
  INV_X1 U7435 ( .A(n10689), .ZN(n10265) );
  NAND2_X1 U7436 ( .A1(n8961), .A2(n8960), .ZN(n9175) );
  CLKBUF_X1 U7437 ( .A(n12829), .Z(n12797) );
  OAI21_X1 U7438 ( .B1(n9060), .B2(P3_D_REG_0__SCAN_IN), .A(n9061), .ZN(n9585)
         );
  INV_X1 U7439 ( .A(n10024), .ZN(n8674) );
  NAND4_X2 U7440 ( .A1(n7502), .A2(n7501), .A3(n7500), .A4(n7499), .ZN(n13721)
         );
  NAND2_X1 U7441 ( .A1(n8216), .A2(n6537), .ZN(n13126) );
  NAND4_X1 U7442 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n12551)
         );
  NAND4_X1 U7443 ( .A1(n9118), .A2(n9117), .A3(n9116), .A4(n9115), .ZN(n12553)
         );
  NAND2_X1 U7444 ( .A1(n7551), .A2(n7550), .ZN(n7568) );
  OAI211_X1 U7445 ( .C1(n11854), .C2(n6739), .A(n7596), .B(n6568), .ZN(n13718)
         );
  INV_X1 U7446 ( .A(n9381), .ZN(n9160) );
  NAND4_X1 U7447 ( .A1(n8164), .A2(n8162), .A3(n8163), .A4(n8161), .ZN(n8668)
         );
  CLKBUF_X1 U7448 ( .A(n8030), .Z(n14167) );
  INV_X2 U7449 ( .A(n6471), .ZN(n6483) );
  OAI21_X1 U7450 ( .B1(n9362), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9032) );
  INV_X1 U7451 ( .A(n10282), .ZN(n11075) );
  BUF_X4 U7452 ( .A(n8206), .Z(n6479) );
  OR2_X1 U7453 ( .A1(n8489), .A2(n6649), .ZN(n8162) );
  INV_X1 U7454 ( .A(n10515), .ZN(n9582) );
  INV_X1 U7455 ( .A(n8489), .ZN(n8614) );
  AND2_X2 U7456 ( .A1(n9094), .A2(n9095), .ZN(n9169) );
  INV_X1 U7457 ( .A(n8004), .ZN(n7561) );
  INV_X1 U7458 ( .A(n12965), .ZN(n9095) );
  INV_X1 U7459 ( .A(n7467), .ZN(n14154) );
  NAND2_X1 U7460 ( .A1(n9039), .A2(n9041), .ZN(n10515) );
  CLKBUF_X2 U7461 ( .A(n8551), .Z(n10282) );
  INV_X1 U7462 ( .A(n8159), .ZN(n8157) );
  NAND2_X1 U7463 ( .A1(n7092), .A2(n7091), .ZN(n12965) );
  NAND2_X1 U7464 ( .A1(n9050), .A2(n9051), .ZN(n11291) );
  NAND2_X1 U7465 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  OAI21_X2 U7466 ( .B1(n8018), .B2(n7432), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7057) );
  NAND2_X1 U7467 ( .A1(n8648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8142) );
  MUX2_X1 U7468 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9047), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9050) );
  INV_X2 U7469 ( .A(n13543), .ZN(n13550) );
  NAND2_X1 U7470 ( .A1(n6838), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U7471 ( .A1(n9092), .A2(n6560), .ZN(n7091) );
  OR2_X1 U7472 ( .A1(n9093), .A2(n12958), .ZN(n9091) );
  INV_X1 U7473 ( .A(n7834), .ZN(n6684) );
  NOR2_X1 U7474 ( .A1(n9053), .A2(n7395), .ZN(n9022) );
  NAND2_X2 U7475 ( .A1(n9735), .A2(P1_U3086), .ZN(n14163) );
  NAND2_X1 U7476 ( .A1(n6679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8167) );
  XNOR2_X1 U7477 ( .A(n7549), .B(SI_3_), .ZN(n7546) );
  NAND2_X1 U7478 ( .A1(n6850), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7016) );
  NAND2_X2 U7479 ( .A1(n7495), .A2(P1_U3086), .ZN(n14166) );
  NOR2_X1 U7480 ( .A1(n9034), .A2(n9033), .ZN(n9038) );
  AND2_X2 U7481 ( .A1(n7604), .A2(n7459), .ZN(n7813) );
  INV_X1 U7482 ( .A(n8266), .ZN(n8123) );
  AND3_X1 U7483 ( .A1(n6583), .A2(n6994), .A3(n9014), .ZN(n7097) );
  NAND2_X1 U7484 ( .A1(n8177), .A2(n8176), .ZN(n14660) );
  INV_X4 U7485 ( .A(n7887), .ZN(n7495) );
  NAND2_X1 U7486 ( .A1(n7433), .A2(n7473), .ZN(n7432) );
  NOR2_X1 U7487 ( .A1(n9033), .A2(n6995), .ZN(n6994) );
  AND2_X1 U7488 ( .A1(n6583), .A2(n9014), .ZN(n6795) );
  NAND2_X1 U7489 ( .A1(n7018), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9023) );
  AND2_X1 U7490 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  AND2_X1 U7491 ( .A1(n7483), .A2(n7455), .ZN(n7505) );
  AND4_X1 U7492 ( .A1(n9013), .A2(n9012), .A3(n9215), .A4(n9196), .ZN(n9014)
         );
  AND3_X1 U7493 ( .A1(n6745), .A2(n6744), .A3(n9011), .ZN(n9144) );
  NAND4_X1 U7494 ( .A1(n9016), .A2(n9017), .A3(n9029), .A4(n9363), .ZN(n9033)
         );
  AND2_X1 U7495 ( .A1(n7406), .A2(n7404), .ZN(n7021) );
  INV_X1 U7496 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9080) );
  INV_X1 U7497 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8220) );
  NOR2_X1 U7498 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7404) );
  NOR2_X1 U7499 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7406) );
  NOR2_X1 U7500 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7405) );
  INV_X4 U7501 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7502 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8036) );
  NOR2_X1 U7503 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n9012) );
  NOR2_X1 U7504 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n9013) );
  INV_X1 U7505 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9029) );
  INV_X1 U7506 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9363) );
  INV_X4 U7507 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7508 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8649) );
  NOR2_X1 U7509 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n9016) );
  NOR2_X1 U7510 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9017) );
  INV_X1 U7511 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8155) );
  INV_X1 U7512 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9037) );
  INV_X1 U7513 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9721) );
  INV_X1 U7514 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9011) );
  NOR2_X1 U7515 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6744) );
  INV_X1 U7516 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9021) );
  INV_X4 U7517 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7518 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7481) );
  INV_X1 U7519 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7479) );
  NOR2_X1 U7520 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8119) );
  NOR2_X1 U7521 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n9020) );
  INV_X1 U7522 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9018) );
  NAND4_X4 U7523 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(n9495)
         );
  XNOR2_X2 U7524 ( .A(n8978), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U7525 ( .A1(n8670), .A2(n8669), .ZN(n8681) );
  AND2_X1 U7526 ( .A1(n8135), .A2(n8137), .ZN(n8139) );
  NOR2_X2 U7527 ( .A1(n11513), .A2(n14472), .ZN(n6891) );
  XNOR2_X2 U7528 ( .A(n8034), .B(P1_IR_REG_21__SCAN_IN), .ZN(n14043) );
  AND2_X4 U7529 ( .A1(n8175), .A2(n8117), .ZN(n8188) );
  NOR2_X1 U7531 ( .A1(n9595), .A2(n9598), .ZN(n10741) );
  AOI21_X2 U7532 ( .B1(n13052), .B2(n13053), .A(n11987), .ZN(n11989) );
  INV_X1 U7533 ( .A(n6471), .ZN(n6481) );
  AOI21_X2 U7534 ( .B1(n13035), .B2(n13034), .A(n6664), .ZN(n13004) );
  OR2_X2 U7535 ( .A1(n8401), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n6513) );
  AOI21_X2 U7536 ( .B1(n7390), .B2(n7389), .A(n7386), .ZN(n12214) );
  NOR2_X1 U7537 ( .A1(n9586), .A2(n12524), .ZN(n6484) );
  OAI21_X2 U7538 ( .B1(n12727), .B2(n12355), .A(n12353), .ZN(n12717) );
  AOI21_X2 U7539 ( .B1(n12539), .B2(n12486), .A(n12743), .ZN(n12727) );
  OAI21_X2 U7540 ( .B1(n12214), .B2(n12213), .A(n9648), .ZN(n12273) );
  NAND2_X2 U7541 ( .A1(n11956), .A2(n9533), .ZN(n9102) );
  OAI21_X2 U7542 ( .B1(n12230), .B2(n9625), .A(n9624), .ZN(n12021) );
  BUF_X8 U7543 ( .A(n9169), .Z(n6486) );
  INV_X1 U7544 ( .A(n9746), .ZN(n6487) );
  NAND2_X1 U7545 ( .A1(n11956), .A2(n9533), .ZN(n6488) );
  NAND2_X1 U7546 ( .A1(n11956), .A2(n9533), .ZN(n6489) );
  CLKBUF_X3 U7547 ( .A(n7540), .Z(n8003) );
  AOI21_X2 U7548 ( .B1(n12706), .B2(n12705), .A(n7005), .ZN(n12693) );
  NOR2_X4 U7549 ( .A1(n10963), .A2(n11748), .ZN(n11082) );
  OR2_X2 U7550 ( .A1(n11037), .A2(n11739), .ZN(n10963) );
  NOR2_X1 U7551 ( .A1(n11813), .A2(n11814), .ZN(n6878) );
  INV_X1 U7552 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8200) );
  NOR2_X2 U7553 ( .A1(n7078), .A2(n12658), .ZN(n7077) );
  INV_X1 U7554 ( .A(n7080), .ZN(n7078) );
  OR3_X1 U7555 ( .A1(n13259), .A2(n8605), .A3(n6831), .ZN(n6828) );
  INV_X1 U7556 ( .A(n6834), .ZN(n6831) );
  OAI21_X1 U7557 ( .B1(n7130), .B2(n8506), .A(n6566), .ZN(n7129) );
  NAND2_X1 U7558 ( .A1(n8833), .A2(n8832), .ZN(n8863) );
  NAND2_X1 U7559 ( .A1(n8830), .A2(n8829), .ZN(n8833) );
  INV_X1 U7560 ( .A(n7300), .ZN(n6820) );
  AOI21_X1 U7561 ( .B1(n7300), .B2(n6819), .A(n6818), .ZN(n6817) );
  AOI21_X1 U7562 ( .B1(n7302), .B2(n7305), .A(n7301), .ZN(n7300) );
  XNOR2_X1 U7564 ( .A(n6642), .B(n12158), .ZN(n10574) );
  NOR2_X1 U7565 ( .A1(n13898), .A2(n7238), .ZN(n7237) );
  INV_X1 U7566 ( .A(n7923), .ZN(n7238) );
  OAI21_X1 U7567 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14198), .A(n14197), .ZN(
        n14251) );
  OR2_X1 U7568 ( .A1(n14528), .A2(n14529), .ZN(n6919) );
  INV_X1 U7569 ( .A(n8765), .ZN(n6658) );
  NOR2_X1 U7570 ( .A1(n6767), .A2(n12447), .ZN(n6766) );
  NOR2_X1 U7571 ( .A1(n6769), .A2(n6768), .ZN(n6767) );
  INV_X1 U7572 ( .A(n12448), .ZN(n6768) );
  AND2_X1 U7573 ( .A1(n7000), .A2(n12444), .ZN(n6769) );
  INV_X1 U7574 ( .A(n11812), .ZN(n7427) );
  NAND2_X1 U7575 ( .A1(n6575), .A2(n6876), .ZN(n6872) );
  NOR2_X1 U7576 ( .A1(n13253), .A2(n6833), .ZN(n6832) );
  INV_X1 U7577 ( .A(n8606), .ZN(n6833) );
  NOR2_X1 U7578 ( .A1(n7037), .A2(n8068), .ZN(n7036) );
  INV_X1 U7579 ( .A(n8067), .ZN(n7037) );
  INV_X1 U7580 ( .A(n7812), .ZN(n6975) );
  NAND2_X1 U7581 ( .A1(n7438), .A2(n7847), .ZN(n7850) );
  NAND2_X1 U7582 ( .A1(n6922), .A2(n14176), .ZN(n14177) );
  NAND2_X1 U7583 ( .A1(n14223), .A2(n14224), .ZN(n6922) );
  NAND2_X1 U7584 ( .A1(n10709), .A2(n9582), .ZN(n9584) );
  NOR2_X1 U7585 ( .A1(n6779), .A2(n6781), .ZN(n6778) );
  NAND2_X1 U7586 ( .A1(n6771), .A2(n6770), .ZN(n6779) );
  NAND2_X1 U7587 ( .A1(n12515), .A2(n12519), .ZN(n6771) );
  NAND2_X1 U7588 ( .A1(n6500), .A2(n12378), .ZN(n6777) );
  OR2_X1 U7589 ( .A1(n12885), .A2(n9640), .ZN(n12474) );
  OR2_X1 U7590 ( .A1(n12948), .A2(n12796), .ZN(n12478) );
  NAND2_X1 U7591 ( .A1(n10872), .A2(n10947), .ZN(n12425) );
  AND2_X1 U7592 ( .A1(n9177), .A2(n6853), .ZN(n6851) );
  INV_X1 U7593 ( .A(n7250), .ZN(n7249) );
  OAI21_X1 U7594 ( .B1(n9240), .B2(n7251), .A(n8974), .ZN(n7250) );
  AND2_X1 U7595 ( .A1(n7246), .A2(n8963), .ZN(n7245) );
  INV_X1 U7596 ( .A(n9191), .ZN(n7246) );
  INV_X1 U7597 ( .A(n13541), .ZN(n8160) );
  OR2_X1 U7598 ( .A1(n8844), .A2(n9861), .ZN(n8170) );
  AND2_X1 U7599 ( .A1(n8121), .A2(n8122), .ZN(n7349) );
  INV_X1 U7600 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U7601 ( .A1(n6942), .A2(n13252), .ZN(n6941) );
  NOR2_X1 U7602 ( .A1(n8850), .A2(n12018), .ZN(n6942) );
  OR2_X1 U7603 ( .A1(n13441), .A2(n6929), .ZN(n6928) );
  INV_X1 U7604 ( .A(n7313), .ZN(n6827) );
  NOR2_X1 U7605 ( .A1(n13096), .A2(n13488), .ZN(n6937) );
  NOR2_X1 U7606 ( .A1(n8357), .A2(n7138), .ZN(n7137) );
  INV_X1 U7607 ( .A(n8340), .ZN(n7138) );
  AND2_X1 U7608 ( .A1(n8912), .A2(n8356), .ZN(n7135) );
  INV_X1 U7609 ( .A(n8607), .ZN(n6835) );
  NOR3_X1 U7610 ( .A1(n13328), .A2(n13010), .A3(n6928), .ZN(n13280) );
  INV_X1 U7611 ( .A(n7468), .ZN(n7466) );
  NOR2_X1 U7612 ( .A1(n7035), .A2(n10648), .ZN(n6718) );
  NAND2_X1 U7613 ( .A1(n7537), .A2(n11686), .ZN(n11892) );
  NAND2_X1 U7614 ( .A1(n6478), .A2(n6646), .ZN(n7537) );
  NAND2_X1 U7615 ( .A1(n7039), .A2(n7040), .ZN(n11518) );
  AOI21_X1 U7616 ( .B1(n7043), .B2(n7045), .A(n7041), .ZN(n7040) );
  AND2_X1 U7617 ( .A1(n11451), .A2(n7044), .ZN(n7043) );
  NAND2_X1 U7618 ( .A1(n7407), .A2(n7412), .ZN(n11890) );
  AND2_X1 U7619 ( .A1(n7494), .A2(n7408), .ZN(n7407) );
  NAND2_X1 U7620 ( .A1(n7999), .A2(n7998), .ZN(n8830) );
  OR2_X1 U7621 ( .A1(n7995), .A2(n7994), .ZN(n7999) );
  INV_X1 U7622 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8032) );
  INV_X1 U7623 ( .A(n6966), .ZN(n6965) );
  AOI21_X1 U7624 ( .B1(n6966), .B2(n6964), .A(n6963), .ZN(n6962) );
  AOI21_X1 U7625 ( .B1(n7194), .B2(n7196), .A(n7769), .ZN(n6966) );
  AOI21_X1 U7626 ( .B1(n7192), .B2(n7190), .A(n7189), .ZN(n7188) );
  NAND2_X1 U7627 ( .A1(n7651), .A2(n6552), .ZN(n6869) );
  INV_X1 U7628 ( .A(n7687), .ZN(n7189) );
  NAND2_X1 U7629 ( .A1(n7379), .A2(n7377), .ZN(n12312) );
  AND2_X1 U7630 ( .A1(n7378), .A2(n12313), .ZN(n7377) );
  NAND2_X1 U7631 ( .A1(n7380), .A2(n12241), .ZN(n7378) );
  AOI21_X1 U7632 ( .B1(n12381), .B2(n12900), .A(n12385), .ZN(n7095) );
  INV_X1 U7633 ( .A(n12391), .ZN(n7272) );
  NAND2_X1 U7634 ( .A1(n12392), .A2(n9044), .ZN(n7273) );
  INV_X1 U7635 ( .A(n6482), .ZN(n9488) );
  NOR2_X1 U7636 ( .A1(n14899), .A2(n6846), .ZN(n14923) );
  AND2_X1 U7637 ( .A1(n10441), .A2(n10459), .ZN(n6846) );
  NAND2_X1 U7638 ( .A1(n6887), .A2(n6886), .ZN(n6885) );
  INV_X1 U7639 ( .A(n10753), .ZN(n6886) );
  AOI21_X1 U7640 ( .B1(n14323), .B2(n12565), .A(n14331), .ZN(n12566) );
  OR2_X1 U7641 ( .A1(n12505), .A2(n12915), .ZN(n7445) );
  NAND2_X1 U7642 ( .A1(n6564), .A2(n7081), .ZN(n7080) );
  AOI22_X2 U7643 ( .A1(n12677), .A2(n12676), .B1(n12536), .B2(n12501), .ZN(
        n12667) );
  INV_X1 U7644 ( .A(n12827), .ZN(n15042) );
  AOI21_X1 U7645 ( .B1(n7281), .B2(n9007), .A(n6624), .ZN(n7280) );
  AND2_X1 U7646 ( .A1(n8968), .A2(n8967), .ZN(n9210) );
  AND4_X1 U7647 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n13079)
         );
  NAND2_X1 U7648 ( .A1(n8157), .A2(n13541), .ZN(n8844) );
  XNOR2_X1 U7649 ( .A(n13218), .B(n12013), .ZN(n8923) );
  AND2_X1 U7650 ( .A1(n13507), .A2(n13280), .ZN(n13266) );
  OR2_X1 U7651 ( .A1(n13259), .A2(n8605), .ZN(n6837) );
  AOI21_X1 U7652 ( .B1(n7304), .B2(n7303), .A(n6576), .ZN(n7302) );
  INV_X1 U7653 ( .A(n11245), .ZN(n7303) );
  AND2_X1 U7654 ( .A1(n8661), .A2(n8670), .ZN(n9953) );
  OR2_X1 U7655 ( .A1(n10282), .A2(n8935), .ZN(n10033) );
  OAI21_X2 U7657 ( .B1(n6513), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8146) );
  INV_X1 U7658 ( .A(n10338), .ZN(n7185) );
  OR2_X1 U7659 ( .A1(n11633), .A2(n7436), .ZN(n7166) );
  INV_X1 U7660 ( .A(n7436), .ZN(n7169) );
  INV_X1 U7661 ( .A(n13627), .ZN(n7159) );
  AOI21_X1 U7662 ( .B1(n13627), .B2(n7158), .A(n7157), .ZN(n7156) );
  INV_X1 U7663 ( .A(n13609), .ZN(n7157) );
  NAND2_X1 U7664 ( .A1(n7411), .A2(n7410), .ZN(n7409) );
  NAND2_X1 U7665 ( .A1(n9932), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U7666 ( .A1(n7408), .A2(n12147), .ZN(n7411) );
  NAND2_X1 U7667 ( .A1(n13611), .A2(n12138), .ZN(n13677) );
  NAND2_X1 U7668 ( .A1(n13677), .A2(n13678), .ZN(n13676) );
  NAND2_X1 U7669 ( .A1(n7467), .A2(n7466), .ZN(n7540) );
  OAI21_X1 U7670 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n13861) );
  INV_X1 U7671 ( .A(n13885), .ZN(n7024) );
  AOI21_X1 U7672 ( .B1(n7025), .B2(n11918), .A(n13873), .ZN(n7022) );
  INV_X1 U7673 ( .A(n7025), .ZN(n7023) );
  INV_X1 U7674 ( .A(n11918), .ZN(n11942) );
  INV_X1 U7675 ( .A(n13703), .ZN(n13603) );
  OR2_X1 U7676 ( .A1(n13928), .A2(n13704), .ZN(n7923) );
  NOR2_X1 U7677 ( .A1(n13914), .A2(n7240), .ZN(n7239) );
  INV_X1 U7678 ( .A(n7910), .ZN(n7240) );
  INV_X1 U7679 ( .A(n11871), .ZN(n7151) );
  OR2_X1 U7680 ( .A1(n12047), .A2(n14462), .ZN(n11784) );
  NAND2_X1 U7681 ( .A1(n11509), .A2(n7767), .ZN(n11590) );
  INV_X1 U7682 ( .A(n9746), .ZN(n7836) );
  NAND2_X1 U7683 ( .A1(n10639), .A2(n7598), .ZN(n11034) );
  NAND2_X1 U7684 ( .A1(n11861), .A2(n8042), .ZN(n14028) );
  NAND2_X1 U7685 ( .A1(n10554), .A2(n7497), .ZN(n10133) );
  INV_X1 U7686 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7459) );
  AOI22_X1 U7687 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14201), .B1(n14251), 
        .B2(n14200), .ZN(n14254) );
  INV_X1 U7688 ( .A(n13194), .ZN(n13196) );
  NAND2_X1 U7689 ( .A1(n7983), .A2(n7982), .ZN(n14070) );
  NAND2_X1 U7690 ( .A1(n6921), .A2(n14530), .ZN(n6920) );
  NAND2_X1 U7691 ( .A1(n14528), .A2(n14529), .ZN(n6921) );
  OAI21_X1 U7692 ( .B1(n10247), .B2(n8666), .A(n8681), .ZN(n8671) );
  NAND2_X1 U7693 ( .A1(n8699), .A2(n6695), .ZN(n6694) );
  INV_X1 U7694 ( .A(n8698), .ZN(n6695) );
  MUX2_X1 U7695 ( .A(n13124), .B(n14803), .S(n8884), .Z(n8708) );
  OAI21_X1 U7696 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n11709) );
  INV_X1 U7697 ( .A(n8730), .ZN(n6665) );
  NAND2_X1 U7698 ( .A1(n11758), .A2(n7419), .ZN(n7418) );
  NAND2_X1 U7699 ( .A1(n8764), .A2(n8763), .ZN(n8766) );
  NOR2_X1 U7700 ( .A1(n11783), .A2(n11782), .ZN(n7401) );
  AOI21_X1 U7701 ( .B1(n7738), .B2(n11860), .A(n6567), .ZN(n11783) );
  OAI21_X1 U7702 ( .B1(n12409), .B2(n6743), .A(n6741), .ZN(n6740) );
  INV_X1 U7703 ( .A(n6742), .ZN(n6741) );
  NAND2_X1 U7704 ( .A1(n10657), .A2(n7004), .ZN(n6743) );
  OAI21_X1 U7705 ( .B1(n15039), .B2(n12405), .A(n12410), .ZN(n6742) );
  INV_X1 U7706 ( .A(n11811), .ZN(n7428) );
  NOR2_X1 U7707 ( .A1(n6882), .A2(n6881), .ZN(n6880) );
  INV_X1 U7708 ( .A(n11814), .ZN(n6881) );
  INV_X1 U7709 ( .A(n11813), .ZN(n6882) );
  AOI21_X1 U7710 ( .B1(n6766), .B2(n6511), .A(n12451), .ZN(n6764) );
  INV_X1 U7711 ( .A(n6766), .ZN(n6765) );
  NAND2_X1 U7712 ( .A1(n7428), .A2(n7427), .ZN(n7426) );
  NAND2_X1 U7713 ( .A1(n6874), .A2(n6880), .ZN(n6871) );
  AND2_X1 U7714 ( .A1(n6879), .A2(n6875), .ZN(n6874) );
  INV_X1 U7715 ( .A(n6878), .ZN(n6875) );
  AOI21_X1 U7716 ( .B1(n11815), .B2(n6878), .A(n6877), .ZN(n6876) );
  INV_X1 U7717 ( .A(n11816), .ZN(n6877) );
  AND2_X1 U7718 ( .A1(n6756), .A2(n6760), .ZN(n6755) );
  NAND2_X1 U7719 ( .A1(n6757), .A2(n6759), .ZN(n6756) );
  NAND2_X1 U7720 ( .A1(n8789), .A2(n8787), .ZN(n7356) );
  AOI21_X1 U7721 ( .B1(n6755), .B2(n6753), .A(n12468), .ZN(n6752) );
  INV_X1 U7722 ( .A(n6757), .ZN(n6753) );
  INV_X1 U7723 ( .A(n6755), .ZN(n6754) );
  INV_X1 U7724 ( .A(n12471), .ZN(n6750) );
  INV_X1 U7725 ( .A(n11825), .ZN(n6868) );
  NAND2_X1 U7726 ( .A1(n11825), .A2(n6866), .ZN(n6865) );
  OR2_X1 U7727 ( .A1(n11830), .A2(n11828), .ZN(n7413) );
  INV_X1 U7728 ( .A(n7881), .ZN(n7883) );
  NAND2_X1 U7729 ( .A1(n12666), .A2(n6787), .ZN(n6786) );
  INV_X1 U7730 ( .A(n12503), .ZN(n6787) );
  NAND2_X1 U7731 ( .A1(n6790), .A2(n12697), .ZN(n6789) );
  NAND2_X1 U7732 ( .A1(n6792), .A2(n6791), .ZN(n6790) );
  NAND2_X1 U7733 ( .A1(n12395), .A2(n6610), .ZN(n6791) );
  NAND2_X1 U7734 ( .A1(n6794), .A2(n6793), .ZN(n6792) );
  NOR2_X1 U7735 ( .A1(n12500), .A2(n12676), .ZN(n6788) );
  INV_X1 U7736 ( .A(n8567), .ZN(n7290) );
  NOR2_X1 U7737 ( .A1(n11006), .A2(n7119), .ZN(n7118) );
  NOR2_X1 U7738 ( .A1(n10884), .A2(n7120), .ZN(n7119) );
  INV_X1 U7739 ( .A(n8293), .ZN(n7120) );
  NAND2_X1 U7740 ( .A1(n7029), .A2(n8075), .ZN(n7028) );
  NOR2_X1 U7741 ( .A1(n6948), .A2(n7980), .ZN(n6947) );
  INV_X1 U7742 ( .A(n6951), .ZN(n6948) );
  AOI21_X1 U7743 ( .B1(n7947), .B2(n6960), .A(n6959), .ZN(n6958) );
  INV_X1 U7744 ( .A(n7961), .ZN(n6959) );
  AOI21_X1 U7745 ( .B1(n7947), .B2(n7946), .A(SI_26_), .ZN(n6957) );
  AOI21_X1 U7746 ( .B1(n7809), .B2(n6974), .A(n6972), .ZN(n6971) );
  INV_X1 U7747 ( .A(n7849), .ZN(n6972) );
  AOI21_X1 U7748 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n7849) );
  INV_X1 U7749 ( .A(n7194), .ZN(n6964) );
  INV_X1 U7750 ( .A(n6858), .ZN(n6857) );
  OAI21_X1 U7751 ( .B1(n7600), .B2(n6859), .A(n7614), .ZN(n6858) );
  INV_X1 U7752 ( .A(n7603), .ZN(n6859) );
  OR2_X1 U7753 ( .A1(n10627), .A2(n6807), .ZN(n6806) );
  NOR2_X1 U7754 ( .A1(n10624), .A2(n10450), .ZN(n6807) );
  NAND2_X1 U7755 ( .A1(n12571), .A2(n6612), .ZN(n12572) );
  OR2_X1 U7756 ( .A1(n12605), .A2(n12604), .ZN(n12607) );
  INV_X1 U7757 ( .A(n14316), .ZN(n6848) );
  INV_X1 U7758 ( .A(n12565), .ZN(n6802) );
  INV_X1 U7759 ( .A(n14324), .ZN(n6800) );
  NAND2_X1 U7760 ( .A1(n12506), .A2(n12505), .ZN(n7081) );
  INV_X1 U7761 ( .A(n9359), .ZN(n7066) );
  OR2_X1 U7762 ( .A1(n12215), .A2(n12275), .ZN(n12481) );
  INV_X1 U7763 ( .A(n9511), .ZN(n7002) );
  INV_X1 U7764 ( .A(n7062), .ZN(n7061) );
  OAI21_X1 U7765 ( .B1(n12358), .B2(n7063), .A(n12435), .ZN(n7062) );
  INV_X1 U7766 ( .A(n12432), .ZN(n7063) );
  INV_X1 U7767 ( .A(n12529), .ZN(n9543) );
  OAI21_X1 U7768 ( .B1(n9414), .B2(n7276), .A(n7274), .ZN(n9001) );
  AOI21_X1 U7769 ( .B1(n7277), .B2(n7275), .A(n6622), .ZN(n7274) );
  INV_X1 U7770 ( .A(n7277), .ZN(n7276) );
  NAND2_X1 U7771 ( .A1(n9380), .A2(n8993), .ZN(n8994) );
  INV_X1 U7772 ( .A(n8973), .ZN(n7251) );
  NAND2_X1 U7773 ( .A1(n13074), .A2(n12004), .ZN(n7329) );
  INV_X1 U7774 ( .A(n13044), .ZN(n7316) );
  INV_X1 U7775 ( .A(n11983), .ZN(n7319) );
  INV_X1 U7776 ( .A(n13024), .ZN(n7338) );
  OAI211_X1 U7777 ( .C1(n8856), .C2(n8855), .A(n8857), .B(n8825), .ZN(n8826)
         );
  INV_X1 U7778 ( .A(n6832), .ZN(n6830) );
  NOR2_X1 U7779 ( .A1(n13377), .A2(n6822), .ZN(n6821) );
  INV_X1 U7780 ( .A(n8591), .ZN(n6822) );
  INV_X1 U7781 ( .A(n7285), .ZN(n7284) );
  OAI21_X1 U7782 ( .B1(n7128), .B2(n7290), .A(n8902), .ZN(n7285) );
  INV_X1 U7783 ( .A(n8561), .ZN(n7294) );
  XNOR2_X1 U7784 ( .A(n13126), .B(n10413), .ZN(n8905) );
  INV_X1 U7785 ( .A(n10306), .ZN(n8904) );
  INV_X1 U7786 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8166) );
  AND3_X1 U7787 ( .A1(n6572), .A2(n8143), .A3(n8129), .ZN(n8632) );
  INV_X1 U7788 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U7789 ( .A1(n8143), .A2(n8129), .ZN(n8130) );
  INV_X1 U7790 ( .A(n12061), .ZN(n7172) );
  INV_X1 U7791 ( .A(n13882), .ZN(n6731) );
  OAI21_X1 U7792 ( .B1(n6736), .B2(n13882), .A(n13883), .ZN(n6735) );
  NOR2_X1 U7793 ( .A1(n13918), .A2(n6733), .ZN(n6732) );
  INV_X1 U7794 ( .A(n8092), .ZN(n6733) );
  AND2_X1 U7795 ( .A1(n14005), .A2(n8084), .ZN(n7056) );
  INV_X1 U7796 ( .A(n7807), .ZN(n7233) );
  INV_X1 U7797 ( .A(n11798), .ZN(n7230) );
  NAND2_X1 U7798 ( .A1(n14507), .A2(n7739), .ZN(n11775) );
  OR2_X1 U7799 ( .A1(n14507), .A2(n7739), .ZN(n11774) );
  NOR2_X1 U7800 ( .A1(n11757), .A2(n14489), .ZN(n6897) );
  INV_X1 U7801 ( .A(n6477), .ZN(n7029) );
  NAND2_X1 U7802 ( .A1(n7033), .A2(n8070), .ZN(n6714) );
  NAND2_X1 U7803 ( .A1(n7053), .A2(n7048), .ZN(n7051) );
  NOR2_X1 U7804 ( .A1(n8064), .A2(n7052), .ZN(n7048) );
  INV_X1 U7805 ( .A(n8062), .ZN(n7052) );
  NAND2_X1 U7806 ( .A1(n14020), .A2(n14024), .ZN(n8085) );
  OAI21_X1 U7807 ( .B1(n8465), .B2(n7898), .A(n7897), .ZN(n7913) );
  XNOR2_X1 U7808 ( .A(n7770), .B(SI_14_), .ZN(n7741) );
  NAND2_X1 U7809 ( .A1(n7690), .A2(n15176), .ZN(n7706) );
  INV_X1 U7810 ( .A(n7193), .ZN(n7192) );
  OAI21_X1 U7811 ( .B1(n6516), .B2(n7650), .A(n7670), .ZN(n7193) );
  NAND2_X1 U7812 ( .A1(n7631), .A2(n7630), .ZN(n6944) );
  NAND2_X1 U7813 ( .A1(n14179), .A2(n14178), .ZN(n14180) );
  OR2_X1 U7814 ( .A1(n14213), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U7815 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n14184), .A(n14183), .ZN(
        n14185) );
  NAND2_X1 U7816 ( .A1(n14235), .A2(n14236), .ZN(n14183) );
  OAI21_X1 U7817 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14954), .A(n14190), .ZN(
        n14192) );
  AOI21_X1 U7818 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14196), .A(n14195), .ZN(
        n14247) );
  NAND2_X1 U7819 ( .A1(n7385), .A2(n9433), .ZN(n7384) );
  INV_X1 U7820 ( .A(n9638), .ZN(n7388) );
  AOI21_X1 U7821 ( .B1(n9677), .B2(n12535), .A(n12173), .ZN(n12176) );
  NOR2_X1 U7822 ( .A1(n12223), .A2(n7375), .ZN(n7374) );
  INV_X1 U7823 ( .A(n7437), .ZN(n7375) );
  AND2_X1 U7824 ( .A1(n12242), .A2(n9667), .ZN(n12265) );
  NAND2_X1 U7825 ( .A1(n9657), .A2(n9656), .ZN(n9658) );
  NOR2_X1 U7826 ( .A1(n7381), .A2(n7382), .ZN(n7380) );
  INV_X1 U7827 ( .A(n9672), .ZN(n7382) );
  NOR2_X1 U7828 ( .A1(n12241), .A2(n12242), .ZN(n7381) );
  NAND2_X1 U7829 ( .A1(n12513), .A2(n6778), .ZN(n6775) );
  NOR2_X1 U7830 ( .A1(n12513), .A2(n6777), .ZN(n6772) );
  AND4_X1 U7831 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(n9640)
         );
  OAI21_X1 U7832 ( .B1(n10182), .B2(n10061), .A(n10062), .ZN(n10165) );
  NAND2_X1 U7833 ( .A1(n10446), .A2(n10445), .ZN(n6805) );
  NOR2_X1 U7834 ( .A1(n6514), .A2(n10462), .ZN(n10623) );
  NOR2_X1 U7835 ( .A1(n10452), .A2(n10451), .ZN(n10627) );
  OR2_X1 U7836 ( .A1(n10623), .A2(n6884), .ZN(n10749) );
  NOR2_X1 U7837 ( .A1(n10624), .A2(n15079), .ZN(n6884) );
  NAND2_X1 U7838 ( .A1(n6885), .A2(n6611), .ZN(n11187) );
  NOR2_X1 U7839 ( .A1(n12556), .A2(n6810), .ZN(n12558) );
  AND2_X1 U7840 ( .A1(n12557), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6810) );
  XNOR2_X1 U7841 ( .A(n12572), .B(n12593), .ZN(n14958) );
  INV_X1 U7842 ( .A(n14973), .ZN(n7100) );
  NOR2_X1 U7843 ( .A1(n14967), .A2(n14966), .ZN(n14965) );
  NAND2_X1 U7844 ( .A1(n14984), .A2(n6843), .ZN(n15001) );
  OR2_X1 U7845 ( .A1(n12595), .A2(n12596), .ZN(n6843) );
  NAND2_X1 U7846 ( .A1(n14303), .A2(n12580), .ZN(n14320) );
  AND2_X1 U7847 ( .A1(n14307), .A2(n14308), .ZN(n14305) );
  NAND2_X1 U7848 ( .A1(n14333), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14332) );
  AOI21_X1 U7849 ( .B1(n7074), .B2(n7076), .A(n7072), .ZN(n7071) );
  NAND2_X1 U7850 ( .A1(n12680), .A2(n7074), .ZN(n7073) );
  INV_X1 U7851 ( .A(n12393), .ZN(n7072) );
  AOI21_X1 U7852 ( .B1(n6525), .B2(n7088), .A(n6495), .ZN(n7084) );
  NAND2_X1 U7853 ( .A1(n6525), .A2(n7083), .ZN(n7082) );
  NAND2_X1 U7854 ( .A1(n9653), .A2(n12538), .ZN(n7006) );
  NAND2_X1 U7855 ( .A1(n6577), .A2(n12487), .ZN(n7088) );
  OR2_X1 U7856 ( .A1(n12355), .A2(n12354), .ZN(n12726) );
  NOR2_X1 U7857 ( .A1(n12738), .A2(n12740), .ZN(n7089) );
  NOR2_X1 U7858 ( .A1(n6522), .A2(n7069), .ZN(n7068) );
  INV_X1 U7859 ( .A(n12478), .ZN(n7069) );
  NAND2_X1 U7860 ( .A1(n12777), .A2(n9359), .ZN(n7070) );
  INV_X1 U7861 ( .A(n12781), .ZN(n7009) );
  AOI21_X1 U7862 ( .B1(n6980), .B2(n6983), .A(n6530), .ZN(n6977) );
  INV_X1 U7863 ( .A(n9514), .ZN(n6983) );
  AOI21_X1 U7864 ( .B1(n10057), .B2(n9102), .A(n12514), .ZN(n12829) );
  CLKBUF_X1 U7865 ( .A(n11491), .Z(n11492) );
  CLKBUF_X1 U7866 ( .A(n11274), .Z(n11275) );
  AND2_X1 U7867 ( .A1(n12438), .A2(n12439), .ZN(n12435) );
  NOR2_X1 U7868 ( .A1(n9135), .A2(n9134), .ZN(n9587) );
  INV_X1 U7869 ( .A(n12829), .ZN(n15040) );
  NOR2_X1 U7870 ( .A1(n9542), .A2(n9541), .ZN(n10809) );
  NAND2_X1 U7871 ( .A1(n7394), .A2(n7393), .ZN(n7392) );
  NOR2_X1 U7872 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n7394) );
  NAND2_X1 U7873 ( .A1(n7393), .A2(n7018), .ZN(n7017) );
  NAND2_X1 U7874 ( .A1(n9006), .A2(n9005), .ZN(n9461) );
  XNOR2_X1 U7875 ( .A(n9056), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U7876 ( .A1(n9038), .A2(n9037), .ZN(n9041) );
  AND2_X1 U7877 ( .A1(n8988), .A2(n8987), .ZN(n9342) );
  NAND2_X1 U7878 ( .A1(n9328), .A2(n8986), .ZN(n9343) );
  NAND2_X1 U7879 ( .A1(n9343), .A2(n9342), .ZN(n9345) );
  NAND2_X1 U7880 ( .A1(n9310), .A2(n8984), .ZN(n9326) );
  AND2_X1 U7881 ( .A1(n8973), .A2(n8972), .ZN(n9240) );
  NAND2_X1 U7882 ( .A1(n9241), .A2(n9240), .ZN(n9243) );
  INV_X1 U7883 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9245) );
  INV_X1 U7884 ( .A(n7243), .ZN(n7242) );
  OAI21_X1 U7885 ( .B1(n7245), .B2(n7244), .A(n9210), .ZN(n7243) );
  INV_X1 U7886 ( .A(n8966), .ZN(n7244) );
  NAND2_X1 U7887 ( .A1(n8964), .A2(n7245), .ZN(n9194) );
  INV_X1 U7888 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9122) );
  AND2_X1 U7889 ( .A1(n11560), .A2(n11558), .ZN(n7348) );
  OR2_X1 U7890 ( .A1(n12969), .A2(n7331), .ZN(n7330) );
  INV_X1 U7891 ( .A(n12004), .ZN(n7331) );
  INV_X1 U7892 ( .A(n12012), .ZN(n7326) );
  AND2_X1 U7893 ( .A1(n11986), .A2(n11985), .ZN(n11987) );
  NAND2_X1 U7894 ( .A1(n7341), .A2(n7340), .ZN(n10503) );
  INV_X1 U7895 ( .A(n10367), .ZN(n7339) );
  INV_X1 U7896 ( .A(n11106), .ZN(n11103) );
  AOI21_X2 U7897 ( .B1(n12990), .B2(n12986), .A(n12988), .ZN(n13043) );
  NAND2_X1 U7898 ( .A1(n13043), .A2(n13044), .ZN(n13042) );
  AND4_X1 U7899 ( .A1(n8516), .A2(n8515), .A3(n8514), .A4(n8513), .ZN(n13005)
         );
  OR2_X1 U7900 ( .A1(n8545), .A2(n8168), .ZN(n8172) );
  OR2_X1 U7901 ( .A1(n8489), .A2(n8169), .ZN(n8171) );
  NOR2_X1 U7902 ( .A1(n13212), .A2(n6941), .ZN(n6940) );
  INV_X1 U7903 ( .A(n8921), .ZN(n13253) );
  NAND2_X1 U7904 ( .A1(n7314), .A2(n8604), .ZN(n13259) );
  NAND2_X1 U7905 ( .A1(n13274), .A2(n8603), .ZN(n7314) );
  NAND2_X1 U7906 ( .A1(n8495), .A2(n6523), .ZN(n13278) );
  NOR2_X1 U7907 ( .A1(n13328), .A2(n6928), .ZN(n13297) );
  AOI21_X1 U7908 ( .B1(n6499), .B2(n6827), .A(n6554), .ZN(n6823) );
  AOI21_X1 U7909 ( .B1(n7313), .B2(n13339), .A(n6561), .ZN(n6826) );
  OR2_X1 U7910 ( .A1(n13343), .A2(n6827), .ZN(n6825) );
  AND2_X1 U7911 ( .A1(n8917), .A2(n8599), .ZN(n7313) );
  OAI21_X1 U7912 ( .B1(n13356), .B2(n8449), .A(n8450), .ZN(n13340) );
  NAND2_X1 U7913 ( .A1(n13343), .A2(n13342), .ZN(n13341) );
  NAND2_X1 U7914 ( .A1(n11667), .A2(n8588), .ZN(n13391) );
  NAND2_X1 U7915 ( .A1(n8582), .A2(n7312), .ZN(n7310) );
  AND2_X1 U7916 ( .A1(n6538), .A2(n8581), .ZN(n7312) );
  AOI21_X1 U7917 ( .B1(n7135), .B2(n7133), .A(n7132), .ZN(n7131) );
  INV_X1 U7918 ( .A(n7135), .ZN(n7134) );
  NAND2_X1 U7919 ( .A1(n8341), .A2(n7137), .ZN(n7136) );
  NAND2_X1 U7920 ( .A1(n7136), .A2(n7135), .ZN(n14405) );
  NAND2_X1 U7921 ( .A1(n8349), .A2(n8348), .ZN(n11431) );
  INV_X1 U7922 ( .A(n8576), .ZN(n7306) );
  NOR2_X1 U7923 ( .A1(n10307), .A2(n7294), .ZN(n7291) );
  OAI21_X1 U7924 ( .B1(n8904), .B2(n7294), .A(n8905), .ZN(n7293) );
  OAI21_X1 U7925 ( .B1(n10249), .B2(n10248), .A(n8678), .ZN(n10267) );
  NAND2_X1 U7926 ( .A1(n8674), .A2(n10683), .ZN(n8179) );
  NAND2_X1 U7927 ( .A1(n10248), .A2(n10244), .ZN(n10243) );
  NAND2_X1 U7928 ( .A1(n13239), .A2(n13238), .ZN(n6634) );
  NAND2_X1 U7929 ( .A1(n6836), .A2(n6834), .ZN(n13236) );
  OR3_X1 U7930 ( .A1(n13266), .A2(n13265), .A3(n13295), .ZN(n13429) );
  NAND2_X1 U7931 ( .A1(n8391), .A2(n8390), .ZN(n13488) );
  OR2_X1 U7932 ( .A1(n8864), .A2(n9711), .ZN(n6632) );
  NAND2_X1 U7933 ( .A1(n7363), .A2(n8166), .ZN(n7362) );
  INV_X1 U7934 ( .A(n7364), .ZN(n7363) );
  NAND2_X1 U7935 ( .A1(n8152), .A2(n8123), .ZN(n8639) );
  AND2_X2 U7936 ( .A1(n8632), .A2(n8151), .ZN(n8152) );
  NOR3_X1 U7937 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n8151) );
  INV_X1 U7938 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7365) );
  CLKBUF_X1 U7939 ( .A(n8639), .Z(n8640) );
  OR2_X1 U7940 ( .A1(n8635), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8637) );
  AND2_X1 U7941 ( .A1(n8120), .A2(n8188), .ZN(n8264) );
  OR2_X1 U7942 ( .A1(n8209), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8219) );
  AND2_X1 U7943 ( .A1(n13626), .A2(n12116), .ZN(n13572) );
  AND2_X1 U7944 ( .A1(n13609), .A2(n12126), .ZN(n13627) );
  NAND2_X1 U7945 ( .A1(n11162), .A2(n7182), .ZN(n7181) );
  NOR2_X1 U7946 ( .A1(n11164), .A2(n7183), .ZN(n7182) );
  INV_X1 U7947 ( .A(n11161), .ZN(n7183) );
  INV_X1 U7948 ( .A(n10335), .ZN(n10233) );
  NAND2_X1 U7949 ( .A1(n12046), .A2(n12045), .ZN(n6675) );
  AND4_X1 U7950 ( .A1(n7878), .A2(n7877), .A3(n7876), .A4(n7875), .ZN(n13656)
         );
  AND2_X1 U7951 ( .A1(n7493), .A2(n7492), .ZN(n7412) );
  NAND2_X1 U7952 ( .A1(n11850), .A2(n11849), .ZN(n11919) );
  OAI21_X1 U7953 ( .B1(n13885), .B2(n11918), .A(n7025), .ZN(n13860) );
  NAND2_X1 U7954 ( .A1(n11941), .A2(n11942), .ZN(n11940) );
  NAND2_X1 U7955 ( .A1(n13885), .A2(n8094), .ZN(n11941) );
  NAND2_X1 U7956 ( .A1(n7916), .A2(n7915), .ZN(n13928) );
  NAND2_X1 U7957 ( .A1(n13987), .A2(n13971), .ZN(n13968) );
  NOR2_X1 U7958 ( .A1(n7198), .A2(n6728), .ZN(n6727) );
  INV_X1 U7959 ( .A(n14024), .ZN(n6728) );
  NAND2_X1 U7960 ( .A1(n8085), .A2(n7056), .ZN(n14004) );
  NAND2_X1 U7961 ( .A1(n11597), .A2(n8081), .ZN(n11648) );
  OR2_X1 U7962 ( .A1(n11648), .A2(n7236), .ZN(n11650) );
  NAND2_X1 U7963 ( .A1(n11518), .A2(n11512), .ZN(n7213) );
  NAND2_X1 U7964 ( .A1(n7213), .A2(n7212), .ZN(n11597) );
  AND2_X1 U7965 ( .A1(n11784), .A2(n11908), .ZN(n7212) );
  INV_X1 U7966 ( .A(n7738), .ZN(n11451) );
  NAND2_X1 U7967 ( .A1(n11319), .A2(n11905), .ZN(n6711) );
  NAND2_X1 U7968 ( .A1(n8074), .A2(n6477), .ZN(n11086) );
  NAND2_X1 U7969 ( .A1(n7666), .A2(n6477), .ZN(n6680) );
  NAND2_X1 U7970 ( .A1(n6703), .A2(n7029), .ZN(n11079) );
  CLKBUF_X1 U7971 ( .A(n11080), .Z(n6703) );
  OAI21_X1 U7972 ( .B1(n10648), .B2(n7035), .A(n7033), .ZN(n10724) );
  INV_X1 U7973 ( .A(n7612), .ZN(n7218) );
  NAND2_X1 U7974 ( .A1(n11034), .A2(n11041), .ZN(n11036) );
  NAND2_X1 U7975 ( .A1(n7038), .A2(n8067), .ZN(n11042) );
  NAND2_X1 U7976 ( .A1(n10648), .A2(n8066), .ZN(n7038) );
  NAND3_X1 U7977 ( .A1(n10640), .A2(n7227), .A3(n7223), .ZN(n10639) );
  OAI21_X1 U7978 ( .B1(n7580), .B2(n7225), .A(n7581), .ZN(n7227) );
  INV_X1 U7979 ( .A(n10391), .ZN(n7225) );
  NAND2_X1 U7980 ( .A1(n10531), .A2(n11895), .ZN(n10530) );
  OR2_X1 U7981 ( .A1(n11852), .A2(n7519), .ZN(n7520) );
  OR2_X1 U7982 ( .A1(n6472), .A2(n7518), .ZN(n7521) );
  NAND2_X1 U7983 ( .A1(n10355), .A2(n11892), .ZN(n7053) );
  INV_X1 U7984 ( .A(n14045), .ZN(n14008) );
  NAND2_X1 U7985 ( .A1(n14126), .A2(n11688), .ZN(n10127) );
  INV_X1 U7986 ( .A(n13723), .ZN(n10565) );
  OR2_X1 U7987 ( .A1(n11872), .A2(n13726), .ZN(n14045) );
  NOR2_X1 U7988 ( .A1(n6895), .A2(n6894), .ZN(n6893) );
  INV_X1 U7989 ( .A(n14509), .ZN(n14126) );
  NAND2_X1 U7990 ( .A1(n7757), .A2(n7756), .ZN(n12047) );
  NAND2_X1 U7991 ( .A1(n10469), .A2(n7965), .ZN(n7757) );
  NAND2_X1 U7992 ( .A1(n11691), .A2(n7151), .ZN(n14509) );
  XNOR2_X1 U7993 ( .A(n8838), .B(n8837), .ZN(n13536) );
  OAI22_X1 U7994 ( .A1(n8863), .A2(n8861), .B1(n8835), .B2(n15215), .ZN(n8838)
         );
  INV_X1 U7995 ( .A(n7433), .ZN(n7431) );
  NAND2_X1 U7996 ( .A1(n6949), .A2(n6951), .ZN(n7981) );
  BUF_X1 U7997 ( .A(n8017), .Z(n8018) );
  XNOR2_X1 U7998 ( .A(n8016), .B(n8015), .ZN(n8030) );
  INV_X1 U7999 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U8000 ( .A(n7913), .B(n7912), .ZN(n7911) );
  XNOR2_X1 U8001 ( .A(n7832), .B(n7831), .ZN(n10952) );
  NAND2_X1 U8002 ( .A1(n6926), .A2(n14237), .ZN(n14240) );
  AOI21_X1 U8003 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14203), .A(n14202), .ZN(
        n14206) );
  AND2_X1 U8004 ( .A1(n9593), .A2(n9495), .ZN(n9595) );
  INV_X1 U8005 ( .A(n12539), .ZN(n12730) );
  NAND2_X1 U8006 ( .A1(n9601), .A2(n12552), .ZN(n7372) );
  NAND2_X1 U8007 ( .A1(n9393), .A2(n9392), .ZN(n12486) );
  AND4_X1 U8008 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n12325)
         );
  AND4_X1 U8009 ( .A1(n9258), .A2(n9257), .A3(n9256), .A4(n9255), .ZN(n12290)
         );
  INV_X1 U8010 ( .A(n14867), .ZN(n12326) );
  AND3_X1 U8011 ( .A1(n10057), .A2(n12504), .A3(n9102), .ZN(n12827) );
  NAND4_X1 U8012 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), .ZN(n12678)
         );
  INV_X1 U8013 ( .A(n12669), .ZN(n12536) );
  INV_X1 U8014 ( .A(n12277), .ZN(n12744) );
  INV_X1 U8015 ( .A(n12290), .ZN(n12544) );
  NAND4_X2 U8016 ( .A1(n9173), .A2(n9172), .A3(n9171), .A4(n9170), .ZN(n12549)
         );
  OAI21_X1 U8017 ( .B1(n14923), .B2(n14920), .A(n10443), .ZN(n10622) );
  AND2_X1 U8018 ( .A1(n10066), .A2(n10058), .ZN(n14355) );
  INV_X1 U8019 ( .A(n14356), .ZN(n7104) );
  AND2_X1 U8020 ( .A1(n10066), .A2(n12586), .ZN(n15014) );
  INV_X1 U8021 ( .A(n9571), .ZN(n7015) );
  OAI21_X1 U8022 ( .B1(n9524), .B2(n6989), .A(n6987), .ZN(n9558) );
  NAND2_X1 U8023 ( .A1(n9367), .A2(n9366), .ZN(n12885) );
  NAND2_X1 U8024 ( .A1(n10810), .A2(n15032), .ZN(n15045) );
  NAND2_X1 U8025 ( .A1(n12337), .A2(n12336), .ZN(n12900) );
  NAND2_X1 U8026 ( .A1(n7014), .A2(n6494), .ZN(n9580) );
  NAND2_X1 U8027 ( .A1(n15076), .A2(n14383), .ZN(n12952) );
  INV_X1 U8028 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9031) );
  CLKBUF_X1 U8029 ( .A(n11262), .Z(n6650) );
  NAND2_X1 U8030 ( .A1(n8452), .A2(n8451), .ZN(n13348) );
  AND2_X1 U8031 ( .A1(n11995), .A2(n11996), .ZN(n6664) );
  NAND2_X1 U8032 ( .A1(n10205), .A2(n7342), .ZN(n7341) );
  NOR2_X1 U8033 ( .A1(n10368), .A2(n7343), .ZN(n7342) );
  INV_X1 U8034 ( .A(n10204), .ZN(n7343) );
  NAND2_X1 U8035 ( .A1(n9960), .A2(n9959), .ZN(n13091) );
  NAND2_X1 U8036 ( .A1(n9954), .A2(n13300), .ZN(n13095) );
  AOI211_X1 U8037 ( .C1(n8929), .C2(n8670), .A(n10282), .B(n8928), .ZN(n8931)
         );
  NAND2_X1 U8038 ( .A1(n6668), .A2(n6667), .ZN(n14666) );
  OR2_X1 U8039 ( .A1(n14660), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U8040 ( .A1(n14660), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6667) );
  INV_X1 U8041 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6698) );
  OR3_X1 U8042 ( .A1(n13248), .A2(n13247), .A3(n13295), .ZN(n13426) );
  NAND2_X1 U8043 ( .A1(n9953), .A2(n14791), .ZN(n13300) );
  AND2_X1 U8044 ( .A1(n6961), .A2(n6626), .ZN(n13218) );
  NAND2_X1 U8045 ( .A1(n13539), .A2(n6474), .ZN(n6961) );
  INV_X1 U8046 ( .A(n13218), .ZN(n8850) );
  NAND2_X1 U8047 ( .A1(n13229), .A2(n13228), .ZN(n13421) );
  NOR2_X1 U8048 ( .A1(n6634), .A2(n6633), .ZN(n7146) );
  INV_X1 U8049 ( .A(n7146), .ZN(n7140) );
  NAND2_X1 U8050 ( .A1(n7143), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7145) );
  OAI21_X1 U8051 ( .B1(n13677), .B2(n12146), .A(n7175), .ZN(n13562) );
  NAND2_X1 U8052 ( .A1(n13676), .A2(n6503), .ZN(n6647) );
  NOR2_X1 U8053 ( .A1(n13569), .A2(n13699), .ZN(n6706) );
  CLKBUF_X1 U8054 ( .A(n11471), .Z(n6682) );
  NAND2_X1 U8055 ( .A1(n6682), .A2(n11470), .ZN(n14482) );
  NAND2_X1 U8056 ( .A1(n10233), .A2(n10337), .ZN(n10338) );
  INV_X1 U8057 ( .A(n10336), .ZN(n10337) );
  AOI21_X1 U8058 ( .B1(n7175), .B2(n12146), .A(n12157), .ZN(n7174) );
  NAND2_X1 U8059 ( .A1(n6708), .A2(n6551), .ZN(n10115) );
  INV_X1 U8060 ( .A(n10114), .ZN(n7150) );
  INV_X1 U8061 ( .A(n13971), .ZN(n14109) );
  AOI21_X1 U8062 ( .B1(n7168), .B2(n7166), .A(n7164), .ZN(n7163) );
  INV_X1 U8063 ( .A(n7166), .ZN(n7165) );
  INV_X1 U8064 ( .A(n11641), .ZN(n7164) );
  AND4_X1 U8065 ( .A1(n7765), .A2(n7764), .A3(n7763), .A4(n7762), .ZN(n14462)
         );
  INV_X1 U8066 ( .A(n13991), .ZN(n14115) );
  AND2_X1 U8067 ( .A1(n13580), .A2(n14124), .ZN(n14490) );
  XNOR2_X1 U8068 ( .A(n10336), .B(n10233), .ZN(n10237) );
  INV_X1 U8069 ( .A(n14467), .ZN(n14483) );
  AND2_X1 U8070 ( .A1(n11884), .A2(n11883), .ZN(n11886) );
  OR2_X1 U8071 ( .A1(n11872), .A2(n8098), .ZN(n14021) );
  NAND3_X2 U8072 ( .A1(n7472), .A2(n6644), .A3(n7471), .ZN(n13722) );
  NAND2_X1 U8073 ( .A1(n7538), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7472) );
  AND2_X1 U8074 ( .A1(n7469), .A2(n7470), .ZN(n6644) );
  AOI21_X1 U8075 ( .B1(n8100), .B2(n14028), .A(n8099), .ZN(n14067) );
  AND2_X1 U8076 ( .A1(n13702), .A2(n14006), .ZN(n8099) );
  INV_X1 U8077 ( .A(n11920), .ZN(n8009) );
  NAND2_X1 U8078 ( .A1(n9746), .A2(n6534), .ZN(n7488) );
  INV_X1 U8079 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7429) );
  INV_X1 U8080 ( .A(n7432), .ZN(n7430) );
  NOR2_X1 U8081 ( .A1(n14524), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U8082 ( .A1(n6918), .A2(n14535), .ZN(n6917) );
  NAND2_X1 U8083 ( .A1(n14534), .A2(n14533), .ZN(n6918) );
  NAND2_X1 U8084 ( .A1(n8674), .A2(n8675), .ZN(n6691) );
  NAND2_X1 U8085 ( .A1(n6669), .A2(n6671), .ZN(n8685) );
  NAND2_X1 U8086 ( .A1(n10265), .A2(n8867), .ZN(n6671) );
  INV_X1 U8087 ( .A(n8699), .ZN(n7367) );
  NAND2_X1 U8088 ( .A1(n8710), .A2(n8708), .ZN(n7360) );
  INV_X1 U8089 ( .A(n8719), .ZN(n7351) );
  OR2_X1 U8090 ( .A1(n7424), .A2(n11723), .ZN(n7423) );
  INV_X1 U8091 ( .A(n11722), .ZN(n7424) );
  INV_X1 U8092 ( .A(n11735), .ZN(n7421) );
  NAND2_X1 U8093 ( .A1(n8736), .A2(n7355), .ZN(n7354) );
  NAND2_X1 U8094 ( .A1(n8754), .A2(n8756), .ZN(n7350) );
  OAI21_X1 U8095 ( .B1(n6685), .B2(n6686), .A(n7352), .ZN(n8775) );
  NAND2_X1 U8096 ( .A1(n8771), .A2(n7353), .ZN(n7352) );
  AOI21_X1 U8097 ( .B1(n8766), .B2(n8767), .A(n6658), .ZN(n6686) );
  NOR2_X1 U8098 ( .A1(n7402), .A2(n7401), .ZN(n7400) );
  OAI21_X1 U8099 ( .B1(n11788), .B2(n11787), .A(n11786), .ZN(n7402) );
  NAND2_X1 U8100 ( .A1(n6740), .A2(n12407), .ZN(n12413) );
  AND2_X1 U8101 ( .A1(n11803), .A2(n14005), .ZN(n6861) );
  INV_X1 U8102 ( .A(n12463), .ZN(n6759) );
  AOI21_X1 U8103 ( .B1(n6764), .B2(n6765), .A(n6763), .ZN(n6762) );
  INV_X1 U8104 ( .A(n12450), .ZN(n6763) );
  AND2_X1 U8105 ( .A1(n12821), .A2(n6758), .ZN(n6757) );
  NAND2_X1 U8106 ( .A1(n6556), .A2(n12463), .ZN(n6758) );
  NOR2_X1 U8107 ( .A1(n6874), .A2(n6876), .ZN(n6873) );
  AND2_X1 U8108 ( .A1(n6872), .A2(n6871), .ZN(n6870) );
  AOI21_X1 U8109 ( .B1(n6751), .B2(n6749), .A(n6748), .ZN(n12473) );
  NOR2_X1 U8110 ( .A1(n6754), .A2(n6750), .ZN(n6749) );
  OAI21_X1 U8111 ( .B1(n6752), .B2(n6750), .A(n6609), .ZN(n6748) );
  NAND2_X1 U8112 ( .A1(n7358), .A2(n8796), .ZN(n7357) );
  AND2_X1 U8113 ( .A1(n11827), .A2(n6868), .ZN(n6867) );
  NOR2_X1 U8114 ( .A1(n12494), .A2(n12705), .ZN(n6793) );
  OR2_X1 U8115 ( .A1(n11692), .A2(n8056), .ZN(n11693) );
  AND2_X1 U8116 ( .A1(n7946), .A2(SI_26_), .ZN(n6960) );
  INV_X1 U8117 ( .A(n7808), .ZN(n7811) );
  INV_X1 U8118 ( .A(n7688), .ZN(n7191) );
  INV_X1 U8119 ( .A(n12512), .ZN(n6783) );
  NOR2_X1 U8120 ( .A1(n12517), .A2(n12518), .ZN(n6785) );
  NAND2_X1 U8121 ( .A1(n12911), .A2(n12670), .ZN(n6993) );
  AND2_X1 U8122 ( .A1(n9020), .A2(n7396), .ZN(n6853) );
  AOI21_X1 U8123 ( .B1(n9413), .B2(n9000), .A(n7278), .ZN(n7277) );
  INV_X1 U8124 ( .A(n9423), .ZN(n7278) );
  INV_X1 U8125 ( .A(n9000), .ZN(n7275) );
  INV_X1 U8126 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9019) );
  INV_X1 U8127 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7391) );
  INV_X1 U8128 ( .A(n8867), .ZN(n6670) );
  INV_X1 U8129 ( .A(n8517), .ZN(n7130) );
  INV_X1 U8130 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U8131 ( .A1(n7415), .A2(n7414), .ZN(n11843) );
  OR2_X1 U8132 ( .A1(n7416), .A2(n11841), .ZN(n7414) );
  OR2_X1 U8133 ( .A1(n6720), .A2(n6717), .ZN(n6713) );
  INV_X1 U8134 ( .A(n8070), .ZN(n6717) );
  NAND2_X1 U8135 ( .A1(n7054), .A2(n6725), .ZN(n6724) );
  INV_X1 U8136 ( .A(n6727), .ZN(n6725) );
  OR2_X1 U8137 ( .A1(n11906), .A2(n7045), .ZN(n7044) );
  INV_X1 U8138 ( .A(n8079), .ZN(n7045) );
  INV_X1 U8139 ( .A(n11774), .ZN(n7041) );
  INV_X1 U8140 ( .A(n6960), .ZN(n6953) );
  INV_X1 U8141 ( .A(n7776), .ZN(n6963) );
  AOI21_X1 U8142 ( .B1(n6574), .B2(n7725), .A(n7195), .ZN(n7194) );
  NOR2_X1 U8143 ( .A1(n7706), .A2(SI_13_), .ZN(n7195) );
  NOR2_X1 U8144 ( .A1(n7725), .A2(n15175), .ZN(n7196) );
  AND2_X1 U8145 ( .A1(n7191), .A2(n6516), .ZN(n7190) );
  AND2_X1 U8146 ( .A1(n9711), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7199) );
  NAND3_X1 U8147 ( .A1(n13201), .A2(n7479), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7206) );
  NOR2_X1 U8148 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7200) );
  NOR2_X1 U8149 ( .A1(n9285), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9298) );
  NOR2_X1 U8150 ( .A1(n9336), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9352) );
  AND2_X1 U8151 ( .A1(n9352), .A2(n12260), .ZN(n9369) );
  NOR2_X1 U8152 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9440), .ZN(n9451) );
  AOI21_X1 U8153 ( .B1(n6789), .B2(n6788), .A(n6786), .ZN(n12510) );
  OAI21_X1 U8154 ( .B1(n12515), .B2(n12378), .A(n12519), .ZN(n6782) );
  NAND2_X1 U8155 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  NAND2_X1 U8156 ( .A1(n9533), .A2(n10168), .ZN(n6840) );
  OR2_X1 U8157 ( .A1(n9533), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8158 ( .A1(n6839), .A2(n10047), .ZN(n10049) );
  AOI21_X1 U8159 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n14902), .A(n14896), .ZN(
        n10448) );
  NAND2_X1 U8160 ( .A1(n14908), .A2(n6557), .ZN(n10460) );
  NOR2_X1 U8161 ( .A1(n11202), .A2(n6811), .ZN(n11204) );
  AND2_X1 U8162 ( .A1(n11203), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U8163 ( .A1(n14975), .A2(n6883), .ZN(n12574) );
  NAND2_X1 U8164 ( .A1(n14981), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8165 ( .A1(n15023), .A2(n12603), .ZN(n12605) );
  NAND2_X1 U8166 ( .A1(n15011), .A2(n12601), .ZN(n12579) );
  NAND2_X1 U8167 ( .A1(n6796), .A2(n12602), .ZN(n12563) );
  AOI21_X1 U8168 ( .B1(n7077), .B2(n7075), .A(n12394), .ZN(n7074) );
  INV_X1 U8169 ( .A(n6527), .ZN(n7075) );
  INV_X1 U8170 ( .A(n7077), .ZN(n7076) );
  AND2_X1 U8171 ( .A1(n6993), .A2(n9523), .ZN(n6992) );
  NAND2_X1 U8172 ( .A1(n6991), .A2(n6993), .ZN(n6990) );
  INV_X1 U8173 ( .A(n12491), .ZN(n7085) );
  OR2_X1 U8174 ( .A1(n12395), .A2(n9433), .ZN(n12497) );
  AND2_X1 U8175 ( .A1(n12454), .A2(n6981), .ZN(n6980) );
  NAND2_X1 U8176 ( .A1(n6982), .A2(n9514), .ZN(n6981) );
  NAND2_X1 U8177 ( .A1(n10867), .A2(n9503), .ZN(n10939) );
  NOR2_X1 U8178 ( .A1(n12333), .A2(n7268), .ZN(n7267) );
  INV_X1 U8179 ( .A(n12188), .ZN(n7268) );
  INV_X1 U8180 ( .A(n9008), .ZN(n7282) );
  INV_X1 U8181 ( .A(n7256), .ZN(n7255) );
  OAI21_X1 U8182 ( .B1(n9342), .B2(n7257), .A(n8990), .ZN(n7256) );
  INV_X1 U8183 ( .A(n8988), .ZN(n7257) );
  AND2_X1 U8184 ( .A1(n8298), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8312) );
  INV_X1 U8185 ( .A(n12009), .ZN(n11975) );
  NOR2_X1 U8186 ( .A1(n8361), .A2(n11566), .ZN(n8374) );
  INV_X1 U8187 ( .A(n8666), .ZN(n10022) );
  OR2_X1 U8188 ( .A1(n8926), .A2(n8860), .ZN(n8879) );
  INV_X1 U8189 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8190 ( .A1(n14708), .A2(n13154), .ZN(n13155) );
  NAND2_X1 U8191 ( .A1(n13519), .A2(n6930), .ZN(n6929) );
  OR2_X1 U8192 ( .A1(n8392), .A2(n13016), .ZN(n8407) );
  INV_X1 U8193 ( .A(n7137), .ZN(n7133) );
  INV_X1 U8194 ( .A(n8899), .ZN(n7301) );
  INV_X1 U8195 ( .A(n7302), .ZN(n6819) );
  INV_X1 U8196 ( .A(n8900), .ZN(n6818) );
  NOR2_X1 U8197 ( .A1(n11263), .A2(n11014), .ZN(n6934) );
  NOR2_X1 U8198 ( .A1(n7299), .A2(n8570), .ZN(n7298) );
  INV_X1 U8199 ( .A(n8569), .ZN(n7299) );
  NAND2_X1 U8200 ( .A1(n11013), .A2(n11151), .ZN(n11014) );
  NAND2_X1 U8201 ( .A1(n7293), .A2(n8563), .ZN(n6815) );
  NAND2_X1 U8202 ( .A1(n8674), .A2(n10246), .ZN(n8678) );
  NAND2_X1 U8203 ( .A1(n11619), .A2(n6498), .ZN(n13399) );
  AOI21_X1 U8204 ( .B1(n7118), .B2(n7120), .A(n6550), .ZN(n7116) );
  NAND2_X1 U8205 ( .A1(n8153), .A2(n7365), .ZN(n7364) );
  CLKBUF_X1 U8206 ( .A(n8294), .Z(n8631) );
  INV_X1 U8207 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8118) );
  INV_X1 U8208 ( .A(n12158), .ZN(n12129) );
  INV_X1 U8209 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7697) );
  INV_X1 U8210 ( .A(n8094), .ZN(n7027) );
  INV_X1 U8211 ( .A(n8095), .ZN(n7026) );
  INV_X1 U8212 ( .A(n13902), .ZN(n7047) );
  INV_X1 U8213 ( .A(n7917), .ZN(n7918) );
  NOR2_X1 U8214 ( .A1(n6904), .A2(n6903), .ZN(n6901) );
  INV_X1 U8215 ( .A(n6721), .ZN(n6720) );
  INV_X1 U8216 ( .A(n7036), .ZN(n7035) );
  AOI21_X1 U8217 ( .B1(n7036), .B2(n7034), .A(n6573), .ZN(n7033) );
  INV_X1 U8218 ( .A(n8066), .ZN(n7034) );
  NOR2_X1 U8219 ( .A1(n7558), .A2(n7228), .ZN(n7226) );
  INV_X1 U8220 ( .A(n7581), .ZN(n7228) );
  NAND2_X1 U8221 ( .A1(n10579), .A2(n10354), .ZN(n11686) );
  NOR2_X1 U8222 ( .A1(n13925), .A2(n14084), .ZN(n13879) );
  NAND2_X1 U8223 ( .A1(n8056), .A2(n11687), .ZN(n11871) );
  NAND3_X1 U8224 ( .A1(n7019), .A2(n7021), .A3(n6521), .ZN(n7020) );
  INV_X1 U8225 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7463) );
  INV_X1 U8226 ( .A(n6947), .ZN(n6946) );
  AOI21_X1 U8227 ( .B1(n6947), .B2(n6956), .A(n6620), .ZN(n6945) );
  AND2_X1 U8228 ( .A1(n7464), .A2(n8019), .ZN(n7433) );
  INV_X1 U8229 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7464) );
  AND2_X1 U8230 ( .A1(n6954), .A2(n6952), .ZN(n6951) );
  NAND2_X1 U8231 ( .A1(n6957), .A2(n6955), .ZN(n6954) );
  NAND2_X1 U8232 ( .A1(n6958), .A2(n6953), .ZN(n6952) );
  INV_X1 U8233 ( .A(n7946), .ZN(n6955) );
  AOI21_X1 U8234 ( .B1(n6971), .B2(n6504), .A(n6969), .ZN(n6968) );
  NAND2_X1 U8235 ( .A1(n6971), .A2(n6607), .ZN(n6970) );
  INV_X1 U8236 ( .A(n7885), .ZN(n6969) );
  INV_X1 U8237 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U8238 ( .A1(n6967), .A2(n6971), .ZN(n7886) );
  NOR2_X1 U8239 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7674) );
  NOR2_X2 U8240 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7748) );
  AOI21_X1 U8241 ( .B1(n6857), .B2(n6859), .A(n6569), .ZN(n6855) );
  INV_X1 U8242 ( .A(n7546), .ZN(n7547) );
  INV_X1 U8243 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U8244 ( .A1(n14174), .A2(n6653), .ZN(n14175) );
  NAND2_X1 U8245 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6654), .ZN(n6653) );
  XNOR2_X1 U8246 ( .A(n14177), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14213) );
  AND2_X1 U8247 ( .A1(n15030), .A2(n6526), .ZN(n9588) );
  OR2_X1 U8248 ( .A1(n9650), .A2(n12730), .ZN(n7437) );
  OR2_X1 U8249 ( .A1(n9268), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9285) );
  AND2_X1 U8250 ( .A1(n12555), .A2(n11678), .ZN(n12400) );
  NOR2_X1 U8251 ( .A1(n9405), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9417) );
  OAI21_X1 U8252 ( .B1(n10047), .B2(n6839), .A(n10049), .ZN(n10176) );
  XNOR2_X1 U8253 ( .A(n6805), .B(n10456), .ZN(n14877) );
  NOR2_X1 U8254 ( .A1(n14884), .A2(n10439), .ZN(n14901) );
  OR2_X1 U8255 ( .A1(n14911), .A2(n14910), .ZN(n14908) );
  XNOR2_X1 U8256 ( .A(n10460), .B(n10447), .ZN(n14929) );
  NAND2_X1 U8257 ( .A1(n14929), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n14928) );
  NAND2_X1 U8258 ( .A1(n7114), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7112) );
  AND2_X1 U8259 ( .A1(n7113), .A2(n7112), .ZN(n10452) );
  INV_X1 U8260 ( .A(n6806), .ZN(n10761) );
  NOR2_X1 U8261 ( .A1(n10767), .A2(n10766), .ZN(n11202) );
  NAND2_X1 U8262 ( .A1(n10750), .A2(n10751), .ZN(n6887) );
  XNOR2_X1 U8263 ( .A(n11204), .B(n14945), .ZN(n14941) );
  AOI21_X1 U8264 ( .B1(n14937), .B2(n14934), .A(n11197), .ZN(n11199) );
  OAI21_X1 U8265 ( .B1(n7107), .B2(n14941), .A(n7106), .ZN(n12556) );
  NAND2_X1 U8266 ( .A1(n7108), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U8267 ( .A1(n11205), .A2(n7108), .ZN(n7106) );
  INV_X1 U8268 ( .A(n11207), .ZN(n7108) );
  NOR2_X1 U8269 ( .A1(n14941), .A2(n14940), .ZN(n14939) );
  NAND2_X1 U8270 ( .A1(n7102), .A2(n6493), .ZN(n7101) );
  NAND2_X1 U8271 ( .A1(n14957), .A2(n12573), .ZN(n14977) );
  NAND2_X1 U8272 ( .A1(n14977), .A2(n14976), .ZN(n14975) );
  XNOR2_X1 U8273 ( .A(n12574), .B(n12599), .ZN(n14994) );
  OR2_X1 U8274 ( .A1(n7100), .A2(n7098), .ZN(n6809) );
  OR2_X1 U8275 ( .A1(n15010), .A2(n15009), .ZN(n6796) );
  XNOR2_X1 U8276 ( .A(n12579), .B(n14299), .ZN(n14304) );
  NAND2_X1 U8277 ( .A1(n14304), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U8278 ( .A1(n6849), .A2(n6847), .ZN(n14336) );
  NAND2_X1 U8279 ( .A1(n14307), .A2(n6512), .ZN(n6849) );
  AOI21_X1 U8280 ( .B1(n12608), .B2(n6623), .A(n6848), .ZN(n6847) );
  OAI211_X1 U8281 ( .C1(n14325), .C2(n6799), .A(n6798), .B(n6797), .ZN(n14339)
         );
  NAND2_X1 U8282 ( .A1(n6800), .A2(n12612), .ZN(n6799) );
  AOI21_X1 U8283 ( .B1(n6801), .B2(n14324), .A(n6803), .ZN(n6798) );
  NAND2_X1 U8284 ( .A1(n14332), .A2(n12583), .ZN(n14348) );
  INV_X1 U8285 ( .A(n12581), .ZN(n12582) );
  AOI21_X1 U8286 ( .B1(n6990), .B2(n6988), .A(n12378), .ZN(n6987) );
  INV_X1 U8287 ( .A(n6992), .ZN(n6988) );
  INV_X1 U8288 ( .A(n6990), .ZN(n6989) );
  NAND2_X1 U8289 ( .A1(n6986), .A2(n6990), .ZN(n9527) );
  NAND2_X1 U8290 ( .A1(n9524), .A2(n6992), .ZN(n6986) );
  INV_X1 U8291 ( .A(n12535), .ZN(n12670) );
  AND2_X1 U8292 ( .A1(n12395), .A2(n12537), .ZN(n7005) );
  AND2_X1 U8293 ( .A1(n12496), .A2(n12495), .ZN(n12697) );
  INV_X1 U8294 ( .A(n6515), .ZN(n7067) );
  AOI21_X1 U8295 ( .B1(n6515), .B2(n7066), .A(n7065), .ZN(n7064) );
  INV_X1 U8296 ( .A(n12474), .ZN(n7065) );
  AND2_X1 U8297 ( .A1(n12464), .A2(n12779), .ZN(n12802) );
  OR2_X1 U8298 ( .A1(n14369), .A2(n12542), .ZN(n12819) );
  NAND2_X1 U8299 ( .A1(n11498), .A2(n6982), .ZN(n7090) );
  OR2_X1 U8300 ( .A1(n9251), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9268) );
  AOI21_X1 U8301 ( .B1(n6999), .B2(n7002), .A(n6531), .ZN(n6996) );
  AOI21_X1 U8302 ( .B1(n7061), .B2(n7063), .A(n7059), .ZN(n7058) );
  INV_X1 U8303 ( .A(n12438), .ZN(n7059) );
  NAND2_X1 U8304 ( .A1(n10994), .A2(n12432), .ZN(n11175) );
  NOR2_X1 U8305 ( .A1(n7447), .A2(n9505), .ZN(n9506) );
  NAND2_X1 U8306 ( .A1(n10995), .A2(n12358), .ZN(n10994) );
  XNOR2_X1 U8307 ( .A(n12550), .B(n10971), .ZN(n12364) );
  INV_X1 U8308 ( .A(n12364), .ZN(n12423) );
  INV_X1 U8309 ( .A(n12553), .ZN(n15039) );
  NAND2_X1 U8310 ( .A1(n6494), .A2(n15085), .ZN(n7013) );
  NAND2_X1 U8311 ( .A1(n9450), .A2(n9449), .ZN(n12501) );
  NAND2_X1 U8312 ( .A1(n9439), .A2(n9438), .ZN(n9664) );
  NAND2_X1 U8313 ( .A1(n9416), .A2(n9415), .ZN(n9653) );
  NAND2_X1 U8314 ( .A1(n9385), .A2(n9384), .ZN(n12215) );
  NAND2_X1 U8315 ( .A1(n9335), .A2(n9334), .ZN(n12470) );
  OR2_X1 U8316 ( .A1(n12683), .A2(n15072), .ZN(n15054) );
  INV_X1 U8317 ( .A(n12335), .ZN(n7264) );
  AOI21_X1 U8318 ( .B1(n7269), .B2(n7267), .A(n7266), .ZN(n7265) );
  NOR2_X1 U8319 ( .A1(n12332), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U8320 ( .A1(n7265), .A2(n7261), .ZN(n7260) );
  NAND2_X1 U8321 ( .A1(n7262), .A2(n7264), .ZN(n7261) );
  INV_X1 U8322 ( .A(n7267), .ZN(n7262) );
  INV_X1 U8323 ( .A(n12186), .ZN(n7269) );
  NAND2_X1 U8324 ( .A1(n9003), .A2(n9002), .ZN(n9437) );
  XNOR2_X1 U8325 ( .A(n9081), .B(n9080), .ZN(n10040) );
  OAI21_X1 U8326 ( .B1(n6519), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U8327 ( .A1(n7254), .A2(n7252), .ZN(n9378) );
  AOI21_X1 U8328 ( .B1(n7255), .B2(n7257), .A(n7253), .ZN(n7252) );
  NAND2_X1 U8329 ( .A1(n9343), .A2(n7255), .ZN(n7254) );
  INV_X1 U8330 ( .A(n8991), .ZN(n7253) );
  AND2_X1 U8331 ( .A1(n8993), .A2(n8992), .ZN(n9377) );
  NAND2_X1 U8332 ( .A1(n9378), .A2(n9377), .ZN(n9380) );
  INV_X1 U8333 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9347) );
  AND2_X1 U8334 ( .A1(n8986), .A2(n8985), .ZN(n9325) );
  NAND2_X1 U8335 ( .A1(n9326), .A2(n9325), .ZN(n9328) );
  INV_X1 U8336 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9312) );
  OAI21_X1 U8337 ( .B1(n9293), .B2(n8981), .A(n8982), .ZN(n9308) );
  AND2_X1 U8338 ( .A1(n10388), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8981) );
  AOI21_X1 U8339 ( .B1(n7249), .B2(n7251), .A(n6613), .ZN(n7247) );
  INV_X1 U8340 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9215) );
  OR2_X1 U8341 ( .A1(n9214), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9217) );
  OR2_X1 U8342 ( .A1(n9217), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9244) );
  INV_X1 U8343 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U8344 ( .A1(n8957), .A2(n8956), .ZN(n9159) );
  NOR2_X1 U8345 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n6747) );
  NOR2_X1 U8346 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n6745) );
  NAND2_X1 U8347 ( .A1(n8950), .A2(n8949), .ZN(n9131) );
  INV_X1 U8348 ( .A(n7328), .ZN(n7327) );
  OAI22_X1 U8349 ( .A1(n12969), .A2(n7329), .B1(n12007), .B2(n12008), .ZN(
        n7328) );
  NAND2_X2 U8350 ( .A1(n10023), .A2(n10022), .ZN(n12009) );
  NAND2_X1 U8351 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  INV_X1 U8352 ( .A(n13023), .ZN(n7337) );
  NAND2_X1 U8353 ( .A1(n13014), .A2(n13013), .ZN(n13025) );
  NOR2_X1 U8354 ( .A1(n8478), .A2(n8477), .ZN(n8488) );
  INV_X1 U8355 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11108) );
  OR2_X1 U8356 ( .A1(n8332), .A2(n8331), .ZN(n8350) );
  INV_X1 U8357 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11442) );
  INV_X1 U8358 ( .A(n8468), .ZN(n8469) );
  NAND2_X1 U8359 ( .A1(n8469), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8478) );
  INV_X1 U8360 ( .A(n7318), .ZN(n7317) );
  AOI21_X1 U8361 ( .B1(n7318), .B2(n7316), .A(n6578), .ZN(n7315) );
  NOR2_X1 U8362 ( .A1(n12995), .A2(n11980), .ZN(n7318) );
  XNOR2_X1 U8363 ( .A(n10246), .B(n12009), .ZN(n10153) );
  NAND2_X1 U8364 ( .A1(n13014), .A2(n6535), .ZN(n7335) );
  AND4_X1 U8365 ( .A1(n8530), .A2(n8529), .A3(n8528), .A4(n8527), .ZN(n13077)
         );
  INV_X1 U8366 ( .A(n8615), .ZN(n8845) );
  INV_X1 U8367 ( .A(n6655), .ZN(n8520) );
  NAND2_X1 U8368 ( .A1(n8614), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6812) );
  AOI21_X1 U8369 ( .B1(n9863), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9994), .ZN(
        n14683) );
  AOI21_X1 U8370 ( .B1(n9880), .B2(P2_REG2_REG_3__SCAN_IN), .A(n14681), .ZN(
        n10096) );
  AOI21_X1 U8371 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10293), .A(n10292), .ZN(
        n10295) );
  CLKBUF_X1 U8372 ( .A(P2_IR_REG_14__SCAN_IN), .Z(n8369) );
  INV_X1 U8373 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U8374 ( .A1(n13185), .A2(n14740), .ZN(n6696) );
  INV_X1 U8375 ( .A(n8923), .ZN(n8608) );
  AOI21_X1 U8376 ( .B1(n6830), .B2(n6834), .A(n6507), .ZN(n6829) );
  INV_X1 U8377 ( .A(n6941), .ZN(n6939) );
  NAND2_X1 U8378 ( .A1(n13248), .A2(n13502), .ZN(n13230) );
  XNOR2_X1 U8379 ( .A(n13010), .B(n13079), .ZN(n13279) );
  AOI21_X1 U8380 ( .B1(n13340), .B2(n13339), .A(n8463), .ZN(n13322) );
  AND2_X1 U8381 ( .A1(n6498), .A2(n6936), .ZN(n6935) );
  NAND2_X1 U8382 ( .A1(n11619), .A2(n14424), .ZN(n11620) );
  NOR2_X1 U8383 ( .A1(n7311), .A2(n8911), .ZN(n7309) );
  OR2_X1 U8384 ( .A1(n11382), .A2(n11431), .ZN(n14411) );
  NAND2_X1 U8385 ( .A1(n6934), .A2(n7308), .ZN(n11382) );
  NAND2_X1 U8386 ( .A1(n7307), .A2(n8576), .ZN(n11216) );
  NAND2_X1 U8387 ( .A1(n11240), .A2(n11245), .ZN(n7307) );
  INV_X1 U8388 ( .A(n6934), .ZN(n11246) );
  INV_X1 U8389 ( .A(n10263), .ZN(n14410) );
  NOR2_X1 U8390 ( .A1(n6539), .A2(n7287), .ZN(n7286) );
  INV_X1 U8391 ( .A(n8901), .ZN(n7287) );
  NAND2_X1 U8392 ( .A1(n10978), .A2(n10980), .ZN(n10979) );
  NAND2_X1 U8393 ( .A1(n7289), .A2(n8567), .ZN(n10856) );
  NAND2_X1 U8394 ( .A1(n10671), .A2(n7128), .ZN(n7289) );
  NAND2_X1 U8395 ( .A1(n10849), .A2(n14813), .ZN(n10985) );
  AND2_X1 U8396 ( .A1(n10666), .A2(n10669), .ZN(n10849) );
  NOR2_X1 U8397 ( .A1(n10523), .A2(n14796), .ZN(n10666) );
  NAND2_X1 U8398 ( .A1(n6932), .A2(n6931), .ZN(n10523) );
  INV_X1 U8399 ( .A(n8920), .ZN(n13233) );
  OR3_X1 U8400 ( .A1(n13281), .A2(n13280), .A3(n13295), .ZN(n13435) );
  NAND2_X1 U8401 ( .A1(n8441), .A2(n8440), .ZN(n13465) );
  NAND2_X1 U8402 ( .A1(n7127), .A2(n8235), .ZN(n10665) );
  INV_X1 U8403 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8153) );
  AND2_X1 U8404 ( .A1(n8210), .A2(n8219), .ZN(n9881) );
  INV_X1 U8405 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8117) );
  INV_X1 U8406 ( .A(n7902), .ZN(n7903) );
  OR2_X1 U8407 ( .A1(n7639), .A2(n11354), .ZN(n7659) );
  INV_X1 U8408 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7658) );
  AND2_X1 U8409 ( .A1(n13563), .A2(n7176), .ZN(n7175) );
  OR2_X1 U8410 ( .A1(n13678), .A2(n12146), .ZN(n7176) );
  OR2_X1 U8411 ( .A1(n7759), .A2(n13691), .ZN(n7784) );
  INV_X1 U8412 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7783) );
  NOR2_X1 U8413 ( .A1(n7784), .A2(n7783), .ZN(n7803) );
  NAND2_X1 U8414 ( .A1(n13574), .A2(n13626), .ZN(n7155) );
  NAND2_X1 U8415 ( .A1(n10574), .A2(n10575), .ZN(n7186) );
  OR2_X1 U8416 ( .A1(n7698), .A2(n7697), .ZN(n7717) );
  NOR2_X1 U8417 ( .A1(n7717), .A2(n13649), .ZN(n7731) );
  INV_X1 U8418 ( .A(n7889), .ZN(n7890) );
  AND2_X1 U8419 ( .A1(n7803), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7821) );
  AND2_X1 U8420 ( .A1(n7171), .A2(n13617), .ZN(n7170) );
  NAND2_X1 U8421 ( .A1(n13616), .A2(n7172), .ZN(n7171) );
  AND3_X1 U8422 ( .A1(n11857), .A2(n11856), .A3(n11855), .ZN(n11877) );
  NAND2_X1 U8423 ( .A1(n7538), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7499) );
  OR2_X1 U8424 ( .A1(n7540), .A2(n10557), .ZN(n7470) );
  AND2_X1 U8425 ( .A1(n7491), .A2(n7490), .ZN(n7494) );
  OR2_X1 U8426 ( .A1(n7540), .A2(n7489), .ZN(n7490) );
  INV_X1 U8427 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n13649) );
  NOR2_X1 U8428 ( .A1(n14075), .A2(n13887), .ZN(n7978) );
  NOR2_X1 U8429 ( .A1(n6505), .A2(n7046), .ZN(n13900) );
  AND2_X1 U8430 ( .A1(n6732), .A2(n6731), .ZN(n6730) );
  INV_X1 U8431 ( .A(n11917), .ZN(n13883) );
  NAND2_X1 U8432 ( .A1(n13987), .A2(n6899), .ZN(n13925) );
  NOR2_X1 U8433 ( .A1(n6900), .A2(n13928), .ZN(n6899) );
  INV_X1 U8434 ( .A(n6901), .ZN(n6900) );
  NAND2_X1 U8435 ( .A1(n13937), .A2(n8092), .ZN(n13919) );
  NAND2_X1 U8436 ( .A1(n13939), .A2(n13938), .ZN(n13937) );
  NAND2_X1 U8437 ( .A1(n13987), .A2(n6901), .ZN(n13942) );
  INV_X1 U8438 ( .A(n7873), .ZN(n7874) );
  AND2_X1 U8439 ( .A1(n7871), .A2(n7870), .ZN(n13971) );
  NAND2_X1 U8440 ( .A1(n14004), .A2(n7197), .ZN(n13982) );
  AND2_X1 U8441 ( .A1(n7821), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7839) );
  INV_X1 U8442 ( .A(n7232), .ZN(n7231) );
  AOI21_X1 U8443 ( .B1(n7232), .B2(n7235), .A(n7230), .ZN(n7229) );
  NOR2_X1 U8444 ( .A1(n11800), .A2(n7233), .ZN(n7232) );
  NAND2_X1 U8445 ( .A1(n6891), .A2(n6890), .ZN(n14031) );
  NAND2_X1 U8446 ( .A1(n11334), .A2(n11906), .ZN(n7042) );
  NAND3_X1 U8447 ( .A1(n13655), .A2(n6491), .A3(n11082), .ZN(n11457) );
  AND2_X1 U8448 ( .A1(n7031), .A2(n6549), .ZN(n7030) );
  NAND2_X1 U8449 ( .A1(n6581), .A2(n8074), .ZN(n6712) );
  NAND2_X1 U8450 ( .A1(n11082), .A2(n14635), .ZN(n11294) );
  NAND2_X1 U8451 ( .A1(n11082), .A2(n6897), .ZN(n11326) );
  NOR2_X1 U8452 ( .A1(n7659), .A2(n7658), .ZN(n7680) );
  NAND2_X1 U8453 ( .A1(n6719), .A2(n6720), .ZN(n6715) );
  INV_X1 U8454 ( .A(n7033), .ZN(n6719) );
  NAND2_X1 U8455 ( .A1(n6718), .A2(n6720), .ZN(n6716) );
  NOR2_X1 U8456 ( .A1(n10642), .A2(n11725), .ZN(n11038) );
  NAND2_X1 U8457 ( .A1(n10535), .A2(n8065), .ZN(n10648) );
  NAND2_X1 U8458 ( .A1(n7051), .A2(n8063), .ZN(n10533) );
  NAND2_X1 U8459 ( .A1(n7049), .A2(n7051), .ZN(n10535) );
  NOR2_X1 U8460 ( .A1(n11895), .A2(n7050), .ZN(n7049) );
  INV_X1 U8461 ( .A(n8063), .ZN(n7050) );
  AND4_X1 U8462 ( .A1(n7545), .A2(n7544), .A3(n7543), .A4(n7542), .ZN(n11714)
         );
  NAND2_X1 U8463 ( .A1(n10352), .A2(n11686), .ZN(n10393) );
  INV_X1 U8464 ( .A(n11892), .ZN(n10356) );
  NOR2_X1 U8465 ( .A1(n10560), .A2(n7516), .ZN(n10353) );
  OAI22_X1 U8466 ( .A1(n8059), .A2(n11890), .B1(n14590), .B2(n13722), .ZN(
        n10135) );
  INV_X1 U8467 ( .A(n9760), .ZN(n6710) );
  INV_X1 U8468 ( .A(n11700), .ZN(n6661) );
  AND2_X1 U8469 ( .A1(n14065), .A2(n14124), .ZN(n6892) );
  NAND2_X1 U8470 ( .A1(n10127), .A2(n9937), .ZN(n14124) );
  INV_X1 U8471 ( .A(n14124), .ZN(n14634) );
  XNOR2_X1 U8472 ( .A(n8863), .B(n8862), .ZN(n11953) );
  XNOR2_X1 U8473 ( .A(n8830), .B(n8829), .ZN(n13539) );
  INV_X1 U8474 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7473) );
  XNOR2_X1 U8475 ( .A(n7948), .B(n7947), .ZN(n13554) );
  AND2_X1 U8476 ( .A1(n7727), .A2(n7714), .ZN(n10587) );
  NAND2_X1 U8477 ( .A1(n7707), .A2(n7706), .ZN(n7726) );
  OR2_X1 U8478 ( .A1(n7693), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7694) );
  XNOR2_X1 U8479 ( .A(n7689), .B(n7688), .ZN(n9964) );
  OR2_X1 U8480 ( .A1(n7554), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7573) );
  CLKBUF_X1 U8481 ( .A(n7505), .Z(n7506) );
  OAI211_X1 U8482 ( .C1(n7887), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n6635), .B(
        SI_0_), .ZN(n7510) );
  NAND2_X1 U8483 ( .A1(n7887), .A2(n6636), .ZN(n6635) );
  CLKBUF_X1 U8484 ( .A(n7483), .Z(n7484) );
  AND2_X1 U8485 ( .A1(n6915), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14218) );
  INV_X1 U8486 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6915) );
  XNOR2_X1 U8487 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14215) );
  XNOR2_X1 U8488 ( .A(n14175), .B(n6923), .ZN(n14223) );
  INV_X1 U8489 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8490 ( .A1(n14232), .A2(n14233), .ZN(n14234) );
  NAND2_X1 U8491 ( .A1(n14182), .A2(n14181), .ZN(n14236) );
  OR2_X1 U8492 ( .A1(n14229), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n14181) );
  OAI21_X1 U8493 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14189), .A(n14188), .ZN(
        n14212) );
  NAND2_X1 U8494 ( .A1(n14194), .A2(n14193), .ZN(n14208) );
  NAND2_X1 U8495 ( .A1(n12312), .A2(n12174), .ZN(n9678) );
  INV_X1 U8496 ( .A(n7384), .ZN(n7383) );
  NAND2_X1 U8497 ( .A1(n7385), .A2(n12264), .ZN(n12206) );
  NAND2_X1 U8498 ( .A1(n11364), .A2(n9615), .ZN(n11575) );
  AND2_X1 U8499 ( .A1(n9646), .A2(n9636), .ZN(n7389) );
  NAND2_X1 U8500 ( .A1(n6580), .A2(n7387), .ZN(n7386) );
  NAND2_X1 U8501 ( .A1(n9646), .A2(n7388), .ZN(n7387) );
  AOI21_X1 U8502 ( .B1(n12312), .B2(n12177), .A(n6496), .ZN(n12179) );
  NAND2_X1 U8503 ( .A1(n7376), .A2(n7437), .ZN(n12222) );
  AND4_X1 U8504 ( .A1(n9446), .A2(n9445), .A3(n9444), .A4(n9443), .ZN(n12708)
         );
  AOI21_X1 U8505 ( .B1(n12240), .B2(n12242), .A(n12241), .ZN(n12244) );
  NAND2_X1 U8506 ( .A1(n7390), .A2(n9636), .ZN(n12251) );
  AND2_X1 U8507 ( .A1(n12526), .A2(n9698), .ZN(n14865) );
  NAND2_X1 U8508 ( .A1(n12251), .A2(n9638), .ZN(n12259) );
  NAND2_X1 U8509 ( .A1(n10740), .A2(n9599), .ZN(n10611) );
  NAND2_X1 U8510 ( .A1(n9686), .A2(n15032), .ZN(n14847) );
  OAI21_X1 U8511 ( .B1(n12240), .B2(n12241), .A(n6639), .ZN(n6638) );
  AND2_X1 U8512 ( .A1(n6640), .A2(n7380), .ZN(n6639) );
  INV_X1 U8513 ( .A(n12313), .ZN(n6640) );
  INV_X1 U8514 ( .A(n12310), .ZN(n14857) );
  OAI211_X1 U8515 ( .C1(n6570), .C2(n7096), .A(n7094), .B(n7270), .ZN(n12525)
         );
  NAND2_X1 U8516 ( .A1(n6528), .A2(n6784), .ZN(n7096) );
  NAND2_X1 U8517 ( .A1(n6570), .A2(n7095), .ZN(n7094) );
  NAND2_X1 U8518 ( .A1(n12523), .A2(n15034), .ZN(n6660) );
  INV_X1 U8519 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14876) );
  OR2_X1 U8520 ( .A1(n10165), .A2(n10046), .ZN(n10167) );
  OAI21_X1 U8521 ( .B1(n10175), .B2(n10054), .A(n10053), .ZN(n14882) );
  AND2_X1 U8522 ( .A1(n14877), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14878) );
  NOR2_X1 U8523 ( .A1(n14878), .A2(n6804), .ZN(n14898) );
  AND2_X1 U8524 ( .A1(n6805), .A2(n14889), .ZN(n6804) );
  NOR2_X1 U8525 ( .A1(n10449), .A2(n7112), .ZN(n14917) );
  AND2_X1 U8526 ( .A1(n10620), .A2(n10624), .ZN(n6845) );
  XNOR2_X1 U8527 ( .A(n10749), .B(n10762), .ZN(n10625) );
  INV_X1 U8528 ( .A(n6885), .ZN(n11185) );
  INV_X1 U8529 ( .A(n6887), .ZN(n10752) );
  NAND2_X1 U8530 ( .A1(n14942), .A2(n11188), .ZN(n11191) );
  NAND2_X1 U8531 ( .A1(n11191), .A2(n11190), .ZN(n12571) );
  INV_X1 U8532 ( .A(n7102), .ZN(n14955) );
  AND2_X1 U8533 ( .A1(n7101), .A2(n7100), .ZN(n14972) );
  INV_X1 U8534 ( .A(n7101), .ZN(n14974) );
  NOR2_X1 U8535 ( .A1(n14965), .A2(n6844), .ZN(n14986) );
  AND2_X1 U8536 ( .A1(n12592), .A2(n12593), .ZN(n6844) );
  NAND2_X1 U8537 ( .A1(n14986), .A2(n14985), .ZN(n14984) );
  INV_X1 U8538 ( .A(n6796), .ZN(n15008) );
  NOR2_X1 U8539 ( .A1(n15000), .A2(n6842), .ZN(n15025) );
  AND2_X1 U8540 ( .A1(n12598), .A2(n12599), .ZN(n6842) );
  NAND2_X1 U8541 ( .A1(n15025), .A2(n15024), .ZN(n15023) );
  NOR2_X1 U8542 ( .A1(n14305), .A2(n12608), .ZN(n14318) );
  INV_X1 U8543 ( .A(n7105), .ZN(n14357) );
  NOR2_X1 U8544 ( .A1(n14346), .A2(n12770), .ZN(n7103) );
  NAND2_X1 U8545 ( .A1(n7079), .A2(n7080), .ZN(n12659) );
  NAND2_X1 U8546 ( .A1(n12680), .A2(n6520), .ZN(n12665) );
  NAND2_X1 U8547 ( .A1(n7086), .A2(n12491), .ZN(n12715) );
  OR2_X1 U8548 ( .A1(n7089), .A2(n7088), .ZN(n7086) );
  INV_X1 U8549 ( .A(n12487), .ZN(n7087) );
  AND2_X1 U8550 ( .A1(n12746), .A2(n12745), .ZN(n12877) );
  NAND2_X1 U8551 ( .A1(n7070), .A2(n7068), .ZN(n12774) );
  NOR2_X1 U8552 ( .A1(n7009), .A2(n7008), .ZN(n12765) );
  INV_X1 U8553 ( .A(n9519), .ZN(n7008) );
  NAND2_X1 U8554 ( .A1(n9316), .A2(n9315), .ZN(n14364) );
  AOI21_X1 U8555 ( .B1(n9774), .B2(n12338), .A(n9284), .ZN(n14376) );
  NAND2_X1 U8556 ( .A1(n11492), .A2(n12367), .ZN(n6979) );
  NAND2_X1 U8557 ( .A1(n6998), .A2(n9511), .ZN(n11252) );
  NAND2_X1 U8558 ( .A1(n11275), .A2(n11276), .ZN(n6998) );
  INV_X1 U8559 ( .A(n15032), .ZN(n12805) );
  AND2_X1 U8560 ( .A1(n9044), .A2(n10515), .ZN(n15034) );
  INV_X1 U8561 ( .A(n7013), .ZN(n7012) );
  INV_X1 U8562 ( .A(n9676), .ZN(n12911) );
  INV_X1 U8563 ( .A(n12506), .ZN(n12915) );
  INV_X1 U8564 ( .A(n12501), .ZN(n12919) );
  INV_X1 U8565 ( .A(n9664), .ZN(n12923) );
  INV_X1 U8566 ( .A(n12486), .ZN(n12939) );
  NAND2_X1 U8567 ( .A1(n9351), .A2(n9350), .ZN(n12948) );
  INV_X1 U8568 ( .A(n12470), .ZN(n12953) );
  AND2_X1 U8569 ( .A1(n9059), .A2(n9058), .ZN(n12954) );
  INV_X1 U8570 ( .A(n9585), .ZN(n12956) );
  AND2_X1 U8571 ( .A1(n10040), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12955) );
  OAI21_X1 U8572 ( .B1(n7265), .B2(n12335), .A(n7260), .ZN(n7259) );
  NAND2_X1 U8573 ( .A1(n7265), .A2(n7264), .ZN(n7263) );
  OAI21_X1 U8574 ( .B1(n12187), .B2(n7269), .A(n12188), .ZN(n12334) );
  NOR2_X1 U8575 ( .A1(n7093), .A2(n9093), .ZN(n7092) );
  NOR2_X1 U8576 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n7093) );
  OAI21_X1 U8577 ( .B1(n9461), .B2(n9007), .A(n9008), .ZN(n9472) );
  INV_X1 U8578 ( .A(SI_25_), .ZN(n15221) );
  NAND2_X1 U8579 ( .A1(n9046), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9047) );
  OAI21_X1 U8580 ( .B1(n9414), .B2(n9413), .A(n9000), .ZN(n9424) );
  XNOR2_X1 U8581 ( .A(n9040), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12529) );
  INV_X1 U8582 ( .A(SI_20_), .ZN(n10513) );
  INV_X1 U8583 ( .A(SI_19_), .ZN(n15160) );
  NAND2_X1 U8584 ( .A1(n9345), .A2(n8988), .ZN(n9361) );
  INV_X1 U8585 ( .A(SI_16_), .ZN(n15194) );
  INV_X1 U8586 ( .A(SI_15_), .ZN(n9915) );
  INV_X1 U8587 ( .A(SI_14_), .ZN(n15127) );
  INV_X1 U8588 ( .A(SI_12_), .ZN(n15176) );
  INV_X1 U8589 ( .A(SI_11_), .ZN(n15213) );
  NAND2_X1 U8590 ( .A1(n9243), .A2(n8973), .ZN(n9260) );
  INV_X1 U8591 ( .A(SI_10_), .ZN(n9754) );
  XNOR2_X1 U8592 ( .A(n9248), .B(n9247), .ZN(n12557) );
  NAND2_X1 U8593 ( .A1(n9194), .A2(n8966), .ZN(n9211) );
  NAND2_X1 U8594 ( .A1(n8964), .A2(n8963), .ZN(n9192) );
  NAND2_X1 U8595 ( .A1(n9112), .A2(n7109), .ZN(n10182) );
  OAI21_X1 U8596 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        n7111), .ZN(n7110) );
  AND2_X1 U8597 ( .A1(n11559), .A2(n11558), .ZN(n11561) );
  NAND2_X1 U8598 ( .A1(n8476), .A2(n8475), .ZN(n13313) );
  NAND2_X1 U8599 ( .A1(n10205), .A2(n10204), .ZN(n10369) );
  NAND2_X1 U8600 ( .A1(n13061), .A2(n6677), .ZN(n12990) );
  NAND2_X1 U8601 ( .A1(n11973), .A2(n6678), .ZN(n6677) );
  INV_X1 U8602 ( .A(n11974), .ZN(n6678) );
  NAND2_X1 U8603 ( .A1(n8426), .A2(n8425), .ZN(n13383) );
  NOR2_X1 U8604 ( .A1(n7330), .A2(n7326), .ZN(n7321) );
  OAI21_X1 U8605 ( .B1(n7327), .B2(n12012), .A(n7323), .ZN(n7322) );
  NAND2_X1 U8606 ( .A1(n7327), .A2(n7324), .ZN(n7323) );
  NAND2_X1 U8607 ( .A1(n7330), .A2(n7326), .ZN(n7324) );
  NAND2_X1 U8608 ( .A1(n7327), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U8609 ( .A1(n13042), .A2(n11981), .ZN(n12996) );
  INV_X1 U8610 ( .A(n7345), .ZN(n7344) );
  INV_X1 U8611 ( .A(n11412), .ZN(n7346) );
  NAND2_X1 U8612 ( .A1(n7333), .A2(n7336), .ZN(n13027) );
  NAND2_X1 U8613 ( .A1(n8487), .A2(n8486), .ZN(n13441) );
  NAND2_X1 U8614 ( .A1(n7332), .A2(n11102), .ZN(n11105) );
  INV_X1 U8615 ( .A(n10034), .ZN(n8554) );
  AND2_X1 U8617 ( .A1(n6650), .A2(n11261), .ZN(n11265) );
  AND2_X1 U8618 ( .A1(n9960), .A2(n9948), .ZN(n13085) );
  NAND2_X1 U8619 ( .A1(n7335), .A2(n7334), .ZN(n13061) );
  AND2_X1 U8620 ( .A1(n13062), .A2(n6501), .ZN(n7334) );
  AND2_X1 U8621 ( .A1(n7333), .A2(n6501), .ZN(n13063) );
  INV_X1 U8622 ( .A(n13091), .ZN(n13060) );
  NAND2_X1 U8623 ( .A1(n10206), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13087) );
  INV_X1 U8624 ( .A(n13078), .ZN(n13064) );
  INV_X1 U8625 ( .A(n13077), .ZN(n13102) );
  NAND2_X1 U8626 ( .A1(n14666), .A2(n6548), .ZN(n14665) );
  OAI21_X1 U8627 ( .B1(n10084), .B2(n9917), .A(n9916), .ZN(n9919) );
  OAI211_X1 U8628 ( .C1(n14726), .C2(n13162), .A(n13161), .B(n13160), .ZN(
        n13183) );
  NOR2_X1 U8629 ( .A1(n13202), .A2(n13295), .ZN(n13412) );
  INV_X1 U8630 ( .A(n6634), .ZN(n13420) );
  AND2_X1 U8631 ( .A1(n8519), .A2(n8518), .ZN(n13252) );
  NAND2_X1 U8632 ( .A1(n6837), .A2(n8606), .ZN(n13244) );
  NAND2_X1 U8633 ( .A1(n13278), .A2(n8506), .ZN(n13264) );
  NAND2_X1 U8634 ( .A1(n6825), .A2(n6826), .ZN(n13307) );
  NAND2_X1 U8635 ( .A1(n13341), .A2(n7313), .ZN(n13326) );
  NAND2_X1 U8636 ( .A1(n13341), .A2(n8599), .ZN(n13324) );
  NAND2_X1 U8637 ( .A1(n7283), .A2(n8591), .ZN(n13376) );
  AND2_X1 U8638 ( .A1(n8385), .A2(n8911), .ZN(n7147) );
  NAND2_X1 U8639 ( .A1(n11611), .A2(n8385), .ZN(n11607) );
  NAND2_X1 U8640 ( .A1(n8582), .A2(n8581), .ZN(n11614) );
  NAND2_X1 U8641 ( .A1(n7136), .A2(n8356), .ZN(n14407) );
  OAI21_X1 U8642 ( .B1(n11240), .B2(n7305), .A(n7302), .ZN(n11375) );
  NAND2_X1 U8643 ( .A1(n8341), .A2(n8340), .ZN(n11380) );
  NAND2_X1 U8644 ( .A1(n7117), .A2(n8293), .ZN(n11007) );
  NAND2_X1 U8645 ( .A1(n10883), .A2(n10884), .ZN(n7117) );
  NAND2_X1 U8646 ( .A1(n6813), .A2(n8563), .ZN(n10518) );
  OR2_X1 U8647 ( .A1(n7293), .A2(n7291), .ZN(n6813) );
  NAND2_X1 U8648 ( .A1(n10243), .A2(n8179), .ZN(n10262) );
  OR2_X1 U8649 ( .A1(n14420), .A2(n10482), .ZN(n13406) );
  INV_X1 U8650 ( .A(n13372), .ZN(n14417) );
  NAND2_X1 U8651 ( .A1(n8665), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6701) );
  INV_X1 U8652 ( .A(n8883), .ZN(n13496) );
  AND2_X1 U8653 ( .A1(n8508), .A2(n8507), .ZN(n13507) );
  INV_X1 U8654 ( .A(n13313), .ZN(n13519) );
  INV_X1 U8655 ( .A(n13383), .ZN(n13532) );
  AND2_X1 U8656 ( .A1(n9951), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14791) );
  CLKBUF_X1 U8657 ( .A(n14769), .Z(n14786) );
  INV_X1 U8658 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6676) );
  OAI21_X2 U8659 ( .B1(n8639), .B2(n7362), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7148) );
  XNOR2_X1 U8660 ( .A(n8643), .B(n7365), .ZN(n13553) );
  INV_X1 U8661 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13556) );
  NAND2_X1 U8662 ( .A1(n8636), .A2(n8637), .ZN(n13558) );
  INV_X1 U8663 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11076) );
  OAI21_X1 U8664 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n8141) );
  NAND2_X1 U8665 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8137), .ZN(n8136) );
  INV_X1 U8666 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11024) );
  INV_X1 U8667 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10423) );
  INV_X1 U8668 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10385) );
  INV_X1 U8669 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10471) );
  INV_X1 U8670 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10214) );
  INV_X1 U8671 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10039) );
  INV_X1 U8672 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9965) );
  INV_X1 U8673 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9911) );
  INV_X1 U8674 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9860) );
  INV_X1 U8675 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9778) );
  INV_X1 U8676 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9768) );
  INV_X1 U8677 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9752) );
  INV_X1 U8678 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9727) );
  INV_X1 U8679 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9723) );
  INV_X1 U8680 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9725) );
  MUX2_X1 U8681 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8174), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8177) );
  INV_X1 U8682 ( .A(n11734), .ZN(n14622) );
  INV_X1 U8683 ( .A(n13718), .ZN(n11062) );
  NOR2_X1 U8684 ( .A1(n14453), .A2(n7178), .ZN(n7177) );
  INV_X1 U8685 ( .A(n12044), .ZN(n7178) );
  NAND2_X1 U8686 ( .A1(n13645), .A2(n12044), .ZN(n14454) );
  INV_X1 U8687 ( .A(n7181), .ZN(n11347) );
  NAND2_X1 U8688 ( .A1(n11162), .A2(n11161), .ZN(n11163) );
  NAND2_X1 U8689 ( .A1(n7162), .A2(n7166), .ZN(n11642) );
  NAND2_X1 U8690 ( .A1(n6682), .A2(n7167), .ZN(n7162) );
  AND2_X1 U8691 ( .A1(n13607), .A2(n7153), .ZN(n7152) );
  NAND2_X1 U8692 ( .A1(n7156), .A2(n7159), .ZN(n7153) );
  NAND2_X1 U8693 ( .A1(n12058), .A2(n13688), .ZN(n14468) );
  AND2_X1 U8694 ( .A1(n11352), .A2(n7180), .ZN(n7179) );
  INV_X1 U8695 ( .A(n7454), .ZN(n7180) );
  NOR2_X1 U8696 ( .A1(n11347), .A2(n7454), .ZN(n11353) );
  AND2_X1 U8697 ( .A1(n14482), .A2(n11633), .ZN(n14485) );
  AND2_X1 U8698 ( .A1(n10345), .A2(n11934), .ZN(n14494) );
  INV_X1 U8699 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13691) );
  CLKBUF_X1 U8700 ( .A(n13687), .Z(n13688) );
  AND2_X1 U8701 ( .A1(n11927), .A2(n11926), .ZN(n11928) );
  INV_X1 U8702 ( .A(n13657), .ZN(n13705) );
  NAND2_X1 U8703 ( .A1(n11870), .A2(n11869), .ZN(n14055) );
  INV_X1 U8704 ( .A(n11919), .ZN(n14060) );
  AND2_X1 U8705 ( .A1(n13868), .A2(n7452), .ZN(n14069) );
  INV_X1 U8706 ( .A(n6895), .ZN(n7452) );
  AOI21_X1 U8707 ( .B1(n13866), .B2(n14028), .A(n13865), .ZN(n14072) );
  NAND2_X1 U8708 ( .A1(n13864), .A2(n13863), .ZN(n13865) );
  NAND2_X1 U8709 ( .A1(n13861), .A2(n7444), .ZN(n13866) );
  AOI21_X1 U8710 ( .B1(n11944), .B2(n14028), .A(n11943), .ZN(n11945) );
  NAND2_X1 U8711 ( .A1(n13917), .A2(n7923), .ZN(n13897) );
  NAND2_X1 U8712 ( .A1(n13934), .A2(n7910), .ZN(n13915) );
  NAND2_X1 U8713 ( .A1(n6726), .A2(n7054), .ZN(n13977) );
  NAND2_X1 U8714 ( .A1(n14020), .A2(n6727), .ZN(n6726) );
  AND2_X1 U8715 ( .A1(n7853), .A2(n7852), .ZN(n13991) );
  NAND2_X1 U8716 ( .A1(n11653), .A2(n7807), .ZN(n14023) );
  NAND2_X1 U8717 ( .A1(n7792), .A2(n7791), .ZN(n11654) );
  NAND2_X1 U8718 ( .A1(n7782), .A2(n7781), .ZN(n14472) );
  NAND2_X1 U8719 ( .A1(n7213), .A2(n11784), .ZN(n11595) );
  NAND2_X2 U8720 ( .A1(n7730), .A2(n7729), .ZN(n14507) );
  NAND2_X1 U8721 ( .A1(n11336), .A2(n7724), .ZN(n11450) );
  NAND2_X1 U8722 ( .A1(n11086), .A2(n8075), .ZN(n11292) );
  OAI21_X1 U8723 ( .B1(n6703), .B2(n7222), .A(n7221), .ZN(n11298) );
  NAND2_X1 U8724 ( .A1(n7666), .A2(n11079), .ZN(n11299) );
  NAND2_X1 U8725 ( .A1(n9910), .A2(n7965), .ZN(n7657) );
  NAND2_X1 U8726 ( .A1(n14047), .A2(n8103), .ZN(n14035) );
  NAND2_X1 U8727 ( .A1(n11036), .A2(n7612), .ZN(n10729) );
  NAND2_X1 U8728 ( .A1(n10530), .A2(n7581), .ZN(n10641) );
  NAND2_X1 U8729 ( .A1(n7053), .A2(n8062), .ZN(n10398) );
  NAND2_X1 U8730 ( .A1(n8057), .A2(n9943), .ZN(n14011) );
  INV_X1 U8731 ( .A(n14035), .ZN(n14049) );
  AND2_X2 U8732 ( .A1(n10144), .A2(n10130), .ZN(n14654) );
  INV_X2 U8733 ( .A(n14639), .ZN(n14641) );
  INV_X1 U8734 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U8735 ( .A1(n6738), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6737) );
  OAI21_X1 U8736 ( .B1(n8017), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7475) );
  XNOR2_X1 U8737 ( .A(n8020), .B(n8019), .ZN(n14160) );
  INV_X1 U8738 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8024) );
  INV_X1 U8739 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11077) );
  INV_X1 U8740 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11936) );
  INV_X1 U8741 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10844) );
  INV_X1 U8742 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10384) );
  INV_X1 U8743 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10470) );
  INV_X1 U8744 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10388) );
  INV_X1 U8745 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10213) );
  INV_X1 U8746 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9912) );
  INV_X1 U8747 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9858) );
  INV_X1 U8748 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9776) );
  INV_X1 U8749 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9765) );
  INV_X1 U8750 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9750) );
  INV_X1 U8751 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9739) );
  XNOR2_X1 U8752 ( .A(n14234), .B(n6927), .ZN(n14276) );
  INV_X1 U8753 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6927) );
  AND2_X1 U8754 ( .A1(n6925), .A2(n6582), .ZN(n14278) );
  OR2_X1 U8755 ( .A1(n15294), .A2(n15295), .ZN(n6925) );
  NAND2_X1 U8756 ( .A1(n14278), .A2(n14279), .ZN(n14277) );
  NAND2_X1 U8757 ( .A1(n6924), .A2(n14277), .ZN(n14282) );
  OAI21_X1 U8758 ( .B1(n14278), .B2(n14279), .A(P2_ADDR_REG_8__SCAN_IN), .ZN(
        n6924) );
  NOR2_X1 U8759 ( .A1(n14249), .A2(n14250), .ZN(n14524) );
  OAI21_X1 U8760 ( .B1(n14538), .B2(n14539), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n6652) );
  AND2_X1 U8761 ( .A1(n14267), .A2(n14266), .ZN(n15088) );
  NAND2_X1 U8762 ( .A1(n14858), .A2(n7372), .ZN(n10831) );
  NOR2_X1 U8763 ( .A1(n14358), .A2(n7103), .ZN(n12570) );
  AND2_X1 U8764 ( .A1(n7014), .A2(n7015), .ZN(n12643) );
  OAI21_X1 U8765 ( .B1(n9580), .B2(n15074), .A(n6619), .ZN(n9581) );
  NOR2_X1 U8766 ( .A1(n9086), .A2(n9088), .ZN(n9539) );
  NAND2_X1 U8767 ( .A1(n7341), .A2(n10367), .ZN(n10377) );
  MUX2_X1 U8768 ( .A(n13198), .B(n13197), .S(n8653), .Z(n13200) );
  OAI22_X1 U8769 ( .A1(n13218), .A2(n13474), .B1(n14842), .B2(n8662), .ZN(
        n8663) );
  NAND2_X1 U8770 ( .A1(n6702), .A2(n6699), .ZN(P2_U3527) );
  INV_X1 U8771 ( .A(n6700), .ZN(n6699) );
  NAND2_X1 U8772 ( .A1(n13501), .A2(n14842), .ZN(n6702) );
  OAI21_X1 U8773 ( .B1(n13502), .B2(n13474), .A(n6701), .ZN(n6700) );
  AND2_X1 U8774 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  AOI21_X1 U8775 ( .B1(n7142), .B2(n7140), .A(n7144), .ZN(n7139) );
  AOI21_X1 U8776 ( .B1(n7146), .B2(n13485), .A(n7143), .ZN(n7142) );
  CLKBUF_X1 U8777 ( .A(n13728), .Z(P1_U4016) );
  NOR2_X1 U8778 ( .A1(n6706), .A2(n6705), .ZN(n6704) );
  INV_X1 U8779 ( .A(n13568), .ZN(n6705) );
  NAND2_X1 U8780 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  INV_X1 U8781 ( .A(n10115), .ZN(n10118) );
  INV_X1 U8782 ( .A(n8115), .ZN(n8116) );
  OAI21_X1 U8783 ( .B1(n14067), .B2(n14041), .A(n8114), .ZN(n8115) );
  INV_X1 U8784 ( .A(n6919), .ZN(n14527) );
  INV_X1 U8785 ( .A(n6916), .ZN(n14532) );
  INV_X1 U8786 ( .A(n6909), .ZN(n14295) );
  INV_X2 U8787 ( .A(n11738), .ZN(n11839) );
  INV_X2 U8788 ( .A(n11738), .ZN(n11860) );
  AND2_X1 U8789 ( .A1(n6897), .A2(n6896), .ZN(n6491) );
  INV_X1 U8790 ( .A(n12740), .ZN(n7083) );
  OR2_X1 U8792 ( .A1(n13328), .A2(n13332), .ZN(n6492) );
  OR2_X1 U8793 ( .A1(n12593), .A2(n12558), .ZN(n6493) );
  AND2_X1 U8794 ( .A1(n9577), .A2(n7015), .ZN(n6494) );
  NOR2_X1 U8795 ( .A1(n9653), .A2(n12729), .ZN(n6495) );
  NOR2_X1 U8796 ( .A1(n12173), .A2(n12176), .ZN(n6496) );
  AND2_X1 U8797 ( .A1(n6889), .A2(n6888), .ZN(n6497) );
  AND2_X1 U8798 ( .A1(n6937), .A2(n13033), .ZN(n6498) );
  AND2_X1 U8799 ( .A1(n6826), .A2(n6543), .ZN(n6499) );
  AND2_X1 U8800 ( .A1(n6785), .A2(n12504), .ZN(n6500) );
  NAND2_X1 U8801 ( .A1(n7373), .A2(n9658), .ZN(n12283) );
  AND2_X1 U8802 ( .A1(n7336), .A2(n6558), .ZN(n6501) );
  AND2_X1 U8803 ( .A1(n7413), .A2(n6865), .ZN(n6502) );
  AND2_X1 U8804 ( .A1(n7900), .A2(n7899), .ZN(n13943) );
  INV_X1 U8805 ( .A(n13943), .ZN(n6904) );
  NOR2_X1 U8806 ( .A1(n13563), .A2(n12146), .ZN(n6503) );
  AND2_X1 U8807 ( .A1(n6973), .A2(n6607), .ZN(n6504) );
  AND2_X1 U8808 ( .A1(n13937), .A2(n6732), .ZN(n6505) );
  INV_X1 U8809 ( .A(n11257), .ZN(n7000) );
  NOR2_X1 U8810 ( .A1(n7362), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n6506) );
  AND2_X1 U8811 ( .A1(n13502), .A2(n13101), .ZN(n6507) );
  AND2_X1 U8812 ( .A1(n11103), .A2(n11102), .ZN(n6508) );
  AND2_X1 U8813 ( .A1(n6493), .A2(n7099), .ZN(n6509) );
  AND2_X1 U8814 ( .A1(n7430), .A2(n7429), .ZN(n6510) );
  INV_X1 U8815 ( .A(n12367), .ZN(n6982) );
  NOR2_X1 U8816 ( .A1(n6957), .A2(n6958), .ZN(n6956) );
  NAND3_X1 U8817 ( .A1(n12440), .A2(n12448), .A3(n7001), .ZN(n6511) );
  NAND2_X1 U8818 ( .A1(n7696), .A2(n7695), .ZN(n11768) );
  INV_X1 U8819 ( .A(n11768), .ZN(n6896) );
  INV_X2 U8820 ( .A(n15074), .ZN(n15076) );
  AND2_X1 U8821 ( .A1(n6623), .A2(n14308), .ZN(n6512) );
  INV_X1 U8822 ( .A(n10413), .ZN(n6931) );
  OAI211_X2 U8823 ( .C1(n9746), .C2(n9795), .A(n7515), .B(n7514), .ZN(n7516)
         );
  AND2_X1 U8824 ( .A1(n10461), .A2(n14928), .ZN(n6514) );
  INV_X1 U8825 ( .A(n11911), .ZN(n7236) );
  AND2_X1 U8826 ( .A1(n7068), .A2(n12372), .ZN(n6515) );
  INV_X1 U8827 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12958) );
  XNOR2_X1 U8828 ( .A(n8037), .B(n8036), .ZN(n8056) );
  MUX2_X1 U8829 ( .A(n14663), .B(n13561), .S(n9868), .Z(n10247) );
  AND2_X1 U8830 ( .A1(n7667), .A2(n9754), .ZN(n6516) );
  OR2_X1 U8831 ( .A1(n13186), .A2(n14738), .ZN(n6517) );
  INV_X1 U8832 ( .A(n10672), .ZN(n7128) );
  AND2_X1 U8833 ( .A1(n7383), .A2(n12264), .ZN(n6518) );
  INV_X2 U8834 ( .A(n12148), .ZN(n12062) );
  OR2_X1 U8835 ( .A1(n9041), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6519) );
  OR2_X1 U8836 ( .A1(n12919), .A2(n12536), .ZN(n6520) );
  AND4_X1 U8837 ( .A1(n8036), .A2(n7816), .A3(n6683), .A4(n7463), .ZN(n6521)
         );
  INV_X1 U8838 ( .A(n7305), .ZN(n7304) );
  OR2_X1 U8839 ( .A1(n8577), .A2(n7306), .ZN(n7305) );
  NAND2_X1 U8840 ( .A1(n6488), .A2(n9735), .ZN(n9165) );
  NOR2_X1 U8841 ( .A1(n12472), .A2(n12779), .ZN(n6522) );
  AND2_X1 U8842 ( .A1(n13279), .A2(n8494), .ZN(n6523) );
  OR2_X1 U8843 ( .A1(n9165), .A2(n9176), .ZN(n6524) );
  NOR2_X1 U8844 ( .A1(n12396), .A2(n7085), .ZN(n6525) );
  NAND2_X1 U8845 ( .A1(n9495), .A2(n15031), .ZN(n6526) );
  MUX2_X1 U8846 ( .A(n13702), .B(n14070), .S(n11839), .Z(n11841) );
  MUX2_X1 U8847 ( .A(n14547), .B(n14170), .S(n9746), .Z(n11694) );
  INV_X1 U8848 ( .A(n13419), .ZN(n6633) );
  AND2_X1 U8849 ( .A1(n7081), .A2(n6520), .ZN(n6527) );
  INV_X1 U8850 ( .A(n7198), .ZN(n7197) );
  NAND2_X1 U8851 ( .A1(n13993), .A2(n8087), .ZN(n7198) );
  AND4_X1 U8852 ( .A1(n12387), .A2(n12398), .A3(n9044), .A4(n12519), .ZN(n6528) );
  OR2_X1 U8853 ( .A1(n15088), .A2(n15086), .ZN(n6529) );
  XNOR2_X1 U8854 ( .A(n9178), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10624) );
  INV_X1 U8855 ( .A(n13502), .ZN(n12018) );
  AND2_X1 U8856 ( .A1(n14376), .A2(n12828), .ZN(n6530) );
  XNOR2_X1 U8857 ( .A(n6737), .B(n7465), .ZN(n7468) );
  AND2_X1 U8858 ( .A1(n12545), .A2(n11316), .ZN(n6531) );
  INV_X1 U8859 ( .A(n12658), .ZN(n6991) );
  AND2_X1 U8860 ( .A1(n11794), .A2(n11911), .ZN(n6532) );
  INV_X1 U8861 ( .A(n11815), .ZN(n6879) );
  NAND2_X1 U8862 ( .A1(n9663), .A2(n9662), .ZN(n12264) );
  NOR2_X1 U8863 ( .A1(n8883), .A2(n13098), .ZN(n6533) );
  AND2_X1 U8864 ( .A1(n9735), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6534) );
  INV_X1 U8865 ( .A(n8737), .ZN(n7355) );
  INV_X1 U8866 ( .A(n11759), .ZN(n7419) );
  INV_X1 U8867 ( .A(n8772), .ZN(n7353) );
  NAND2_X1 U8868 ( .A1(n12393), .A2(n9574), .ZN(n12511) );
  AND2_X1 U8869 ( .A1(n7338), .A2(n13013), .ZN(n6535) );
  INV_X1 U8870 ( .A(n8916), .ZN(n13398) );
  NAND2_X1 U8871 ( .A1(n8373), .A2(n8372), .ZN(n13096) );
  AND2_X1 U8872 ( .A1(n7019), .A2(n7021), .ZN(n6536) );
  AND2_X1 U8873 ( .A1(n8497), .A2(n8496), .ZN(n13511) );
  INV_X1 U8874 ( .A(n13511), .ZN(n13010) );
  INV_X1 U8875 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8137) );
  AND3_X1 U8876 ( .A1(n8214), .A2(n8215), .A3(n6812), .ZN(n6537) );
  OR2_X1 U8877 ( .A1(n13096), .A2(n8583), .ZN(n6538) );
  AND2_X1 U8878 ( .A1(n14169), .A2(n9746), .ZN(n14104) );
  INV_X1 U8879 ( .A(n14104), .ZN(n13957) );
  AND2_X1 U8880 ( .A1(n7536), .A2(n7535), .ZN(n10354) );
  INV_X1 U8881 ( .A(n10354), .ZN(n6646) );
  AND2_X1 U8882 ( .A1(n8902), .A2(n7290), .ZN(n6539) );
  OR2_X1 U8883 ( .A1(n12162), .A2(n12160), .ZN(n6540) );
  OR2_X1 U8884 ( .A1(n9868), .A2(n14660), .ZN(n6541) );
  AND3_X1 U8885 ( .A1(n11781), .A2(n11776), .A3(n11778), .ZN(n6542) );
  OR2_X1 U8886 ( .A1(n13313), .A2(n11988), .ZN(n6543) );
  AND2_X1 U8887 ( .A1(n7523), .A2(n7522), .ZN(n6544) );
  AND2_X1 U8888 ( .A1(n9043), .A2(n6519), .ZN(n12398) );
  AND2_X1 U8889 ( .A1(n6523), .A2(n8517), .ZN(n6545) );
  INV_X1 U8890 ( .A(n11827), .ZN(n6866) );
  OR2_X1 U8891 ( .A1(n7509), .A2(n9712), .ZN(n6546) );
  AND2_X1 U8892 ( .A1(n7425), .A2(n7426), .ZN(n6547) );
  AND2_X1 U8893 ( .A1(n14663), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6548) );
  OR2_X1 U8894 ( .A1(n14489), .A2(n8077), .ZN(n6549) );
  AND2_X1 U8895 ( .A1(n11133), .A2(n13119), .ZN(n6550) );
  NAND2_X1 U8896 ( .A1(n10107), .A2(n12158), .ZN(n6551) );
  INV_X1 U8897 ( .A(n7235), .ZN(n7234) );
  NAND2_X1 U8898 ( .A1(n7236), .A2(n7791), .ZN(n7235) );
  AND2_X1 U8899 ( .A1(n7192), .A2(n7191), .ZN(n6552) );
  NOR2_X1 U8900 ( .A1(n14364), .A2(n12254), .ZN(n6553) );
  INV_X1 U8901 ( .A(n13212), .ZN(n13500) );
  NAND2_X1 U8902 ( .A1(n8866), .A2(n8865), .ZN(n13212) );
  AND2_X1 U8903 ( .A1(n13313), .A2(n11988), .ZN(n6554) );
  OR2_X1 U8904 ( .A1(n13328), .A2(n6929), .ZN(n6555) );
  NAND2_X1 U8905 ( .A1(n8405), .A2(n8404), .ZN(n13482) );
  NAND2_X1 U8906 ( .A1(n12826), .A2(n12460), .ZN(n6556) );
  OR2_X1 U8907 ( .A1(n10459), .A2(n10458), .ZN(n6557) );
  NAND2_X1 U8908 ( .A1(n11972), .A2(n11971), .ZN(n6558) );
  NOR2_X1 U8909 ( .A1(n11739), .A2(n13716), .ZN(n6559) );
  AND2_X1 U8910 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n6560) );
  NOR2_X1 U8911 ( .A1(n13332), .A2(n12981), .ZN(n6561) );
  AND2_X1 U8912 ( .A1(n12931), .A2(n12729), .ZN(n6562) );
  INV_X1 U8913 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6636) );
  INV_X1 U8914 ( .A(n8075), .ZN(n7032) );
  INV_X1 U8915 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U8916 ( .A1(n7461), .A2(n7460), .ZN(n6563) );
  AND2_X1 U8917 ( .A1(n12915), .A2(n12678), .ZN(n6564) );
  INV_X1 U8918 ( .A(n12522), .ZN(n6784) );
  NOR2_X1 U8919 ( .A1(n9557), .A2(n12655), .ZN(n6565) );
  NAND2_X1 U8920 ( .A1(n13507), .A2(n13005), .ZN(n6566) );
  AND2_X1 U8921 ( .A1(n11779), .A2(n11780), .ZN(n6567) );
  INV_X1 U8922 ( .A(n6903), .ZN(n6902) );
  NAND2_X1 U8923 ( .A1(n13971), .A2(n13957), .ZN(n6903) );
  INV_X1 U8924 ( .A(n7046), .ZN(n6736) );
  NAND2_X1 U8925 ( .A1(n13898), .A2(n7047), .ZN(n7046) );
  AND2_X1 U8926 ( .A1(n7597), .A2(n7595), .ZN(n6568) );
  AND2_X1 U8927 ( .A1(n7616), .A2(SI_7_), .ZN(n6569) );
  NAND2_X1 U8928 ( .A1(n7396), .A2(n9021), .ZN(n7395) );
  INV_X1 U8929 ( .A(n7395), .ZN(n7393) );
  AND2_X1 U8930 ( .A1(n12347), .A2(n12516), .ZN(n6570) );
  AND2_X1 U8931 ( .A1(n11793), .A2(n11792), .ZN(n6571) );
  AND4_X1 U8932 ( .A1(n8150), .A2(n8149), .A3(n8137), .A4(n8649), .ZN(n6572)
         );
  NAND2_X1 U8933 ( .A1(n7155), .A2(n13627), .ZN(n13606) );
  NOR2_X1 U8934 ( .A1(n11055), .A2(n11734), .ZN(n6573) );
  NAND2_X1 U8935 ( .A1(n7706), .A2(SI_13_), .ZN(n6574) );
  OR2_X1 U8936 ( .A1(n6880), .A2(n6879), .ZN(n6575) );
  INV_X1 U8937 ( .A(n7168), .ZN(n7167) );
  NAND2_X1 U8938 ( .A1(n7169), .A2(n11470), .ZN(n7168) );
  INV_X1 U8939 ( .A(n7666), .ZN(n7222) );
  AND2_X1 U8940 ( .A1(n7308), .A2(n13117), .ZN(n6576) );
  AND2_X1 U8941 ( .A1(n12474), .A2(n12477), .ZN(n12372) );
  INV_X1 U8942 ( .A(n12372), .ZN(n12773) );
  OR2_X1 U8943 ( .A1(n12731), .A2(n12277), .ZN(n6577) );
  AND2_X1 U8944 ( .A1(n11982), .A2(n7319), .ZN(n6578) );
  NAND2_X1 U8945 ( .A1(n7716), .A2(n7715), .ZN(n12040) );
  NAND2_X1 U8946 ( .A1(n9600), .A2(n15039), .ZN(n6579) );
  OR2_X1 U8947 ( .A1(n12301), .A2(n9645), .ZN(n6580) );
  INV_X1 U8948 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7018) );
  AND2_X1 U8949 ( .A1(n8076), .A2(n7028), .ZN(n6581) );
  OR2_X1 U8950 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14240), .ZN(n6582) );
  AND2_X1 U8951 ( .A1(n9015), .A2(n7391), .ZN(n6583) );
  NOR2_X1 U8952 ( .A1(n14489), .A2(n13713), .ZN(n6584) );
  INV_X1 U8953 ( .A(n7055), .ZN(n7054) );
  OR2_X1 U8954 ( .A1(n12062), .A2(n10579), .ZN(n6585) );
  INV_X1 U8955 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6746) );
  AND2_X1 U8956 ( .A1(n8495), .A2(n8494), .ZN(n6586) );
  AND2_X1 U8957 ( .A1(n7738), .A2(n7724), .ZN(n6587) );
  NAND2_X1 U8958 ( .A1(n12009), .A2(n10034), .ZN(n6588) );
  AND2_X1 U8959 ( .A1(n9616), .A2(n9615), .ZN(n6589) );
  AND2_X1 U8960 ( .A1(n8085), .A2(n8084), .ZN(n6590) );
  OR2_X1 U8961 ( .A1(n7353), .A2(n8771), .ZN(n6591) );
  OR2_X1 U8962 ( .A1(n11724), .A2(n11722), .ZN(n6592) );
  AND2_X1 U8963 ( .A1(n12773), .A2(n9519), .ZN(n6593) );
  OR2_X1 U8964 ( .A1(n8789), .A2(n8787), .ZN(n6594) );
  AND2_X1 U8965 ( .A1(n14004), .A2(n8087), .ZN(n6595) );
  OR2_X1 U8966 ( .A1(n8736), .A2(n7355), .ZN(n6596) );
  OR2_X1 U8967 ( .A1(n8756), .A2(n8754), .ZN(n6597) );
  OR2_X1 U8968 ( .A1(n7419), .A2(n11758), .ZN(n6598) );
  OR2_X1 U8969 ( .A1(n8719), .A2(n8721), .ZN(n6599) );
  OR2_X1 U8970 ( .A1(n7421), .A2(n11736), .ZN(n6600) );
  OR2_X1 U8971 ( .A1(n7351), .A2(n8720), .ZN(n6601) );
  OR2_X1 U8972 ( .A1(n11735), .A2(n11737), .ZN(n6602) );
  OR2_X1 U8973 ( .A1(n9276), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n6603) );
  INV_X1 U8974 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7396) );
  INV_X1 U8975 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8019) );
  AND2_X1 U8976 ( .A1(n11828), .A2(n11830), .ZN(n6604) );
  OR2_X1 U8977 ( .A1(n7428), .A2(n7427), .ZN(n6605) );
  NAND2_X1 U8978 ( .A1(n11841), .A2(n7416), .ZN(n6606) );
  INV_X1 U8979 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6683) );
  INV_X2 U8980 ( .A(n12062), .ZN(n12132) );
  XNOR2_X1 U8981 ( .A(n9032), .B(n9031), .ZN(n12623) );
  INV_X1 U8982 ( .A(n11276), .ZN(n7001) );
  NAND2_X1 U8983 ( .A1(n7792), .A2(n7234), .ZN(n11653) );
  NAND2_X1 U8984 ( .A1(n7070), .A2(n6515), .ZN(n12772) );
  AND2_X1 U8985 ( .A1(n7451), .A2(n7453), .ZN(n6607) );
  CLKBUF_X1 U8986 ( .A(n9591), .Z(n12404) );
  AND2_X1 U8987 ( .A1(n13987), .A2(n6902), .ZN(n6608) );
  INV_X1 U8988 ( .A(n7538), .ZN(n11852) );
  OR3_X1 U8989 ( .A1(n12470), .A2(n12469), .A3(n12514), .ZN(n6609) );
  NAND2_X1 U8990 ( .A1(n6711), .A2(n8078), .ZN(n11334) );
  NAND2_X1 U8991 ( .A1(n7090), .A2(n12457), .ZN(n11501) );
  NAND2_X1 U8992 ( .A1(n7042), .A2(n8079), .ZN(n11452) );
  OAI21_X1 U8993 ( .B1(n11240), .B2(n6820), .A(n6817), .ZN(n14396) );
  NAND2_X1 U8994 ( .A1(n6712), .A2(n7030), .ZN(n11319) );
  NAND2_X1 U8995 ( .A1(n6979), .A2(n9514), .ZN(n11502) );
  NAND2_X1 U8996 ( .A1(n14468), .A2(n12061), .ZN(n13615) );
  INV_X1 U8997 ( .A(n13626), .ZN(n7158) );
  NAND2_X1 U8998 ( .A1(n8002), .A2(n8001), .ZN(n14065) );
  NAND2_X1 U8999 ( .A1(n9177), .A2(n9014), .ZN(n9276) );
  AND4_X1 U9000 ( .A1(n8542), .A2(n8541), .A3(n8540), .A4(n8539), .ZN(n12971)
         );
  INV_X1 U9001 ( .A(n12971), .ZN(n13101) );
  NOR2_X1 U9002 ( .A1(n12537), .A2(n12514), .ZN(n6610) );
  INV_X1 U9003 ( .A(n12647), .ZN(n9557) );
  NAND2_X1 U9004 ( .A1(n9027), .A2(n9026), .ZN(n12647) );
  NAND2_X1 U9005 ( .A1(n11619), .A2(n6937), .ZN(n6938) );
  OR2_X1 U9006 ( .A1(n11186), .A2(n15081), .ZN(n6611) );
  INV_X1 U9007 ( .A(n8797), .ZN(n7358) );
  INV_X1 U9008 ( .A(n6889), .ZN(n14030) );
  NOR2_X1 U9009 ( .A1(n14031), .A2(n14125), .ZN(n6889) );
  OR2_X1 U9010 ( .A1(n12590), .A2(n11189), .ZN(n6612) );
  INV_X1 U9011 ( .A(n6891), .ZN(n11655) );
  INV_X1 U9012 ( .A(n8584), .ZN(n7311) );
  AND2_X1 U9013 ( .A1(n9967), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6613) );
  OAI21_X1 U9014 ( .B1(n13502), .B2(n13531), .A(n7145), .ZN(n7144) );
  AND2_X1 U9015 ( .A1(n12459), .A2(n12457), .ZN(n6614) );
  INV_X1 U9016 ( .A(n6974), .ZN(n6973) );
  NOR2_X1 U9017 ( .A1(n7850), .A2(n6975), .ZN(n6974) );
  OR2_X1 U9018 ( .A1(n7358), .A2(n8796), .ZN(n6615) );
  AND2_X1 U9019 ( .A1(n7310), .A2(n8584), .ZN(n6616) );
  NAND2_X1 U9020 ( .A1(n8467), .A2(n8466), .ZN(n13332) );
  INV_X1 U9021 ( .A(n13332), .ZN(n6930) );
  NAND2_X1 U9022 ( .A1(n8414), .A2(n8413), .ZN(n13477) );
  INV_X1 U9023 ( .A(n13477), .ZN(n6936) );
  NAND2_X1 U9024 ( .A1(n7802), .A2(n7801), .ZN(n13623) );
  INV_X1 U9025 ( .A(n13623), .ZN(n6890) );
  NAND2_X1 U9026 ( .A1(n7347), .A2(n6650), .ZN(n11410) );
  INV_X1 U9027 ( .A(n14439), .ZN(n7308) );
  NAND2_X1 U9028 ( .A1(n7060), .A2(n7058), .ZN(n11273) );
  INV_X1 U9029 ( .A(n14119), .ZN(n6888) );
  AND2_X1 U9030 ( .A1(n12340), .A2(SI_30_), .ZN(n6617) );
  NOR2_X1 U9031 ( .A1(n14939), .A2(n11205), .ZN(n6618) );
  INV_X1 U9032 ( .A(n14404), .ZN(n7132) );
  OR2_X1 U9033 ( .A1(n15076), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6619) );
  INV_X1 U9034 ( .A(n7099), .ZN(n7098) );
  NAND2_X1 U9035 ( .A1(n14981), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7099) );
  AND2_X1 U9036 ( .A1(n7979), .A2(SI_27_), .ZN(n6620) );
  NOR2_X1 U9037 ( .A1(n15085), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U9038 ( .A1(n11082), .A2(n6491), .ZN(n6898) );
  OAI21_X1 U9039 ( .B1(n10393), .B2(n7558), .A(n10391), .ZN(n10529) );
  AND2_X1 U9040 ( .A1(n11393), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6622) );
  INV_X1 U9041 ( .A(SI_26_), .ZN(n15186) );
  INV_X1 U9042 ( .A(n9956), .ZN(n10263) );
  INV_X1 U9043 ( .A(n12832), .ZN(n15038) );
  INV_X1 U9044 ( .A(n14836), .ZN(n7143) );
  INV_X1 U9045 ( .A(n11112), .ZN(n7297) );
  AND2_X1 U9046 ( .A1(n10023), .A2(n14805), .ZN(n13485) );
  INV_X1 U9047 ( .A(n10408), .ZN(n6932) );
  OR2_X1 U9048 ( .A1(n9588), .A2(n12404), .ZN(n10656) );
  AND2_X1 U9049 ( .A1(n12529), .A2(n12398), .ZN(n12504) );
  NAND2_X1 U9050 ( .A1(n12585), .A2(n12610), .ZN(n6623) );
  NOR2_X1 U9051 ( .A1(n12565), .A2(n14331), .ZN(n6803) );
  NAND2_X1 U9052 ( .A1(n6526), .A2(n7004), .ZN(n10736) );
  AND2_X1 U9053 ( .A1(n14155), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6624) );
  AND2_X1 U9054 ( .A1(n7267), .A2(n12335), .ZN(n6625) );
  OR2_X1 U9055 ( .A1(n6681), .A2(n13540), .ZN(n6626) );
  OR2_X1 U9056 ( .A1(n9044), .A2(n12398), .ZN(n6627) );
  NOR2_X1 U9057 ( .A1(n9009), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U9058 ( .A1(n12623), .A2(n10515), .ZN(n9547) );
  INV_X1 U9059 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7211) );
  INV_X1 U9060 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7210) );
  INV_X1 U9061 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6654) );
  INV_X1 U9062 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6739) );
  AND2_X1 U9063 ( .A1(n9931), .A2(n9730), .ZN(n9943) );
  NOR2_X1 U9064 ( .A1(n6802), .A2(n12612), .ZN(n6801) );
  XNOR2_X1 U9065 ( .A(n12581), .B(n12612), .ZN(n14333) );
  XNOR2_X1 U9066 ( .A(n11263), .B(n6637), .ZN(n11407) );
  INV_X2 U9067 ( .A(n8871), .ZN(n8867) );
  NAND3_X1 U9068 ( .A1(n6631), .A2(n6594), .A3(n6630), .ZN(n6689) );
  NAND3_X1 U9069 ( .A1(n8707), .A2(n7359), .A3(n8706), .ZN(n6656) );
  NAND2_X1 U9070 ( .A1(n6628), .A2(n7350), .ZN(n8759) );
  NAND3_X1 U9071 ( .A1(n8753), .A2(n6597), .A3(n8752), .ZN(n6628) );
  NAND2_X1 U9072 ( .A1(n6629), .A2(n7357), .ZN(n8800) );
  NAND3_X1 U9073 ( .A1(n6673), .A2(n6615), .A3(n6672), .ZN(n6629) );
  NAND2_X1 U9074 ( .A1(n8786), .A2(n8785), .ZN(n6630) );
  NAND2_X1 U9075 ( .A1(n8782), .A2(n8781), .ZN(n6631) );
  AND3_X4 U9076 ( .A1(n8191), .A2(n8192), .A3(n7448), .ZN(n10689) );
  NAND2_X2 U9077 ( .A1(n8160), .A2(n8159), .ZN(n8489) );
  NAND3_X1 U9078 ( .A1(n8697), .A2(n6694), .A3(n8696), .ZN(n6693) );
  NAND3_X1 U9079 ( .A1(n8718), .A2(n6599), .A3(n8717), .ZN(n6690) );
  INV_X1 U9080 ( .A(n8684), .ZN(n8687) );
  NAND4_X1 U9081 ( .A1(n8680), .A2(n6691), .A3(n8679), .A4(n6692), .ZN(n8684)
         );
  NAND3_X2 U9082 ( .A1(n8178), .A2(n6632), .A3(n6541), .ZN(n10246) );
  XNOR2_X2 U9083 ( .A(n10683), .B(n13129), .ZN(n10248) );
  INV_X1 U9084 ( .A(n7142), .ZN(n7141) );
  NAND2_X1 U9085 ( .A1(n13374), .A2(n8594), .ZN(n13364) );
  NAND2_X1 U9086 ( .A1(n6824), .A2(n6823), .ZN(n13289) );
  NAND2_X1 U9087 ( .A1(n6836), .A2(n8607), .ZN(n13234) );
  NAND2_X1 U9088 ( .A1(n7291), .A2(n8563), .ZN(n6814) );
  NAND2_X1 U9089 ( .A1(n14396), .A2(n8579), .ZN(n8582) );
  NAND2_X1 U9090 ( .A1(n6816), .A2(n8565), .ZN(n10671) );
  AOI21_X1 U9091 ( .B1(n6502), .B2(n6867), .A(n6604), .ZN(n6863) );
  NAND2_X1 U9092 ( .A1(n6864), .A2(n6863), .ZN(n11833) );
  XNOR2_X1 U9093 ( .A(n7927), .B(SI_24_), .ZN(n7924) );
  INV_X1 U9094 ( .A(n6735), .ZN(n6734) );
  NAND2_X1 U9095 ( .A1(n7530), .A2(n7529), .ZN(n7548) );
  NAND2_X1 U9096 ( .A1(n10504), .A2(n10505), .ZN(n10546) );
  NAND2_X1 U9097 ( .A1(n7332), .A2(n6508), .ZN(n11141) );
  NOR2_X1 U9098 ( .A1(n13089), .A2(n13092), .ZN(n13090) );
  INV_X1 U9099 ( .A(n9046), .ZN(n9049) );
  NAND2_X1 U9100 ( .A1(n11027), .A2(n11026), .ZN(n11025) );
  NAND2_X1 U9101 ( .A1(n11231), .A2(n11230), .ZN(n11229) );
  NAND2_X1 U9102 ( .A1(n12273), .A2(n12274), .ZN(n7376) );
  AND2_X1 U9103 ( .A1(n7372), .A2(n7369), .ZN(n7368) );
  XNOR2_X1 U9104 ( .A(n11962), .B(n11963), .ZN(n13089) );
  NAND2_X1 U9105 ( .A1(n10503), .A2(n10502), .ZN(n10504) );
  NAND2_X1 U9106 ( .A1(n11440), .A2(n11439), .ZN(n11559) );
  NAND2_X1 U9107 ( .A1(n11101), .A2(n11100), .ZN(n7332) );
  NAND2_X1 U9108 ( .A1(n11141), .A2(n11140), .ZN(n11262) );
  XNOR2_X1 U9109 ( .A(n10153), .B(n10154), .ZN(n10028) );
  NOR2_X2 U9111 ( .A1(n13090), .A2(n7439), .ZN(n13014) );
  OAI21_X2 U9112 ( .B1(n11262), .B2(n7346), .A(n7344), .ZN(n11430) );
  NOR2_X1 U9113 ( .A1(n10376), .A2(n7339), .ZN(n7340) );
  NAND2_X1 U9114 ( .A1(n10027), .A2(n10028), .ZN(n10157) );
  OR2_X2 U9115 ( .A1(n13075), .A2(n13074), .ZN(n13072) );
  NAND2_X1 U9116 ( .A1(n6638), .A2(n12312), .ZN(n12314) );
  NAND2_X1 U9117 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  NAND2_X1 U9118 ( .A1(n7097), .A2(n9177), .ZN(n9046) );
  OAI21_X1 U9119 ( .B1(n12323), .B2(n12254), .A(n12321), .ZN(n9635) );
  INV_X4 U9120 ( .A(n10246), .ZN(n10683) );
  XNOR2_X2 U9121 ( .A(n8010), .B(n8009), .ZN(n14068) );
  NAND2_X1 U9122 ( .A1(n11338), .A2(n11337), .ZN(n11336) );
  NOR2_X2 U9123 ( .A1(n11939), .A2(n11942), .ZN(n11938) );
  NAND2_X1 U9124 ( .A1(n10957), .A2(n11902), .ZN(n10956) );
  NAND2_X1 U9125 ( .A1(n14001), .A2(n8086), .ZN(n13992) );
  NAND2_X1 U9126 ( .A1(n11448), .A2(n7740), .ZN(n11511) );
  NAND2_X1 U9127 ( .A1(n7601), .A2(n7600), .ZN(n6856) );
  NAND2_X1 U9128 ( .A1(n6856), .A2(n7603), .ZN(n7615) );
  NOR2_X1 U9129 ( .A1(n11041), .A2(n7218), .ZN(n7217) );
  AOI21_X1 U9130 ( .B1(n7216), .B2(n7218), .A(n6559), .ZN(n7215) );
  NAND2_X1 U9131 ( .A1(n11320), .A2(n7704), .ZN(n11338) );
  NAND2_X1 U9132 ( .A1(n13874), .A2(n13873), .ZN(n13872) );
  NAND2_X2 U9133 ( .A1(n13667), .A2(n13668), .ZN(n13583) );
  NAND2_X2 U9134 ( .A1(n7160), .A2(n12097), .ZN(n13593) );
  NAND2_X2 U9135 ( .A1(n12117), .A2(n13572), .ZN(n13574) );
  NAND2_X1 U9136 ( .A1(n6585), .A2(n10333), .ZN(n6642) );
  NAND2_X1 U9137 ( .A1(n13954), .A2(n13959), .ZN(n13953) );
  NAND3_X1 U9138 ( .A1(n7203), .A2(n7204), .A3(n7207), .ZN(n7509) );
  OAI22_X1 U9139 ( .A1(n13878), .A2(n13883), .B1(n13603), .B2(n13892), .ZN(
        n11939) );
  NOR2_X1 U9140 ( .A1(n11938), .A2(n7978), .ZN(n13874) );
  NOR4_X1 U9141 ( .A1(n12658), .A2(n12676), .A3(n12376), .A4(n12375), .ZN(
        n12377) );
  NAND2_X1 U9142 ( .A1(n7154), .A2(n7152), .ZN(n13611) );
  AOI21_X1 U9143 ( .B1(n12525), .B2(n9582), .A(n6659), .ZN(n12532) );
  NAND2_X1 U9144 ( .A1(n13562), .A2(n6647), .ZN(n13564) );
  OR2_X1 U9145 ( .A1(n12392), .A2(n6627), .ZN(n7271) );
  NAND2_X2 U9146 ( .A1(n8160), .A2(n8157), .ZN(n8545) );
  OAI21_X1 U9147 ( .B1(n12523), .B2(n9547), .A(n6660), .ZN(n6659) );
  OAI21_X2 U9148 ( .B1(n13967), .B2(n8089), .A(n7879), .ZN(n13954) );
  NAND2_X1 U9149 ( .A1(n10350), .A2(n10356), .ZN(n10352) );
  AND3_X2 U9150 ( .A1(n7520), .A2(n7521), .A3(n6544), .ZN(n10579) );
  INV_X4 U9151 ( .A(n8614), .ZN(n8842) );
  NAND2_X1 U9152 ( .A1(n7766), .A2(n11910), .ZN(n11509) );
  NAND2_X1 U9153 ( .A1(n6670), .A2(n13128), .ZN(n6669) );
  NAND2_X1 U9154 ( .A1(n11336), .A2(n6587), .ZN(n11448) );
  XNOR2_X1 U9155 ( .A(n14240), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15294) );
  NAND2_X1 U9156 ( .A1(n14276), .A2(n14275), .ZN(n6926) );
  NOR2_X1 U9157 ( .A1(n14282), .A2(n14283), .ZN(n14244) );
  INV_X1 U9158 ( .A(n14520), .ZN(n6908) );
  NAND2_X1 U9159 ( .A1(n14537), .A2(n6652), .ZN(n14543) );
  NAND2_X1 U9160 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  NAND2_X1 U9161 ( .A1(n10546), .A2(n10545), .ZN(n10716) );
  XNOR2_X1 U9162 ( .A(n6529), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  OAI21_X2 U9163 ( .B1(n10716), .B2(n10715), .A(n10714), .ZN(n10917) );
  NAND2_X1 U9164 ( .A1(n6656), .A2(n7360), .ZN(n8713) );
  NAND2_X1 U9165 ( .A1(n6657), .A2(n7170), .ZN(n13667) );
  NAND3_X1 U9166 ( .A1(n12058), .A2(n13687), .A3(n13616), .ZN(n6657) );
  INV_X1 U9167 ( .A(n10108), .ZN(n6708) );
  NAND2_X1 U9168 ( .A1(n12781), .A2(n6593), .ZN(n12764) );
  INV_X1 U9169 ( .A(n10939), .ZN(n9504) );
  NAND2_X1 U9170 ( .A1(n6976), .A2(n9507), .ZN(n11176) );
  OAI21_X2 U9171 ( .B1(n12811), .B2(n6553), .A(n9517), .ZN(n12793) );
  AOI21_X2 U9172 ( .B1(n7007), .B2(n7006), .A(n6562), .ZN(n12706) );
  NAND2_X1 U9173 ( .A1(n10063), .A2(n10064), .ZN(n10446) );
  NOR2_X1 U9174 ( .A1(n14301), .A2(n12816), .ZN(n14300) );
  INV_X1 U9175 ( .A(n7110), .ZN(n7109) );
  XNOR2_X1 U9176 ( .A(n6806), .B(n10754), .ZN(n10629) );
  NOR2_X1 U9177 ( .A1(n14990), .A2(n12561), .ZN(n15010) );
  OAI21_X1 U9178 ( .B1(n6687), .B2(n6688), .A(n7354), .ZN(n8740) );
  NAND2_X1 U9179 ( .A1(n8735), .A2(n6596), .ZN(n6687) );
  NAND2_X1 U9180 ( .A1(n9402), .A2(n8997), .ZN(n8999) );
  OR2_X2 U9181 ( .A1(n9308), .A2(n9307), .ZN(n9310) );
  NAND2_X1 U9182 ( .A1(n6776), .A2(n6775), .ZN(n6780) );
  OAI211_X1 U9183 ( .C1(n6777), .C2(n12512), .A(n6774), .B(n6784), .ZN(n6773)
         );
  OAI21_X1 U9184 ( .B1(n14068), .B2(n14583), .A(n6662), .ZN(n14135) );
  XNOR2_X2 U9185 ( .A(n13722), .B(n6661), .ZN(n10556) );
  NAND2_X1 U9186 ( .A1(n6663), .A2(n8946), .ZN(n9120) );
  NAND2_X1 U9187 ( .A1(n8945), .A2(n9111), .ZN(n6663) );
  NAND2_X1 U9188 ( .A1(n6780), .A2(n12521), .ZN(n12523) );
  INV_X1 U9189 ( .A(n6785), .ZN(n6781) );
  NAND2_X1 U9190 ( .A1(n10956), .A2(n7645), .ZN(n11080) );
  NAND2_X1 U9191 ( .A1(n6778), .A2(n6782), .ZN(n6774) );
  NAND2_X1 U9192 ( .A1(n9448), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U9193 ( .A1(n13227), .A2(n13233), .ZN(n13229) );
  NAND2_X1 U9194 ( .A1(n13395), .A2(n8422), .ZN(n13373) );
  NAND2_X1 U9195 ( .A1(n10405), .A2(n8217), .ZN(n10516) );
  NAND2_X1 U9196 ( .A1(n11662), .A2(n11664), .ZN(n11661) );
  OAI21_X1 U9197 ( .B1(n13317), .B2(n8485), .A(n8897), .ZN(n13293) );
  OAI22_X1 U9198 ( .A1(n11244), .A2(n8321), .B1(n13118), .B2(n11263), .ZN(
        n11213) );
  AOI211_X2 U9199 ( .C1(n14816), .C2(n13216), .A(n13223), .B(n13217), .ZN(
        n8944) );
  XNOR2_X1 U9200 ( .A(n6933), .B(n8166), .ZN(n8612) );
  NAND2_X1 U9201 ( .A1(n11559), .A2(n7348), .ZN(n11961) );
  NAND2_X1 U9202 ( .A1(n8684), .A2(n8685), .ZN(n8683) );
  AOI21_X1 U9203 ( .B1(n8731), .B2(n8732), .A(n6665), .ZN(n6688) );
  XNOR2_X1 U9204 ( .A(n11986), .B(n11984), .ZN(n13052) );
  NAND2_X1 U9205 ( .A1(n9655), .A2(n9654), .ZN(n7373) );
  NAND2_X1 U9206 ( .A1(n14845), .A2(n14844), .ZN(n14843) );
  INV_X1 U9207 ( .A(n10832), .ZN(n7369) );
  NOR2_X1 U9208 ( .A1(n9633), .A2(n9631), .ZN(n12323) );
  NAND2_X1 U9209 ( .A1(n7370), .A2(n7371), .ZN(n14858) );
  NAND2_X1 U9210 ( .A1(n10611), .A2(n10612), .ZN(n7370) );
  NAND2_X1 U9211 ( .A1(n9331), .A2(n9347), .ZN(n9362) );
  AOI21_X1 U9212 ( .B1(n9919), .B2(n9865), .A(n9864), .ZN(n9969) );
  NAND2_X1 U9213 ( .A1(n6697), .A2(n6696), .ZN(n14739) );
  NOR2_X1 U9214 ( .A1(n14683), .A2(n14682), .ZN(n14681) );
  NOR2_X1 U9215 ( .A1(n10096), .A2(n10095), .ZN(n10094) );
  NOR2_X1 U9216 ( .A1(n10086), .A2(n10085), .ZN(n10084) );
  NAND2_X1 U9217 ( .A1(n10996), .A2(n12436), .ZN(n6976) );
  INV_X1 U9218 ( .A(n11678), .ZN(n10636) );
  OAI22_X2 U9219 ( .A1(n12693), .A2(n9522), .B1(n12708), .B2(n12923), .ZN(
        n12677) );
  NAND2_X1 U9220 ( .A1(n9500), .A2(n9499), .ZN(n11094) );
  NAND2_X1 U9221 ( .A1(n7003), .A2(n9496), .ZN(n10659) );
  INV_X1 U9222 ( .A(n12717), .ZN(n7007) );
  INV_X1 U9223 ( .A(n8185), .ZN(n8206) );
  NAND2_X1 U9224 ( .A1(n8795), .A2(n8794), .ZN(n6672) );
  NAND2_X1 U9225 ( .A1(n8791), .A2(n8790), .ZN(n6673) );
  INV_X1 U9226 ( .A(n7361), .ZN(n7359) );
  NAND2_X1 U9227 ( .A1(n6674), .A2(n10115), .ZN(n10235) );
  INV_X1 U9228 ( .A(n10117), .ZN(n6674) );
  NAND2_X1 U9229 ( .A1(n10234), .A2(n7149), .ZN(n10117) );
  OAI22_X2 U9230 ( .A1(n14046), .A2(n10334), .B1(n12109), .B2(n14590), .ZN(
        n10112) );
  AND2_X4 U9231 ( .A1(n9931), .A2(n9930), .ZN(n12147) );
  NAND2_X2 U9232 ( .A1(n9868), .A2(n7495), .ZN(n8864) );
  NAND2_X2 U9233 ( .A1(n8612), .A2(n13547), .ZN(n9868) );
  NAND2_X1 U9234 ( .A1(n6693), .A2(n7366), .ZN(n8702) );
  NAND2_X1 U9235 ( .A1(n6689), .A2(n7356), .ZN(n8792) );
  NAND2_X1 U9236 ( .A1(n6690), .A2(n6601), .ZN(n8724) );
  NAND2_X1 U9237 ( .A1(n8780), .A2(n8779), .ZN(n8783) );
  NAND2_X1 U9238 ( .A1(n8689), .A2(n8688), .ZN(n8692) );
  NAND3_X1 U9239 ( .A1(n10683), .A2(n13129), .A3(n8884), .ZN(n6692) );
  XNOR2_X2 U9240 ( .A(n7148), .B(n6676), .ZN(n13541) );
  AND3_X2 U9241 ( .A1(n8126), .A2(n8124), .A3(n8125), .ZN(n8143) );
  NAND2_X1 U9242 ( .A1(n13072), .A2(n12004), .ZN(n12970) );
  NAND2_X1 U9243 ( .A1(n11430), .A2(n11429), .ZN(n11437) );
  XNOR2_X1 U9244 ( .A(n13155), .B(n13171), .ZN(n14717) );
  NAND2_X1 U9245 ( .A1(n14716), .A2(n13156), .ZN(n14729) );
  NAND2_X1 U9246 ( .A1(n14698), .A2(n14697), .ZN(n14696) );
  INV_X1 U9247 ( .A(n13186), .ZN(n6697) );
  AOI21_X1 U9248 ( .B1(n7221), .B2(n7222), .A(n6584), .ZN(n7219) );
  XNOR2_X1 U9249 ( .A(n7509), .B(n9712), .ZN(n7511) );
  AOI21_X2 U9250 ( .B1(n12657), .B2(n12832), .A(n12656), .ZN(n12849) );
  NAND2_X1 U9251 ( .A1(n10736), .A2(n9596), .ZN(n7003) );
  NAND2_X1 U9252 ( .A1(n9516), .A2(n9515), .ZN(n12811) );
  INV_X1 U9253 ( .A(n9591), .ZN(n7004) );
  NAND2_X1 U9254 ( .A1(n6997), .A2(n6996), .ZN(n11394) );
  NAND2_X1 U9255 ( .A1(n6978), .A2(n6977), .ZN(n12825) );
  NAND3_X1 U9256 ( .A1(n8152), .A2(n7365), .A3(n8123), .ZN(n6679) );
  NAND2_X2 U9257 ( .A1(n11590), .A2(n7790), .ZN(n7792) );
  NAND2_X2 U9258 ( .A1(n13934), .A2(n7239), .ZN(n13917) );
  NAND2_X1 U9259 ( .A1(n7220), .A2(n7219), .ZN(n11322) );
  OAI21_X2 U9260 ( .B1(n8994), .B2(P1_DATAO_REG_20__SCAN_IN), .A(n8995), .ZN(
        n9391) );
  NAND2_X1 U9261 ( .A1(n7248), .A2(n7247), .ZN(n9275) );
  NAND2_X1 U9262 ( .A1(n9213), .A2(n8968), .ZN(n9222) );
  NAND2_X1 U9263 ( .A1(n7073), .A2(n7071), .ZN(n12346) );
  AND2_X4 U9264 ( .A1(n9929), .A2(n9931), .ZN(n12148) );
  OAI21_X2 U9265 ( .B1(n8035), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8034) );
  AOI21_X2 U9266 ( .B1(n8888), .B2(n8887), .A(n8886), .ZN(n8929) );
  NAND2_X1 U9267 ( .A1(n8792), .A2(n8793), .ZN(n8791) );
  NAND2_X1 U9268 ( .A1(n8759), .A2(n8760), .ZN(n8758) );
  NAND2_X1 U9269 ( .A1(n8713), .A2(n8714), .ZN(n8712) );
  NAND2_X1 U9270 ( .A1(n8724), .A2(n8725), .ZN(n8723) );
  NAND2_X1 U9271 ( .A1(n8770), .A2(n6591), .ZN(n6685) );
  NAND2_X1 U9272 ( .A1(n8805), .A2(n8804), .ZN(n8808) );
  NAND2_X1 U9273 ( .A1(n8745), .A2(n8744), .ZN(n8748) );
  NAND2_X1 U9274 ( .A1(n8800), .A2(n8801), .ZN(n8799) );
  NAND2_X1 U9275 ( .A1(n14717), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14716) );
  NAND2_X1 U9276 ( .A1(n14709), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14708) );
  CLKBUF_X2 U9277 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n14663) );
  AOI21_X1 U9278 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(n8880) );
  INV_X2 U9279 ( .A(n8681), .ZN(n8884) );
  NAND2_X1 U9280 ( .A1(n7127), .A2(n7125), .ZN(n10663) );
  OAI21_X2 U9281 ( .B1(n7792), .B2(n7231), .A(n7229), .ZN(n14001) );
  NAND2_X2 U9282 ( .A1(n7909), .A2(n7908), .ZN(n13934) );
  NOR2_X2 U9283 ( .A1(n13896), .A2(n7945), .ZN(n13878) );
  NAND2_X1 U9284 ( .A1(n11322), .A2(n11321), .ZN(n11320) );
  NAND2_X1 U9285 ( .A1(n7205), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7208) );
  NAND2_X2 U9286 ( .A1(n7587), .A2(n7586), .ZN(n7601) );
  NOR2_X1 U9287 ( .A1(n11900), .A2(n7217), .ZN(n7216) );
  AOI22_X2 U9288 ( .A1(n10785), .A2(n10784), .B1(n10782), .B2(n10783), .ZN(
        n10894) );
  XNOR2_X2 U9289 ( .A(n10781), .B(n10782), .ZN(n10785) );
  INV_X1 U9290 ( .A(n9933), .ZN(n9934) );
  NAND2_X1 U9291 ( .A1(n6707), .A2(n6704), .ZN(P1_U3214) );
  NAND2_X1 U9292 ( .A1(n13564), .A2(n14483), .ZN(n6707) );
  NAND3_X2 U9293 ( .A1(n7487), .A2(n6709), .A3(n7488), .ZN(n11700) );
  NAND2_X1 U9294 ( .A1(n7571), .A2(n6710), .ZN(n6709) );
  NOR2_X2 U9295 ( .A1(n8017), .A2(n7431), .ZN(n7476) );
  OAI21_X1 U9296 ( .B1(n6718), .B2(n6714), .A(n6713), .ZN(n8072) );
  NAND3_X1 U9297 ( .A1(n6716), .A2(n8070), .A3(n6715), .ZN(n10960) );
  INV_X1 U9298 ( .A(n11900), .ZN(n6721) );
  NAND3_X1 U9299 ( .A1(n14020), .A2(n6724), .A3(n8089), .ZN(n6723) );
  NAND3_X1 U9300 ( .A1(n6723), .A2(n6722), .A3(n8090), .ZN(n13960) );
  NAND3_X1 U9301 ( .A1(n6724), .A2(n7055), .A3(n8089), .ZN(n6722) );
  NAND2_X1 U9302 ( .A1(n13937), .A2(n6730), .ZN(n6729) );
  NAND2_X1 U9303 ( .A1(n7241), .A2(n7813), .ZN(n8017) );
  NAND3_X1 U9304 ( .A1(n7241), .A2(n7813), .A3(n6510), .ZN(n6738) );
  NAND3_X1 U9305 ( .A1(n6747), .A2(n9011), .A3(n6746), .ZN(n9145) );
  INV_X1 U9306 ( .A(n12461), .ZN(n6751) );
  INV_X1 U9307 ( .A(n12465), .ZN(n6760) );
  NAND2_X1 U9308 ( .A1(n6761), .A2(n6762), .ZN(n12452) );
  NAND2_X1 U9309 ( .A1(n12441), .A2(n6764), .ZN(n6761) );
  NAND3_X1 U9310 ( .A1(n12378), .A2(n12519), .A3(n6783), .ZN(n6770) );
  NOR2_X1 U9311 ( .A1(n6773), .A2(n6772), .ZN(n6776) );
  NAND3_X1 U9312 ( .A1(n12493), .A2(n12492), .A3(n12714), .ZN(n6794) );
  NAND2_X1 U9313 ( .A1(n9177), .A2(n6795), .ZN(n9034) );
  INV_X1 U9314 ( .A(n9034), .ZN(n9028) );
  NAND2_X1 U9315 ( .A1(n14325), .A2(n6801), .ZN(n6797) );
  NOR2_X1 U9316 ( .A1(n14339), .A2(n14340), .ZN(n14341) );
  OR2_X1 U9317 ( .A1(n14325), .A2(n14324), .ZN(n14323) );
  NAND2_X1 U9318 ( .A1(n7102), .A2(n6509), .ZN(n6808) );
  NAND2_X1 U9319 ( .A1(n6808), .A2(n6809), .ZN(n12560) );
  XNOR2_X1 U9320 ( .A(n12560), .B(n12599), .ZN(n14991) );
  NAND3_X1 U9321 ( .A1(n6815), .A2(n10517), .A3(n6814), .ZN(n6816) );
  NAND2_X1 U9322 ( .A1(n7284), .A2(n10671), .ZN(n7288) );
  NAND2_X1 U9323 ( .A1(n7283), .A2(n6821), .ZN(n13374) );
  NAND2_X1 U9324 ( .A1(n13343), .A2(n6499), .ZN(n6824) );
  NAND2_X1 U9325 ( .A1(n6828), .A2(n6829), .ZN(n8609) );
  NAND2_X1 U9326 ( .A1(n6837), .A2(n6832), .ZN(n6836) );
  NAND3_X1 U9327 ( .A1(n8152), .A2(n8123), .A3(n6506), .ZN(n6838) );
  NOR2_X1 U9328 ( .A1(n14336), .A2(n14335), .ZN(n14334) );
  AND2_X1 U9329 ( .A1(n9177), .A2(n9020), .ZN(n6852) );
  NAND2_X1 U9330 ( .A1(n7097), .A2(n6851), .ZN(n6850) );
  NAND4_X1 U9331 ( .A1(n7210), .A2(n13201), .A3(n7479), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7201) );
  MUX2_X1 U9332 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7495), .Z(n7549) );
  NAND2_X1 U9333 ( .A1(n7601), .A2(n6857), .ZN(n6854) );
  NAND2_X1 U9334 ( .A1(n6860), .A2(n11805), .ZN(n11808) );
  OAI21_X1 U9335 ( .B1(n6571), .B2(n6862), .A(n6861), .ZN(n6860) );
  OAI21_X1 U9336 ( .B1(n11791), .B2(n11790), .A(n6532), .ZN(n6862) );
  NAND2_X1 U9337 ( .A1(n11826), .A2(n6502), .ZN(n6864) );
  OAI21_X1 U9338 ( .B1(n6547), .B2(n6873), .A(n6870), .ZN(n11819) );
  NOR2_X2 U9339 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10060) );
  NAND2_X1 U9340 ( .A1(n10060), .A2(n9122), .ZN(n9132) );
  XNOR2_X2 U9341 ( .A(n7474), .B(n7473), .ZN(n8098) );
  NOR3_X4 U9342 ( .A1(n13867), .A2(n14070), .A3(n14065), .ZN(n13855) );
  NOR2_X1 U9343 ( .A1(n13867), .A2(n14070), .ZN(n6895) );
  INV_X1 U9344 ( .A(n14065), .ZN(n6894) );
  INV_X1 U9345 ( .A(n6898), .ZN(n11339) );
  NAND2_X1 U9346 ( .A1(n6908), .A2(n6905), .ZN(n14249) );
  NAND2_X1 U9347 ( .A1(n6907), .A2(n6906), .ZN(n6905) );
  INV_X1 U9348 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U9349 ( .A1(n14521), .A2(n14522), .ZN(n6907) );
  NAND2_X1 U9350 ( .A1(n6910), .A2(n6909), .ZN(n14267) );
  NAND2_X1 U9351 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  INV_X1 U9352 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U9353 ( .A1(n14297), .A2(n14296), .ZN(n6912) );
  OR2_X1 U9354 ( .A1(n14543), .A2(n14542), .ZN(n6913) );
  NAND2_X1 U9355 ( .A1(n14541), .A2(n14255), .ZN(n6914) );
  NAND2_X1 U9356 ( .A1(n14543), .A2(n14542), .ZN(n14541) );
  OAI21_X2 U9357 ( .B1(n8639), .B2(n7364), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6933) );
  NOR2_X2 U9358 ( .A1(n10986), .A2(n11112), .ZN(n11013) );
  NAND2_X1 U9359 ( .A1(n6935), .A2(n11619), .ZN(n13400) );
  INV_X1 U9360 ( .A(n6938), .ZN(n11670) );
  AND2_X1 U9361 ( .A1(n13266), .A2(n6939), .ZN(n13208) );
  AND2_X1 U9362 ( .A1(n13266), .A2(n13252), .ZN(n13248) );
  NAND2_X1 U9363 ( .A1(n13266), .A2(n6940), .ZN(n13209) );
  NAND2_X1 U9364 ( .A1(n7584), .A2(n7583), .ZN(n7587) );
  NAND2_X1 U9365 ( .A1(n7568), .A2(n7567), .ZN(n6943) );
  INV_X1 U9366 ( .A(n7948), .ZN(n6950) );
  OAI21_X1 U9367 ( .B1(n7948), .B2(n7947), .A(n7946), .ZN(n7962) );
  OAI21_X1 U9368 ( .B1(n7707), .B2(n6965), .A(n6962), .ZN(n7794) );
  OAI21_X1 U9369 ( .B1(n7810), .B2(n7809), .A(n7812), .ZN(n7851) );
  NAND2_X1 U9370 ( .A1(n7810), .A2(n6974), .ZN(n6967) );
  OAI211_X1 U9371 ( .C1(n10996), .C2(n12436), .A(n6976), .B(n12832), .ZN(
        n10999) );
  NAND2_X1 U9372 ( .A1(n11491), .A2(n6980), .ZN(n6978) );
  NAND2_X1 U9373 ( .A1(n9524), .A2(n6987), .ZN(n6984) );
  NAND2_X1 U9374 ( .A1(n6984), .A2(n6985), .ZN(n9566) );
  NAND2_X1 U9375 ( .A1(n9524), .A2(n9523), .ZN(n12653) );
  NAND4_X1 U9376 ( .A1(n9018), .A2(n9019), .A3(n9037), .A4(n9080), .ZN(n6995)
         );
  NAND2_X1 U9377 ( .A1(n11274), .A2(n6999), .ZN(n6997) );
  AOI21_X1 U9378 ( .B1(n7001), .B2(n9511), .A(n7000), .ZN(n6999) );
  NOR2_X2 U9379 ( .A1(n9495), .A2(n15031), .ZN(n9591) );
  NAND2_X1 U9380 ( .A1(n12764), .A2(n9520), .ZN(n12753) );
  OR2_X1 U9381 ( .A1(n9572), .A2(n7013), .ZN(n7010) );
  NAND2_X1 U9382 ( .A1(n9572), .A2(n12832), .ZN(n7014) );
  NAND2_X1 U9383 ( .A1(n7010), .A2(n7011), .ZN(n9579) );
  NAND2_X2 U9384 ( .A1(n9025), .A2(n9092), .ZN(n11956) );
  OR2_X2 U9385 ( .A1(n9053), .A2(n7017), .ZN(n9092) );
  NAND2_X1 U9386 ( .A1(n11650), .A2(n8082), .ZN(n14020) );
  INV_X1 U9387 ( .A(n7020), .ZN(n8011) );
  NOR2_X2 U9388 ( .A1(n7020), .A2(n6563), .ZN(n7241) );
  NAND3_X1 U9389 ( .A1(n8076), .A2(n7028), .A3(n7032), .ZN(n7031) );
  NAND2_X1 U9390 ( .A1(n11334), .A2(n7043), .ZN(n7039) );
  OAI21_X1 U9391 ( .B1(n7056), .B2(n7198), .A(n8088), .ZN(n7055) );
  NAND2_X1 U9392 ( .A1(n8072), .A2(n8071), .ZN(n10958) );
  NAND2_X1 U9393 ( .A1(n7206), .A2(n7210), .ZN(n7209) );
  OAI21_X1 U9394 ( .B1(n13960), .B2(n13959), .A(n8091), .ZN(n13939) );
  OR2_X2 U9395 ( .A1(n7476), .A2(n7588), .ZN(n7474) );
  OR2_X1 U9396 ( .A1(n10539), .A2(n11721), .ZN(n10642) );
  NAND2_X1 U9397 ( .A1(n10995), .A2(n7061), .ZN(n7060) );
  OAI21_X1 U9398 ( .B1(n12777), .B2(n7067), .A(n7064), .ZN(n12752) );
  NAND2_X1 U9399 ( .A1(n12680), .A2(n6527), .ZN(n7079) );
  OAI21_X1 U9400 ( .B1(n12738), .B2(n7082), .A(n7084), .ZN(n12704) );
  INV_X1 U9401 ( .A(n7089), .ZN(n12737) );
  OR2_X1 U9402 ( .A1(n7089), .A2(n7087), .ZN(n12725) );
  NAND2_X1 U9403 ( .A1(n7090), .A2(n6614), .ZN(n9291) );
  NAND3_X1 U9404 ( .A1(n9231), .A2(n7000), .A3(n9230), .ZN(n11256) );
  NAND2_X1 U9405 ( .A1(n11256), .A2(n12446), .ZN(n11398) );
  NAND2_X1 U9406 ( .A1(n9231), .A2(n9230), .ZN(n11258) );
  NOR2_X2 U9407 ( .A1(n14300), .A2(n12564), .ZN(n14325) );
  XNOR2_X1 U9408 ( .A(n12563), .B(n12604), .ZN(n14301) );
  OR2_X2 U9409 ( .A1(n14956), .A2(n9253), .ZN(n7102) );
  AND2_X2 U9410 ( .A1(n7105), .A2(n7104), .ZN(n14358) );
  NAND3_X1 U9411 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U9412 ( .A1(n7113), .A2(n7114), .ZN(n14918) );
  INV_X1 U9413 ( .A(n10449), .ZN(n7113) );
  NAND2_X1 U9414 ( .A1(n10448), .A2(n10447), .ZN(n7114) );
  NAND2_X1 U9415 ( .A1(n10881), .A2(n7118), .ZN(n7115) );
  INV_X1 U9416 ( .A(n8179), .ZN(n7124) );
  AND2_X1 U9417 ( .A1(n7121), .A2(n10266), .ZN(n7123) );
  NAND2_X1 U9418 ( .A1(n7122), .A2(n8179), .ZN(n7121) );
  INV_X1 U9419 ( .A(n10244), .ZN(n7122) );
  OAI21_X1 U9420 ( .B1(n10248), .B2(n7124), .A(n7123), .ZN(n10261) );
  NAND2_X1 U9421 ( .A1(n10516), .A2(n8234), .ZN(n7127) );
  NOR2_X1 U9422 ( .A1(n7128), .A2(n7126), .ZN(n7125) );
  INV_X1 U9423 ( .A(n8235), .ZN(n7126) );
  OAI21_X1 U9424 ( .B1(n8341), .B2(n7134), .A(n7131), .ZN(n8368) );
  OAI21_X1 U9425 ( .B1(n13421), .B2(n13485), .A(n7146), .ZN(n13501) );
  OAI21_X1 U9426 ( .B1(n13421), .B2(n7141), .A(n7139), .ZN(P2_U3495) );
  NAND2_X1 U9427 ( .A1(n13490), .A2(n8400), .ZN(n11662) );
  INV_X1 U9428 ( .A(n10112), .ZN(n10113) );
  NAND2_X1 U9429 ( .A1(n7150), .A2(n10112), .ZN(n7149) );
  NAND3_X1 U9430 ( .A1(n11691), .A2(n7151), .A3(n13843), .ZN(n14013) );
  NAND2_X1 U9431 ( .A1(n13574), .A2(n7156), .ZN(n7154) );
  INV_X1 U9432 ( .A(n13596), .ZN(n7160) );
  NAND2_X1 U9433 ( .A1(n7161), .A2(n12091), .ZN(n13596) );
  NAND2_X1 U9434 ( .A1(n13637), .A2(n13638), .ZN(n7161) );
  OAI21_X2 U9435 ( .B1(n11471), .B2(n7165), .A(n7163), .ZN(n12037) );
  NAND2_X1 U9436 ( .A1(n13677), .A2(n7175), .ZN(n7173) );
  NAND2_X1 U9437 ( .A1(n7173), .A2(n7174), .ZN(n12166) );
  NAND2_X1 U9438 ( .A1(n13645), .A2(n7177), .ZN(n14456) );
  XNOR2_X1 U9439 ( .A(n10574), .B(n10575), .ZN(n10341) );
  NOR2_X1 U9440 ( .A1(n10341), .A2(n7185), .ZN(n7184) );
  AND2_X2 U9441 ( .A1(n7187), .A2(n7186), .ZN(n10781) );
  NAND2_X1 U9442 ( .A1(n7184), .A2(n10339), .ZN(n7187) );
  INV_X1 U9443 ( .A(n7187), .ZN(n10573) );
  NAND2_X1 U9444 ( .A1(n7205), .A2(n7199), .ZN(n7204) );
  NAND3_X1 U9445 ( .A1(n7480), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n7481), .ZN(
        n7205) );
  NAND2_X1 U9446 ( .A1(n7206), .A2(n7200), .ZN(n7207) );
  AND2_X2 U9447 ( .A1(n7202), .A2(n7201), .ZN(n7887) );
  NAND4_X1 U9448 ( .A1(n7480), .A2(n7481), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7202) );
  NAND3_X1 U9449 ( .A1(n7208), .A2(n7209), .A3(n7211), .ZN(n7203) );
  INV_X1 U9450 ( .A(n10556), .ZN(n11893) );
  NAND2_X1 U9451 ( .A1(n10555), .A2(n10556), .ZN(n10554) );
  OAI21_X1 U9452 ( .B1(n11034), .B2(n7218), .A(n7216), .ZN(n10728) );
  NAND2_X1 U9453 ( .A1(n7215), .A2(n7214), .ZN(n10957) );
  NAND2_X1 U9454 ( .A1(n11034), .A2(n7216), .ZN(n7214) );
  NAND2_X1 U9455 ( .A1(n11080), .A2(n7221), .ZN(n7220) );
  NAND2_X1 U9456 ( .A1(n7226), .A2(n7224), .ZN(n7223) );
  INV_X1 U9457 ( .A(n10393), .ZN(n7224) );
  AND2_X2 U9458 ( .A1(n13917), .A2(n7237), .ZN(n13896) );
  NAND2_X2 U9459 ( .A1(n7478), .A2(n7477), .ZN(n14157) );
  NOR2_X2 U9460 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7483) );
  NAND2_X1 U9461 ( .A1(n9241), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U9462 ( .A1(n12187), .A2(n6625), .ZN(n7258) );
  OAI211_X1 U9463 ( .C1(n12187), .C2(n7263), .A(n7258), .B(n7259), .ZN(n12957)
         );
  NAND3_X1 U9464 ( .A1(n7273), .A2(n7272), .A3(n7271), .ZN(n7270) );
  NAND2_X1 U9465 ( .A1(n9461), .A2(n7281), .ZN(n7279) );
  OAI21_X2 U9466 ( .B1(n9437), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9003), .ZN(
        n9448) );
  OAI21_X2 U9467 ( .B1(n9391), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8995), .ZN(
        n9402) );
  NAND2_X1 U9468 ( .A1(n13391), .A2(n8589), .ZN(n7283) );
  NAND2_X1 U9469 ( .A1(n7288), .A2(n7286), .ZN(n10978) );
  NAND2_X1 U9470 ( .A1(n7292), .A2(n8561), .ZN(n10409) );
  NAND2_X1 U9471 ( .A1(n10307), .A2(n8904), .ZN(n7292) );
  NAND2_X1 U9472 ( .A1(n8571), .A2(n7295), .ZN(n11009) );
  INV_X1 U9473 ( .A(n7296), .ZN(n7295) );
  AOI21_X1 U9474 ( .B1(n10979), .B2(n7298), .A(n7297), .ZN(n7296) );
  NAND2_X1 U9475 ( .A1(n10979), .A2(n8569), .ZN(n10885) );
  NAND2_X1 U9476 ( .A1(n11009), .A2(n11006), .ZN(n8574) );
  NAND2_X1 U9477 ( .A1(n7310), .A2(n7309), .ZN(n11665) );
  NAND2_X1 U9478 ( .A1(n13075), .A2(n7321), .ZN(n7320) );
  OAI211_X1 U9479 ( .C1(n13075), .C2(n7325), .A(n7322), .B(n7320), .ZN(n12020)
         );
  CLKBUF_X1 U9480 ( .A(n7335), .Z(n7333) );
  NAND2_X1 U9481 ( .A1(n10158), .A2(n10159), .ZN(n10205) );
  OAI21_X1 U9482 ( .B1(n7347), .B2(n7346), .A(n11411), .ZN(n7345) );
  NAND3_X2 U9483 ( .A1(n8120), .A2(n8188), .A3(n7349), .ZN(n8294) );
  NAND3_X1 U9484 ( .A1(n8120), .A2(n8188), .A3(n8121), .ZN(n8266) );
  NOR2_X1 U9485 ( .A1(n8710), .A2(n8708), .ZN(n7361) );
  NAND2_X1 U9486 ( .A1(n8698), .A2(n7367), .ZN(n7366) );
  XNOR2_X1 U9487 ( .A(n9601), .B(n9602), .ZN(n14859) );
  AND2_X1 U9488 ( .A1(n7370), .A2(n6579), .ZN(n14860) );
  AND2_X1 U9489 ( .A1(n14859), .A2(n6579), .ZN(n7371) );
  NAND3_X1 U9490 ( .A1(n7373), .A2(n9658), .A3(n12729), .ZN(n12284) );
  NAND2_X1 U9491 ( .A1(n7376), .A2(n7374), .ZN(n12220) );
  NAND2_X1 U9492 ( .A1(n12240), .A2(n7380), .ZN(n7379) );
  NAND2_X1 U9493 ( .A1(n7384), .A2(n12264), .ZN(n9668) );
  NAND2_X1 U9494 ( .A1(n11364), .A2(n6589), .ZN(n11573) );
  NOR2_X2 U9495 ( .A1(n9053), .A2(n7392), .ZN(n9093) );
  NAND2_X1 U9496 ( .A1(n7397), .A2(n6542), .ZN(n7403) );
  NAND2_X1 U9497 ( .A1(n15308), .A2(n7398), .ZN(n7397) );
  NAND2_X1 U9498 ( .A1(n11770), .A2(n11769), .ZN(n7398) );
  NAND2_X1 U9500 ( .A1(n7403), .A2(n7400), .ZN(n11791) );
  NAND2_X1 U9501 ( .A1(n7412), .A2(n7494), .ZN(n13723) );
  AOI21_X1 U9502 ( .B1(n13723), .B2(n12148), .A(n7409), .ZN(n10107) );
  NAND3_X1 U9503 ( .A1(n11838), .A2(n11837), .A3(n6606), .ZN(n7415) );
  INV_X1 U9504 ( .A(n11840), .ZN(n7416) );
  NAND2_X1 U9505 ( .A1(n7417), .A2(n7418), .ZN(n11762) );
  NAND3_X1 U9506 ( .A1(n11756), .A2(n6598), .A3(n11755), .ZN(n7417) );
  NAND2_X1 U9507 ( .A1(n7420), .A2(n6600), .ZN(n11742) );
  NAND3_X1 U9508 ( .A1(n11733), .A2(n6602), .A3(n11732), .ZN(n7420) );
  NAND2_X1 U9509 ( .A1(n7422), .A2(n7423), .ZN(n11728) );
  NAND3_X1 U9510 ( .A1(n11720), .A2(n11719), .A3(n6592), .ZN(n7422) );
  NAND3_X1 U9511 ( .A1(n11810), .A2(n11809), .A3(n6605), .ZN(n7425) );
  INV_X1 U9512 ( .A(n11946), .ZN(n14077) );
  OAI21_X1 U9513 ( .B1(n14078), .B2(n14025), .A(n11945), .ZN(n11946) );
  NAND2_X1 U9514 ( .A1(n14154), .A2(n7468), .ZN(n7517) );
  OR2_X2 U9515 ( .A1(n13293), .A2(n8600), .ZN(n8495) );
  OR2_X1 U9516 ( .A1(n9746), .A2(n9856), .ZN(n7487) );
  CLKBUF_X1 U9517 ( .A(n10881), .Z(n10883) );
  CLKBUF_X1 U9518 ( .A(n10776), .Z(n10937) );
  NAND2_X1 U9519 ( .A1(n9153), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9138) );
  NAND2_X4 U9520 ( .A1(n9930), .A2(n11689), .ZN(n12158) );
  INV_X1 U9521 ( .A(n8648), .ZN(n8133) );
  INV_X1 U9522 ( .A(n11511), .ZN(n7766) );
  NAND2_X1 U9523 ( .A1(n8139), .A2(n8149), .ZN(n8648) );
  OR3_X1 U9524 ( .A1(n8139), .A2(n8154), .A3(n8149), .ZN(n8132) );
  OR2_X1 U9525 ( .A1(n8545), .A2(n10283), .ZN(n8164) );
  INV_X1 U9526 ( .A(n10480), .ZN(n8653) );
  INV_X1 U9527 ( .A(n8552), .ZN(n8148) );
  OAI21_X1 U9528 ( .B1(n10334), .B2(n10565), .A(n9934), .ZN(n9935) );
  AND2_X1 U9529 ( .A1(n6513), .A2(n8403), .ZN(n13177) );
  CLKBUF_X1 U9530 ( .A(n8612), .Z(n9873) );
  NAND2_X1 U9531 ( .A1(n11890), .A2(n11878), .ZN(n11696) );
  OAI22_X2 U9532 ( .A1(n13004), .A2(n13003), .B1(n12000), .B2(n11999), .ZN(
        n13075) );
  NAND2_X1 U9533 ( .A1(n12284), .A2(n9658), .ZN(n9663) );
  INV_X1 U9534 ( .A(n12363), .ZN(n10657) );
  NOR2_X2 U9535 ( .A1(n12555), .A2(n11678), .ZN(n15030) );
  OAI22_X2 U9536 ( .A1(n13373), .A2(n8439), .B1(n13532), .B2(n8592), .ZN(
        n13356) );
  INV_X1 U9537 ( .A(n13879), .ZN(n13907) );
  INV_X1 U9538 ( .A(n12447), .ZN(n9266) );
  INV_X1 U9539 ( .A(n11910), .ZN(n11512) );
  NAND2_X1 U9540 ( .A1(n10939), .A2(n10938), .ZN(n7434) );
  INV_X1 U9541 ( .A(n12898), .ZN(n9554) );
  OR3_X1 U9542 ( .A1(n10048), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n7435) );
  AND2_X1 U9543 ( .A1(n11636), .A2(n11635), .ZN(n7436) );
  OR2_X1 U9544 ( .A1(n7843), .A2(n10259), .ZN(n7438) );
  AND2_X1 U9545 ( .A1(n11965), .A2(n11964), .ZN(n7439) );
  AND2_X1 U9546 ( .A1(n11923), .A2(n11875), .ZN(n7440) );
  OR2_X1 U9547 ( .A1(n14068), .A2(n14019), .ZN(n7441) );
  OR2_X1 U9548 ( .A1(n12637), .A2(n12898), .ZN(n7442) );
  OR2_X1 U9549 ( .A1(n12637), .A2(n12952), .ZN(n7443) );
  OR2_X1 U9550 ( .A1(n13860), .A2(n13859), .ZN(n7444) );
  NOR2_X1 U9551 ( .A1(n9557), .A2(n12952), .ZN(n9086) );
  INV_X1 U9552 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9015) );
  INV_X1 U9553 ( .A(n7513), .ZN(n7571) );
  AND2_X1 U9554 ( .A1(n7706), .A2(n7692), .ZN(n7446) );
  AND2_X1 U9555 ( .A1(n12549), .A2(n10947), .ZN(n7447) );
  OR2_X1 U9556 ( .A1(n9868), .A2(n10004), .ZN(n7448) );
  INV_X1 U9557 ( .A(n12538), .ZN(n12729) );
  NAND2_X2 U9558 ( .A1(n8109), .A2(n14011), .ZN(n14047) );
  XNOR2_X1 U9559 ( .A(n12620), .B(n12619), .ZN(n7449) );
  OR2_X2 U9560 ( .A1(n12793), .A2(n12802), .ZN(n7450) );
  INV_X1 U9561 ( .A(n6490), .ZN(n9044) );
  OR2_X1 U9562 ( .A1(n7880), .A2(SI_20_), .ZN(n7451) );
  NAND2_X1 U9563 ( .A1(n8890), .A2(n8610), .ZN(n14399) );
  OR2_X1 U9564 ( .A1(n7883), .A2(SI_21_), .ZN(n7453) );
  INV_X1 U9565 ( .A(n13531), .ZN(n8940) );
  INV_X1 U9566 ( .A(n14842), .ZN(n8665) );
  AND2_X1 U9567 ( .A1(n11346), .A2(n11345), .ZN(n7454) );
  INV_X1 U9568 ( .A(n13887), .ZN(n7977) );
  INV_X1 U9569 ( .A(n8671), .ZN(n8672) );
  INV_X1 U9570 ( .A(n8685), .ZN(n8686) );
  NOR2_X1 U9571 ( .A1(n13722), .A2(n11839), .ZN(n11701) );
  OAI21_X1 U9572 ( .B1(n11718), .B2(n11717), .A(n11716), .ZN(n11720) );
  AND2_X1 U9573 ( .A1(n11784), .A2(n11774), .ZN(n11781) );
  INV_X1 U9574 ( .A(n8809), .ZN(n8810) );
  NAND2_X1 U9575 ( .A1(n12398), .A2(n10515), .ZN(n9583) );
  NAND2_X1 U9576 ( .A1(n10866), .A2(n12364), .ZN(n10867) );
  INV_X1 U9577 ( .A(n11902), .ZN(n8071) );
  OAI21_X1 U9578 ( .B1(n9585), .B2(n9584), .A(n9583), .ZN(n9586) );
  INV_X1 U9579 ( .A(n11576), .ZN(n9616) );
  AOI21_X1 U9580 ( .B1(n12613), .B2(n12612), .A(n14334), .ZN(n12615) );
  INV_X1 U9581 ( .A(n10867), .ZN(n10868) );
  NAND2_X1 U9582 ( .A1(n6476), .A2(n9504), .ZN(n10941) );
  XNOR2_X1 U9583 ( .A(n12553), .B(n10905), .ZN(n12363) );
  INV_X1 U9584 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8975) );
  AND2_X1 U9585 ( .A1(n8498), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8509) );
  AND2_X1 U9586 ( .A1(n8509), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8522) );
  INV_X1 U9587 ( .A(n8911), .ZN(n8585) );
  NOR2_X1 U9588 ( .A1(n8287), .A2(n11108), .ZN(n8298) );
  INV_X1 U9589 ( .A(n13595), .ZN(n12097) );
  INV_X1 U9590 ( .A(n13938), .ZN(n7908) );
  NAND2_X1 U9591 ( .A1(n7854), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7873) );
  INV_X1 U9592 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7480) );
  OAI21_X1 U9593 ( .B1(n7511), .B2(n7510), .A(n6546), .ZN(n7512) );
  NOR2_X1 U9594 ( .A1(n14209), .A2(n14208), .ZN(n14195) );
  INV_X1 U9595 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15195) );
  OR2_X1 U9596 ( .A1(n9317), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9336) );
  AND2_X1 U9597 ( .A1(n9203), .A2(n9202), .ZN(n9234) );
  OR2_X1 U9598 ( .A1(n9475), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U9599 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  INV_X1 U9600 ( .A(n12607), .ZN(n12608) );
  OR2_X1 U9601 ( .A1(n12506), .A2(n12678), .ZN(n9523) );
  OR2_X1 U9602 ( .A1(n14364), .A2(n12830), .ZN(n12466) );
  XNOR2_X1 U9603 ( .A(n10689), .B(n12009), .ZN(n10148) );
  NOR2_X1 U9604 ( .A1(n8407), .A2(n8406), .ZN(n8431) );
  OAI21_X1 U9605 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8888) );
  AND2_X1 U9606 ( .A1(n8431), .A2(n8430), .ZN(n8442) );
  OR2_X1 U9607 ( .A1(n8350), .A2(n11442), .ZN(n8361) );
  AND2_X1 U9608 ( .A1(n8522), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8534) );
  OR2_X1 U9609 ( .A1(n8272), .A2(n8271), .ZN(n8287) );
  OAI22_X1 U9610 ( .A1(n12971), .A2(n13078), .B1(n13204), .B2(n8619), .ZN(
        n8620) );
  INV_X1 U9611 ( .A(n11613), .ZN(n8384) );
  INV_X1 U9612 ( .A(n11619), .ZN(n14413) );
  INV_X1 U9613 ( .A(n10033), .ZN(n8661) );
  NAND2_X1 U9614 ( .A1(n7903), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7917) );
  INV_X1 U9615 ( .A(n13702), .ZN(n12160) );
  INV_X1 U9616 ( .A(n12034), .ZN(n12035) );
  NAND2_X1 U9617 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n7918), .ZN(n7937) );
  NAND2_X1 U9618 ( .A1(n7890), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U9619 ( .A1(n7874), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U9620 ( .A1(n11456), .A2(n13700), .ZN(n11513) );
  OR2_X1 U9621 ( .A1(n7622), .A2(n7621), .ZN(n7639) );
  INV_X1 U9622 ( .A(n11713), .ZN(n11715) );
  OR2_X1 U9623 ( .A1(n14167), .A2(P1_B_REG_SCAN_IN), .ZN(n8022) );
  NAND2_X1 U9624 ( .A1(n7829), .A2(SI_19_), .ZN(n7847) );
  NAND2_X1 U9625 ( .A1(n7671), .A2(n15213), .ZN(n7687) );
  INV_X1 U9626 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15192) );
  OR2_X1 U9627 ( .A1(n9427), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U9628 ( .A1(n9369), .A2(n9368), .ZN(n9395) );
  OR2_X1 U9629 ( .A1(n9395), .A2(n9394), .ZN(n9405) );
  INV_X1 U9630 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15219) );
  AND2_X1 U9631 ( .A1(n9167), .A2(n9166), .ZN(n9181) );
  INV_X1 U9632 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14173) );
  INV_X1 U9633 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15191) );
  AND2_X1 U9634 ( .A1(n10044), .A2(n10072), .ZN(n10066) );
  AND2_X1 U9635 ( .A1(n9151), .A2(n15191), .ZN(n9167) );
  NOR2_X1 U9636 ( .A1(n9683), .A2(n15068), .ZN(n9685) );
  INV_X1 U9637 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9087) );
  INV_X1 U9638 ( .A(n14848), .ZN(n11304) );
  INV_X1 U9639 ( .A(n15054), .ZN(n14372) );
  NAND2_X1 U9640 ( .A1(n9057), .A2(n9084), .ZN(n9060) );
  NAND2_X1 U9641 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  AND2_X1 U9642 ( .A1(n8952), .A2(n8951), .ZN(n9130) );
  INV_X1 U9643 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11566) );
  INV_X1 U9644 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U9645 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  INV_X1 U9646 ( .A(n11438), .ZN(n11439) );
  OR2_X1 U9647 ( .A1(n11075), .A2(n8148), .ZN(n9958) );
  AND2_X1 U9648 ( .A1(n8442), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8453) );
  NOR2_X1 U9649 ( .A1(n13400), .A2(n13383), .ZN(n13381) );
  OR2_X1 U9650 ( .A1(n14420), .A2(n6641), .ZN(n14415) );
  NAND2_X1 U9651 ( .A1(n8841), .A2(n8840), .ZN(n8883) );
  NAND2_X1 U9652 ( .A1(n8661), .A2(n8933), .ZN(n14828) );
  XNOR2_X1 U9653 ( .A(n13127), .B(n8204), .ZN(n10306) );
  INV_X1 U9654 ( .A(n14399), .ZN(n13393) );
  AOI21_X1 U9655 ( .B1(n14754), .B2(n8656), .A(n8655), .ZN(n9947) );
  NAND2_X1 U9656 ( .A1(n11052), .A2(n11051), .ZN(n11053) );
  INV_X1 U9657 ( .A(n13673), .ZN(n14477) );
  AND2_X1 U9658 ( .A1(n7839), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7854) );
  INV_X1 U9659 ( .A(n7517), .ZN(n7498) );
  INV_X1 U9660 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11354) );
  OR2_X1 U9661 ( .A1(n10188), .A2(n10189), .ZN(n14554) );
  OR2_X1 U9662 ( .A1(n10591), .A2(n10592), .ZN(n11528) );
  OR2_X1 U9663 ( .A1(n13830), .A2(n11538), .ZN(n11540) );
  AOI21_X1 U9664 ( .B1(n14063), .B2(n13999), .A(n8113), .ZN(n8114) );
  NAND2_X1 U9665 ( .A1(n13879), .A2(n13892), .ZN(n13880) );
  OR2_X1 U9666 ( .A1(n10134), .A2(n11688), .ZN(n14025) );
  INV_X1 U9667 ( .A(n11908), .ZN(n11594) );
  NAND2_X1 U9668 ( .A1(n8035), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8037) );
  OR2_X1 U9669 ( .A1(n7779), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n7799) );
  INV_X1 U9670 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14224) );
  OAI21_X1 U9671 ( .B1(n12911), .B2(n14856), .A(n9702), .ZN(n9703) );
  INV_X1 U9672 ( .A(n12276), .ZN(n12315) );
  AND4_X1 U9673 ( .A1(n12345), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(n12348)
         );
  AND4_X1 U9674 ( .A1(n9459), .A2(n9458), .A3(n9457), .A4(n9456), .ZN(n12669)
         );
  AND4_X1 U9675 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n12277)
         );
  AND4_X1 U9676 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(n12254)
         );
  INV_X1 U9677 ( .A(n15003), .ZN(n15022) );
  INV_X1 U9678 ( .A(n15018), .ZN(n14944) );
  NAND2_X1 U9679 ( .A1(n9526), .A2(n9525), .ZN(n12832) );
  AND2_X1 U9680 ( .A1(n15045), .A2(n15044), .ZN(n12841) );
  NAND2_X1 U9681 ( .A1(n9685), .A2(n15034), .ZN(n15032) );
  AND2_X1 U9682 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  AND2_X1 U9683 ( .A1(n15034), .A2(n9543), .ZN(n15072) );
  AND2_X1 U9684 ( .A1(n12955), .A2(n9709), .ZN(n10043) );
  OR2_X1 U9685 ( .A1(n9060), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9059) );
  AND2_X1 U9686 ( .A1(n8970), .A2(n8969), .ZN(n9221) );
  INV_X1 U9687 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9161) );
  INV_X1 U9688 ( .A(n13076), .ZN(n13065) );
  INV_X1 U9689 ( .A(n13087), .ZN(n13068) );
  NOR2_X1 U9690 ( .A1(n9949), .A2(n14788), .ZN(n9960) );
  AND3_X1 U9691 ( .A1(n8848), .A2(n8847), .A3(n8846), .ZN(n13203) );
  OR2_X1 U9692 ( .A1(n9886), .A2(n9885), .ZN(n14668) );
  OR2_X1 U9693 ( .A1(n10224), .A2(n10223), .ZN(n10290) );
  INV_X1 U9694 ( .A(n14668), .ZN(n14743) );
  OR2_X1 U9695 ( .A1(n13227), .A2(n13233), .ZN(n13228) );
  INV_X1 U9696 ( .A(n8917), .ZN(n13323) );
  INV_X1 U9697 ( .A(n8913), .ZN(n11664) );
  INV_X1 U9698 ( .A(n13406), .ZN(n14403) );
  INV_X1 U9699 ( .A(n14415), .ZN(n13402) );
  INV_X1 U9700 ( .A(n14828), .ZN(n14819) );
  AND2_X1 U9701 ( .A1(n14409), .A2(n14408), .ZN(n14433) );
  INV_X1 U9702 ( .A(n13485), .ZN(n14816) );
  NOR2_X1 U9703 ( .A1(n10276), .A2(n9953), .ZN(n8939) );
  AND2_X1 U9704 ( .A1(n8645), .A2(n8644), .ZN(n14754) );
  AND2_X1 U9705 ( .A1(n9867), .A2(n9706), .ZN(n9951) );
  AND2_X1 U9706 ( .A1(n8328), .A2(n8342), .ZN(n13144) );
  NOR2_X1 U9707 ( .A1(n9941), .A2(n11931), .ZN(n13658) );
  OR2_X1 U9708 ( .A1(n8003), .A2(n13871), .ZN(n7990) );
  AND4_X1 U9709 ( .A1(n7907), .A2(n7906), .A3(n7905), .A4(n7904), .ZN(n13657)
         );
  AND2_X1 U9710 ( .A1(n7862), .A2(n7861), .ZN(n13598) );
  AND4_X1 U9711 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), .ZN(n7739)
         );
  AND2_X1 U9712 ( .A1(n14556), .A2(n10328), .ZN(n10330) );
  INV_X1 U9713 ( .A(n11530), .ZN(n14574) );
  INV_X1 U9714 ( .A(n11539), .ZN(n14575) );
  INV_X1 U9715 ( .A(n14579), .ZN(n14560) );
  INV_X1 U9716 ( .A(n14021), .ZN(n14006) );
  AND2_X1 U9717 ( .A1(n8101), .A2(n13843), .ZN(n13999) );
  AND2_X1 U9718 ( .A1(n8029), .A2(n8028), .ZN(n10130) );
  AND2_X1 U9719 ( .A1(n14025), .A2(n14130), .ZN(n14583) );
  INV_X1 U9720 ( .A(n14583), .ZN(n14638) );
  AND2_X1 U9721 ( .A1(n7780), .A2(n7799), .ZN(n11534) );
  AND2_X1 U9722 ( .A1(n7555), .A2(n7573), .ZN(n13762) );
  AND2_X1 U9723 ( .A1(n14249), .A2(n14250), .ZN(n14525) );
  AND2_X1 U9724 ( .A1(n10073), .A2(n10072), .ZN(n15021) );
  AND2_X1 U9725 ( .A1(n10613), .A2(n12531), .ZN(n14867) );
  NAND2_X1 U9726 ( .A1(n9681), .A2(n10043), .ZN(n12310) );
  INV_X1 U9727 ( .A(n14847), .ZN(n14856) );
  AND4_X1 U9728 ( .A1(n9493), .A2(n9492), .A3(n9491), .A4(n9490), .ZN(n12655)
         );
  INV_X1 U9729 ( .A(n12254), .ZN(n12830) );
  INV_X1 U9730 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14954) );
  INV_X1 U9731 ( .A(n14355), .ZN(n15028) );
  OR2_X1 U9732 ( .A1(n10810), .A2(n10904), .ZN(n12807) );
  INV_X1 U9733 ( .A(n12900), .ZN(n12846) );
  NAND2_X1 U9734 ( .A1(n15085), .A2(n14383), .ZN(n12898) );
  AND2_X2 U9735 ( .A1(n10809), .A2(n9551), .ZN(n15085) );
  NAND2_X1 U9736 ( .A1(n9552), .A2(n15076), .ZN(n9538) );
  INV_X1 U9737 ( .A(n9653), .ZN(n12931) );
  NAND2_X1 U9738 ( .A1(n9085), .A2(n10043), .ZN(n15074) );
  NAND2_X1 U9739 ( .A1(n9060), .A2(n12955), .ZN(n9968) );
  INV_X1 U9740 ( .A(SI_18_), .ZN(n10259) );
  INV_X1 U9741 ( .A(SI_13_), .ZN(n15175) );
  INV_X1 U9742 ( .A(n10931), .ZN(n12967) );
  AND2_X1 U9743 ( .A1(n9707), .A2(n9867), .ZN(n9866) );
  INV_X1 U9744 ( .A(n13085), .ZN(n13066) );
  INV_X1 U9745 ( .A(n12013), .ZN(n13100) );
  INV_X1 U9746 ( .A(P2_U3947), .ZN(n13121) );
  INV_X1 U9747 ( .A(n14741), .ZN(n14694) );
  OR2_X1 U9748 ( .A1(n9874), .A2(P2_U3088), .ZN(n14752) );
  INV_X1 U9749 ( .A(n13336), .ZN(n14420) );
  OR2_X1 U9750 ( .A1(n14420), .A2(n10476), .ZN(n13372) );
  INV_X1 U9751 ( .A(n13336), .ZN(n13411) );
  NAND2_X1 U9752 ( .A1(n14842), .A2(n14819), .ZN(n13474) );
  AND2_X2 U9753 ( .A1(n8660), .A2(n8939), .ZN(n14842) );
  NAND2_X1 U9754 ( .A1(n14836), .A2(n14819), .ZN(n13531) );
  AND2_X1 U9755 ( .A1(n14444), .A2(n14443), .ZN(n14451) );
  AND2_X2 U9756 ( .A1(n10277), .A2(n8939), .ZN(n14836) );
  NOR2_X1 U9757 ( .A1(n14754), .A2(n14788), .ZN(n14769) );
  INV_X1 U9758 ( .A(n14791), .ZN(n14788) );
  INV_X1 U9759 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11174) );
  INV_X1 U9760 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10389) );
  INV_X1 U9761 ( .A(n11757), .ZN(n14635) );
  NAND2_X1 U9762 ( .A1(n9940), .A2(n9939), .ZN(n14467) );
  INV_X1 U9763 ( .A(n12040), .ZN(n13655) );
  INV_X1 U9764 ( .A(n14490), .ZN(n13699) );
  NAND4_X1 U9765 ( .A1(n7975), .A2(n7974), .A3(n7973), .A4(n7972), .ZN(n13887)
         );
  INV_X1 U9766 ( .A(n13656), .ZN(n13983) );
  INV_X1 U9767 ( .A(n7739), .ZN(n13710) );
  NOR2_X2 U9768 ( .A1(n9931), .A2(n9708), .ZN(n13728) );
  OR2_X1 U9769 ( .A1(n14550), .A2(n14546), .ZN(n11539) );
  INV_X1 U9770 ( .A(n14570), .ZN(n14566) );
  NAND2_X1 U9771 ( .A1(n14047), .A2(n8058), .ZN(n14019) );
  INV_X1 U9772 ( .A(n14654), .ZN(n14651) );
  NAND2_X1 U9773 ( .A1(n10144), .A2(n10143), .ZN(n14639) );
  AND2_X1 U9774 ( .A1(n9743), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9730) );
  INV_X1 U9775 ( .A(n11687), .ZN(n14168) );
  INV_X1 U9776 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10421) );
  INV_X1 U9777 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9967) );
  AND2_X1 U9778 ( .A1(n12955), .A2(n9710), .ZN(P3_U3897) );
  NAND2_X1 U9779 ( .A1(n9539), .A2(n9538), .ZN(P3_U3455) );
  AND2_X1 U9780 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9866), .ZN(P2_U3947) );
  NAND2_X1 U9781 ( .A1(n7441), .A2(n8116), .ZN(P1_U3356) );
  NOR2_X1 U9782 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n7457) );
  NOR2_X1 U9783 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7456) );
  AND2_X1 U9784 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  AND2_X2 U9785 ( .A1(n7505), .A2(n7458), .ZN(n7604) );
  NOR2_X1 U9786 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n7461) );
  NOR2_X1 U9787 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7460) );
  NOR2_X1 U9788 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7462) );
  AND2_X4 U9789 ( .A1(n7466), .A2(n14154), .ZN(n7538) );
  AND2_X4 U9790 ( .A1(n7467), .A2(n7468), .ZN(n8004) );
  NAND2_X1 U9791 ( .A1(n8004), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7471) );
  INV_X1 U9792 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U9793 ( .A1(n7498), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7469) );
  MUX2_X1 U9794 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7475), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n7478) );
  INV_X1 U9795 ( .A(n7476), .ZN(n7477) );
  NAND2_X1 U9796 ( .A1(n9746), .A2(n7495), .ZN(n7513) );
  XNOR2_X1 U9797 ( .A(n7511), .B(n7510), .ZN(n9760) );
  NAND2_X1 U9798 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7482) );
  MUX2_X1 U9799 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7482), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7486) );
  INV_X1 U9800 ( .A(n7484), .ZN(n7485) );
  NAND2_X1 U9801 ( .A1(n7486), .A2(n7485), .ZN(n9856) );
  NAND2_X1 U9802 ( .A1(n7498), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7491) );
  INV_X1 U9803 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7489) );
  NAND2_X1 U9804 ( .A1(n7538), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U9805 ( .A1(n8004), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7492) );
  INV_X1 U9806 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14547) );
  INV_X1 U9807 ( .A(SI_0_), .ZN(n9758) );
  NOR2_X1 U9808 ( .A1(n9735), .A2(n9758), .ZN(n7496) );
  XNOR2_X1 U9809 ( .A(n7496), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14170) );
  NAND2_X1 U9810 ( .A1(n13723), .A2(n7408), .ZN(n10555) );
  INV_X1 U9811 ( .A(n11700), .ZN(n14590) );
  NAND2_X1 U9812 ( .A1(n14046), .A2(n14590), .ZN(n7497) );
  INV_X1 U9813 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13730) );
  OR2_X1 U9814 ( .A1(n7540), .A2(n13730), .ZN(n7502) );
  NAND2_X1 U9815 ( .A1(n7498), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7501) );
  NAND2_X1 U9816 ( .A1(n8004), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7500) );
  NOR2_X1 U9817 ( .A1(n7484), .A2(n7588), .ZN(n7503) );
  MUX2_X1 U9818 ( .A(n7588), .B(n7503), .S(P1_IR_REG_2__SCAN_IN), .Z(n7504) );
  INV_X1 U9819 ( .A(n7504), .ZN(n7508) );
  INV_X1 U9820 ( .A(n7506), .ZN(n7507) );
  NAND2_X1 U9821 ( .A1(n7508), .A2(n7507), .ZN(n9795) );
  INV_X1 U9822 ( .A(SI_1_), .ZN(n9712) );
  INV_X1 U9823 ( .A(n7512), .ZN(n7527) );
  XNOR2_X1 U9824 ( .A(n7527), .B(SI_2_), .ZN(n7526) );
  INV_X1 U9825 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9741) );
  MUX2_X1 U9826 ( .A(n9741), .B(n9721), .S(n7777), .Z(n7524) );
  XNOR2_X1 U9827 ( .A(n7526), .B(n7524), .ZN(n9720) );
  NAND2_X1 U9828 ( .A1(n9720), .A2(n7571), .ZN(n7515) );
  NAND2_X1 U9829 ( .A1(n7531), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7514) );
  INV_X1 U9830 ( .A(n11891), .ZN(n10132) );
  NAND2_X1 U9831 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  INV_X1 U9832 ( .A(n13721), .ZN(n10566) );
  INV_X1 U9833 ( .A(n7516), .ZN(n10425) );
  NAND2_X1 U9834 ( .A1(n10566), .A2(n10425), .ZN(n11706) );
  NAND2_X1 U9835 ( .A1(n10131), .A2(n11706), .ZN(n10350) );
  INV_X1 U9836 ( .A(n7517), .ZN(n7984) );
  NAND2_X1 U9837 ( .A1(n7984), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7523) );
  OR2_X1 U9838 ( .A1(n7540), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7522) );
  INV_X1 U9839 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7518) );
  INV_X1 U9840 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7519) );
  INV_X1 U9841 ( .A(n7524), .ZN(n7525) );
  NAND2_X1 U9842 ( .A1(n7526), .A2(n7525), .ZN(n7530) );
  INV_X1 U9843 ( .A(n7527), .ZN(n7528) );
  NAND2_X1 U9844 ( .A1(n7528), .A2(SI_2_), .ZN(n7529) );
  XNOR2_X1 U9845 ( .A(n7548), .B(n7546), .ZN(n9724) );
  NAND2_X1 U9846 ( .A1(n9724), .A2(n7571), .ZN(n7536) );
  BUF_X4 U9847 ( .A(n7531), .Z(n8000) );
  NOR2_X1 U9848 ( .A1(n7506), .A2(n7588), .ZN(n7532) );
  MUX2_X1 U9849 ( .A(n7588), .B(n7532), .S(P1_IR_REG_3__SCAN_IN), .Z(n7534) );
  INV_X1 U9850 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7533) );
  AND2_X1 U9851 ( .A1(n7506), .A2(n7533), .ZN(n7552) );
  NOR2_X1 U9852 ( .A1(n7534), .A2(n7552), .ZN(n13750) );
  AOI22_X1 U9853 ( .A1(n7531), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6487), .B2(
        n13750), .ZN(n7535) );
  NAND2_X1 U9854 ( .A1(n7538), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7545) );
  INV_X1 U9855 ( .A(n7984), .ZN(n11854) );
  INV_X1 U9856 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7539) );
  OR2_X1 U9857 ( .A1(n11854), .A2(n7539), .ZN(n7544) );
  NAND2_X1 U9858 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7559) );
  OAI21_X1 U9859 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7559), .ZN(n10583) );
  OR2_X1 U9860 ( .A1(n8003), .A2(n10583), .ZN(n7543) );
  INV_X1 U9861 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7541) );
  OR2_X1 U9862 ( .A1(n7561), .A2(n7541), .ZN(n7542) );
  NAND2_X1 U9863 ( .A1(n7548), .A2(n7547), .ZN(n7551) );
  NAND2_X1 U9864 ( .A1(n7549), .A2(SI_3_), .ZN(n7550) );
  MUX2_X1 U9865 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7777), .Z(n7569) );
  XNOR2_X1 U9866 ( .A(n7569), .B(SI_4_), .ZN(n7566) );
  XNOR2_X1 U9867 ( .A(n7568), .B(n7566), .ZN(n9722) );
  NAND2_X1 U9868 ( .A1(n9722), .A2(n7965), .ZN(n7557) );
  INV_X1 U9869 ( .A(n7552), .ZN(n7554) );
  NAND2_X1 U9870 ( .A1(n7554), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7553) );
  MUX2_X1 U9871 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7553), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7555) );
  AOI22_X1 U9872 ( .A1(n8000), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7836), .B2(
        n13762), .ZN(n7556) );
  OR2_X1 U9873 ( .A1(n13720), .A2(n11715), .ZN(n10392) );
  INV_X1 U9874 ( .A(n10392), .ZN(n7558) );
  NAND2_X1 U9875 ( .A1(n11715), .A2(n13720), .ZN(n10391) );
  NAND2_X1 U9876 ( .A1(n7538), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7565) );
  INV_X1 U9877 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10797) );
  AND2_X1 U9878 ( .A1(n7559), .A2(n10797), .ZN(n7560) );
  NOR2_X1 U9879 ( .A1(n7559), .A2(n10797), .ZN(n7593) );
  OR2_X1 U9880 ( .A1(n7560), .A2(n7593), .ZN(n10796) );
  OR2_X1 U9881 ( .A1(n8003), .A2(n10796), .ZN(n7564) );
  INV_X1 U9882 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9805) );
  OR2_X1 U9883 ( .A1(n6472), .A2(n9805), .ZN(n7563) );
  NAND2_X1 U9884 ( .A1(n7984), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7562) );
  NAND4_X1 U9885 ( .A1(n7565), .A2(n7564), .A3(n7563), .A4(n7562), .ZN(n13719)
         );
  INV_X1 U9886 ( .A(n13719), .ZN(n10580) );
  INV_X1 U9887 ( .A(n7566), .ZN(n7567) );
  NAND2_X1 U9888 ( .A1(n7569), .A2(SI_4_), .ZN(n7570) );
  MUX2_X1 U9889 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7777), .Z(n7585) );
  XNOR2_X1 U9890 ( .A(n7585), .B(SI_5_), .ZN(n7582) );
  XNOR2_X1 U9891 ( .A(n7584), .B(n7582), .ZN(n9726) );
  NAND2_X1 U9892 ( .A1(n9726), .A2(n7571), .ZN(n7579) );
  NAND2_X1 U9893 ( .A1(n7573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7572) );
  MUX2_X1 U9894 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7572), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7576) );
  INV_X1 U9895 ( .A(n7573), .ZN(n7575) );
  INV_X1 U9896 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U9897 ( .A1(n7575), .A2(n7574), .ZN(n7589) );
  NAND2_X1 U9898 ( .A1(n7576), .A2(n7589), .ZN(n9816) );
  INV_X1 U9899 ( .A(n9816), .ZN(n7577) );
  AOI22_X1 U9900 ( .A1(n8000), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7836), .B2(
        n7577), .ZN(n7578) );
  NAND2_X1 U9901 ( .A1(n7579), .A2(n7578), .ZN(n11721) );
  XNOR2_X1 U9902 ( .A(n10580), .B(n11721), .ZN(n11895) );
  INV_X1 U9903 ( .A(n11895), .ZN(n7580) );
  OR2_X1 U9904 ( .A1(n11721), .A2(n13719), .ZN(n7581) );
  INV_X1 U9905 ( .A(n7582), .ZN(n7583) );
  NAND2_X1 U9906 ( .A1(n7585), .A2(SI_5_), .ZN(n7586) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7777), .Z(n7602) );
  XNOR2_X1 U9908 ( .A(n7602), .B(SI_6_), .ZN(n7599) );
  XNOR2_X1 U9909 ( .A(n7601), .B(n7599), .ZN(n9749) );
  NAND2_X1 U9910 ( .A1(n9749), .A2(n7965), .ZN(n7592) );
  NAND2_X1 U9911 ( .A1(n7589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7590) );
  XNOR2_X1 U9912 ( .A(n7590), .B(P1_IR_REG_6__SCAN_IN), .ZN(n13778) );
  AOI22_X1 U9913 ( .A1(n8000), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7836), .B2(
        n13778), .ZN(n7591) );
  NAND2_X1 U9914 ( .A1(n7592), .A2(n7591), .ZN(n11725) );
  NAND2_X1 U9915 ( .A1(n7538), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U9916 ( .A1(n7593), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7622) );
  OR2_X1 U9917 ( .A1(n7593), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9918 ( .A1(n7622), .A2(n7594), .ZN(n10899) );
  OR2_X1 U9919 ( .A1(n8003), .A2(n10899), .ZN(n7596) );
  NAND2_X1 U9920 ( .A1(n8004), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7595) );
  XNOR2_X1 U9921 ( .A(n11725), .B(n13718), .ZN(n11897) );
  INV_X1 U9922 ( .A(n11897), .ZN(n10640) );
  OR2_X1 U9923 ( .A1(n11725), .A2(n13718), .ZN(n7598) );
  INV_X1 U9924 ( .A(n7599), .ZN(n7600) );
  NAND2_X1 U9925 ( .A1(n7602), .A2(SI_6_), .ZN(n7603) );
  MUX2_X1 U9926 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7777), .Z(n7616) );
  XNOR2_X1 U9927 ( .A(n7616), .B(SI_7_), .ZN(n7613) );
  NAND2_X1 U9928 ( .A1(n9764), .A2(n7965), .ZN(n7607) );
  OR2_X1 U9929 ( .A1(n7604), .A2(n7588), .ZN(n7605) );
  XNOR2_X1 U9930 ( .A(n7605), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U9931 ( .A1(n8000), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7836), .B2(
        n9818), .ZN(n7606) );
  NAND2_X1 U9932 ( .A1(n7984), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U9933 ( .A1(n8004), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7610) );
  INV_X1 U9934 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7620) );
  XNOR2_X1 U9935 ( .A(n7622), .B(n7620), .ZN(n11039) );
  OR2_X1 U9936 ( .A1(n8003), .A2(n11039), .ZN(n7609) );
  NAND2_X1 U9937 ( .A1(n7538), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7608) );
  NAND4_X1 U9938 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n13717)
         );
  XNOR2_X1 U9939 ( .A(n11734), .B(n13717), .ZN(n11898) );
  INV_X1 U9940 ( .A(n11898), .ZN(n11041) );
  OR2_X1 U9941 ( .A1(n11734), .A2(n13717), .ZN(n7612) );
  INV_X1 U9942 ( .A(n7613), .ZN(n7614) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n7777), .Z(n7632) );
  XNOR2_X1 U9944 ( .A(n7632), .B(SI_8_), .ZN(n7629) );
  NAND2_X1 U9945 ( .A1(n9775), .A2(n7965), .ZN(n7618) );
  INV_X1 U9946 ( .A(n7813), .ZN(n7750) );
  NAND2_X1 U9947 ( .A1(n7750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7635) );
  XNOR2_X1 U9948 ( .A(n7635), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U9949 ( .A1(n8000), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7836), .B2(
        n9901), .ZN(n7617) );
  NAND2_X1 U9950 ( .A1(n7538), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7628) );
  INV_X1 U9951 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7619) );
  OAI21_X1 U9952 ( .B1(n7622), .B2(n7620), .A(n7619), .ZN(n7623) );
  NAND2_X1 U9953 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n7621) );
  NAND2_X1 U9954 ( .A1(n7623), .A2(n7639), .ZN(n11168) );
  OR2_X1 U9955 ( .A1(n8003), .A2(n11168), .ZN(n7627) );
  INV_X1 U9956 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7624) );
  OR2_X1 U9957 ( .A1(n7561), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U9958 ( .A1(n8105), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7625) );
  NAND4_X1 U9959 ( .A1(n7628), .A2(n7627), .A3(n7626), .A4(n7625), .ZN(n13716)
         );
  XNOR2_X1 U9960 ( .A(n11739), .B(n13716), .ZN(n11900) );
  INV_X1 U9961 ( .A(n7629), .ZN(n7630) );
  NAND2_X1 U9962 ( .A1(n7632), .A2(SI_8_), .ZN(n7633) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n7777), .Z(n7649) );
  XNOR2_X1 U9964 ( .A(n7649), .B(SI_9_), .ZN(n7646) );
  XNOR2_X1 U9965 ( .A(n7648), .B(n7646), .ZN(n9857) );
  NAND2_X1 U9966 ( .A1(n9857), .A2(n7965), .ZN(n7638) );
  INV_X1 U9967 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9968 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U9969 ( .A1(n7636), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7677) );
  XNOR2_X1 U9970 ( .A(n7677), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U9971 ( .A1(n8000), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7836), .B2(
        n10183), .ZN(n7637) );
  NAND2_X1 U9972 ( .A1(n7538), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9973 ( .A1(n7639), .A2(n11354), .ZN(n7640) );
  NAND2_X1 U9974 ( .A1(n7659), .A2(n7640), .ZN(n10964) );
  OR2_X1 U9975 ( .A1(n8003), .A2(n10964), .ZN(n7643) );
  INV_X1 U9976 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9900) );
  OR2_X1 U9977 ( .A1(n7561), .A2(n9900), .ZN(n7642) );
  NAND2_X1 U9978 ( .A1(n8105), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7641) );
  NAND4_X1 U9979 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n13715)
         );
  INV_X1 U9980 ( .A(n13715), .ZN(n11474) );
  XNOR2_X1 U9981 ( .A(n11748), .B(n11474), .ZN(n11902) );
  OR2_X1 U9982 ( .A1(n11748), .A2(n13715), .ZN(n7645) );
  INV_X1 U9983 ( .A(n7646), .ZN(n7647) );
  NAND2_X1 U9984 ( .A1(n7649), .A2(SI_9_), .ZN(n7650) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n7777), .Z(n7669) );
  XNOR2_X1 U9986 ( .A(n7669), .B(SI_10_), .ZN(n7652) );
  INV_X1 U9987 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U9988 ( .A1(n7677), .A2(n7653), .ZN(n7654) );
  NAND2_X1 U9989 ( .A1(n7654), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7655) );
  XNOR2_X1 U9990 ( .A(n7655), .B(P1_IR_REG_10__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U9991 ( .A1(n8000), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7836), .B2(
        n13788), .ZN(n7656) );
  NAND2_X2 U9992 ( .A1(n7657), .A2(n7656), .ZN(n11757) );
  NAND2_X1 U9993 ( .A1(n7538), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U9994 ( .A1(n8105), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7664) );
  INV_X1 U9995 ( .A(n7680), .ZN(n7661) );
  NAND2_X1 U9996 ( .A1(n7659), .A2(n7658), .ZN(n7660) );
  NAND2_X1 U9997 ( .A1(n7661), .A2(n7660), .ZN(n11472) );
  OR2_X1 U9998 ( .A1(n8003), .A2(n11472), .ZN(n7663) );
  NAND2_X1 U9999 ( .A1(n8004), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7662) );
  NAND4_X1 U10000 ( .A1(n7665), .A2(n7664), .A3(n7663), .A4(n7662), .ZN(n13714) );
  INV_X1 U10001 ( .A(n13714), .ZN(n14476) );
  XNOR2_X1 U10002 ( .A(n11757), .B(n14476), .ZN(n11903) );
  OR2_X1 U10003 ( .A1(n11757), .A2(n13714), .ZN(n7666) );
  INV_X1 U10004 ( .A(n7669), .ZN(n7667) );
  NAND2_X1 U10005 ( .A1(n7669), .A2(SI_10_), .ZN(n7670) );
  MUX2_X1 U10006 ( .A(n9967), .B(n9965), .S(n7777), .Z(n7671) );
  INV_X1 U10007 ( .A(n7671), .ZN(n7672) );
  NAND2_X1 U10008 ( .A1(n7672), .A2(SI_11_), .ZN(n7673) );
  NAND2_X1 U10009 ( .A1(n7687), .A2(n7673), .ZN(n7688) );
  NAND2_X1 U10010 ( .A1(n9964), .A2(n7965), .ZN(n7679) );
  INV_X1 U10011 ( .A(n7674), .ZN(n7675) );
  NAND2_X1 U10012 ( .A1(n7675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U10013 ( .A1(n7677), .A2(n7676), .ZN(n7693) );
  INV_X1 U10014 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7746) );
  XNOR2_X1 U10015 ( .A(n7693), .B(n7746), .ZN(n10324) );
  AOI22_X1 U10016 ( .A1(n8000), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7836), 
        .B2(n10324), .ZN(n7678) );
  NAND2_X2 U10017 ( .A1(n7679), .A2(n7678), .ZN(n14489) );
  NAND2_X1 U10018 ( .A1(n7680), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7698) );
  OR2_X1 U10019 ( .A1(n7680), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U10020 ( .A1(n7698), .A2(n7681), .ZN(n14493) );
  OR2_X1 U10021 ( .A1(n8003), .A2(n14493), .ZN(n7686) );
  NAND2_X1 U10022 ( .A1(n7984), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7685) );
  INV_X1 U10023 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7682) );
  OR2_X1 U10024 ( .A1(n7561), .A2(n7682), .ZN(n7684) );
  NAND2_X1 U10025 ( .A1(n7538), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7683) );
  NAND4_X1 U10026 ( .A1(n7686), .A2(n7685), .A3(n7684), .A4(n7683), .ZN(n13713) );
  INV_X1 U10027 ( .A(n13713), .ZN(n8077) );
  XNOR2_X1 U10028 ( .A(n14489), .B(n8077), .ZN(n11904) );
  MUX2_X1 U10029 ( .A(n8975), .B(n10039), .S(n7777), .Z(n7690) );
  INV_X1 U10030 ( .A(n7690), .ZN(n7691) );
  NAND2_X1 U10031 ( .A1(n7691), .A2(SI_12_), .ZN(n7692) );
  NAND2_X1 U10032 ( .A1(n10020), .A2(n7965), .ZN(n7696) );
  NAND2_X1 U10033 ( .A1(n7694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7710) );
  XNOR2_X1 U10034 ( .A(n7710), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U10035 ( .A1(n8000), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7836), 
        .B2(n14562), .ZN(n7695) );
  NAND2_X1 U10036 ( .A1(n7538), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U10037 ( .A1(n8105), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U10038 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  NAND2_X1 U10039 ( .A1(n7717), .A2(n7699), .ZN(n11328) );
  OR2_X1 U10040 ( .A1(n8003), .A2(n11328), .ZN(n7701) );
  NAND2_X1 U10041 ( .A1(n8004), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7700) );
  NAND4_X1 U10042 ( .A1(n7703), .A2(n7702), .A3(n7701), .A4(n7700), .ZN(n13712) );
  XNOR2_X1 U10043 ( .A(n11768), .B(n13712), .ZN(n11905) );
  INV_X1 U10044 ( .A(n11905), .ZN(n11321) );
  OR2_X1 U10045 ( .A1(n11768), .A2(n13712), .ZN(n7704) );
  MUX2_X1 U10046 ( .A(n10213), .B(n10214), .S(n7777), .Z(n7725) );
  XNOR2_X1 U10047 ( .A(n7725), .B(SI_13_), .ZN(n7708) );
  XNOR2_X1 U10048 ( .A(n7726), .B(n7708), .ZN(n10212) );
  NAND2_X1 U10049 ( .A1(n10212), .A2(n7965), .ZN(n7716) );
  INV_X1 U10050 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U10051 ( .A1(n7710), .A2(n7709), .ZN(n7711) );
  NAND2_X1 U10052 ( .A1(n7711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7713) );
  INV_X1 U10053 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U10054 ( .A1(n7713), .A2(n7712), .ZN(n7727) );
  OR2_X1 U10055 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  AOI22_X1 U10056 ( .A1(n8000), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10587), 
        .B2(n7836), .ZN(n7715) );
  NAND2_X1 U10057 ( .A1(n7538), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U10058 ( .A1(n8105), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7722) );
  INV_X1 U10059 ( .A(n7731), .ZN(n7719) );
  NAND2_X1 U10060 ( .A1(n7717), .A2(n13649), .ZN(n7718) );
  NAND2_X1 U10061 ( .A1(n7719), .A2(n7718), .ZN(n13648) );
  OR2_X1 U10062 ( .A1(n8003), .A2(n13648), .ZN(n7721) );
  NAND2_X1 U10063 ( .A1(n8004), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7720) );
  NAND4_X1 U10064 ( .A1(n7723), .A2(n7722), .A3(n7721), .A4(n7720), .ZN(n13711) );
  XNOR2_X1 U10065 ( .A(n12040), .B(n13711), .ZN(n11906) );
  INV_X1 U10066 ( .A(n11906), .ZN(n11337) );
  OR2_X1 U10067 ( .A1(n12040), .A2(n13711), .ZN(n7724) );
  MUX2_X1 U10068 ( .A(n10388), .B(n10389), .S(n7777), .Z(n7771) );
  NAND2_X1 U10069 ( .A1(n10387), .A2(n7965), .ZN(n7730) );
  NAND2_X1 U10070 ( .A1(n7727), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7728) );
  XNOR2_X1 U10071 ( .A(n7728), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U10072 ( .A1(n11526), .A2(n7836), .B1(n8000), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U10073 ( .A1(n7984), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10074 ( .A1(n7731), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7759) );
  OR2_X1 U10075 ( .A1(n7731), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U10076 ( .A1(n7759), .A2(n7732), .ZN(n14461) );
  OR2_X1 U10077 ( .A1(n8003), .A2(n14461), .ZN(n7736) );
  INV_X1 U10078 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7733) );
  OR2_X1 U10079 ( .A1(n7561), .A2(n7733), .ZN(n7735) );
  INV_X1 U10080 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11548) );
  OR2_X1 U10081 ( .A1(n11852), .A2(n11548), .ZN(n7734) );
  NAND2_X1 U10082 ( .A1(n14507), .A2(n13710), .ZN(n7740) );
  NAND2_X1 U10083 ( .A1(n7741), .A2(n7771), .ZN(n7743) );
  NAND2_X1 U10084 ( .A1(n7770), .A2(n15127), .ZN(n7742) );
  NAND2_X1 U10085 ( .A1(n7743), .A2(n7742), .ZN(n7745) );
  MUX2_X1 U10086 ( .A(n10470), .B(n10471), .S(n7777), .Z(n7773) );
  XNOR2_X1 U10087 ( .A(n7773), .B(SI_15_), .ZN(n7744) );
  NOR2_X1 U10088 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7747) );
  NAND4_X1 U10089 ( .A1(n7748), .A2(n7674), .A3(n7747), .A4(n7746), .ZN(n7749)
         );
  OR2_X1 U10090 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  NAND2_X1 U10091 ( .A1(n7752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7751) );
  MUX2_X1 U10092 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7751), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n7755) );
  INV_X1 U10093 ( .A(n7752), .ZN(n7754) );
  INV_X1 U10094 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10095 ( .A1(n7754), .A2(n7753), .ZN(n7779) );
  NAND2_X1 U10096 ( .A1(n7755), .A2(n7779), .ZN(n11530) );
  AOI22_X1 U10097 ( .A1(n8000), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6487), 
        .B2(n14574), .ZN(n7756) );
  NAND2_X1 U10098 ( .A1(n7984), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7765) );
  INV_X1 U10099 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7758) );
  OR2_X1 U10100 ( .A1(n7561), .A2(n7758), .ZN(n7764) );
  NAND2_X1 U10101 ( .A1(n7759), .A2(n13691), .ZN(n7760) );
  NAND2_X1 U10102 ( .A1(n7784), .A2(n7760), .ZN(n11515) );
  OR2_X1 U10103 ( .A1(n8003), .A2(n11515), .ZN(n7763) );
  INV_X1 U10104 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7761) );
  OR2_X1 U10105 ( .A1(n11852), .A2(n7761), .ZN(n7762) );
  NAND2_X1 U10106 ( .A1(n12047), .A2(n14462), .ZN(n11785) );
  NAND2_X1 U10107 ( .A1(n11784), .A2(n11785), .ZN(n11910) );
  INV_X1 U10108 ( .A(n14462), .ZN(n13709) );
  OR2_X1 U10109 ( .A1(n12047), .A2(n13709), .ZN(n7767) );
  INV_X1 U10110 ( .A(n7773), .ZN(n7768) );
  NAND2_X1 U10111 ( .A1(n7768), .A2(SI_15_), .ZN(n7774) );
  OAI21_X1 U10112 ( .B1(n15127), .B2(n7771), .A(n7774), .ZN(n7769) );
  INV_X1 U10113 ( .A(n7771), .ZN(n7772) );
  NOR2_X1 U10114 ( .A1(n7772), .A2(SI_14_), .ZN(n7775) );
  AOI22_X1 U10115 ( .A1(n7775), .A2(n7774), .B1(n7773), .B2(n9915), .ZN(n7776)
         );
  MUX2_X1 U10116 ( .A(n10384), .B(n10385), .S(n7777), .Z(n7795) );
  XNOR2_X1 U10117 ( .A(n7795), .B(SI_16_), .ZN(n7793) );
  XNOR2_X1 U10118 ( .A(n7794), .B(n7793), .ZN(n10383) );
  NAND2_X1 U10119 ( .A1(n10383), .A2(n7965), .ZN(n7782) );
  NAND2_X1 U10120 ( .A1(n7779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7778) );
  MUX2_X1 U10121 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7778), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n7780) );
  AOI22_X1 U10122 ( .A1(n8000), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7836), 
        .B2(n11534), .ZN(n7781) );
  AND2_X1 U10123 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  OR2_X1 U10124 ( .A1(n7785), .A2(n7803), .ZN(n14475) );
  NAND2_X1 U10125 ( .A1(n8105), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10126 ( .A1(n7538), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7786) );
  AND2_X1 U10127 ( .A1(n7787), .A2(n7786), .ZN(n7789) );
  NAND2_X1 U10128 ( .A1(n8004), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7788) );
  OAI211_X1 U10129 ( .C1(n8003), .C2(n14475), .A(n7789), .B(n7788), .ZN(n13708) );
  NAND2_X1 U10130 ( .A1(n14472), .A2(n13708), .ZN(n7790) );
  OR2_X1 U10131 ( .A1(n14472), .A2(n13708), .ZN(n7791) );
  NAND2_X1 U10132 ( .A1(n7794), .A2(n7793), .ZN(n7797) );
  NAND2_X1 U10133 ( .A1(n7795), .A2(n15194), .ZN(n7796) );
  MUX2_X1 U10134 ( .A(n10421), .B(n10423), .S(n9735), .Z(n7808) );
  XNOR2_X1 U10135 ( .A(n7808), .B(SI_17_), .ZN(n7798) );
  XNOR2_X1 U10136 ( .A(n7810), .B(n7798), .ZN(n10420) );
  NAND2_X1 U10137 ( .A1(n10420), .A2(n7965), .ZN(n7802) );
  NAND2_X1 U10138 ( .A1(n7799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U10139 ( .A(n7800), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U10140 ( .A1(n8000), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6487), 
        .B2(n11545), .ZN(n7801) );
  NOR2_X1 U10141 ( .A1(n7803), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7804) );
  OR2_X1 U10142 ( .A1(n7821), .A2(n7804), .ZN(n13621) );
  AOI22_X1 U10143 ( .A1(n7538), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n7984), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U10144 ( .A1(n8004), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7805) );
  OAI211_X1 U10145 ( .C1(n13621), .C2(n8003), .A(n7806), .B(n7805), .ZN(n13707) );
  XNOR2_X1 U10146 ( .A(n13623), .B(n13707), .ZN(n11911) );
  NAND2_X1 U10147 ( .A1(n13623), .A2(n13707), .ZN(n7807) );
  NOR2_X1 U10148 ( .A1(n7811), .A2(SI_17_), .ZN(n7809) );
  NAND2_X1 U10149 ( .A1(n7811), .A2(SI_17_), .ZN(n7812) );
  XNOR2_X1 U10150 ( .A(n7851), .B(SI_18_), .ZN(n7825) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9735), .Z(n7844) );
  XNOR2_X1 U10152 ( .A(n7825), .B(n7844), .ZN(n10843) );
  NAND2_X1 U10153 ( .A1(n10843), .A2(n7965), .ZN(n7820) );
  AND2_X2 U10154 ( .A1(n7813), .A2(n6536), .ZN(n7817) );
  INV_X1 U10155 ( .A(n7817), .ZN(n7814) );
  NAND2_X1 U10156 ( .A1(n7814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7815) );
  MUX2_X1 U10157 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7815), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n7818) );
  NAND2_X1 U10158 ( .A1(n7818), .A2(n7834), .ZN(n11554) );
  INV_X1 U10159 ( .A(n11554), .ZN(n13833) );
  AOI22_X1 U10160 ( .A1(n8000), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6487), 
        .B2(n13833), .ZN(n7819) );
  NOR2_X1 U10161 ( .A1(n7821), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7822) );
  OR2_X1 U10162 ( .A1(n7839), .A2(n7822), .ZN(n14032) );
  AOI22_X1 U10163 ( .A1(n7538), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n8105), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10164 ( .A1(n8004), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7823) );
  OAI211_X1 U10165 ( .C1(n14032), .C2(n8003), .A(n7824), .B(n7823), .ZN(n14007) );
  NAND2_X1 U10166 ( .A1(n14125), .A2(n14007), .ZN(n11789) );
  INV_X1 U10167 ( .A(n11789), .ZN(n11800) );
  OR2_X1 U10168 ( .A1(n14125), .A2(n14007), .ZN(n11798) );
  INV_X1 U10169 ( .A(n7825), .ZN(n7826) );
  NAND2_X1 U10170 ( .A1(n7826), .A2(n7844), .ZN(n7828) );
  NAND2_X1 U10171 ( .A1(n7851), .A2(SI_18_), .ZN(n7827) );
  NAND2_X1 U10172 ( .A1(n7828), .A2(n7827), .ZN(n7832) );
  MUX2_X1 U10173 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9735), .Z(n7829) );
  INV_X1 U10174 ( .A(n7829), .ZN(n7830) );
  NAND2_X1 U10175 ( .A1(n7830), .A2(n15160), .ZN(n7845) );
  NAND2_X1 U10176 ( .A1(n7847), .A2(n7845), .ZN(n7831) );
  NAND2_X1 U10177 ( .A1(n10952), .A2(n7965), .ZN(n7838) );
  NAND2_X1 U10178 ( .A1(n7834), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7833) );
  MUX2_X1 U10179 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7833), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n7835) );
  NAND2_X2 U10180 ( .A1(n8035), .A2(n7835), .ZN(n13843) );
  AOI22_X1 U10181 ( .A1(n8000), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11688), 
        .B2(n6487), .ZN(n7837) );
  NOR2_X1 U10182 ( .A1(n7839), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7840) );
  OR2_X1 U10183 ( .A1(n7854), .A2(n7840), .ZN(n14012) );
  AOI22_X1 U10184 ( .A1(n8004), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n7984), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U10185 ( .A1(n7538), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7841) );
  OAI211_X1 U10186 ( .C1(n14012), .C2(n8003), .A(n7842), .B(n7841), .ZN(n13984) );
  XNOR2_X1 U10187 ( .A(n14119), .B(n13984), .ZN(n14005) );
  INV_X1 U10188 ( .A(n14005), .ZN(n8086) );
  NOR2_X1 U10189 ( .A1(n14119), .A2(n13984), .ZN(n13994) );
  INV_X1 U10190 ( .A(n13994), .ZN(n7863) );
  INV_X1 U10191 ( .A(n7844), .ZN(n7843) );
  NOR2_X1 U10192 ( .A1(n7844), .A2(SI_18_), .ZN(n7848) );
  INV_X1 U10193 ( .A(n7845), .ZN(n7846) );
  XNOR2_X1 U10194 ( .A(n7886), .B(SI_20_), .ZN(n7867) );
  MUX2_X1 U10195 ( .A(n11936), .B(n11024), .S(n9735), .Z(n7882) );
  XNOR2_X1 U10196 ( .A(n7867), .B(n7882), .ZN(n11022) );
  NAND2_X1 U10197 ( .A1(n11022), .A2(n7965), .ZN(n7853) );
  NAND2_X1 U10198 ( .A1(n8000), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7852) );
  OR2_X1 U10199 ( .A1(n7854), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7855) );
  AND2_X1 U10200 ( .A1(n7855), .A2(n7873), .ZN(n13989) );
  INV_X1 U10201 ( .A(n8003), .ZN(n7856) );
  NAND2_X1 U10202 ( .A1(n13989), .A2(n7856), .ZN(n7862) );
  INV_X1 U10203 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10204 ( .A1(n8105), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10205 ( .A1(n7538), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7857) );
  OAI211_X1 U10206 ( .C1(n7859), .C2(n7561), .A(n7858), .B(n7857), .ZN(n7860)
         );
  INV_X1 U10207 ( .A(n7860), .ZN(n7861) );
  XNOR2_X1 U10208 ( .A(n14115), .B(n13598), .ZN(n11914) );
  AND2_X1 U10209 ( .A1(n7863), .A2(n11914), .ZN(n7864) );
  OR2_X1 U10210 ( .A1(n13991), .A2(n13598), .ZN(n7865) );
  INV_X1 U10211 ( .A(n7882), .ZN(n7880) );
  NOR2_X1 U10212 ( .A1(n7886), .A2(n10513), .ZN(n7866) );
  AOI21_X1 U10213 ( .B1(n7867), .B2(n7880), .A(n7866), .ZN(n7869) );
  MUX2_X1 U10214 ( .A(n11077), .B(n11076), .S(n9735), .Z(n7881) );
  XNOR2_X1 U10215 ( .A(n7881), .B(SI_21_), .ZN(n7868) );
  XNOR2_X1 U10216 ( .A(n7869), .B(n7868), .ZN(n11074) );
  NAND2_X1 U10217 ( .A1(n11074), .A2(n7965), .ZN(n7871) );
  NAND2_X1 U10218 ( .A1(n8000), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10219 ( .A1(n8105), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7878) );
  INV_X1 U10220 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7872) );
  OR2_X1 U10221 ( .A1(n7561), .A2(n7872), .ZN(n7877) );
  OAI21_X1 U10222 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n7874), .A(n7889), .ZN(
        n13972) );
  OR2_X1 U10223 ( .A1(n8003), .A2(n13972), .ZN(n7876) );
  INV_X1 U10224 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n13973) );
  OR2_X1 U10225 ( .A1(n11852), .A2(n13973), .ZN(n7875) );
  XNOR2_X1 U10226 ( .A(n14109), .B(n13656), .ZN(n13976) );
  INV_X1 U10227 ( .A(n13976), .ZN(n8089) );
  NAND2_X1 U10228 ( .A1(n13971), .A2(n13656), .ZN(n7879) );
  NOR2_X1 U10229 ( .A1(n7882), .A2(n10513), .ZN(n7884) );
  AOI22_X1 U10230 ( .A1(n7884), .A2(n7453), .B1(n7883), .B2(SI_21_), .ZN(n7885) );
  OR2_X1 U10231 ( .A1(n8465), .A2(n9735), .ZN(n7888) );
  XNOR2_X1 U10232 ( .A(n7888), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14169) );
  NAND2_X1 U10233 ( .A1(n8105), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10234 ( .A1(n8004), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7893) );
  OAI21_X1 U10235 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n7890), .A(n7902), .ZN(
        n13963) );
  OR2_X1 U10236 ( .A1(n8003), .A2(n13963), .ZN(n7892) );
  NAND2_X1 U10237 ( .A1(n7538), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7891) );
  NAND4_X1 U10238 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n13706) );
  XNOR2_X1 U10239 ( .A(n13957), .B(n13706), .ZN(n13959) );
  OR2_X1 U10240 ( .A1(n14104), .A2(n13706), .ZN(n7895) );
  NAND2_X1 U10241 ( .A1(n13953), .A2(n7895), .ZN(n13936) );
  INV_X1 U10242 ( .A(n13936), .ZN(n7909) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9735), .Z(n8464) );
  INV_X1 U10244 ( .A(n8464), .ZN(n7898) );
  NAND2_X1 U10245 ( .A1(n7896), .A2(SI_22_), .ZN(n7897) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9735), .Z(n7912) );
  XNOR2_X1 U10247 ( .A(n7911), .B(SI_23_), .ZN(n11390) );
  NAND2_X1 U10248 ( .A1(n11390), .A2(n7965), .ZN(n7900) );
  NAND2_X1 U10249 ( .A1(n8000), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U10250 ( .A1(n8105), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7907) );
  INV_X1 U10251 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7901) );
  OR2_X1 U10252 ( .A1(n7561), .A2(n7901), .ZN(n7906) );
  OAI21_X1 U10253 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n7903), .A(n7917), .ZN(
        n13944) );
  OR2_X1 U10254 ( .A1(n8003), .A2(n13944), .ZN(n7905) );
  INV_X1 U10255 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13945) );
  OR2_X1 U10256 ( .A1(n11852), .A2(n13945), .ZN(n7904) );
  XNOR2_X1 U10257 ( .A(n6904), .B(n13705), .ZN(n13938) );
  OR2_X1 U10258 ( .A1(n13943), .A2(n13657), .ZN(n7910) );
  NAND2_X1 U10259 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  MUX2_X1 U10260 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9735), .Z(n7925) );
  XNOR2_X1 U10261 ( .A(n7924), .B(n7925), .ZN(n13557) );
  NAND2_X1 U10262 ( .A1(n13557), .A2(n7965), .ZN(n7916) );
  NAND2_X1 U10263 ( .A1(n8000), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10264 ( .A1(n7538), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10265 ( .A1(n7984), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7921) );
  OAI21_X1 U10266 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7918), .A(n7937), .ZN(
        n13631) );
  OR2_X1 U10267 ( .A1(n8003), .A2(n13631), .ZN(n7920) );
  NAND2_X1 U10268 ( .A1(n8004), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7919) );
  NAND4_X1 U10269 ( .A1(n7922), .A2(n7921), .A3(n7920), .A4(n7919), .ZN(n13704) );
  XNOR2_X1 U10270 ( .A(n13928), .B(n13704), .ZN(n13914) );
  INV_X1 U10271 ( .A(n7924), .ZN(n7926) );
  NAND2_X1 U10272 ( .A1(n7926), .A2(n7925), .ZN(n7929) );
  NAND2_X1 U10273 ( .A1(n7927), .A2(SI_24_), .ZN(n7928) );
  INV_X1 U10274 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14161) );
  MUX2_X1 U10275 ( .A(n14161), .B(n13556), .S(n9735), .Z(n7930) );
  NAND2_X1 U10276 ( .A1(n7930), .A2(n15221), .ZN(n7946) );
  INV_X1 U10277 ( .A(n7930), .ZN(n7931) );
  NAND2_X1 U10278 ( .A1(n7931), .A2(SI_25_), .ZN(n7932) );
  NAND2_X1 U10279 ( .A1(n7946), .A2(n7932), .ZN(n7947) );
  NAND2_X1 U10280 ( .A1(n13554), .A2(n7965), .ZN(n7934) );
  NAND2_X1 U10281 ( .A1(n8000), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7933) );
  NAND2_X2 U10282 ( .A1(n7934), .A2(n7933), .ZN(n14084) );
  NAND2_X1 U10283 ( .A1(n7538), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10284 ( .A1(n7984), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7941) );
  INV_X1 U10285 ( .A(n7937), .ZN(n7935) );
  NAND2_X1 U10286 ( .A1(n7935), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7954) );
  INV_X1 U10287 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10288 ( .A1(n7937), .A2(n7936), .ZN(n7938) );
  NAND2_X1 U10289 ( .A1(n7954), .A2(n7938), .ZN(n13908) );
  OR2_X1 U10290 ( .A1(n8003), .A2(n13908), .ZN(n7940) );
  NAND2_X1 U10291 ( .A1(n8004), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7939) );
  NAND4_X1 U10292 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .ZN(n13886) );
  NAND2_X1 U10293 ( .A1(n14084), .A2(n13886), .ZN(n7944) );
  OR2_X1 U10294 ( .A1(n14084), .A2(n13886), .ZN(n7943) );
  NAND2_X1 U10295 ( .A1(n7944), .A2(n7943), .ZN(n13898) );
  INV_X1 U10296 ( .A(n7944), .ZN(n7945) );
  INV_X1 U10297 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14158) );
  INV_X1 U10298 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13551) );
  MUX2_X1 U10299 ( .A(n14158), .B(n13551), .S(n9735), .Z(n7961) );
  XNOR2_X1 U10300 ( .A(n7961), .B(SI_26_), .ZN(n7949) );
  XNOR2_X1 U10301 ( .A(n7962), .B(n7949), .ZN(n13549) );
  NAND2_X1 U10302 ( .A1(n13549), .A2(n7965), .ZN(n7951) );
  NAND2_X1 U10303 ( .A1(n8000), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10304 ( .A1(n7984), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10305 ( .A1(n8004), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7958) );
  INV_X1 U10306 ( .A(n7954), .ZN(n7952) );
  NAND2_X1 U10307 ( .A1(n7952), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7970) );
  INV_X1 U10308 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U10309 ( .A1(n7954), .A2(n7953), .ZN(n7955) );
  NAND2_X1 U10310 ( .A1(n7970), .A2(n7955), .ZN(n13680) );
  OR2_X1 U10311 ( .A1(n8003), .A2(n13680), .ZN(n7957) );
  NAND2_X1 U10312 ( .A1(n7538), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7956) );
  NAND4_X1 U10313 ( .A1(n7959), .A2(n7958), .A3(n7957), .A4(n7956), .ZN(n13703) );
  NAND2_X1 U10314 ( .A1(n14079), .A2(n13603), .ZN(n8094) );
  OR2_X1 U10315 ( .A1(n14079), .A2(n13603), .ZN(n7960) );
  NAND2_X1 U10316 ( .A1(n8094), .A2(n7960), .ZN(n11917) );
  INV_X1 U10317 ( .A(n14079), .ZN(n13892) );
  MUX2_X1 U10318 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9735), .Z(n7979) );
  INV_X1 U10319 ( .A(n7979), .ZN(n7963) );
  XNOR2_X1 U10320 ( .A(n7963), .B(SI_27_), .ZN(n7964) );
  XNOR2_X1 U10321 ( .A(n7981), .B(n7964), .ZN(n13546) );
  NAND2_X1 U10322 ( .A1(n13546), .A2(n7965), .ZN(n7967) );
  NAND2_X1 U10323 ( .A1(n8000), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7966) );
  NAND2_X2 U10324 ( .A1(n7967), .A2(n7966), .ZN(n14075) );
  NAND2_X1 U10325 ( .A1(n8105), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U10326 ( .A1(n8004), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7974) );
  INV_X1 U10327 ( .A(n7970), .ZN(n7968) );
  NAND2_X1 U10328 ( .A1(n7968), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7987) );
  INV_X1 U10329 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10330 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  NAND2_X1 U10331 ( .A1(n7987), .A2(n7971), .ZN(n11948) );
  OR2_X1 U10332 ( .A1(n8003), .A2(n11948), .ZN(n7973) );
  NAND2_X1 U10333 ( .A1(n7538), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10334 ( .A1(n14075), .A2(n7977), .ZN(n8095) );
  OR2_X1 U10335 ( .A1(n14075), .A2(n7977), .ZN(n7976) );
  NAND2_X1 U10336 ( .A1(n8095), .A2(n7976), .ZN(n11918) );
  INV_X1 U10337 ( .A(n14075), .ZN(n13569) );
  NOR2_X1 U10338 ( .A1(n7979), .A2(SI_27_), .ZN(n7980) );
  MUX2_X1 U10339 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9735), .Z(n7996) );
  XNOR2_X1 U10340 ( .A(n7996), .B(SI_28_), .ZN(n7994) );
  NAND2_X1 U10341 ( .A1(n11684), .A2(n7965), .ZN(n7983) );
  NAND2_X1 U10342 ( .A1(n8000), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10343 ( .A1(n7538), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10344 ( .A1(n8105), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7991) );
  INV_X1 U10345 ( .A(n7987), .ZN(n7985) );
  NAND2_X1 U10346 ( .A1(n7985), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8104) );
  INV_X1 U10347 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10348 ( .A1(n7987), .A2(n7986), .ZN(n7988) );
  NAND2_X1 U10349 ( .A1(n8104), .A2(n7988), .ZN(n13871) );
  NAND2_X1 U10350 ( .A1(n8004), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7989) );
  NAND4_X1 U10351 ( .A1(n7992), .A2(n7991), .A3(n7990), .A4(n7989), .ZN(n13702) );
  NAND2_X1 U10352 ( .A1(n14070), .A2(n12160), .ZN(n8096) );
  OR2_X1 U10353 ( .A1(n14070), .A2(n12160), .ZN(n7993) );
  NAND2_X1 U10354 ( .A1(n8096), .A2(n7993), .ZN(n13873) );
  INV_X1 U10355 ( .A(n14070), .ZN(n12162) );
  NAND2_X1 U10356 ( .A1(n13872), .A2(n6540), .ZN(n8010) );
  INV_X1 U10357 ( .A(n7996), .ZN(n7997) );
  INV_X1 U10358 ( .A(SI_28_), .ZN(n15184) );
  NAND2_X1 U10359 ( .A1(n7997), .A2(n15184), .ZN(n7998) );
  INV_X1 U10360 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14152) );
  INV_X1 U10361 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13540) );
  MUX2_X1 U10362 ( .A(n14152), .B(n13540), .S(n9735), .Z(n8831) );
  XNOR2_X1 U10363 ( .A(n8831), .B(SI_29_), .ZN(n8829) );
  NAND2_X1 U10364 ( .A1(n13539), .A2(n7965), .ZN(n8002) );
  NAND2_X1 U10365 ( .A1(n8000), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10366 ( .A1(n7538), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10367 ( .A1(n8105), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8007) );
  OR2_X1 U10368 ( .A1(n8003), .A2(n8104), .ZN(n8006) );
  NAND2_X1 U10369 ( .A1(n8004), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8005) );
  NAND4_X1 U10370 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n13862) );
  XNOR2_X1 U10371 ( .A(n14065), .B(n13862), .ZN(n11920) );
  NAND2_X1 U10372 ( .A1(n7813), .A2(n8011), .ZN(n8038) );
  INV_X1 U10373 ( .A(n8038), .ZN(n8013) );
  NAND2_X1 U10374 ( .A1(n8013), .A2(n8012), .ZN(n8040) );
  INV_X1 U10375 ( .A(n8040), .ZN(n8014) );
  NAND2_X1 U10376 ( .A1(n8014), .A2(n8032), .ZN(n8023) );
  NAND2_X1 U10377 ( .A1(n8023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10378 ( .A1(n8018), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8020) );
  INV_X1 U10379 ( .A(n14160), .ZN(n8021) );
  AND2_X1 U10380 ( .A1(n8022), .A2(n8021), .ZN(n8027) );
  NAND3_X1 U10381 ( .A1(n8031), .A2(P1_B_REG_SCAN_IN), .A3(n14167), .ZN(n8026)
         );
  NAND2_X1 U10382 ( .A1(n8027), .A2(n8026), .ZN(n10125) );
  OR2_X1 U10383 ( .A1(n10125), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10384 ( .A1(n14167), .A2(n14160), .ZN(n8028) );
  INV_X1 U10385 ( .A(n10130), .ZN(n10143) );
  OR3_X4 U10386 ( .A1(n8031), .A2(n14160), .A3(n8030), .ZN(n9931) );
  NAND2_X1 U10387 ( .A1(n8040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U10388 ( .A(n8033), .B(n8032), .ZN(n9743) );
  INV_X1 U10389 ( .A(n8056), .ZN(n8102) );
  NAND2_X1 U10390 ( .A1(n14043), .A2(n8102), .ZN(n11861) );
  NAND2_X1 U10391 ( .A1(n8038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8039) );
  MUX2_X1 U10392 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8039), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8041) );
  NAND2_X1 U10393 ( .A1(n8041), .A2(n8040), .ZN(n11687) );
  NAND2_X1 U10394 ( .A1(n11688), .A2(n14168), .ZN(n8042) );
  NAND2_X1 U10395 ( .A1(n14043), .A2(n14168), .ZN(n11872) );
  INV_X1 U10396 ( .A(n11872), .ZN(n8043) );
  NAND2_X1 U10397 ( .A1(n14028), .A2(n8043), .ZN(n10342) );
  NAND2_X1 U10398 ( .A1(n9943), .A2(n10342), .ZN(n11931) );
  INV_X1 U10399 ( .A(n11931), .ZN(n9942) );
  NOR4_X1 U10400 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8047) );
  NOR4_X1 U10401 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8046) );
  NOR4_X1 U10402 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8045) );
  NOR4_X1 U10403 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8044) );
  NAND4_X1 U10404 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8053)
         );
  NOR2_X1 U10405 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n8051) );
  NOR4_X1 U10406 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8050) );
  NOR4_X1 U10407 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8049) );
  NOR4_X1 U10408 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8048) );
  NAND4_X1 U10409 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n8052)
         );
  NOR2_X1 U10410 ( .A1(n8053), .A2(n8052), .ZN(n10124) );
  AND2_X1 U10411 ( .A1(n10124), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8054) );
  OR2_X1 U10412 ( .A1(n10125), .A2(n8054), .ZN(n8055) );
  NAND2_X1 U10413 ( .A1(n8031), .A2(n14160), .ZN(n10123) );
  AND2_X1 U10414 ( .A1(n8055), .A2(n10123), .ZN(n9936) );
  NAND3_X1 U10415 ( .A1(n10143), .A2(n9942), .A3(n9936), .ZN(n8109) );
  INV_X1 U10416 ( .A(n10127), .ZN(n8057) );
  NAND2_X2 U10417 ( .A1(n14043), .A2(n8056), .ZN(n9930) );
  OR2_X1 U10418 ( .A1(n9930), .A2(n11689), .ZN(n14042) );
  NAND2_X1 U10419 ( .A1(n14042), .A2(n12158), .ZN(n10134) );
  INV_X1 U10420 ( .A(n10134), .ZN(n8058) );
  AND2_X1 U10421 ( .A1(n13722), .A2(n14590), .ZN(n8059) );
  NAND2_X1 U10422 ( .A1(n10135), .A2(n11891), .ZN(n8061) );
  NAND2_X1 U10423 ( .A1(n10566), .A2(n7516), .ZN(n8060) );
  NAND2_X1 U10424 ( .A1(n8061), .A2(n8060), .ZN(n10355) );
  NAND2_X1 U10425 ( .A1(n6646), .A2(n10579), .ZN(n8062) );
  NOR2_X1 U10426 ( .A1(n11713), .A2(n13720), .ZN(n8064) );
  NAND2_X1 U10427 ( .A1(n11713), .A2(n13720), .ZN(n8063) );
  NAND2_X1 U10428 ( .A1(n11721), .A2(n10580), .ZN(n8065) );
  OR2_X1 U10429 ( .A1(n11725), .A2(n11062), .ZN(n8066) );
  NAND2_X1 U10430 ( .A1(n11725), .A2(n11062), .ZN(n8067) );
  INV_X1 U10431 ( .A(n13717), .ZN(n11055) );
  AND2_X1 U10432 ( .A1(n11734), .A2(n11055), .ZN(n8068) );
  INV_X1 U10433 ( .A(n13716), .ZN(n8069) );
  OR2_X1 U10434 ( .A1(n11739), .A2(n8069), .ZN(n8070) );
  NAND2_X1 U10435 ( .A1(n11748), .A2(n11474), .ZN(n8073) );
  NAND2_X1 U10436 ( .A1(n10958), .A2(n8073), .ZN(n11085) );
  INV_X1 U10437 ( .A(n11085), .ZN(n8074) );
  OR2_X1 U10438 ( .A1(n11757), .A2(n14476), .ZN(n8075) );
  INV_X1 U10439 ( .A(n11904), .ZN(n8076) );
  INV_X1 U10440 ( .A(n13712), .ZN(n14479) );
  OR2_X1 U10441 ( .A1(n11768), .A2(n14479), .ZN(n8078) );
  INV_X1 U10442 ( .A(n13711), .ZN(n14452) );
  OR2_X1 U10443 ( .A1(n12040), .A2(n14452), .ZN(n8079) );
  XNOR2_X1 U10444 ( .A(n14472), .B(n13708), .ZN(n11908) );
  INV_X1 U10445 ( .A(n13708), .ZN(n8080) );
  NAND2_X1 U10446 ( .A1(n14472), .A2(n8080), .ZN(n8081) );
  INV_X1 U10447 ( .A(n13707), .ZN(n14463) );
  OR2_X1 U10448 ( .A1(n13623), .A2(n14463), .ZN(n8082) );
  NAND2_X1 U10449 ( .A1(n11798), .A2(n11789), .ZN(n14024) );
  INV_X1 U10450 ( .A(n14007), .ZN(n8083) );
  OR2_X1 U10451 ( .A1(n14125), .A2(n8083), .ZN(n8084) );
  INV_X1 U10452 ( .A(n13984), .ZN(n14022) );
  NAND2_X1 U10453 ( .A1(n14119), .A2(n14022), .ZN(n8087) );
  INV_X1 U10454 ( .A(n11914), .ZN(n13993) );
  INV_X1 U10455 ( .A(n13598), .ZN(n14009) );
  NAND2_X1 U10456 ( .A1(n13991), .A2(n14009), .ZN(n8088) );
  NAND2_X1 U10457 ( .A1(n13971), .A2(n13983), .ZN(n8090) );
  INV_X1 U10458 ( .A(n13706), .ZN(n13597) );
  NAND2_X1 U10459 ( .A1(n14104), .A2(n13597), .ZN(n8091) );
  OR2_X1 U10460 ( .A1(n13943), .A2(n13705), .ZN(n8092) );
  INV_X1 U10461 ( .A(n13914), .ZN(n13918) );
  INV_X1 U10462 ( .A(n13898), .ZN(n13901) );
  INV_X1 U10463 ( .A(n13704), .ZN(n13604) );
  NOR2_X1 U10464 ( .A1(n13928), .A2(n13604), .ZN(n13902) );
  INV_X1 U10465 ( .A(n14084), .ZN(n8093) );
  NOR2_X1 U10466 ( .A1(n8093), .A2(n13886), .ZN(n13882) );
  INV_X1 U10467 ( .A(n13873), .ZN(n13859) );
  NAND2_X1 U10468 ( .A1(n13861), .A2(n8096), .ZN(n8097) );
  XNOR2_X1 U10469 ( .A(n8097), .B(n11920), .ZN(n8100) );
  NAND2_X1 U10470 ( .A1(n14590), .A2(n11694), .ZN(n10560) );
  NAND2_X1 U10471 ( .A1(n10353), .A2(n10354), .ZN(n10394) );
  OR2_X1 U10472 ( .A1(n10394), .A2(n11715), .ZN(n10539) );
  NAND2_X1 U10473 ( .A1(n11038), .A2(n14622), .ZN(n11037) );
  NOR2_X2 U10474 ( .A1(n11457), .A2(n14507), .ZN(n11456) );
  AND2_X2 U10475 ( .A1(n6497), .A2(n13991), .ZN(n13987) );
  OR2_X2 U10476 ( .A1(n14075), .A2(n13880), .ZN(n13867) );
  INV_X1 U10477 ( .A(n8109), .ZN(n8101) );
  INV_X1 U10478 ( .A(n14043), .ZN(n11691) );
  NAND2_X1 U10479 ( .A1(n11691), .A2(n8102), .ZN(n11925) );
  OR2_X1 U10480 ( .A1(n11925), .A2(n14168), .ZN(n9937) );
  INV_X1 U10481 ( .A(n9937), .ZN(n8103) );
  NOR2_X1 U10482 ( .A1(n14011), .A2(n8104), .ZN(n8111) );
  INV_X1 U10483 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8107) );
  AOI22_X1 U10484 ( .A1(n7538), .A2(P1_REG2_REG_30__SCAN_IN), .B1(n8105), .B2(
        P1_REG0_REG_30__SCAN_IN), .ZN(n8106) );
  OAI21_X1 U10485 ( .B1(n7561), .B2(n8107), .A(n8106), .ZN(n13701) );
  INV_X1 U10486 ( .A(n13701), .ZN(n14062) );
  INV_X1 U10487 ( .A(P1_B_REG_SCAN_IN), .ZN(n8108) );
  INV_X1 U10488 ( .A(n8098), .ZN(n13726) );
  OAI21_X1 U10489 ( .B1(n14157), .B2(n8108), .A(n14008), .ZN(n14061) );
  NOR3_X1 U10490 ( .A1(n14062), .A2(n14061), .A3(n8109), .ZN(n8110) );
  AOI211_X1 U10491 ( .C1(n14041), .C2(P1_REG2_REG_29__SCAN_IN), .A(n8111), .B(
        n8110), .ZN(n8112) );
  OAI21_X1 U10492 ( .B1(n6894), .B2(n14035), .A(n8112), .ZN(n8113) );
  NOR2_X4 U10493 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8175) );
  AND4_X2 U10494 ( .A1(n8119), .A2(n8118), .A3(n8200), .A4(n8220), .ZN(n8120)
         );
  NOR2_X2 U10495 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n8126) );
  NOR2_X2 U10496 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8125) );
  NOR2_X2 U10497 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8124) );
  NOR2_X1 U10498 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8128) );
  NOR2_X1 U10499 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8127) );
  NOR2_X2 U10500 ( .A1(n8294), .A2(n8130), .ZN(n8135) );
  NAND2_X1 U10501 ( .A1(n8154), .A2(n8149), .ZN(n8131) );
  NAND2_X1 U10502 ( .A1(n8132), .A2(n8131), .ZN(n8134) );
  NOR2_X1 U10503 ( .A1(n8135), .A2(n8154), .ZN(n8138) );
  INV_X1 U10504 ( .A(n8139), .ZN(n8140) );
  XNOR2_X1 U10505 ( .A(n8148), .B(n8666), .ZN(n8147) );
  INV_X1 U10506 ( .A(n8143), .ZN(n8144) );
  NOR2_X2 U10507 ( .A1(n8294), .A2(n8144), .ZN(n8386) );
  NAND2_X1 U10508 ( .A1(n8386), .A2(n8145), .ZN(n8401) );
  XNOR2_X2 U10509 ( .A(n8146), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10480) );
  AND2_X2 U10510 ( .A1(n10480), .A2(n11023), .ZN(n8670) );
  NAND2_X1 U10511 ( .A1(n8670), .A2(n8148), .ZN(n14805) );
  XNOR2_X2 U10512 ( .A(n8156), .B(n8155), .ZN(n8159) );
  INV_X1 U10513 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10283) );
  INV_X1 U10514 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8158) );
  AND2_X2 U10515 ( .A1(n8159), .A2(n13541), .ZN(n8456) );
  NAND2_X1 U10516 ( .A1(n8456), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U10517 ( .A1(n9735), .A2(SI_0_), .ZN(n8165) );
  XNOR2_X1 U10518 ( .A(n8165), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13561) );
  XNOR2_X2 U10519 ( .A(n8167), .B(n8153), .ZN(n13547) );
  NAND2_X1 U10520 ( .A1(n13131), .A2(n8554), .ZN(n10244) );
  NAND2_X1 U10521 ( .A1(n8456), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8173) );
  INV_X1 U10522 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8168) );
  INV_X1 U10523 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8169) );
  INV_X1 U10524 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9861) );
  NAND4_X1 U10525 ( .A1(n8173), .A2(n8172), .A3(n8171), .A4(n8170), .ZN(n10024) );
  NAND2_X1 U10526 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n14663), .ZN(n8174) );
  INV_X1 U10527 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U10528 ( .A1(n9868), .A2(n9735), .ZN(n8185) );
  OR2_X1 U10529 ( .A1(n8185), .A2(n9760), .ZN(n8178) );
  INV_X1 U10530 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9711) );
  INV_X1 U10531 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10690) );
  OR2_X1 U10532 ( .A1(n8545), .A2(n10690), .ZN(n8184) );
  NAND2_X1 U10533 ( .A1(n8456), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8183) );
  INV_X1 U10534 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9877) );
  OR2_X1 U10535 ( .A1(n8489), .A2(n9877), .ZN(n8182) );
  INV_X1 U10536 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8180) );
  OR2_X1 U10537 ( .A1(n8844), .A2(n8180), .ZN(n8181) );
  NAND4_X2 U10538 ( .A1(n8184), .A2(n8183), .A3(n8182), .A4(n8181), .ZN(n13128) );
  OR2_X1 U10539 ( .A1(n8864), .A2(n9721), .ZN(n8192) );
  NAND2_X1 U10540 ( .A1(n9720), .A2(n8206), .ZN(n8191) );
  NOR2_X1 U10541 ( .A1(n8175), .A2(n8154), .ZN(n8186) );
  MUX2_X1 U10542 ( .A(n8154), .B(n8186), .S(P2_IR_REG_2__SCAN_IN), .Z(n8187)
         );
  INV_X1 U10543 ( .A(n8187), .ZN(n8190) );
  INV_X1 U10544 ( .A(n8188), .ZN(n8189) );
  NAND2_X1 U10545 ( .A1(n8190), .A2(n8189), .ZN(n10004) );
  INV_X1 U10546 ( .A(n13128), .ZN(n8557) );
  NAND2_X1 U10547 ( .A1(n8557), .A2(n10689), .ZN(n8193) );
  NAND2_X1 U10548 ( .A1(n10261), .A2(n8193), .ZN(n10302) );
  NAND2_X1 U10549 ( .A1(n8456), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8198) );
  OR2_X1 U10550 ( .A1(n8545), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8197) );
  INV_X1 U10551 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9879) );
  OR2_X1 U10552 ( .A1(n8489), .A2(n9879), .ZN(n8196) );
  INV_X1 U10553 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8194) );
  OR2_X1 U10554 ( .A1(n8844), .A2(n8194), .ZN(n8195) );
  NAND4_X1 U10555 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(n13127) );
  NAND2_X1 U10556 ( .A1(n9724), .A2(n6474), .ZN(n8203) );
  INV_X2 U10557 ( .A(n8864), .ZN(n8424) );
  INV_X2 U10558 ( .A(n9868), .ZN(n8423) );
  NOR2_X1 U10559 ( .A1(n8188), .A2(n8154), .ZN(n8199) );
  MUX2_X1 U10560 ( .A(n8154), .B(n8199), .S(P2_IR_REG_3__SCAN_IN), .Z(n8201)
         );
  AND2_X1 U10561 ( .A1(n8188), .A2(n8200), .ZN(n8207) );
  AOI22_X1 U10562 ( .A1(n8424), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8423), .B2(
        n9880), .ZN(n8202) );
  NAND2_X1 U10563 ( .A1(n10302), .A2(n10306), .ZN(n10301) );
  INV_X1 U10564 ( .A(n13127), .ZN(n8560) );
  NAND2_X1 U10565 ( .A1(n8204), .A2(n8560), .ZN(n8205) );
  NAND2_X1 U10566 ( .A1(n10301), .A2(n8205), .ZN(n10406) );
  NAND2_X1 U10567 ( .A1(n9722), .A2(n6479), .ZN(n8212) );
  INV_X1 U10568 ( .A(n8207), .ZN(n8209) );
  NAND2_X1 U10569 ( .A1(n8209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8208) );
  MUX2_X1 U10570 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8208), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8210) );
  AOI22_X1 U10571 ( .A1(n8424), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8423), .B2(
        n9881), .ZN(n8211) );
  NAND2_X1 U10572 ( .A1(n8615), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8216) );
  INV_X1 U10573 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10479) );
  OR2_X1 U10574 ( .A1(n8844), .A2(n10479), .ZN(n8215) );
  AND2_X1 U10575 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8225) );
  INV_X1 U10576 ( .A(n8225), .ZN(n8227) );
  OAI21_X1 U10577 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8227), .ZN(n10483) );
  OR2_X1 U10578 ( .A1(n8545), .A2(n10483), .ZN(n8214) );
  INV_X1 U10579 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8213) );
  INV_X1 U10580 ( .A(n8905), .ZN(n10410) );
  NAND2_X1 U10581 ( .A1(n10406), .A2(n10410), .ZN(n10405) );
  OR2_X1 U10582 ( .A1(n10413), .A2(n13126), .ZN(n8217) );
  NAND2_X1 U10583 ( .A1(n9726), .A2(n6479), .ZN(n8224) );
  NAND2_X1 U10584 ( .A1(n8219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U10585 ( .A(n8218), .B(P2_IR_REG_31__SCAN_IN), .S(n8220), .Z(n8222)
         );
  INV_X1 U10586 ( .A(n8219), .ZN(n8221) );
  NAND2_X1 U10587 ( .A1(n8221), .A2(n8220), .ZN(n8248) );
  NAND2_X1 U10588 ( .A1(n8222), .A2(n8248), .ZN(n10093) );
  INV_X1 U10589 ( .A(n10093), .ZN(n9882) );
  AOI22_X1 U10590 ( .A1(n8424), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8423), .B2(
        n9882), .ZN(n8223) );
  NAND2_X1 U10591 ( .A1(n8224), .A2(n8223), .ZN(n14796) );
  NAND2_X1 U10592 ( .A1(n8615), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8233) );
  INV_X1 U10593 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10522) );
  OR2_X1 U10594 ( .A1(n6655), .A2(n10522), .ZN(n8232) );
  NAND2_X1 U10595 ( .A1(n8225), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8240) );
  INV_X1 U10596 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10597 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  NAND2_X1 U10598 ( .A1(n8240), .A2(n8228), .ZN(n10524) );
  OR2_X1 U10599 ( .A1(n6666), .A2(n10524), .ZN(n8231) );
  INV_X1 U10600 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8229) );
  OR2_X1 U10601 ( .A1(n8842), .A2(n8229), .ZN(n8230) );
  NAND4_X1 U10602 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8230), .ZN(n13125) );
  NAND2_X1 U10603 ( .A1(n14796), .A2(n13125), .ZN(n8234) );
  OR2_X1 U10604 ( .A1(n14796), .A2(n13125), .ZN(n8235) );
  NAND2_X1 U10605 ( .A1(n9749), .A2(n6479), .ZN(n8238) );
  NAND2_X1 U10606 ( .A1(n8248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8236) );
  XNOR2_X1 U10607 ( .A(n8236), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U10608 ( .A1(n8424), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8423), .B2(
        n9883), .ZN(n8237) );
  NAND2_X1 U10609 ( .A1(n8615), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8246) );
  INV_X1 U10610 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10676) );
  OR2_X1 U10611 ( .A1(n6655), .A2(n10676), .ZN(n8245) );
  INV_X1 U10612 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8239) );
  NOR2_X1 U10613 ( .A1(n8240), .A2(n8239), .ZN(n8253) );
  INV_X1 U10614 ( .A(n8253), .ZN(n8255) );
  NAND2_X1 U10615 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U10616 ( .A1(n8255), .A2(n8241), .ZN(n10668) );
  OR2_X1 U10617 ( .A1(n6666), .A2(n10668), .ZN(n8244) );
  INV_X1 U10618 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8242) );
  OR2_X1 U10619 ( .A1(n8842), .A2(n8242), .ZN(n8243) );
  NAND4_X1 U10620 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n13124) );
  INV_X1 U10621 ( .A(n13124), .ZN(n8566) );
  XNOR2_X1 U10622 ( .A(n14803), .B(n8566), .ZN(n10672) );
  NAND2_X1 U10623 ( .A1(n14803), .A2(n13124), .ZN(n8247) );
  NAND2_X1 U10624 ( .A1(n10663), .A2(n8247), .ZN(n10848) );
  NAND2_X1 U10625 ( .A1(n9764), .A2(n6479), .ZN(n8251) );
  OAI21_X1 U10626 ( .B1(n8248), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U10627 ( .A(n8249), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U10628 ( .A1(n8424), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8423), .B2(
        n9971), .ZN(n8250) );
  NAND2_X1 U10629 ( .A1(n8251), .A2(n8250), .ZN(n10852) );
  NAND2_X1 U10630 ( .A1(n8615), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8260) );
  INV_X1 U10631 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8252) );
  OR2_X1 U10632 ( .A1(n6655), .A2(n8252), .ZN(n8259) );
  NAND2_X1 U10633 ( .A1(n8253), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8272) );
  INV_X1 U10634 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10635 ( .A1(n8255), .A2(n8254), .ZN(n8256) );
  NAND2_X1 U10636 ( .A1(n8272), .A2(n8256), .ZN(n10850) );
  OR2_X1 U10637 ( .A1(n6666), .A2(n10850), .ZN(n8258) );
  INV_X1 U10638 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9884) );
  OR2_X1 U10639 ( .A1(n8842), .A2(n9884), .ZN(n8257) );
  NAND4_X1 U10640 ( .A1(n8260), .A2(n8259), .A3(n8258), .A4(n8257), .ZN(n13123) );
  OR2_X1 U10641 ( .A1(n10852), .A2(n13123), .ZN(n8261) );
  NAND2_X1 U10642 ( .A1(n10848), .A2(n8261), .ZN(n8263) );
  NAND2_X1 U10643 ( .A1(n10852), .A2(n13123), .ZN(n8262) );
  NAND2_X1 U10644 ( .A1(n8263), .A2(n8262), .ZN(n10977) );
  NAND2_X1 U10645 ( .A1(n9775), .A2(n6479), .ZN(n8269) );
  NOR2_X1 U10646 ( .A1(n8264), .A2(n8154), .ZN(n8265) );
  MUX2_X1 U10647 ( .A(n8154), .B(n8265), .S(P2_IR_REG_8__SCAN_IN), .Z(n8267)
         );
  NOR2_X1 U10648 ( .A1(n8267), .A2(n8123), .ZN(n9972) );
  AOI22_X1 U10649 ( .A1(n8424), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8423), .B2(
        n9972), .ZN(n8268) );
  NAND2_X1 U10650 ( .A1(n8520), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8278) );
  INV_X1 U10651 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8270) );
  OR2_X1 U10652 ( .A1(n8845), .A2(n8270), .ZN(n8277) );
  INV_X1 U10653 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U10654 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  NAND2_X1 U10655 ( .A1(n8287), .A2(n8273), .ZN(n10988) );
  OR2_X1 U10656 ( .A1(n6666), .A2(n10988), .ZN(n8276) );
  INV_X1 U10657 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8274) );
  OR2_X1 U10658 ( .A1(n8842), .A2(n8274), .ZN(n8275) );
  NAND4_X1 U10659 ( .A1(n8278), .A2(n8277), .A3(n8276), .A4(n8275), .ZN(n13122) );
  INV_X1 U10660 ( .A(n13122), .ZN(n8279) );
  NAND2_X1 U10661 ( .A1(n14820), .A2(n8279), .ZN(n8569) );
  OR2_X1 U10662 ( .A1(n14820), .A2(n8279), .ZN(n8280) );
  NAND2_X1 U10663 ( .A1(n8569), .A2(n8280), .ZN(n8908) );
  NAND2_X1 U10664 ( .A1(n10977), .A2(n8908), .ZN(n8282) );
  NAND2_X1 U10665 ( .A1(n14820), .A2(n13122), .ZN(n8281) );
  NAND2_X1 U10666 ( .A1(n8282), .A2(n8281), .ZN(n10881) );
  NAND2_X1 U10667 ( .A1(n9857), .A2(n6479), .ZN(n8285) );
  NAND2_X1 U10668 ( .A1(n8266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8283) );
  XNOR2_X1 U10669 ( .A(n8283), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U10670 ( .A1(n8424), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8423), .B2(
        n10221), .ZN(n8284) );
  NAND2_X2 U10671 ( .A1(n8285), .A2(n8284), .ZN(n11112) );
  NAND2_X1 U10672 ( .A1(n8520), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8292) );
  INV_X1 U10673 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8286) );
  OR2_X1 U10674 ( .A1(n8845), .A2(n8286), .ZN(n8291) );
  INV_X1 U10675 ( .A(n8298), .ZN(n8300) );
  NAND2_X1 U10676 ( .A1(n8287), .A2(n11108), .ZN(n8288) );
  NAND2_X1 U10677 ( .A1(n8300), .A2(n8288), .ZN(n11107) );
  OR2_X1 U10678 ( .A1(n6666), .A2(n11107), .ZN(n8290) );
  INV_X1 U10679 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9975) );
  OR2_X1 U10680 ( .A1(n8842), .A2(n9975), .ZN(n8289) );
  NAND4_X1 U10681 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n13120) );
  XNOR2_X1 U10682 ( .A(n11112), .B(n13120), .ZN(n10882) );
  INV_X1 U10683 ( .A(n10882), .ZN(n10884) );
  NAND2_X1 U10684 ( .A1(n11112), .A2(n13120), .ZN(n8293) );
  NAND2_X1 U10685 ( .A1(n9910), .A2(n6479), .ZN(n8297) );
  NAND2_X1 U10686 ( .A1(n8631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8295) );
  XNOR2_X1 U10687 ( .A(n8295), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U10688 ( .A1(n8424), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8423), 
        .B2(n10293), .ZN(n8296) );
  NAND2_X1 U10689 ( .A1(n8615), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8306) );
  INV_X1 U10690 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11016) );
  OR2_X1 U10691 ( .A1(n6655), .A2(n11016), .ZN(n8305) );
  INV_X1 U10692 ( .A(n8312), .ZN(n8314) );
  INV_X1 U10693 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10694 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  NAND2_X1 U10695 ( .A1(n8314), .A2(n8301), .ZN(n11144) );
  OR2_X1 U10696 ( .A1(n6666), .A2(n11144), .ZN(n8304) );
  INV_X1 U10697 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8302) );
  OR2_X1 U10698 ( .A1(n8842), .A2(n8302), .ZN(n8303) );
  NAND4_X1 U10699 ( .A1(n8306), .A2(n8305), .A3(n8304), .A4(n8303), .ZN(n13119) );
  XNOR2_X1 U10700 ( .A(n11133), .B(n13119), .ZN(n11006) );
  INV_X1 U10701 ( .A(n11006), .ZN(n11008) );
  NAND2_X1 U10702 ( .A1(n9964), .A2(n6479), .ZN(n8310) );
  NOR2_X1 U10703 ( .A1(n8631), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8323) );
  INV_X1 U10704 ( .A(n8323), .ZN(n8307) );
  NAND2_X1 U10705 ( .A1(n8307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8308) );
  XNOR2_X1 U10706 ( .A(n8308), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U10707 ( .A1(n8424), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8423), 
        .B2(n13143), .ZN(n8309) );
  NAND2_X1 U10708 ( .A1(n8520), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8320) );
  INV_X1 U10709 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8311) );
  OR2_X1 U10710 ( .A1(n8845), .A2(n8311), .ZN(n8319) );
  NAND2_X1 U10711 ( .A1(n8312), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8332) );
  INV_X1 U10712 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U10713 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U10714 ( .A1(n8332), .A2(n8315), .ZN(n11267) );
  OR2_X1 U10715 ( .A1(n6666), .A2(n11267), .ZN(n8318) );
  INV_X1 U10716 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8316) );
  OR2_X1 U10717 ( .A1(n8842), .A2(n8316), .ZN(n8317) );
  NAND4_X1 U10718 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(n13118) );
  AND2_X1 U10719 ( .A1(n11263), .A2(n13118), .ZN(n8321) );
  NAND2_X1 U10720 ( .A1(n10020), .A2(n6479), .ZN(n8330) );
  INV_X1 U10721 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8322) );
  AND2_X1 U10722 ( .A1(n8323), .A2(n8322), .ZN(n8327) );
  INV_X1 U10723 ( .A(n8327), .ZN(n8324) );
  NAND2_X1 U10724 ( .A1(n8324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8325) );
  MUX2_X1 U10725 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8325), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8328) );
  INV_X1 U10726 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8326) );
  AND2_X1 U10727 ( .A1(n8327), .A2(n8326), .ZN(n8345) );
  INV_X1 U10728 ( .A(n8345), .ZN(n8342) );
  AOI22_X1 U10729 ( .A1(n8424), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8423), 
        .B2(n13144), .ZN(n8329) );
  NAND2_X2 U10730 ( .A1(n8330), .A2(n8329), .ZN(n14439) );
  NAND2_X1 U10731 ( .A1(n8615), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8338) );
  INV_X1 U10732 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13134) );
  OR2_X1 U10733 ( .A1(n6655), .A2(n13134), .ZN(n8337) );
  INV_X1 U10734 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10735 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  NAND2_X1 U10736 ( .A1(n8350), .A2(n8333), .ZN(n11406) );
  OR2_X1 U10737 ( .A1(n6666), .A2(n11406), .ZN(n8336) );
  INV_X1 U10738 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8334) );
  OR2_X1 U10739 ( .A1(n8842), .A2(n8334), .ZN(n8335) );
  NAND4_X1 U10740 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n13117) );
  NOR2_X1 U10741 ( .A1(n14439), .A2(n13117), .ZN(n8339) );
  OR2_X2 U10742 ( .A1(n11213), .A2(n8339), .ZN(n8341) );
  NAND2_X1 U10743 ( .A1(n14439), .A2(n13117), .ZN(n8340) );
  NAND2_X1 U10744 ( .A1(n10212), .A2(n6479), .ZN(n8349) );
  NAND2_X1 U10745 ( .A1(n8342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8343) );
  MUX2_X1 U10746 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8343), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8346) );
  INV_X1 U10747 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U10748 ( .A1(n8345), .A2(n8344), .ZN(n8370) );
  NAND2_X1 U10749 ( .A1(n8346), .A2(n8370), .ZN(n14693) );
  INV_X1 U10750 ( .A(n14693), .ZN(n8347) );
  AOI22_X1 U10751 ( .A1(n8424), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8347), 
        .B2(n8423), .ZN(n8348) );
  NAND2_X1 U10752 ( .A1(n8615), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8355) );
  INV_X1 U10753 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13152) );
  OR2_X1 U10754 ( .A1(n6655), .A2(n13152), .ZN(n8354) );
  NAND2_X1 U10755 ( .A1(n8350), .A2(n11442), .ZN(n8351) );
  NAND2_X1 U10756 ( .A1(n8361), .A2(n8351), .ZN(n11443) );
  OR2_X1 U10757 ( .A1(n6666), .A2(n11443), .ZN(n8353) );
  INV_X1 U10758 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13168) );
  OR2_X1 U10759 ( .A1(n8842), .A2(n13168), .ZN(n8352) );
  NAND4_X1 U10760 ( .A1(n8355), .A2(n8354), .A3(n8353), .A4(n8352), .ZN(n13116) );
  AND2_X1 U10761 ( .A1(n11431), .A2(n13116), .ZN(n8357) );
  OR2_X1 U10762 ( .A1(n11431), .A2(n13116), .ZN(n8356) );
  NAND2_X1 U10763 ( .A1(n10387), .A2(n6479), .ZN(n8360) );
  NAND2_X1 U10764 ( .A1(n8370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8358) );
  XNOR2_X1 U10765 ( .A(n8358), .B(n8369), .ZN(n14710) );
  AOI22_X1 U10766 ( .A1(n8424), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n14710), 
        .B2(n8423), .ZN(n8359) );
  NAND2_X1 U10767 ( .A1(n8615), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8367) );
  INV_X1 U10768 ( .A(n8374), .ZN(n8376) );
  NAND2_X1 U10769 ( .A1(n8361), .A2(n11566), .ZN(n8362) );
  NAND2_X1 U10770 ( .A1(n8376), .A2(n8362), .ZN(n11563) );
  OR2_X1 U10771 ( .A1(n6666), .A2(n11563), .ZN(n8366) );
  INV_X1 U10772 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13169) );
  OR2_X1 U10773 ( .A1(n8842), .A2(n13169), .ZN(n8365) );
  INV_X1 U10774 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8363) );
  OR2_X1 U10775 ( .A1(n6655), .A2(n8363), .ZN(n8364) );
  NAND4_X1 U10776 ( .A1(n8367), .A2(n8366), .A3(n8365), .A4(n8364), .ZN(n13115) );
  OR2_X1 U10777 ( .A1(n14412), .A2(n13115), .ZN(n8912) );
  NAND2_X1 U10778 ( .A1(n14412), .A2(n13115), .ZN(n14404) );
  INV_X1 U10779 ( .A(n8368), .ZN(n11612) );
  NAND2_X1 U10780 ( .A1(n10469), .A2(n6479), .ZN(n8373) );
  OAI21_X1 U10781 ( .B1(n8370), .B2(n8369), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8371) );
  XNOR2_X1 U10782 ( .A(n8371), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14715) );
  AOI22_X1 U10783 ( .A1(n14715), .A2(n8423), .B1(n8424), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10784 ( .A1(n8374), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8392) );
  INV_X1 U10785 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10786 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  NAND2_X1 U10787 ( .A1(n8392), .A2(n8377), .ZN(n13088) );
  OR2_X1 U10788 ( .A1(n13088), .A2(n6666), .ZN(n8383) );
  INV_X1 U10789 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11618) );
  OR2_X1 U10790 ( .A1(n6655), .A2(n11618), .ZN(n8382) );
  INV_X1 U10791 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8378) );
  OR2_X1 U10792 ( .A1(n8845), .A2(n8378), .ZN(n8381) );
  INV_X1 U10793 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8379) );
  OR2_X1 U10794 ( .A1(n8842), .A2(n8379), .ZN(n8380) );
  NAND4_X1 U10795 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n13114) );
  XNOR2_X1 U10796 ( .A(n13096), .B(n13114), .ZN(n11613) );
  OR2_X1 U10797 ( .A1(n13096), .A2(n13114), .ZN(n8385) );
  NAND2_X1 U10798 ( .A1(n10383), .A2(n6479), .ZN(n8391) );
  INV_X1 U10799 ( .A(n8386), .ZN(n8387) );
  NAND2_X1 U10800 ( .A1(n8387), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8388) );
  MUX2_X1 U10801 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8388), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8389) );
  AND2_X1 U10802 ( .A1(n8401), .A2(n8389), .ZN(n14725) );
  AOI22_X1 U10803 ( .A1(n8424), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8423), 
        .B2(n14725), .ZN(n8390) );
  NAND2_X1 U10804 ( .A1(n8392), .A2(n13016), .ZN(n8393) );
  NAND2_X1 U10805 ( .A1(n8407), .A2(n8393), .ZN(n11604) );
  INV_X1 U10806 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8394) );
  OR2_X1 U10807 ( .A1(n6655), .A2(n8394), .ZN(n8397) );
  INV_X1 U10808 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8395) );
  OR2_X1 U10809 ( .A1(n8845), .A2(n8395), .ZN(n8396) );
  AND2_X1 U10810 ( .A1(n8397), .A2(n8396), .ZN(n8399) );
  NAND2_X1 U10811 ( .A1(n8614), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8398) );
  OAI211_X1 U10812 ( .C1(n11604), .C2(n6666), .A(n8399), .B(n8398), .ZN(n13113) );
  INV_X1 U10813 ( .A(n13113), .ZN(n11966) );
  XNOR2_X1 U10814 ( .A(n13488), .B(n11966), .ZN(n8911) );
  NAND2_X1 U10815 ( .A1(n13488), .A2(n13113), .ZN(n8400) );
  NAND2_X1 U10816 ( .A1(n10420), .A2(n6474), .ZN(n8405) );
  NAND2_X1 U10817 ( .A1(n8401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8402) );
  MUX2_X1 U10818 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8402), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8403) );
  AOI22_X1 U10819 ( .A1(n8424), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8423), 
        .B2(n13177), .ZN(n8404) );
  INV_X1 U10820 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13188) );
  INV_X1 U10821 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8406) );
  INV_X1 U10822 ( .A(n8431), .ZN(n8429) );
  NAND2_X1 U10823 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  NAND2_X1 U10824 ( .A1(n8429), .A2(n8408), .ZN(n11672) );
  OR2_X1 U10825 ( .A1(n11672), .A2(n6666), .ZN(n8410) );
  AOI22_X1 U10826 ( .A1(n8520), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8456), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8409) );
  OAI211_X1 U10827 ( .C1(n8842), .C2(n13188), .A(n8410), .B(n8409), .ZN(n13112) );
  XNOR2_X1 U10828 ( .A(n13482), .B(n13112), .ZN(n8913) );
  NAND2_X1 U10829 ( .A1(n13482), .A2(n13112), .ZN(n8411) );
  NAND2_X1 U10830 ( .A1(n11661), .A2(n8411), .ZN(n13397) );
  INV_X1 U10831 ( .A(n13397), .ZN(n8421) );
  NAND2_X1 U10832 ( .A1(n10843), .A2(n6479), .ZN(n8414) );
  NAND2_X1 U10833 ( .A1(n6513), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8412) );
  XNOR2_X1 U10834 ( .A(n8412), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14740) );
  AOI22_X1 U10835 ( .A1(n8424), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8423), 
        .B2(n14740), .ZN(n8413) );
  XNOR2_X1 U10836 ( .A(n8429), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13403) );
  INV_X1 U10837 ( .A(n6666), .ZN(n8455) );
  NAND2_X1 U10838 ( .A1(n13403), .A2(n8455), .ZN(n8420) );
  INV_X1 U10839 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10840 ( .A1(n8520), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10841 ( .A1(n8456), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8415) );
  OAI211_X1 U10842 ( .C1(n8417), .C2(n8842), .A(n8416), .B(n8415), .ZN(n8418)
         );
  INV_X1 U10843 ( .A(n8418), .ZN(n8419) );
  NAND2_X1 U10844 ( .A1(n8420), .A2(n8419), .ZN(n13111) );
  INV_X1 U10845 ( .A(n13111), .ZN(n8590) );
  XNOR2_X1 U10846 ( .A(n13477), .B(n8590), .ZN(n8916) );
  NAND2_X1 U10847 ( .A1(n8421), .A2(n8916), .ZN(n13395) );
  OR2_X1 U10848 ( .A1(n13477), .A2(n13111), .ZN(n8422) );
  NAND2_X1 U10849 ( .A1(n10952), .A2(n6474), .ZN(n8426) );
  AOI22_X1 U10850 ( .A1(n8424), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6641), 
        .B2(n8423), .ZN(n8425) );
  INV_X1 U10851 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8428) );
  INV_X1 U10852 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8427) );
  OAI21_X1 U10853 ( .B1(n8429), .B2(n8428), .A(n8427), .ZN(n8433) );
  AND2_X1 U10854 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8430) );
  INV_X1 U10855 ( .A(n8442), .ZN(n8432) );
  AND2_X1 U10856 ( .A1(n8433), .A2(n8432), .ZN(n13384) );
  NAND2_X1 U10857 ( .A1(n13384), .A2(n8455), .ZN(n8438) );
  INV_X1 U10858 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13472) );
  NAND2_X1 U10859 ( .A1(n8520), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10860 ( .A1(n8615), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8434) );
  OAI211_X1 U10861 ( .C1(n13472), .C2(n8842), .A(n8435), .B(n8434), .ZN(n8436)
         );
  INV_X1 U10862 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U10863 ( .A1(n8438), .A2(n8437), .ZN(n13110) );
  NOR2_X1 U10864 ( .A1(n13383), .A2(n13110), .ZN(n8439) );
  INV_X1 U10865 ( .A(n13110), .ZN(n8592) );
  NAND2_X1 U10866 ( .A1(n11022), .A2(n6474), .ZN(n8441) );
  OR2_X1 U10867 ( .A1(n6681), .A2(n11024), .ZN(n8440) );
  NOR2_X1 U10868 ( .A1(n8442), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8443) );
  OR2_X1 U10869 ( .A1(n8453), .A2(n8443), .ZN(n13046) );
  INV_X1 U10870 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10871 ( .A1(n8456), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10872 ( .A1(n8614), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8444) );
  OAI211_X1 U10873 ( .C1(n6655), .C2(n8446), .A(n8445), .B(n8444), .ZN(n8447)
         );
  INV_X1 U10874 ( .A(n8447), .ZN(n8448) );
  OAI21_X1 U10875 ( .B1(n13046), .B2(n6666), .A(n8448), .ZN(n13109) );
  AND2_X1 U10876 ( .A1(n13465), .A2(n13109), .ZN(n8449) );
  OR2_X1 U10877 ( .A1(n13465), .A2(n13109), .ZN(n8450) );
  NAND2_X1 U10878 ( .A1(n11074), .A2(n6479), .ZN(n8452) );
  OR2_X1 U10879 ( .A1(n6681), .A2(n11076), .ZN(n8451) );
  OR2_X1 U10880 ( .A1(n8453), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10881 ( .A1(n8453), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8468) );
  AND2_X1 U10882 ( .A1(n8454), .A2(n8468), .ZN(n13349) );
  NAND2_X1 U10883 ( .A1(n13349), .A2(n8455), .ZN(n8462) );
  INV_X1 U10884 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10885 ( .A1(n8614), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10886 ( .A1(n8615), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8457) );
  OAI211_X1 U10887 ( .C1(n6655), .C2(n8459), .A(n8458), .B(n8457), .ZN(n8460)
         );
  INV_X1 U10888 ( .A(n8460), .ZN(n8461) );
  NAND2_X1 U10889 ( .A1(n8462), .A2(n8461), .ZN(n13108) );
  XNOR2_X1 U10890 ( .A(n13348), .B(n13108), .ZN(n13342) );
  INV_X1 U10891 ( .A(n13342), .ZN(n13339) );
  NOR2_X1 U10892 ( .A1(n13348), .A2(n13108), .ZN(n8463) );
  XNOR2_X1 U10893 ( .A(n8465), .B(n8464), .ZN(n11172) );
  NAND2_X1 U10894 ( .A1(n11172), .A2(n6474), .ZN(n8467) );
  OR2_X1 U10895 ( .A1(n6681), .A2(n11174), .ZN(n8466) );
  NAND2_X1 U10896 ( .A1(n8520), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8473) );
  INV_X1 U10897 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13521) );
  OR2_X1 U10898 ( .A1(n8845), .A2(n13521), .ZN(n8472) );
  OAI21_X1 U10899 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8469), .A(n8478), .ZN(
        n13330) );
  OR2_X1 U10900 ( .A1(n6666), .A2(n13330), .ZN(n8471) );
  INV_X1 U10901 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13457) );
  OR2_X1 U10902 ( .A1(n8842), .A2(n13457), .ZN(n8470) );
  NAND4_X1 U10903 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(n13107) );
  XNOR2_X1 U10904 ( .A(n13332), .B(n13107), .ZN(n8917) );
  NAND2_X1 U10905 ( .A1(n13322), .A2(n13323), .ZN(n13321) );
  NAND2_X1 U10906 ( .A1(n13332), .A2(n13107), .ZN(n8474) );
  NAND2_X1 U10907 ( .A1(n11390), .A2(n6479), .ZN(n8476) );
  INV_X1 U10908 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11393) );
  OR2_X1 U10909 ( .A1(n6681), .A2(n11393), .ZN(n8475) );
  NAND2_X1 U10910 ( .A1(n8520), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8484) );
  INV_X1 U10911 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13517) );
  OR2_X1 U10912 ( .A1(n8845), .A2(n13517), .ZN(n8483) );
  INV_X1 U10913 ( .A(n8478), .ZN(n8480) );
  INV_X1 U10914 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8477) );
  INV_X1 U10915 ( .A(n8488), .ZN(n8479) );
  OAI21_X1 U10916 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8480), .A(n8479), .ZN(
        n13306) );
  OR2_X1 U10917 ( .A1(n6666), .A2(n13306), .ZN(n8482) );
  INV_X1 U10918 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13451) );
  OR2_X1 U10919 ( .A1(n8842), .A2(n13451), .ZN(n8481) );
  NAND4_X1 U10920 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n13106) );
  NAND2_X1 U10921 ( .A1(n13313), .A2(n13106), .ZN(n8896) );
  INV_X1 U10922 ( .A(n8896), .ZN(n8485) );
  OR2_X1 U10923 ( .A1(n13313), .A2(n13106), .ZN(n8897) );
  NAND2_X1 U10924 ( .A1(n13557), .A2(n6474), .ZN(n8487) );
  INV_X1 U10925 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13560) );
  OR2_X1 U10926 ( .A1(n6681), .A2(n13560), .ZN(n8486) );
  NAND2_X1 U10927 ( .A1(n8520), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8493) );
  INV_X1 U10928 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13513) );
  OR2_X1 U10929 ( .A1(n8845), .A2(n13513), .ZN(n8492) );
  NAND2_X1 U10930 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8488), .ZN(n8500) );
  OAI21_X1 U10931 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8488), .A(n8500), .ZN(
        n13299) );
  OR2_X1 U10932 ( .A1(n6666), .A2(n13299), .ZN(n8491) );
  INV_X1 U10933 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13446) );
  OR2_X1 U10934 ( .A1(n8842), .A2(n13446), .ZN(n8490) );
  NAND4_X1 U10935 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), .ZN(n13105) );
  INV_X1 U10936 ( .A(n13105), .ZN(n12980) );
  XNOR2_X1 U10937 ( .A(n13441), .B(n12980), .ZN(n13294) );
  INV_X1 U10938 ( .A(n13294), .ZN(n8600) );
  NAND2_X1 U10939 ( .A1(n13441), .A2(n13105), .ZN(n8494) );
  NAND2_X1 U10940 ( .A1(n13554), .A2(n6479), .ZN(n8497) );
  OR2_X1 U10941 ( .A1(n6681), .A2(n13556), .ZN(n8496) );
  NAND2_X1 U10942 ( .A1(n8520), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8505) );
  INV_X1 U10943 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13509) );
  OR2_X1 U10944 ( .A1(n8845), .A2(n13509), .ZN(n8504) );
  INV_X1 U10945 ( .A(n8500), .ZN(n8498) );
  INV_X1 U10946 ( .A(n8509), .ZN(n8511) );
  INV_X1 U10947 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10948 ( .A1(n8500), .A2(n8499), .ZN(n8501) );
  NAND2_X1 U10949 ( .A1(n8511), .A2(n8501), .ZN(n13282) );
  OR2_X1 U10950 ( .A1(n6666), .A2(n13282), .ZN(n8503) );
  INV_X1 U10951 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13439) );
  OR2_X1 U10952 ( .A1(n8842), .A2(n13439), .ZN(n8502) );
  NAND2_X1 U10953 ( .A1(n13511), .A2(n13079), .ZN(n8506) );
  NAND2_X1 U10954 ( .A1(n13549), .A2(n6479), .ZN(n8508) );
  OR2_X1 U10955 ( .A1(n6681), .A2(n13551), .ZN(n8507) );
  NAND2_X1 U10956 ( .A1(n8520), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8516) );
  INV_X1 U10957 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n13505) );
  OR2_X1 U10958 ( .A1(n8845), .A2(n13505), .ZN(n8515) );
  INV_X1 U10959 ( .A(n8522), .ZN(n8524) );
  INV_X1 U10960 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U10961 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  NAND2_X1 U10962 ( .A1(n8524), .A2(n8512), .ZN(n13267) );
  OR2_X1 U10963 ( .A1(n6666), .A2(n13267), .ZN(n8514) );
  INV_X1 U10964 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13433) );
  OR2_X1 U10965 ( .A1(n8842), .A2(n13433), .ZN(n8513) );
  OR2_X1 U10966 ( .A1(n13507), .A2(n13005), .ZN(n8517) );
  NAND2_X1 U10967 ( .A1(n13546), .A2(n6474), .ZN(n8519) );
  INV_X1 U10968 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13548) );
  OR2_X1 U10969 ( .A1(n6681), .A2(n13548), .ZN(n8518) );
  NAND2_X1 U10970 ( .A1(n8520), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8530) );
  INV_X1 U10971 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8521) );
  OR2_X1 U10972 ( .A1(n8845), .A2(n8521), .ZN(n8529) );
  INV_X1 U10973 ( .A(n8534), .ZN(n8536) );
  INV_X1 U10974 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10975 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  NAND2_X1 U10976 ( .A1(n8536), .A2(n8525), .ZN(n13249) );
  OR2_X1 U10977 ( .A1(n6666), .A2(n13249), .ZN(n8528) );
  INV_X1 U10978 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8526) );
  OR2_X1 U10979 ( .A1(n8842), .A2(n8526), .ZN(n8527) );
  XNOR2_X1 U10980 ( .A(n13424), .B(n13102), .ZN(n8921) );
  OR2_X1 U10981 ( .A1(n13252), .A2(n13077), .ZN(n8531) );
  NAND2_X1 U10982 ( .A1(n13422), .A2(n8531), .ZN(n13227) );
  NAND2_X1 U10983 ( .A1(n11684), .A2(n6474), .ZN(n8533) );
  INV_X1 U10984 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9559) );
  OR2_X1 U10985 ( .A1(n6681), .A2(n9559), .ZN(n8532) );
  AND2_X2 U10986 ( .A1(n8533), .A2(n8532), .ZN(n13502) );
  NAND2_X1 U10987 ( .A1(n8615), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8542) );
  INV_X1 U10988 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13231) );
  OR2_X1 U10989 ( .A1(n6655), .A2(n13231), .ZN(n8541) );
  NAND2_X1 U10990 ( .A1(n8534), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13219) );
  INV_X1 U10991 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10992 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  NAND2_X1 U10993 ( .A1(n13219), .A2(n8537), .ZN(n13240) );
  OR2_X1 U10994 ( .A1(n6666), .A2(n13240), .ZN(n8540) );
  INV_X1 U10995 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8538) );
  OR2_X1 U10996 ( .A1(n8842), .A2(n8538), .ZN(n8539) );
  NAND2_X1 U10997 ( .A1(n12018), .A2(n13101), .ZN(n8544) );
  OR2_X1 U10998 ( .A1(n12018), .A2(n13101), .ZN(n8543) );
  NAND2_X1 U10999 ( .A1(n8544), .A2(n8543), .ZN(n8920) );
  NAND2_X1 U11000 ( .A1(n13229), .A2(n8544), .ZN(n8550) );
  NAND2_X1 U11001 ( .A1(n8615), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8549) );
  INV_X1 U11002 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13220) );
  OR2_X1 U11003 ( .A1(n6655), .A2(n13220), .ZN(n8548) );
  OR2_X1 U11004 ( .A1(n6666), .A2(n13219), .ZN(n8547) );
  INV_X1 U11005 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8662) );
  OR2_X1 U11006 ( .A1(n8842), .A2(n8662), .ZN(n8546) );
  AND4_X1 U11007 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n12013)
         );
  INV_X1 U11008 ( .A(n11133), .ZN(n11151) );
  INV_X1 U11009 ( .A(n10852), .ZN(n14813) );
  INV_X1 U11010 ( .A(n14803), .ZN(n10669) );
  OR2_X1 U11011 ( .A1(n10246), .A2(n8554), .ZN(n10264) );
  NAND2_X1 U11012 ( .A1(n10303), .A2(n8204), .ZN(n10408) );
  OR2_X1 U11013 ( .A1(n10985), .A2(n14820), .ZN(n10986) );
  INV_X1 U11014 ( .A(n13482), .ZN(n13033) );
  INV_X1 U11015 ( .A(n13465), .ZN(n13362) );
  NAND2_X1 U11016 ( .A1(n13381), .A2(n13362), .ZN(n13357) );
  OR2_X1 U11017 ( .A1(n13357), .A2(n13348), .ZN(n13328) );
  INV_X1 U11018 ( .A(n11023), .ZN(n8553) );
  AOI211_X1 U11019 ( .C1(n8850), .C2(n13230), .A(n13295), .B(n13208), .ZN(
        n13223) );
  INV_X1 U11020 ( .A(n13131), .ZN(n8555) );
  INV_X1 U11021 ( .A(n10266), .ZN(n8556) );
  NAND2_X1 U11022 ( .A1(n10267), .A2(n8556), .ZN(n8559) );
  NAND2_X1 U11023 ( .A1(n8557), .A2(n10265), .ZN(n8558) );
  NAND2_X1 U11024 ( .A1(n8559), .A2(n8558), .ZN(n10307) );
  NAND2_X1 U11025 ( .A1(n8560), .A2(n10305), .ZN(n8561) );
  INV_X1 U11026 ( .A(n13126), .ZN(n8562) );
  NAND2_X1 U11027 ( .A1(n10413), .A2(n8562), .ZN(n8563) );
  XNOR2_X1 U11028 ( .A(n14796), .B(n13125), .ZN(n10517) );
  INV_X1 U11029 ( .A(n13125), .ZN(n8564) );
  NAND2_X1 U11030 ( .A1(n14796), .A2(n8564), .ZN(n8565) );
  NAND2_X1 U11031 ( .A1(n14803), .A2(n8566), .ZN(n8567) );
  INV_X1 U11032 ( .A(n13123), .ZN(n8568) );
  OR2_X1 U11033 ( .A1(n10852), .A2(n8568), .ZN(n8902) );
  NAND2_X1 U11034 ( .A1(n10852), .A2(n8568), .ZN(n8901) );
  INV_X1 U11035 ( .A(n8908), .ZN(n10980) );
  INV_X1 U11036 ( .A(n13120), .ZN(n8570) );
  NAND2_X1 U11037 ( .A1(n10885), .A2(n8570), .ZN(n8571) );
  INV_X1 U11038 ( .A(n13119), .ZN(n8572) );
  NAND2_X1 U11039 ( .A1(n11133), .A2(n8572), .ZN(n8573) );
  NAND2_X1 U11040 ( .A1(n8574), .A2(n8573), .ZN(n11240) );
  XNOR2_X1 U11041 ( .A(n11263), .B(n13118), .ZN(n11245) );
  INV_X1 U11042 ( .A(n13118), .ZN(n8575) );
  NAND2_X1 U11043 ( .A1(n11263), .A2(n8575), .ZN(n8576) );
  INV_X1 U11044 ( .A(n13117), .ZN(n8898) );
  AND2_X1 U11045 ( .A1(n14439), .A2(n8898), .ZN(n8577) );
  INV_X1 U11046 ( .A(n13116), .ZN(n8578) );
  NAND2_X1 U11047 ( .A1(n11431), .A2(n8578), .ZN(n8899) );
  OR2_X1 U11048 ( .A1(n11431), .A2(n8578), .ZN(n8900) );
  INV_X1 U11049 ( .A(n13115), .ZN(n8580) );
  NAND2_X1 U11050 ( .A1(n14412), .A2(n8580), .ZN(n8579) );
  OR2_X1 U11051 ( .A1(n14412), .A2(n8580), .ZN(n8581) );
  INV_X1 U11052 ( .A(n13114), .ZN(n8583) );
  NAND2_X1 U11053 ( .A1(n13096), .A2(n8583), .ZN(n8584) );
  OR2_X1 U11054 ( .A1(n13488), .A2(n11966), .ZN(n11663) );
  NAND2_X1 U11055 ( .A1(n11665), .A2(n11663), .ZN(n8586) );
  NAND2_X1 U11056 ( .A1(n8586), .A2(n8913), .ZN(n11667) );
  INV_X1 U11057 ( .A(n13112), .ZN(n8587) );
  OR2_X1 U11058 ( .A1(n13482), .A2(n8587), .ZN(n8588) );
  NAND2_X1 U11059 ( .A1(n13477), .A2(n8590), .ZN(n8589) );
  OR2_X1 U11060 ( .A1(n13477), .A2(n8590), .ZN(n8591) );
  NAND2_X1 U11061 ( .A1(n13383), .A2(n8592), .ZN(n8594) );
  OR2_X1 U11062 ( .A1(n13383), .A2(n8592), .ZN(n8593) );
  NAND2_X1 U11063 ( .A1(n8594), .A2(n8593), .ZN(n13377) );
  INV_X1 U11064 ( .A(n13109), .ZN(n8595) );
  NAND2_X1 U11065 ( .A1(n13465), .A2(n8595), .ZN(n8597) );
  OR2_X1 U11066 ( .A1(n13465), .A2(n8595), .ZN(n8596) );
  NAND2_X1 U11067 ( .A1(n8597), .A2(n8596), .ZN(n13355) );
  INV_X1 U11068 ( .A(n13355), .ZN(n13365) );
  NAND2_X1 U11069 ( .A1(n13364), .A2(n13365), .ZN(n13363) );
  NAND2_X1 U11070 ( .A1(n13363), .A2(n8597), .ZN(n13343) );
  INV_X1 U11071 ( .A(n13108), .ZN(n8598) );
  NAND2_X1 U11072 ( .A1(n13348), .A2(n8598), .ZN(n8599) );
  INV_X1 U11073 ( .A(n13107), .ZN(n12981) );
  INV_X1 U11074 ( .A(n13106), .ZN(n11988) );
  NAND2_X1 U11075 ( .A1(n13289), .A2(n8600), .ZN(n8602) );
  NAND2_X1 U11076 ( .A1(n13441), .A2(n12980), .ZN(n8601) );
  NAND2_X1 U11077 ( .A1(n8602), .A2(n8601), .ZN(n13274) );
  INV_X1 U11078 ( .A(n13279), .ZN(n8603) );
  INV_X1 U11079 ( .A(n13079), .ZN(n13104) );
  OR2_X1 U11080 ( .A1(n13511), .A2(n13104), .ZN(n8604) );
  INV_X1 U11081 ( .A(n13005), .ZN(n13103) );
  NOR2_X1 U11082 ( .A1(n13507), .A2(n13103), .ZN(n8605) );
  NAND2_X1 U11083 ( .A1(n13507), .A2(n13103), .ZN(n8606) );
  OR2_X1 U11084 ( .A1(n13252), .A2(n13102), .ZN(n8607) );
  XNOR2_X1 U11085 ( .A(n8609), .B(n8608), .ZN(n8611) );
  OR2_X1 U11086 ( .A1(n11075), .A2(n11023), .ZN(n8890) );
  NAND2_X1 U11087 ( .A1(n6641), .A2(n8935), .ZN(n8610) );
  NAND2_X1 U11088 ( .A1(n8611), .A2(n14399), .ZN(n8622) );
  OR2_X1 U11089 ( .A1(n9958), .A2(n9873), .ZN(n13078) );
  INV_X1 U11090 ( .A(P2_B_REG_SCAN_IN), .ZN(n8613) );
  INV_X1 U11091 ( .A(n9958), .ZN(n8654) );
  NAND2_X1 U11092 ( .A1(n8654), .A2(n9873), .ZN(n13076) );
  OAI21_X1 U11093 ( .B1(n13547), .B2(n8613), .A(n13065), .ZN(n13204) );
  INV_X1 U11094 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11095 ( .A1(n8614), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U11096 ( .A1(n8615), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8616) );
  OAI211_X1 U11097 ( .C1(n6655), .C2(n8618), .A(n8617), .B(n8616), .ZN(n13099)
         );
  INV_X1 U11098 ( .A(n13099), .ZN(n8619) );
  INV_X1 U11099 ( .A(n8620), .ZN(n8621) );
  NAND2_X1 U11100 ( .A1(n8622), .A2(n8621), .ZN(n13217) );
  NOR4_X1 U11101 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8626) );
  NOR4_X1 U11102 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8625) );
  NOR4_X1 U11103 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8624) );
  NOR4_X1 U11104 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8623) );
  NAND4_X1 U11105 ( .A1(n8626), .A2(n8625), .A3(n8624), .A4(n8623), .ZN(n8647)
         );
  NOR2_X1 U11106 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8630) );
  NOR4_X1 U11107 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8629) );
  NOR4_X1 U11108 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8628) );
  NOR4_X1 U11109 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8627) );
  NAND4_X1 U11110 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n8646)
         );
  INV_X1 U11111 ( .A(n8631), .ZN(n8633) );
  NAND2_X1 U11112 ( .A1(n8633), .A2(n8632), .ZN(n8635) );
  NAND2_X1 U11113 ( .A1(n8635), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8634) );
  MUX2_X1 U11114 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8634), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8636) );
  XNOR2_X1 U11115 ( .A(n13558), .B(P2_B_REG_SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11116 ( .A1(n8637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8638) );
  MUX2_X1 U11117 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8638), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8641) );
  NAND2_X1 U11118 ( .A1(n8641), .A2(n8640), .ZN(n13555) );
  NAND2_X1 U11119 ( .A1(n8642), .A2(n13555), .ZN(n8645) );
  NAND2_X1 U11120 ( .A1(n8640), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8643) );
  INV_X1 U11121 ( .A(n13553), .ZN(n8644) );
  OAI21_X1 U11122 ( .B1(n8647), .B2(n8646), .A(n14754), .ZN(n9946) );
  OAI21_X1 U11123 ( .B1(n8648), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8650) );
  XNOR2_X1 U11124 ( .A(n8650), .B(n8649), .ZN(n9867) );
  INV_X1 U11125 ( .A(n13555), .ZN(n8652) );
  NOR2_X1 U11126 ( .A1(n13558), .A2(n13553), .ZN(n8651) );
  NAND2_X1 U11127 ( .A1(n8652), .A2(n8651), .ZN(n9706) );
  NAND2_X1 U11128 ( .A1(n8653), .A2(n11023), .ZN(n8933) );
  NAND2_X1 U11129 ( .A1(n8654), .A2(n8933), .ZN(n9950) );
  NAND3_X1 U11130 ( .A1(n9946), .A2(n14791), .A3(n9950), .ZN(n8938) );
  INV_X1 U11131 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11132 ( .A1(n13558), .A2(n13553), .ZN(n14787) );
  INV_X1 U11133 ( .A(n14787), .ZN(n8655) );
  INV_X1 U11134 ( .A(n9947), .ZN(n8657) );
  NOR2_X1 U11135 ( .A1(n8938), .A2(n8657), .ZN(n8660) );
  INV_X1 U11136 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14789) );
  NAND2_X1 U11137 ( .A1(n14754), .A2(n14789), .ZN(n8659) );
  NAND2_X1 U11138 ( .A1(n13555), .A2(n13553), .ZN(n8658) );
  NAND2_X1 U11139 ( .A1(n8659), .A2(n8658), .ZN(n14790) );
  INV_X1 U11140 ( .A(n14790), .ZN(n10276) );
  INV_X1 U11141 ( .A(n8663), .ZN(n8664) );
  OAI21_X1 U11142 ( .B1(n8944), .B2(n8665), .A(n8664), .ZN(P2_U3528) );
  NAND2_X1 U11143 ( .A1(n10247), .A2(n8666), .ZN(n8667) );
  NAND2_X1 U11144 ( .A1(n8668), .A2(n8667), .ZN(n8673) );
  NOR2_X1 U11145 ( .A1(n11075), .A2(n8552), .ZN(n8669) );
  NAND2_X1 U11146 ( .A1(n8673), .A2(n8672), .ZN(n8676) );
  INV_X1 U11147 ( .A(n8676), .ZN(n8675) );
  OAI21_X1 U11148 ( .B1(n8884), .B2(n10024), .A(n8676), .ZN(n8677) );
  NAND2_X1 U11149 ( .A1(n8677), .A2(n10246), .ZN(n8680) );
  INV_X1 U11150 ( .A(n10247), .ZN(n10034) );
  AND2_X1 U11151 ( .A1(n8668), .A2(n10034), .ZN(n8903) );
  NAND3_X1 U11152 ( .A1(n8678), .A2(n8884), .A3(n8903), .ZN(n8679) );
  INV_X1 U11153 ( .A(n8681), .ZN(n8871) );
  NAND2_X1 U11154 ( .A1(n8683), .A2(n8682), .ZN(n8689) );
  NAND2_X1 U11155 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  MUX2_X1 U11156 ( .A(n13127), .B(n10305), .S(n8884), .Z(n8693) );
  NAND2_X1 U11157 ( .A1(n8692), .A2(n8693), .ZN(n8691) );
  MUX2_X1 U11158 ( .A(n13127), .B(n10305), .S(n8867), .Z(n8690) );
  NAND2_X1 U11159 ( .A1(n8691), .A2(n8690), .ZN(n8697) );
  INV_X1 U11160 ( .A(n8692), .ZN(n8695) );
  INV_X1 U11161 ( .A(n8693), .ZN(n8694) );
  NAND2_X1 U11162 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  MUX2_X1 U11163 ( .A(n13126), .B(n10413), .S(n8867), .Z(n8699) );
  MUX2_X1 U11164 ( .A(n13126), .B(n10413), .S(n8884), .Z(n8698) );
  MUX2_X1 U11165 ( .A(n13125), .B(n14796), .S(n6645), .Z(n8703) );
  NAND2_X1 U11166 ( .A1(n8702), .A2(n8703), .ZN(n8701) );
  MUX2_X1 U11167 ( .A(n13125), .B(n14796), .S(n8867), .Z(n8700) );
  NAND2_X1 U11168 ( .A1(n8701), .A2(n8700), .ZN(n8707) );
  INV_X1 U11169 ( .A(n8702), .ZN(n8705) );
  INV_X1 U11170 ( .A(n8703), .ZN(n8704) );
  NAND2_X1 U11171 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  MUX2_X1 U11172 ( .A(n13124), .B(n14803), .S(n8867), .Z(n8709) );
  INV_X1 U11173 ( .A(n8709), .ZN(n8710) );
  MUX2_X1 U11174 ( .A(n13123), .B(n10852), .S(n6645), .Z(n8714) );
  MUX2_X1 U11175 ( .A(n13123), .B(n10852), .S(n8867), .Z(n8711) );
  NAND2_X1 U11176 ( .A1(n8712), .A2(n8711), .ZN(n8718) );
  INV_X1 U11177 ( .A(n8713), .ZN(n8716) );
  INV_X1 U11178 ( .A(n8714), .ZN(n8715) );
  NAND2_X1 U11179 ( .A1(n8716), .A2(n8715), .ZN(n8717) );
  MUX2_X1 U11180 ( .A(n13122), .B(n14820), .S(n8867), .Z(n8720) );
  MUX2_X1 U11181 ( .A(n13122), .B(n14820), .S(n8849), .Z(n8719) );
  INV_X1 U11182 ( .A(n8720), .ZN(n8721) );
  MUX2_X1 U11183 ( .A(n13120), .B(n11112), .S(n6645), .Z(n8725) );
  MUX2_X1 U11184 ( .A(n13120), .B(n11112), .S(n6643), .Z(n8722) );
  NAND2_X1 U11185 ( .A1(n8723), .A2(n8722), .ZN(n8729) );
  INV_X1 U11186 ( .A(n8724), .ZN(n8727) );
  INV_X1 U11187 ( .A(n8725), .ZN(n8726) );
  NAND2_X1 U11188 ( .A1(n8727), .A2(n8726), .ZN(n8728) );
  NAND2_X1 U11189 ( .A1(n8729), .A2(n8728), .ZN(n8731) );
  MUX2_X1 U11190 ( .A(n13119), .B(n11133), .S(n6643), .Z(n8732) );
  MUX2_X1 U11191 ( .A(n13119), .B(n11133), .S(n8849), .Z(n8730) );
  INV_X1 U11192 ( .A(n8731), .ZN(n8734) );
  INV_X1 U11193 ( .A(n8732), .ZN(n8733) );
  NAND2_X1 U11194 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  MUX2_X1 U11195 ( .A(n13118), .B(n11263), .S(n6645), .Z(n8737) );
  MUX2_X1 U11196 ( .A(n13118), .B(n11263), .S(n6643), .Z(n8736) );
  MUX2_X1 U11197 ( .A(n13117), .B(n14439), .S(n6643), .Z(n8741) );
  NAND2_X1 U11198 ( .A1(n8740), .A2(n8741), .ZN(n8739) );
  MUX2_X1 U11199 ( .A(n13117), .B(n14439), .S(n6645), .Z(n8738) );
  NAND2_X1 U11200 ( .A1(n8739), .A2(n8738), .ZN(n8745) );
  INV_X1 U11201 ( .A(n8740), .ZN(n8743) );
  INV_X1 U11202 ( .A(n8741), .ZN(n8742) );
  NAND2_X1 U11203 ( .A1(n8743), .A2(n8742), .ZN(n8744) );
  MUX2_X1 U11204 ( .A(n13116), .B(n11431), .S(n6645), .Z(n8749) );
  NAND2_X1 U11205 ( .A1(n8748), .A2(n8749), .ZN(n8747) );
  MUX2_X1 U11206 ( .A(n13116), .B(n11431), .S(n6643), .Z(n8746) );
  NAND2_X1 U11207 ( .A1(n8747), .A2(n8746), .ZN(n8753) );
  INV_X1 U11208 ( .A(n8748), .ZN(n8751) );
  INV_X1 U11209 ( .A(n8749), .ZN(n8750) );
  NAND2_X1 U11210 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  MUX2_X1 U11211 ( .A(n13115), .B(n14412), .S(n6643), .Z(n8755) );
  MUX2_X1 U11212 ( .A(n13115), .B(n14412), .S(n6645), .Z(n8754) );
  INV_X1 U11213 ( .A(n8755), .ZN(n8756) );
  MUX2_X1 U11214 ( .A(n13114), .B(n13096), .S(n6645), .Z(n8760) );
  MUX2_X1 U11215 ( .A(n13114), .B(n13096), .S(n6643), .Z(n8757) );
  NAND2_X1 U11216 ( .A1(n8758), .A2(n8757), .ZN(n8764) );
  INV_X1 U11217 ( .A(n8759), .ZN(n8762) );
  INV_X1 U11218 ( .A(n8760), .ZN(n8761) );
  NAND2_X1 U11219 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  MUX2_X1 U11220 ( .A(n13113), .B(n13488), .S(n6643), .Z(n8767) );
  MUX2_X1 U11221 ( .A(n13113), .B(n13488), .S(n8849), .Z(n8765) );
  INV_X1 U11222 ( .A(n8766), .ZN(n8769) );
  INV_X1 U11223 ( .A(n8767), .ZN(n8768) );
  NAND2_X1 U11224 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  MUX2_X1 U11225 ( .A(n13112), .B(n13482), .S(n8849), .Z(n8772) );
  MUX2_X1 U11226 ( .A(n13112), .B(n13482), .S(n6643), .Z(n8771) );
  MUX2_X1 U11227 ( .A(n13111), .B(n13477), .S(n6643), .Z(n8776) );
  NAND2_X1 U11228 ( .A1(n8775), .A2(n8776), .ZN(n8774) );
  INV_X1 U11229 ( .A(n8867), .ZN(n8849) );
  MUX2_X1 U11230 ( .A(n13111), .B(n13477), .S(n8849), .Z(n8773) );
  NAND2_X1 U11231 ( .A1(n8774), .A2(n8773), .ZN(n8780) );
  INV_X1 U11232 ( .A(n8775), .ZN(n8778) );
  INV_X1 U11233 ( .A(n8776), .ZN(n8777) );
  NAND2_X1 U11234 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  MUX2_X1 U11235 ( .A(n13110), .B(n13383), .S(n8849), .Z(n8784) );
  NAND2_X1 U11236 ( .A1(n8783), .A2(n8784), .ZN(n8782) );
  MUX2_X1 U11237 ( .A(n13110), .B(n13383), .S(n6643), .Z(n8781) );
  INV_X1 U11238 ( .A(n8783), .ZN(n8786) );
  INV_X1 U11239 ( .A(n8784), .ZN(n8785) );
  MUX2_X1 U11240 ( .A(n13109), .B(n13465), .S(n6643), .Z(n8788) );
  MUX2_X1 U11241 ( .A(n13109), .B(n13465), .S(n8849), .Z(n8787) );
  INV_X1 U11242 ( .A(n8788), .ZN(n8789) );
  MUX2_X1 U11243 ( .A(n13108), .B(n13348), .S(n8849), .Z(n8793) );
  MUX2_X1 U11244 ( .A(n13108), .B(n13348), .S(n6643), .Z(n8790) );
  INV_X1 U11245 ( .A(n8792), .ZN(n8795) );
  INV_X1 U11246 ( .A(n8793), .ZN(n8794) );
  MUX2_X1 U11247 ( .A(n13107), .B(n13332), .S(n6643), .Z(n8797) );
  MUX2_X1 U11248 ( .A(n13107), .B(n13332), .S(n8849), .Z(n8796) );
  MUX2_X1 U11249 ( .A(n13106), .B(n13313), .S(n8849), .Z(n8801) );
  MUX2_X1 U11250 ( .A(n13106), .B(n13313), .S(n6643), .Z(n8798) );
  NAND2_X1 U11251 ( .A1(n8799), .A2(n8798), .ZN(n8805) );
  INV_X1 U11252 ( .A(n8800), .ZN(n8803) );
  INV_X1 U11253 ( .A(n8801), .ZN(n8802) );
  NAND2_X1 U11254 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  MUX2_X1 U11255 ( .A(n13105), .B(n13441), .S(n6643), .Z(n8809) );
  NAND2_X1 U11256 ( .A1(n8808), .A2(n8809), .ZN(n8807) );
  MUX2_X1 U11257 ( .A(n13105), .B(n13441), .S(n8849), .Z(n8806) );
  NAND2_X1 U11258 ( .A1(n8807), .A2(n8806), .ZN(n8813) );
  INV_X1 U11259 ( .A(n8808), .ZN(n8811) );
  NAND2_X1 U11260 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  NAND2_X1 U11261 ( .A1(n8813), .A2(n8812), .ZN(n8828) );
  MUX2_X1 U11262 ( .A(n13005), .B(n13507), .S(n8849), .Z(n8820) );
  INV_X1 U11263 ( .A(n13507), .ZN(n13082) );
  MUX2_X1 U11264 ( .A(n13103), .B(n13082), .S(n6643), .Z(n8819) );
  NAND2_X1 U11265 ( .A1(n8820), .A2(n8819), .ZN(n8824) );
  MUX2_X1 U11266 ( .A(n13104), .B(n13010), .S(n8849), .Z(n8817) );
  INV_X1 U11267 ( .A(n8817), .ZN(n8815) );
  MUX2_X1 U11268 ( .A(n13079), .B(n13511), .S(n6643), .Z(n8818) );
  INV_X1 U11269 ( .A(n8818), .ZN(n8814) );
  NAND2_X1 U11270 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  AND2_X1 U11271 ( .A1(n8824), .A2(n8816), .ZN(n8827) );
  MUX2_X1 U11272 ( .A(n13077), .B(n13252), .S(n8849), .Z(n8856) );
  MUX2_X1 U11273 ( .A(n13102), .B(n13424), .S(n6643), .Z(n8855) );
  MUX2_X1 U11274 ( .A(n12971), .B(n13502), .S(n6643), .Z(n8852) );
  MUX2_X1 U11275 ( .A(n13101), .B(n12018), .S(n8849), .Z(n8851) );
  NAND2_X1 U11276 ( .A1(n8852), .A2(n8851), .ZN(n8857) );
  AND2_X1 U11277 ( .A1(n8818), .A2(n8817), .ZN(n8823) );
  INV_X1 U11278 ( .A(n8819), .ZN(n8822) );
  INV_X1 U11279 ( .A(n8820), .ZN(n8821) );
  AOI22_X1 U11280 ( .A1(n8824), .A2(n8823), .B1(n8822), .B2(n8821), .ZN(n8825)
         );
  INV_X1 U11281 ( .A(SI_29_), .ZN(n15211) );
  NAND2_X1 U11282 ( .A1(n8831), .A2(n15211), .ZN(n8832) );
  MUX2_X1 U11283 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9735), .Z(n8834) );
  XNOR2_X1 U11284 ( .A(n8834), .B(SI_30_), .ZN(n8861) );
  INV_X1 U11285 ( .A(n8834), .ZN(n8835) );
  INV_X1 U11286 ( .A(SI_30_), .ZN(n15215) );
  MUX2_X1 U11287 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9735), .Z(n8836) );
  XNOR2_X1 U11288 ( .A(n8836), .B(SI_31_), .ZN(n8837) );
  NAND2_X1 U11289 ( .A1(n13536), .A2(n6474), .ZN(n8841) );
  INV_X1 U11290 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8839) );
  OR2_X1 U11291 ( .A1(n6681), .A2(n8839), .ZN(n8840) );
  INV_X1 U11292 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13413) );
  OR2_X1 U11293 ( .A1(n8842), .A2(n13413), .ZN(n8848) );
  INV_X1 U11294 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8843) );
  OR2_X1 U11295 ( .A1(n6655), .A2(n8843), .ZN(n8847) );
  INV_X1 U11296 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13494) );
  OR2_X1 U11297 ( .A1(n8845), .A2(n13494), .ZN(n8846) );
  XNOR2_X1 U11298 ( .A(n8883), .B(n13203), .ZN(n8926) );
  MUX2_X1 U11299 ( .A(n12013), .B(n13218), .S(n6643), .Z(n8873) );
  MUX2_X1 U11300 ( .A(n13100), .B(n8850), .S(n8849), .Z(n8872) );
  INV_X1 U11301 ( .A(n8851), .ZN(n8854) );
  INV_X1 U11302 ( .A(n8852), .ZN(n8853) );
  NAND2_X1 U11303 ( .A1(n8854), .A2(n8853), .ZN(n8859) );
  NAND3_X1 U11304 ( .A1(n8857), .A2(n8856), .A3(n8855), .ZN(n8858) );
  OAI211_X1 U11305 ( .C1(n8873), .C2(n8872), .A(n8859), .B(n8858), .ZN(n8860)
         );
  INV_X1 U11306 ( .A(n8861), .ZN(n8862) );
  NAND2_X1 U11307 ( .A1(n11953), .A2(n6479), .ZN(n8866) );
  INV_X1 U11308 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12189) );
  OR2_X1 U11309 ( .A1(n6681), .A2(n12189), .ZN(n8865) );
  MUX2_X1 U11310 ( .A(n13099), .B(n13212), .S(n6643), .Z(n8882) );
  INV_X1 U11311 ( .A(n13203), .ZN(n13098) );
  NAND2_X1 U11312 ( .A1(n13098), .A2(n6643), .ZN(n8868) );
  INV_X1 U11313 ( .A(n8670), .ZN(n10280) );
  OR2_X1 U11314 ( .A1(n10280), .A2(n8148), .ZN(n8889) );
  NAND4_X1 U11315 ( .A1(n8868), .A2(n10282), .A3(n8889), .A4(n8933), .ZN(n8869) );
  AND2_X1 U11316 ( .A1(n8869), .A2(n13099), .ZN(n8870) );
  AOI21_X1 U11317 ( .B1(n13212), .B2(n6670), .A(n8870), .ZN(n8881) );
  INV_X1 U11318 ( .A(n8872), .ZN(n8875) );
  INV_X1 U11319 ( .A(n8873), .ZN(n8874) );
  OAI22_X1 U11320 ( .A1(n8882), .A2(n8881), .B1(n8875), .B2(n8874), .ZN(n8877)
         );
  INV_X1 U11321 ( .A(n8926), .ZN(n8876) );
  NAND2_X1 U11322 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  NAND2_X1 U11323 ( .A1(n8882), .A2(n8881), .ZN(n8887) );
  MUX2_X1 U11324 ( .A(n13098), .B(n8883), .S(n6645), .Z(n8885) );
  NOR2_X1 U11325 ( .A1(n6533), .A2(n8885), .ZN(n8886) );
  OAI21_X1 U11326 ( .B1(n8890), .B2(n8653), .A(n8889), .ZN(n8891) );
  INV_X1 U11327 ( .A(n8891), .ZN(n8895) );
  NAND2_X1 U11328 ( .A1(n10282), .A2(n8653), .ZN(n8892) );
  OAI211_X1 U11329 ( .C1(n10022), .C2(n8935), .A(n8933), .B(n8892), .ZN(n8893)
         );
  NAND2_X1 U11330 ( .A1(n8929), .A2(n8893), .ZN(n8894) );
  OAI21_X1 U11331 ( .B1(n8929), .B2(n8895), .A(n8894), .ZN(n8932) );
  XNOR2_X1 U11332 ( .A(n13500), .B(n13099), .ZN(n8925) );
  XNOR2_X1 U11333 ( .A(n13082), .B(n13005), .ZN(n13263) );
  NAND2_X1 U11334 ( .A1(n8897), .A2(n8896), .ZN(n13316) );
  XNOR2_X1 U11335 ( .A(n14439), .B(n8898), .ZN(n11214) );
  NAND2_X1 U11336 ( .A1(n8900), .A2(n8899), .ZN(n11381) );
  NAND2_X1 U11337 ( .A1(n8902), .A2(n8901), .ZN(n10854) );
  INV_X1 U11338 ( .A(n8903), .ZN(n9955) );
  NAND2_X1 U11339 ( .A1(n9955), .A2(n10249), .ZN(n10285) );
  NOR4_X1 U11340 ( .A1(n10248), .A2(n10285), .A3(n10266), .A4(n11023), .ZN(
        n8906) );
  NAND4_X1 U11341 ( .A1(n8906), .A2(n10517), .A3(n8905), .A4(n8904), .ZN(n8907) );
  NOR4_X1 U11342 ( .A1(n8908), .A2(n10854), .A3(n8907), .A4(n10672), .ZN(n8909) );
  NAND4_X1 U11343 ( .A1(n11245), .A2(n8909), .A3(n11006), .A4(n10882), .ZN(
        n8910) );
  NOR4_X1 U11344 ( .A1(n8911), .A2(n11214), .A3(n11381), .A4(n8910), .ZN(n8914) );
  NAND2_X1 U11345 ( .A1(n8912), .A2(n14404), .ZN(n14406) );
  NAND4_X1 U11346 ( .A1(n8914), .A2(n11613), .A3(n8913), .A4(n14406), .ZN(
        n8915) );
  NOR4_X1 U11347 ( .A1(n13355), .A2(n13377), .A3(n8916), .A4(n8915), .ZN(n8918) );
  NAND4_X1 U11348 ( .A1(n13316), .A2(n8918), .A3(n8917), .A4(n13342), .ZN(
        n8919) );
  NOR4_X1 U11349 ( .A1(n13263), .A2(n13279), .A3(n13294), .A4(n8919), .ZN(
        n8922) );
  NAND4_X1 U11350 ( .A1(n8923), .A2(n8922), .A3(n8921), .A4(n8920), .ZN(n8924)
         );
  NOR3_X1 U11351 ( .A1(n8926), .A2(n8925), .A3(n8924), .ZN(n8927) );
  XNOR2_X1 U11352 ( .A(n6641), .B(n8927), .ZN(n8928) );
  OR2_X1 U11353 ( .A1(n9867), .A2(P2_U3088), .ZN(n11391) );
  INV_X1 U11354 ( .A(n11391), .ZN(n8930) );
  OAI21_X1 U11355 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n8937) );
  INV_X1 U11356 ( .A(n13547), .ZN(n9885) );
  INV_X1 U11357 ( .A(n8933), .ZN(n9948) );
  NAND4_X1 U11358 ( .A1(n14791), .A2(n9885), .A3(n9948), .A4(n13064), .ZN(
        n8934) );
  OAI211_X1 U11359 ( .C1(n8935), .C2(n11391), .A(n8934), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8936) );
  NAND2_X1 U11360 ( .A1(n8937), .A2(n8936), .ZN(P2_U3328) );
  NOR2_X1 U11361 ( .A1(n8938), .A2(n9947), .ZN(n10277) );
  NAND2_X1 U11362 ( .A1(n8850), .A2(n8940), .ZN(n8942) );
  NAND2_X1 U11363 ( .A1(n7143), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8941) );
  OAI21_X1 U11364 ( .B1(n8944), .B2(n7143), .A(n8943), .ZN(P2_U3496) );
  NAND2_X1 U11365 ( .A1(n6636), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9110) );
  INV_X1 U11366 ( .A(n9110), .ZN(n8945) );
  NAND2_X1 U11367 ( .A1(n9711), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U11368 ( .A1(n9721), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11369 ( .A1(n9741), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U11370 ( .A1(n8949), .A2(n8947), .ZN(n9119) );
  INV_X1 U11371 ( .A(n9119), .ZN(n8948) );
  NAND2_X1 U11372 ( .A1(n9120), .A2(n8948), .ZN(n8950) );
  NAND2_X1 U11373 ( .A1(n9725), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8952) );
  INV_X1 U11374 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U11375 ( .A1(n9761), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U11376 ( .A1(n9131), .A2(n9130), .ZN(n8953) );
  NAND2_X1 U11377 ( .A1(n8953), .A2(n8952), .ZN(n9143) );
  NAND2_X1 U11378 ( .A1(n9723), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8956) );
  INV_X1 U11379 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U11380 ( .A1(n9736), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11381 ( .A1(n8956), .A2(n8954), .ZN(n9142) );
  INV_X1 U11382 ( .A(n9142), .ZN(n8955) );
  NAND2_X1 U11383 ( .A1(n9143), .A2(n8955), .ZN(n8957) );
  NAND2_X1 U11384 ( .A1(n9727), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U11385 ( .A1(n9739), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11386 ( .A1(n8960), .A2(n8958), .ZN(n9158) );
  INV_X1 U11387 ( .A(n9158), .ZN(n8959) );
  NAND2_X1 U11388 ( .A1(n9159), .A2(n8959), .ZN(n8961) );
  NAND2_X1 U11389 ( .A1(n9750), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11390 ( .A1(n9752), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11391 ( .A1(n9765), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11392 ( .A1(n9768), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U11393 ( .A1(n8966), .A2(n8965), .ZN(n9191) );
  NAND2_X1 U11394 ( .A1(n9776), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U11395 ( .A1(n9778), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U11396 ( .A1(n9858), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11397 ( .A1(n9860), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U11398 ( .A1(n9222), .A2(n9221), .ZN(n8971) );
  NAND2_X1 U11399 ( .A1(n8971), .A2(n8970), .ZN(n9241) );
  NAND2_X1 U11400 ( .A1(n9912), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U11401 ( .A1(n9911), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U11402 ( .A1(n9965), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8974) );
  XNOR2_X1 U11403 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9274) );
  NAND2_X1 U11404 ( .A1(n9275), .A2(n9274), .ZN(n8977) );
  NAND2_X1 U11405 ( .A1(n8975), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U11406 ( .A1(n9282), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U11407 ( .A1(n8978), .A2(n10213), .ZN(n8979) );
  NAND2_X1 U11408 ( .A1(n10389), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11409 ( .A1(n10470), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U11410 ( .A1(n10471), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11411 ( .A1(n8984), .A2(n8983), .ZN(n9307) );
  NAND2_X1 U11412 ( .A1(n10384), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11413 ( .A1(n10385), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11414 ( .A1(n10421), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11415 ( .A1(n10423), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8987) );
  NAND2_X1 U11416 ( .A1(n10844), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8991) );
  INV_X1 U11417 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U11418 ( .A1(n10847), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11419 ( .A1(n8991), .A2(n8989), .ZN(n9360) );
  INV_X1 U11420 ( .A(n9360), .ZN(n8990) );
  INV_X1 U11421 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U11422 ( .A1(n10954), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8993) );
  INV_X1 U11423 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U11424 ( .A1(n10953), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U11425 ( .A1(n11077), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U11426 ( .A1(n11076), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U11427 ( .A1(n8998), .A2(n8996), .ZN(n9401) );
  INV_X1 U11428 ( .A(n9401), .ZN(n8997) );
  XNOR2_X1 U11429 ( .A(n11174), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11430 ( .A1(n11174), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9000) );
  XNOR2_X1 U11431 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9423) );
  NAND2_X1 U11432 ( .A1(n9001), .A2(n13560), .ZN(n9002) );
  NAND2_X1 U11433 ( .A1(n13556), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11434 ( .A1(n14161), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9005) );
  AND2_X1 U11435 ( .A1(n14158), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11436 ( .A1(n13551), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9008) );
  AND2_X1 U11437 ( .A1(n13548), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9009) );
  INV_X1 U11438 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14155) );
  XNOR2_X1 U11439 ( .A(n9559), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9010) );
  XNOR2_X1 U11440 ( .A(n9562), .B(n9010), .ZN(n11954) );
  AND2_X2 U11441 ( .A1(n9144), .A2(n9161), .ZN(n9177) );
  OAI21_X1 U11442 ( .B1(n9022), .B2(n12958), .A(P3_IR_REG_28__SCAN_IN), .ZN(
        n9024) );
  NAND2_X1 U11443 ( .A1(n11954), .A2(n12338), .ZN(n9027) );
  NAND2_X1 U11444 ( .A1(n12340), .A2(SI_28_), .ZN(n9026) );
  NAND2_X1 U11445 ( .A1(n9028), .A2(n9029), .ZN(n9311) );
  INV_X1 U11446 ( .A(n9311), .ZN(n9030) );
  NAND2_X1 U11447 ( .A1(n9030), .A2(n9312), .ZN(n9329) );
  INV_X1 U11448 ( .A(n9038), .ZN(n9035) );
  NAND2_X1 U11449 ( .A1(n9035), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9036) );
  MUX2_X1 U11450 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9036), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9039) );
  NAND2_X1 U11451 ( .A1(n6519), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U11452 ( .A1(n9041), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9042) );
  MUX2_X1 U11453 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9042), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9043) );
  AND2_X1 U11454 ( .A1(n12524), .A2(n12504), .ZN(n10606) );
  AND3_X1 U11455 ( .A1(n12529), .A2(n9582), .A3(n10709), .ZN(n9045) );
  AND2_X1 U11456 ( .A1(n9044), .A2(n9045), .ZN(n9689) );
  INV_X1 U11457 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11458 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  XNOR2_X1 U11459 ( .A(n11291), .B(P3_B_REG_SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11460 ( .A1(n9051), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9052) );
  MUX2_X1 U11461 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9052), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9054) );
  NAND2_X1 U11462 ( .A1(n9054), .A2(n9053), .ZN(n11682) );
  NAND2_X1 U11463 ( .A1(n9055), .A2(n11682), .ZN(n9057) );
  NAND2_X1 U11464 ( .A1(n9053), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9056) );
  INV_X1 U11465 ( .A(n9084), .ZN(n11362) );
  NAND2_X1 U11466 ( .A1(n11362), .A2(n11682), .ZN(n9058) );
  NAND2_X1 U11467 ( .A1(n11362), .A2(n11291), .ZN(n9061) );
  NOR2_X1 U11468 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9065) );
  NOR4_X1 U11469 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9064) );
  NOR4_X1 U11470 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9063) );
  NOR4_X1 U11471 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9062) );
  NAND4_X1 U11472 ( .A1(n9065), .A2(n9064), .A3(n9063), .A4(n9062), .ZN(n9071)
         );
  NOR4_X1 U11473 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9069) );
  NOR4_X1 U11474 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9068) );
  NOR4_X1 U11475 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9067) );
  NOR4_X1 U11476 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9066) );
  NAND4_X1 U11477 ( .A1(n9069), .A2(n9068), .A3(n9067), .A4(n9066), .ZN(n9070)
         );
  NOR2_X1 U11478 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  OR2_X1 U11479 ( .A1(n9060), .A2(n9072), .ZN(n9540) );
  NAND3_X1 U11480 ( .A1(n12954), .A2(n12956), .A3(n9540), .ZN(n9688) );
  INV_X1 U11481 ( .A(n9688), .ZN(n9684) );
  OAI21_X1 U11482 ( .B1(n10606), .B2(n9689), .A(n9684), .ZN(n9079) );
  INV_X1 U11483 ( .A(n12954), .ZN(n10803) );
  NAND3_X1 U11484 ( .A1(n9585), .A2(n10803), .A3(n9540), .ZN(n9694) );
  INV_X1 U11485 ( .A(n9694), .ZN(n9698) );
  NAND2_X1 U11486 ( .A1(n12529), .A2(n10515), .ZN(n9073) );
  NAND2_X1 U11487 ( .A1(n9044), .A2(n9073), .ZN(n9074) );
  NAND2_X1 U11488 ( .A1(n9074), .A2(n10709), .ZN(n9077) );
  NAND2_X1 U11489 ( .A1(n10709), .A2(n10515), .ZN(n9075) );
  NAND2_X1 U11490 ( .A1(n9543), .A2(n9075), .ZN(n9076) );
  NAND2_X1 U11491 ( .A1(n9077), .A2(n9076), .ZN(n9687) );
  NAND2_X1 U11492 ( .A1(n9698), .A2(n9687), .ZN(n9078) );
  NAND2_X1 U11493 ( .A1(n9079), .A2(n9078), .ZN(n9085) );
  INV_X1 U11494 ( .A(n11291), .ZN(n9083) );
  INV_X1 U11495 ( .A(n11682), .ZN(n9082) );
  NAND3_X1 U11496 ( .A1(n9084), .A2(n9083), .A3(n9082), .ZN(n9709) );
  NAND2_X1 U11497 ( .A1(n9543), .A2(n10709), .ZN(n15068) );
  INV_X1 U11498 ( .A(n15068), .ZN(n14383) );
  NOR2_X1 U11499 ( .A1(n15076), .A2(n9087), .ZN(n9088) );
  NAND3_X1 U11500 ( .A1(n9687), .A2(n12524), .A3(n15068), .ZN(n9090) );
  NAND2_X1 U11501 ( .A1(n12529), .A2(n9582), .ZN(n9089) );
  OR2_X1 U11502 ( .A1(n9044), .A2(n9089), .ZN(n9548) );
  NAND2_X1 U11503 ( .A1(n9090), .A2(n9548), .ZN(n12683) );
  INV_X1 U11504 ( .A(n9094), .ZN(n12192) );
  INV_X1 U11505 ( .A(n9093), .ZN(n12959) );
  AND2_X2 U11506 ( .A1(n12192), .A2(n9095), .ZN(n9201) );
  NAND2_X1 U11507 ( .A1(n9201), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9099) );
  AND2_X2 U11508 ( .A1(n12192), .A2(n12965), .ZN(n9153) );
  NAND2_X1 U11509 ( .A1(n9153), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11510 ( .A1(n6486), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11511 ( .A1(n6483), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9096) );
  OR2_X1 U11512 ( .A1(n9165), .A2(n9758), .ZN(n9105) );
  INV_X1 U11513 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11514 ( .A1(n9100), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U11515 ( .A1(n9110), .A2(n9101), .ZN(n9757) );
  NAND2_X1 U11516 ( .A1(n9160), .A2(n9757), .ZN(n9104) );
  NAND2_X1 U11517 ( .A1(n9279), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11518 ( .A1(n9169), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11519 ( .A1(n6481), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11520 ( .A1(n9201), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9106) );
  XNOR2_X1 U11521 ( .A(n9111), .B(n9110), .ZN(n9713) );
  INV_X1 U11522 ( .A(n10060), .ZN(n9112) );
  OAI22_X1 U11523 ( .A1(n9381), .A2(n9713), .B1(n9102), .B2(n10182), .ZN(n9114) );
  NOR2_X1 U11524 ( .A1(n9165), .A2(n9712), .ZN(n9113) );
  NOR2_X2 U11525 ( .A1(n9114), .A2(n9113), .ZN(n15031) );
  NAND2_X1 U11526 ( .A1(n9201), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U11527 ( .A1(n6483), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11528 ( .A1(n6486), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U11529 ( .A1(n9153), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9115) );
  XNOR2_X1 U11530 ( .A(n9120), .B(n9119), .ZN(n9771) );
  INV_X1 U11531 ( .A(n9771), .ZN(n9121) );
  OR2_X1 U11532 ( .A1(n9381), .A2(n9121), .ZN(n9125) );
  XNOR2_X2 U11533 ( .A(n9123), .B(n9122), .ZN(n10444) );
  NAND2_X1 U11534 ( .A1(n9279), .A2(n10444), .ZN(n9124) );
  OAI211_X1 U11535 ( .C1(SI_2_), .C2(n9165), .A(n9125), .B(n9124), .ZN(n10905)
         );
  NAND2_X1 U11536 ( .A1(n10656), .A2(n10657), .ZN(n10658) );
  INV_X1 U11537 ( .A(n10905), .ZN(n12405) );
  NAND2_X1 U11538 ( .A1(n15039), .A2(n12405), .ZN(n12406) );
  NAND2_X1 U11539 ( .A1(n10658), .A2(n12406), .ZN(n11097) );
  BUF_X2 U11540 ( .A(n9201), .Z(n9483) );
  NAND2_X1 U11541 ( .A1(n9483), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U11542 ( .A1(n6482), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U11543 ( .A1(n6486), .A2(n14885), .ZN(n9127) );
  NAND2_X1 U11544 ( .A1(n9153), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9126) );
  INV_X1 U11545 ( .A(n12552), .ZN(n9602) );
  XNOR2_X1 U11546 ( .A(n9131), .B(n9130), .ZN(n9733) );
  NAND2_X1 U11547 ( .A1(n9132), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9133) );
  XNOR2_X1 U11548 ( .A(n9133), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10456) );
  OAI22_X1 U11549 ( .A1(n9381), .A2(n9733), .B1(n10456), .B2(n9102), .ZN(n9135) );
  NOR2_X1 U11550 ( .A1(n9165), .A2(SI_3_), .ZN(n9134) );
  NAND2_X1 U11551 ( .A1(n9602), .A2(n9587), .ZN(n12407) );
  INV_X1 U11552 ( .A(n9587), .ZN(n15052) );
  NAND2_X1 U11553 ( .A1(n15052), .A2(n12552), .ZN(n12410) );
  NAND2_X1 U11554 ( .A1(n11097), .A2(n12357), .ZN(n9136) );
  NAND2_X1 U11555 ( .A1(n9136), .A2(n12407), .ZN(n10774) );
  NAND2_X1 U11556 ( .A1(n9201), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U11557 ( .A1(n6483), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9140) );
  AND2_X1 U11558 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9137) );
  NOR2_X1 U11559 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9151) );
  OR2_X1 U11560 ( .A1(n9137), .A2(n9151), .ZN(n10837) );
  NAND2_X1 U11561 ( .A1(n6486), .A2(n10837), .ZN(n9139) );
  XNOR2_X1 U11562 ( .A(n9143), .B(n9142), .ZN(n9772) );
  NAND2_X1 U11563 ( .A1(n9160), .A2(n9772), .ZN(n9150) );
  INV_X1 U11564 ( .A(n9144), .ZN(n9148) );
  NAND2_X1 U11565 ( .A1(n9145), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9146) );
  MUX2_X1 U11566 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9146), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9147) );
  NAND2_X1 U11567 ( .A1(n9148), .A2(n9147), .ZN(n14902) );
  NAND2_X1 U11568 ( .A1(n9279), .A2(n14902), .ZN(n9149) );
  OAI211_X1 U11569 ( .C1(SI_4_), .C2(n9165), .A(n9150), .B(n9149), .ZN(n10821)
         );
  NAND2_X1 U11570 ( .A1(n11093), .A2(n10833), .ZN(n12416) );
  NAND2_X1 U11571 ( .A1(n12551), .A2(n10821), .ZN(n12422) );
  INV_X1 U11572 ( .A(n12414), .ZN(n12359) );
  NAND2_X1 U11573 ( .A1(n10774), .A2(n12359), .ZN(n10775) );
  NAND2_X1 U11574 ( .A1(n10775), .A2(n12416), .ZN(n10864) );
  NAND2_X1 U11575 ( .A1(n6483), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U11576 ( .A1(n9201), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9156) );
  NOR2_X1 U11577 ( .A1(n9151), .A2(n15191), .ZN(n9152) );
  OR2_X1 U11578 ( .A1(n9167), .A2(n9152), .ZN(n11153) );
  NAND2_X1 U11579 ( .A1(n6486), .A2(n11153), .ZN(n9155) );
  NAND2_X1 U11580 ( .A1(n9153), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9154) );
  NAND4_X2 U11581 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(n12550) );
  XNOR2_X1 U11582 ( .A(n9159), .B(n9158), .ZN(n9769) );
  NAND2_X1 U11583 ( .A1(n9160), .A2(n9769), .ZN(n9164) );
  OR2_X1 U11584 ( .A1(n9144), .A2(n12958), .ZN(n9162) );
  XNOR2_X1 U11585 ( .A(n9162), .B(n9161), .ZN(n14924) );
  NAND2_X1 U11586 ( .A1(n9279), .A2(n14924), .ZN(n9163) );
  NAND2_X1 U11587 ( .A1(n10864), .A2(n12423), .ZN(n10863) );
  INV_X1 U11588 ( .A(n12550), .ZN(n12419) );
  INV_X1 U11589 ( .A(n10971), .ZN(n12418) );
  NAND2_X1 U11590 ( .A1(n12419), .A2(n12418), .ZN(n12424) );
  NAND2_X1 U11591 ( .A1(n10863), .A2(n12424), .ZN(n10935) );
  NAND2_X1 U11592 ( .A1(n6482), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U11593 ( .A1(n9483), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9172) );
  INV_X1 U11594 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n9166) );
  NOR2_X1 U11595 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  OR2_X1 U11596 ( .A1(n9181), .A2(n9168), .ZN(n11031) );
  NAND2_X1 U11597 ( .A1(n6486), .A2(n11031), .ZN(n9171) );
  NAND2_X1 U11598 ( .A1(n9153), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9170) );
  INV_X1 U11599 ( .A(n12549), .ZN(n10872) );
  XNOR2_X1 U11600 ( .A(n9752), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9174) );
  XNOR2_X1 U11601 ( .A(n9175), .B(n9174), .ZN(n9763) );
  INV_X1 U11602 ( .A(SI_6_), .ZN(n9176) );
  OR2_X1 U11603 ( .A1(n9177), .A2(n12958), .ZN(n9178) );
  NAND2_X1 U11604 ( .A1(n9279), .A2(n10624), .ZN(n9179) );
  INV_X1 U11605 ( .A(n10947), .ZN(n15057) );
  NAND2_X1 U11606 ( .A1(n12549), .A2(n15057), .ZN(n12428) );
  NAND2_X1 U11607 ( .A1(n10935), .A2(n12356), .ZN(n9180) );
  NAND2_X1 U11608 ( .A1(n9180), .A2(n12425), .ZN(n10995) );
  NAND2_X1 U11609 ( .A1(n9483), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U11610 ( .A1(n9181), .A2(n15192), .ZN(n9204) );
  INV_X1 U11611 ( .A(n9181), .ZN(n9182) );
  NAND2_X1 U11612 ( .A1(n9182), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9183) );
  AND2_X1 U11613 ( .A1(n9204), .A2(n9183), .ZN(n14855) );
  INV_X1 U11614 ( .A(n14855), .ZN(n9184) );
  NAND2_X1 U11615 ( .A1(n6486), .A2(n9184), .ZN(n9189) );
  INV_X1 U11616 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9185) );
  OR2_X1 U11617 ( .A1(n9488), .A2(n9185), .ZN(n9188) );
  INV_X1 U11618 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n9186) );
  OR2_X1 U11619 ( .A1(n9489), .A2(n9186), .ZN(n9187) );
  INV_X1 U11620 ( .A(SI_7_), .ZN(n9717) );
  NAND2_X1 U11621 ( .A1(n12340), .A2(n9717), .ZN(n9200) );
  NAND2_X1 U11622 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  NAND2_X1 U11623 ( .A1(n9194), .A2(n9193), .ZN(n9716) );
  NAND2_X1 U11624 ( .A1(n12338), .A2(n9716), .ZN(n9199) );
  INV_X1 U11625 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11626 ( .A1(n9177), .A2(n9195), .ZN(n9214) );
  NAND2_X1 U11627 ( .A1(n9214), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9197) );
  XNOR2_X1 U11628 ( .A(n9197), .B(n9196), .ZN(n10754) );
  NAND2_X1 U11629 ( .A1(n9279), .A2(n10754), .ZN(n9198) );
  NAND2_X1 U11630 ( .A1(n11232), .A2(n14848), .ZN(n12432) );
  NAND2_X1 U11631 ( .A1(n12548), .A2(n11304), .ZN(n12433) );
  NAND2_X1 U11632 ( .A1(n12432), .A2(n12433), .ZN(n12436) );
  INV_X1 U11633 ( .A(n12436), .ZN(n12358) );
  NAND2_X1 U11634 ( .A1(n9529), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U11635 ( .A1(n9153), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9208) );
  INV_X1 U11636 ( .A(n9204), .ZN(n9203) );
  INV_X1 U11637 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9202) );
  INV_X1 U11638 ( .A(n9234), .ZN(n9232) );
  NAND2_X1 U11639 ( .A1(n9204), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11640 ( .A1(n9232), .A2(n9205), .ZN(n11228) );
  NAND2_X1 U11641 ( .A1(n6486), .A2(n11228), .ZN(n9207) );
  NAND2_X1 U11642 ( .A1(n6483), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9206) );
  NAND4_X1 U11643 ( .A1(n9209), .A2(n9208), .A3(n9207), .A4(n9206), .ZN(n12547) );
  INV_X1 U11644 ( .A(n12547), .ZN(n11278) );
  OR2_X1 U11645 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  NAND2_X1 U11646 ( .A1(n9213), .A2(n9212), .ZN(n9715) );
  NAND2_X1 U11647 ( .A1(n12340), .A2(SI_8_), .ZN(n9220) );
  NAND2_X1 U11648 ( .A1(n9217), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9216) );
  MUX2_X1 U11649 ( .A(n9216), .B(P3_IR_REG_31__SCAN_IN), .S(n9215), .Z(n9218)
         );
  NAND2_X1 U11650 ( .A1(n9218), .A2(n9244), .ZN(n11203) );
  INV_X1 U11651 ( .A(n11203), .ZN(n11186) );
  NAND2_X1 U11652 ( .A1(n9279), .A2(n11186), .ZN(n9219) );
  OAI211_X1 U11653 ( .C1(n9381), .C2(n9715), .A(n9220), .B(n9219), .ZN(n11236)
         );
  NAND2_X1 U11654 ( .A1(n11278), .A2(n11236), .ZN(n12438) );
  INV_X1 U11655 ( .A(n11236), .ZN(n15062) );
  NAND2_X1 U11656 ( .A1(n12547), .A2(n15062), .ZN(n12439) );
  XNOR2_X1 U11657 ( .A(n9222), .B(n9221), .ZN(n9719) );
  NAND2_X1 U11658 ( .A1(n12338), .A2(n9719), .ZN(n9225) );
  NAND2_X1 U11659 ( .A1(n9244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9223) );
  XNOR2_X1 U11660 ( .A(n9223), .B(n9245), .ZN(n11195) );
  NAND2_X1 U11661 ( .A1(n9279), .A2(n11195), .ZN(n9224) );
  OAI211_X1 U11662 ( .C1(SI_9_), .C2(n9382), .A(n9225), .B(n9224), .ZN(n15069)
         );
  INV_X1 U11663 ( .A(n15069), .ZN(n12443) );
  NAND2_X1 U11664 ( .A1(n9529), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11665 ( .A1(n12341), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9228) );
  XNOR2_X1 U11666 ( .A(n9232), .B(P3_REG3_REG_9__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U11667 ( .A1(n6486), .A2(n11370), .ZN(n9227) );
  NAND2_X1 U11668 ( .A1(n6483), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9226) );
  NAND4_X1 U11669 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(n12546) );
  INV_X1 U11670 ( .A(n12546), .ZN(n11233) );
  OAI21_X1 U11671 ( .B1(n11273), .B2(n12443), .A(n11233), .ZN(n9231) );
  NAND2_X1 U11672 ( .A1(n11273), .A2(n12443), .ZN(n9230) );
  NAND2_X1 U11673 ( .A1(n9483), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11674 ( .A1(n6482), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9238) );
  OAI21_X1 U11675 ( .B1(n9232), .B2(P3_REG3_REG_9__SCAN_IN), .A(
        P3_REG3_REG_10__SCAN_IN), .ZN(n9235) );
  NOR2_X1 U11676 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_REG3_REG_10__SCAN_IN), 
        .ZN(n9233) );
  NAND2_X1 U11677 ( .A1(n9234), .A2(n9233), .ZN(n9251) );
  NAND2_X1 U11678 ( .A1(n9235), .A2(n9251), .ZN(n11579) );
  NAND2_X1 U11679 ( .A1(n6486), .A2(n11579), .ZN(n9237) );
  NAND2_X1 U11680 ( .A1(n12341), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9236) );
  NAND4_X1 U11681 ( .A1(n9239), .A2(n9238), .A3(n9237), .A4(n9236), .ZN(n12545) );
  INV_X1 U11682 ( .A(n12545), .ZN(n11277) );
  OR2_X1 U11683 ( .A1(n9241), .A2(n9240), .ZN(n9242) );
  NAND2_X1 U11684 ( .A1(n9243), .A2(n9242), .ZN(n9753) );
  NAND2_X1 U11685 ( .A1(n12338), .A2(n9753), .ZN(n9250) );
  INV_X1 U11686 ( .A(n9244), .ZN(n9246) );
  NAND2_X1 U11687 ( .A1(n9246), .A2(n9245), .ZN(n9261) );
  NAND2_X1 U11688 ( .A1(n9261), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9248) );
  INV_X1 U11689 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11690 ( .A1(n9279), .A2(n12557), .ZN(n9249) );
  OAI211_X1 U11691 ( .C1(SI_10_), .C2(n9382), .A(n9250), .B(n9249), .ZN(n11572) );
  INV_X1 U11692 ( .A(n11572), .ZN(n11316) );
  NAND2_X1 U11693 ( .A1(n11277), .A2(n11316), .ZN(n12445) );
  NAND2_X1 U11694 ( .A1(n12545), .A2(n11572), .ZN(n12446) );
  NAND2_X1 U11695 ( .A1(n12445), .A2(n12446), .ZN(n11257) );
  INV_X1 U11696 ( .A(n11398), .ZN(n9267) );
  NAND2_X1 U11697 ( .A1(n9483), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9258) );
  NAND2_X1 U11698 ( .A1(n9251), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11699 ( .A1(n9268), .A2(n9252), .ZN(n12296) );
  NAND2_X1 U11700 ( .A1(n6486), .A2(n12296), .ZN(n9257) );
  INV_X1 U11701 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9253) );
  OR2_X1 U11702 ( .A1(n9488), .A2(n9253), .ZN(n9256) );
  INV_X1 U11703 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9254) );
  OR2_X1 U11704 ( .A1(n9489), .A2(n9254), .ZN(n9255) );
  XNOR2_X1 U11705 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9259) );
  XNOR2_X1 U11706 ( .A(n9260), .B(n9259), .ZN(n9755) );
  NAND2_X1 U11707 ( .A1(n12338), .A2(n9755), .ZN(n9265) );
  OAI21_X1 U11708 ( .B1(n9261), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9263) );
  INV_X1 U11709 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9262) );
  XNOR2_X1 U11710 ( .A(n9263), .B(n9262), .ZN(n14962) );
  NAND2_X1 U11711 ( .A1(n9279), .A2(n14962), .ZN(n9264) );
  OAI211_X1 U11712 ( .C1(SI_11_), .C2(n9382), .A(n9265), .B(n9264), .ZN(n12294) );
  NAND2_X1 U11713 ( .A1(n12544), .A2(n12294), .ZN(n12397) );
  INV_X1 U11714 ( .A(n12294), .ZN(n14384) );
  NAND2_X1 U11715 ( .A1(n12290), .A2(n14384), .ZN(n12449) );
  NAND2_X1 U11716 ( .A1(n12397), .A2(n12449), .ZN(n12447) );
  NAND2_X1 U11717 ( .A1(n9267), .A2(n9266), .ZN(n11400) );
  NAND2_X1 U11718 ( .A1(n11400), .A2(n12449), .ZN(n11498) );
  NAND2_X1 U11719 ( .A1(n9529), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11720 ( .A1(n12341), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11721 ( .A1(n9268), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11722 ( .A1(n9285), .A2(n9269), .ZN(n12237) );
  NAND2_X1 U11723 ( .A1(n6486), .A2(n12237), .ZN(n9271) );
  NAND2_X1 U11724 ( .A1(n6482), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9270) );
  NAND4_X1 U11725 ( .A1(n9273), .A2(n9272), .A3(n9271), .A4(n9270), .ZN(n12543) );
  INV_X1 U11726 ( .A(n12543), .ZN(n11504) );
  XNOR2_X1 U11727 ( .A(n9275), .B(n9274), .ZN(n9756) );
  NAND2_X1 U11728 ( .A1(n12340), .A2(SI_12_), .ZN(n9281) );
  NAND2_X1 U11729 ( .A1(n9276), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9277) );
  MUX2_X1 U11730 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9277), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9278) );
  AND2_X1 U11731 ( .A1(n9278), .A2(n6603), .ZN(n12596) );
  NAND2_X1 U11732 ( .A1(n9279), .A2(n12596), .ZN(n9280) );
  OAI211_X1 U11733 ( .C1(n9756), .C2(n9381), .A(n9281), .B(n9280), .ZN(n11497)
         );
  NAND2_X1 U11734 ( .A1(n11504), .A2(n11497), .ZN(n12457) );
  INV_X1 U11735 ( .A(n11497), .ZN(n14379) );
  NAND2_X1 U11736 ( .A1(n12543), .A2(n14379), .ZN(n12450) );
  NAND2_X1 U11737 ( .A1(n12457), .A2(n12450), .ZN(n12367) );
  XNOR2_X1 U11738 ( .A(n9282), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U11739 ( .A1(n6603), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9283) );
  XNOR2_X1 U11740 ( .A(n9283), .B(n9015), .ZN(n14997) );
  INV_X1 U11741 ( .A(n14997), .ZN(n12599) );
  OAI22_X1 U11742 ( .A1(n9382), .A2(SI_13_), .B1(n12599), .B2(n9102), .ZN(
        n9284) );
  NAND2_X1 U11743 ( .A1(n6483), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11744 ( .A1(n9529), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9289) );
  INV_X1 U11745 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U11746 ( .A1(n9285), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11747 ( .A1(n9299), .A2(n9286), .ZN(n12024) );
  NAND2_X1 U11748 ( .A1(n6486), .A2(n12024), .ZN(n9288) );
  NAND2_X1 U11749 ( .A1(n12341), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9287) );
  NAND4_X1 U11750 ( .A1(n9290), .A2(n9289), .A3(n9288), .A4(n9287), .ZN(n12828) );
  INV_X1 U11751 ( .A(n12828), .ZN(n12201) );
  NAND2_X1 U11752 ( .A1(n14376), .A2(n12201), .ZN(n12459) );
  OR2_X1 U11753 ( .A1(n14376), .A2(n12201), .ZN(n12458) );
  NAND2_X1 U11754 ( .A1(n9291), .A2(n12458), .ZN(n12840) );
  INV_X1 U11755 ( .A(n12840), .ZN(n9306) );
  XNOR2_X1 U11756 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9292) );
  XNOR2_X1 U11757 ( .A(n9293), .B(n9292), .ZN(n9779) );
  NAND2_X1 U11758 ( .A1(n9779), .A2(n12338), .ZN(n9297) );
  OR2_X1 U11759 ( .A1(n9028), .A2(n12958), .ZN(n9294) );
  XNOR2_X1 U11760 ( .A(n9294), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12578) );
  OAI22_X1 U11761 ( .A1(n9382), .A2(SI_14_), .B1(n12578), .B2(n9102), .ZN(
        n9295) );
  INV_X1 U11762 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U11763 ( .A1(n9297), .A2(n9296), .ZN(n14369) );
  NAND2_X1 U11764 ( .A1(n9529), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U11765 ( .A1(n9298), .A2(n15195), .ZN(n9317) );
  NAND2_X1 U11766 ( .A1(n9299), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11767 ( .A1(n9317), .A2(n9300), .ZN(n12833) );
  NAND2_X1 U11768 ( .A1(n6486), .A2(n12833), .ZN(n9304) );
  INV_X1 U11769 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12835) );
  OR2_X1 U11770 ( .A1(n9488), .A2(n12835), .ZN(n9303) );
  INV_X1 U11771 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11772 ( .A1(n9489), .A2(n9301), .ZN(n9302) );
  INV_X1 U11773 ( .A(n12325), .ZN(n12542) );
  NAND2_X1 U11774 ( .A1(n14369), .A2(n12542), .ZN(n12462) );
  NAND2_X1 U11775 ( .A1(n9306), .A2(n12462), .ZN(n12820) );
  NAND2_X1 U11776 ( .A1(n9308), .A2(n9307), .ZN(n9309) );
  NAND2_X1 U11777 ( .A1(n9310), .A2(n9309), .ZN(n9914) );
  NAND2_X1 U11778 ( .A1(n9914), .A2(n12338), .ZN(n9316) );
  NAND2_X1 U11779 ( .A1(n9311), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11780 ( .A(n9313), .B(n9312), .ZN(n12604) );
  INV_X1 U11781 ( .A(n12604), .ZN(n14299) );
  OAI22_X1 U11782 ( .A1(n9382), .A2(SI_15_), .B1(n14299), .B2(n9102), .ZN(
        n9314) );
  INV_X1 U11783 ( .A(n9314), .ZN(n9315) );
  NAND2_X1 U11784 ( .A1(n9483), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11785 ( .A1(n9317), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11786 ( .A1(n9336), .A2(n9318), .ZN(n12814) );
  NAND2_X1 U11787 ( .A1(n6486), .A2(n12814), .ZN(n9322) );
  INV_X1 U11788 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n9319) );
  OR2_X1 U11789 ( .A1(n9489), .A2(n9319), .ZN(n9321) );
  INV_X1 U11790 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12816) );
  OR2_X1 U11791 ( .A1(n9488), .A2(n12816), .ZN(n9320) );
  AND2_X1 U11792 ( .A1(n12819), .A2(n12466), .ZN(n9324) );
  NAND2_X1 U11793 ( .A1(n12820), .A2(n9324), .ZN(n12777) );
  OR2_X1 U11794 ( .A1(n9326), .A2(n9325), .ZN(n9327) );
  NAND2_X1 U11795 ( .A1(n9328), .A2(n9327), .ZN(n9990) );
  OR2_X1 U11796 ( .A1(n9990), .A2(n9381), .ZN(n9335) );
  NAND2_X1 U11797 ( .A1(n9329), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9330) );
  MUX2_X1 U11798 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9330), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9332) );
  INV_X1 U11799 ( .A(n9331), .ZN(n9346) );
  NAND2_X1 U11800 ( .A1(n9332), .A2(n9346), .ZN(n12610) );
  OAI22_X1 U11801 ( .A1(n9382), .A2(n15194), .B1(n9102), .B2(n12610), .ZN(
        n9333) );
  INV_X1 U11802 ( .A(n9333), .ZN(n9334) );
  NAND2_X1 U11803 ( .A1(n6482), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11804 ( .A1(n9529), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9340) );
  INV_X1 U11805 ( .A(n9352), .ZN(n9353) );
  NAND2_X1 U11806 ( .A1(n9336), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U11807 ( .A1(n9353), .A2(n9337), .ZN(n12804) );
  NAND2_X1 U11808 ( .A1(n6486), .A2(n12804), .ZN(n9339) );
  NAND2_X1 U11809 ( .A1(n12341), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9338) );
  NAND4_X1 U11810 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n12541) );
  INV_X1 U11811 ( .A(n12541), .ZN(n12469) );
  OR2_X1 U11812 ( .A1(n12470), .A2(n12469), .ZN(n12464) );
  NAND2_X1 U11813 ( .A1(n12470), .A2(n12469), .ZN(n12779) );
  NAND2_X1 U11814 ( .A1(n14364), .A2(n12830), .ZN(n12800) );
  AND2_X1 U11815 ( .A1(n12802), .A2(n12800), .ZN(n12778) );
  OR2_X1 U11816 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  NAND2_X1 U11817 ( .A1(n9345), .A2(n9344), .ZN(n10079) );
  NAND2_X1 U11818 ( .A1(n10079), .A2(n12338), .ZN(n9351) );
  NAND2_X1 U11819 ( .A1(n9346), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9348) );
  XNOR2_X1 U11820 ( .A(n9348), .B(n9347), .ZN(n12612) );
  INV_X1 U11821 ( .A(n12612), .ZN(n14331) );
  OAI22_X1 U11822 ( .A1(n9382), .A2(SI_17_), .B1(n14331), .B2(n9102), .ZN(
        n9349) );
  INV_X1 U11823 ( .A(n9349), .ZN(n9350) );
  NAND2_X1 U11824 ( .A1(n6483), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11825 ( .A1(n9529), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9357) );
  INV_X1 U11826 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12260) );
  INV_X1 U11827 ( .A(n9369), .ZN(n9370) );
  NAND2_X1 U11828 ( .A1(n9353), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11829 ( .A1(n9370), .A2(n9354), .ZN(n12787) );
  NAND2_X1 U11830 ( .A1(n6486), .A2(n12787), .ZN(n9356) );
  NAND2_X1 U11831 ( .A1(n12341), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9355) );
  NAND4_X1 U11832 ( .A1(n9358), .A2(n9357), .A3(n9356), .A4(n9355), .ZN(n12796) );
  NAND2_X1 U11833 ( .A1(n12948), .A2(n12796), .ZN(n12475) );
  NAND2_X1 U11834 ( .A1(n12478), .A2(n12475), .ZN(n12472) );
  INV_X1 U11835 ( .A(n12472), .ZN(n12783) );
  AND2_X1 U11836 ( .A1(n12778), .A2(n12783), .ZN(n9359) );
  XNOR2_X1 U11837 ( .A(n9361), .B(n9360), .ZN(n10258) );
  NAND2_X1 U11838 ( .A1(n10258), .A2(n12338), .ZN(n9367) );
  NAND2_X1 U11839 ( .A1(n9362), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9364) );
  XNOR2_X1 U11840 ( .A(n9364), .B(n9363), .ZN(n12614) );
  OAI22_X1 U11841 ( .A1(n9382), .A2(n10259), .B1(n9102), .B2(n12614), .ZN(
        n9365) );
  INV_X1 U11842 ( .A(n9365), .ZN(n9366) );
  NAND2_X1 U11843 ( .A1(n9483), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9376) );
  INV_X1 U11844 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11845 ( .A1(n9370), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11846 ( .A1(n9395), .A2(n9371), .ZN(n12768) );
  NAND2_X1 U11847 ( .A1(n6486), .A2(n12768), .ZN(n9375) );
  INV_X1 U11848 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12770) );
  OR2_X1 U11849 ( .A1(n9488), .A2(n12770), .ZN(n9374) );
  INV_X1 U11850 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n9372) );
  OR2_X1 U11851 ( .A1(n9489), .A2(n9372), .ZN(n9373) );
  NAND2_X1 U11852 ( .A1(n12885), .A2(n9640), .ZN(n12477) );
  OR2_X1 U11853 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  NAND2_X1 U11854 ( .A1(n9380), .A2(n9379), .ZN(n12031) );
  OR2_X1 U11855 ( .A1(n12031), .A2(n9381), .ZN(n9385) );
  OAI22_X1 U11856 ( .A1(n9382), .A2(n15160), .B1(n6490), .B2(n9102), .ZN(n9383) );
  INV_X1 U11857 ( .A(n9383), .ZN(n9384) );
  NAND2_X1 U11858 ( .A1(n6482), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11859 ( .A1(n9529), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9388) );
  XNOR2_X1 U11860 ( .A(n9395), .B(P3_REG3_REG_19__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U11861 ( .A1(n6486), .A2(n12759), .ZN(n9387) );
  NAND2_X1 U11862 ( .A1(n12341), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9386) );
  NAND4_X1 U11863 ( .A1(n9389), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n12766) );
  INV_X1 U11864 ( .A(n12766), .ZN(n12275) );
  INV_X1 U11865 ( .A(n12481), .ZN(n9390) );
  NAND2_X1 U11866 ( .A1(n12215), .A2(n12275), .ZN(n12482) );
  OAI21_X1 U11867 ( .B1(n12752), .B2(n9390), .A(n12482), .ZN(n12738) );
  XNOR2_X1 U11868 ( .A(n9391), .B(n11936), .ZN(n10512) );
  NAND2_X1 U11869 ( .A1(n10512), .A2(n12338), .ZN(n9393) );
  NAND2_X1 U11870 ( .A1(n12340), .A2(SI_20_), .ZN(n9392) );
  NAND2_X1 U11871 ( .A1(n6483), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U11872 ( .A1(n9529), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9399) );
  OAI21_X1 U11873 ( .B1(n9395), .B2(P3_REG3_REG_19__SCAN_IN), .A(
        P3_REG3_REG_20__SCAN_IN), .ZN(n9396) );
  INV_X1 U11874 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15270) );
  INV_X1 U11875 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15251) );
  NAND2_X1 U11876 ( .A1(n15270), .A2(n15251), .ZN(n9394) );
  NAND2_X1 U11877 ( .A1(n9396), .A2(n9405), .ZN(n12747) );
  NAND2_X1 U11878 ( .A1(n6486), .A2(n12747), .ZN(n9398) );
  NAND2_X1 U11879 ( .A1(n12341), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9397) );
  NAND4_X1 U11880 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n12539) );
  XNOR2_X1 U11881 ( .A(n12486), .B(n12730), .ZN(n12740) );
  NAND2_X1 U11882 ( .A1(n12939), .A2(n12539), .ZN(n12487) );
  XNOR2_X1 U11883 ( .A(n9402), .B(n9401), .ZN(n10706) );
  NAND2_X1 U11884 ( .A1(n10706), .A2(n12338), .ZN(n9404) );
  NAND2_X1 U11885 ( .A1(n12340), .A2(SI_21_), .ZN(n9403) );
  NAND2_X1 U11886 ( .A1(n9529), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9412) );
  INV_X1 U11887 ( .A(n9417), .ZN(n9407) );
  NAND2_X1 U11888 ( .A1(n9405), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U11889 ( .A1(n9407), .A2(n9406), .ZN(n12732) );
  NAND2_X1 U11890 ( .A1(n6486), .A2(n12732), .ZN(n9411) );
  INV_X1 U11891 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9408) );
  OR2_X1 U11892 ( .A1(n9488), .A2(n9408), .ZN(n9410) );
  INV_X1 U11893 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12933) );
  OR2_X1 U11894 ( .A1(n9489), .A2(n12933), .ZN(n9409) );
  NAND2_X1 U11895 ( .A1(n12731), .A2(n12277), .ZN(n12491) );
  XNOR2_X1 U11896 ( .A(n9414), .B(n9413), .ZN(n10817) );
  NAND2_X1 U11897 ( .A1(n10817), .A2(n12338), .ZN(n9416) );
  NAND2_X1 U11898 ( .A1(n12340), .A2(SI_22_), .ZN(n9415) );
  NAND2_X1 U11899 ( .A1(n6482), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11900 ( .A1(n9483), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11901 ( .A1(n9417), .A2(n15219), .ZN(n9427) );
  OR2_X1 U11902 ( .A1(n9417), .A2(n15219), .ZN(n9418) );
  NAND2_X1 U11903 ( .A1(n9427), .A2(n9418), .ZN(n12720) );
  NAND2_X1 U11904 ( .A1(n6486), .A2(n12720), .ZN(n9420) );
  NAND2_X1 U11905 ( .A1(n12341), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9419) );
  NAND4_X1 U11906 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n12538) );
  AND2_X1 U11907 ( .A1(n9653), .A2(n12729), .ZN(n12396) );
  XNOR2_X1 U11908 ( .A(n9424), .B(n9423), .ZN(n10932) );
  NAND2_X1 U11909 ( .A1(n10932), .A2(n12338), .ZN(n9426) );
  NAND2_X1 U11910 ( .A1(n12340), .A2(SI_23_), .ZN(n9425) );
  NAND2_X1 U11911 ( .A1(n9427), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11912 ( .A1(n9428), .A2(n9440), .ZN(n12709) );
  NAND2_X1 U11913 ( .A1(n12709), .A2(n6486), .ZN(n9432) );
  NAND2_X1 U11914 ( .A1(n6483), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U11915 ( .A1(n9529), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U11916 ( .A1(n12341), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9429) );
  NAND4_X1 U11917 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(n12537) );
  INV_X1 U11918 ( .A(n12537), .ZN(n9433) );
  NAND2_X1 U11919 ( .A1(n12395), .A2(n9433), .ZN(n9434) );
  NAND2_X1 U11920 ( .A1(n12497), .A2(n9434), .ZN(n12705) );
  INV_X1 U11921 ( .A(n12705), .ZN(n9436) );
  INV_X1 U11922 ( .A(n12497), .ZN(n9435) );
  AOI21_X1 U11923 ( .B1(n12704), .B2(n9436), .A(n9435), .ZN(n12698) );
  INV_X1 U11924 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14164) );
  XNOR2_X1 U11925 ( .A(n9437), .B(n14164), .ZN(n11288) );
  NAND2_X1 U11926 ( .A1(n11288), .A2(n12338), .ZN(n9439) );
  NAND2_X1 U11927 ( .A1(n12340), .A2(SI_24_), .ZN(n9438) );
  NAND2_X1 U11928 ( .A1(n9529), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11929 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9440), .ZN(n9441) );
  INV_X1 U11930 ( .A(n9451), .ZN(n9453) );
  NAND2_X1 U11931 ( .A1(n9441), .A2(n9453), .ZN(n12699) );
  NAND2_X1 U11932 ( .A1(n6486), .A2(n12699), .ZN(n9445) );
  INV_X1 U11933 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n9442) );
  OR2_X1 U11934 ( .A1(n9488), .A2(n9442), .ZN(n9444) );
  INV_X1 U11935 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12921) );
  OR2_X1 U11936 ( .A1(n9489), .A2(n12921), .ZN(n9443) );
  OR2_X1 U11937 ( .A1(n9664), .A2(n12708), .ZN(n12496) );
  NAND2_X1 U11938 ( .A1(n9664), .A2(n12708), .ZN(n12495) );
  NAND2_X1 U11939 ( .A1(n12698), .A2(n12697), .ZN(n12696) );
  NAND2_X1 U11940 ( .A1(n12696), .A2(n12495), .ZN(n12682) );
  XNOR2_X1 U11941 ( .A(n13556), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9447) );
  XNOR2_X1 U11942 ( .A(n9448), .B(n9447), .ZN(n11681) );
  NAND2_X1 U11943 ( .A1(n11681), .A2(n12338), .ZN(n9450) );
  NAND2_X1 U11944 ( .A1(n12340), .A2(SI_25_), .ZN(n9449) );
  NAND2_X1 U11945 ( .A1(n9529), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9459) );
  INV_X1 U11946 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U11947 ( .A1(n9452), .A2(n9451), .ZN(n9465) );
  NAND2_X1 U11948 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n9453), .ZN(n9454) );
  NAND2_X1 U11949 ( .A1(n9465), .A2(n9454), .ZN(n12687) );
  NAND2_X1 U11950 ( .A1(n6486), .A2(n12687), .ZN(n9458) );
  INV_X1 U11951 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n9455) );
  OR2_X1 U11952 ( .A1(n9488), .A2(n9455), .ZN(n9457) );
  INV_X1 U11953 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12917) );
  OR2_X1 U11954 ( .A1(n9489), .A2(n12917), .ZN(n9456) );
  XNOR2_X1 U11955 ( .A(n12501), .B(n12669), .ZN(n12676) );
  INV_X1 U11956 ( .A(n12676), .ZN(n12681) );
  XNOR2_X1 U11957 ( .A(n13551), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9460) );
  XNOR2_X1 U11958 ( .A(n9461), .B(n9460), .ZN(n11361) );
  NAND2_X1 U11959 ( .A1(n11361), .A2(n12338), .ZN(n9463) );
  NAND2_X1 U11960 ( .A1(n12340), .A2(SI_26_), .ZN(n9462) );
  NAND2_X1 U11961 ( .A1(n6482), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11962 ( .A1(n9529), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9469) );
  INV_X1 U11963 ( .A(n9465), .ZN(n9464) );
  INV_X1 U11964 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U11965 ( .A1(n9464), .A2(n15222), .ZN(n9475) );
  NAND2_X1 U11966 ( .A1(n9465), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U11967 ( .A1(n9475), .A2(n9466), .ZN(n12671) );
  NAND2_X1 U11968 ( .A1(n6486), .A2(n12671), .ZN(n9468) );
  NAND2_X1 U11969 ( .A1(n12341), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9467) );
  INV_X1 U11970 ( .A(n12678), .ZN(n12505) );
  XNOR2_X1 U11971 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9471) );
  XNOR2_X1 U11972 ( .A(n9472), .B(n9471), .ZN(n11488) );
  NAND2_X1 U11973 ( .A1(n11488), .A2(n12338), .ZN(n9474) );
  NAND2_X1 U11974 ( .A1(n12340), .A2(SI_27_), .ZN(n9473) );
  NAND2_X1 U11975 ( .A1(n9483), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U11976 ( .A1(n6483), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U11977 ( .A1(n9475), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U11978 ( .A1(n9486), .A2(n9476), .ZN(n12660) );
  NAND2_X1 U11979 ( .A1(n6486), .A2(n12660), .ZN(n9478) );
  NAND2_X1 U11980 ( .A1(n12341), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9477) );
  NAND4_X1 U11981 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(n12535) );
  NAND2_X1 U11982 ( .A1(n9676), .A2(n12670), .ZN(n9573) );
  OR2_X1 U11983 ( .A1(n9676), .A2(n12670), .ZN(n9481) );
  INV_X1 U11984 ( .A(n9573), .ZN(n9482) );
  NOR2_X1 U11985 ( .A1(n9575), .A2(n9482), .ZN(n9494) );
  NAND2_X1 U11986 ( .A1(n9483), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9493) );
  INV_X1 U11987 ( .A(n9486), .ZN(n9485) );
  INV_X1 U11988 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U11989 ( .A1(n9485), .A2(n9484), .ZN(n9528) );
  NAND2_X1 U11990 ( .A1(n9486), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U11991 ( .A1(n9528), .A2(n9487), .ZN(n12180) );
  NAND2_X1 U11992 ( .A1(n6486), .A2(n12180), .ZN(n9492) );
  INV_X1 U11993 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12645) );
  OR2_X1 U11994 ( .A1(n9488), .A2(n12645), .ZN(n9491) );
  OR2_X1 U11995 ( .A1(n9489), .A2(n9087), .ZN(n9490) );
  NAND2_X1 U11996 ( .A1(n12647), .A2(n12655), .ZN(n9574) );
  XNOR2_X1 U11997 ( .A(n9494), .B(n12378), .ZN(n12648) );
  NAND2_X1 U11998 ( .A1(n12555), .A2(n10636), .ZN(n9596) );
  INV_X1 U11999 ( .A(n9495), .ZN(n9592) );
  NAND2_X1 U12000 ( .A1(n9592), .A2(n15031), .ZN(n9496) );
  NAND2_X1 U12001 ( .A1(n10659), .A2(n12363), .ZN(n9498) );
  NAND2_X1 U12002 ( .A1(n15039), .A2(n10905), .ZN(n9497) );
  NAND2_X1 U12003 ( .A1(n9498), .A2(n9497), .ZN(n11092) );
  INV_X1 U12004 ( .A(n11092), .ZN(n9500) );
  INV_X1 U12005 ( .A(n12357), .ZN(n9499) );
  NAND2_X1 U12006 ( .A1(n12552), .A2(n9587), .ZN(n9501) );
  NAND2_X1 U12007 ( .A1(n11094), .A2(n9501), .ZN(n10776) );
  NAND2_X1 U12008 ( .A1(n12419), .A2(n10971), .ZN(n9503) );
  AND2_X1 U12009 ( .A1(n12414), .A2(n9503), .ZN(n10936) );
  AND2_X1 U12010 ( .A1(n6476), .A2(n10936), .ZN(n9502) );
  NAND2_X1 U12011 ( .A1(n10776), .A2(n9502), .ZN(n10940) );
  NAND2_X1 U12012 ( .A1(n12551), .A2(n10833), .ZN(n10866) );
  INV_X1 U12013 ( .A(n10941), .ZN(n9505) );
  NAND2_X1 U12014 ( .A1(n10940), .A2(n9506), .ZN(n10996) );
  NAND2_X1 U12015 ( .A1(n12548), .A2(n14848), .ZN(n9507) );
  NAND2_X1 U12016 ( .A1(n11278), .A2(n15062), .ZN(n9508) );
  NAND2_X1 U12017 ( .A1(n11176), .A2(n9508), .ZN(n9510) );
  NAND2_X1 U12018 ( .A1(n12547), .A2(n11236), .ZN(n9509) );
  NAND2_X1 U12019 ( .A1(n9510), .A2(n9509), .ZN(n11274) );
  XNOR2_X1 U12020 ( .A(n12546), .B(n15069), .ZN(n11276) );
  NAND2_X1 U12021 ( .A1(n12546), .A2(n12443), .ZN(n9511) );
  NAND2_X1 U12022 ( .A1(n11394), .A2(n12447), .ZN(n9513) );
  NAND2_X1 U12023 ( .A1(n12544), .A2(n14384), .ZN(n9512) );
  NAND2_X1 U12024 ( .A1(n9513), .A2(n9512), .ZN(n11491) );
  NAND2_X1 U12025 ( .A1(n12543), .A2(n11497), .ZN(n9514) );
  NAND2_X1 U12026 ( .A1(n12458), .A2(n12459), .ZN(n12454) );
  NAND2_X1 U12027 ( .A1(n12819), .A2(n12462), .ZN(n12839) );
  NAND2_X1 U12028 ( .A1(n12825), .A2(n12839), .ZN(n9516) );
  OR2_X1 U12029 ( .A1(n14369), .A2(n12325), .ZN(n9515) );
  NAND2_X1 U12030 ( .A1(n14364), .A2(n12254), .ZN(n9517) );
  NAND2_X1 U12031 ( .A1(n12470), .A2(n12541), .ZN(n12782) );
  NAND2_X1 U12032 ( .A1(n7450), .A2(n12782), .ZN(n9518) );
  NAND2_X1 U12033 ( .A1(n9518), .A2(n12472), .ZN(n12781) );
  INV_X1 U12034 ( .A(n12796), .ZN(n12307) );
  OR2_X1 U12035 ( .A1(n12948), .A2(n12307), .ZN(n9519) );
  NAND2_X1 U12036 ( .A1(n12481), .A2(n12482), .ZN(n12754) );
  INV_X1 U12037 ( .A(n9640), .ZN(n12540) );
  OR2_X1 U12038 ( .A1(n12885), .A2(n12540), .ZN(n12755) );
  AND2_X1 U12039 ( .A1(n12754), .A2(n12755), .ZN(n9520) );
  NAND2_X1 U12040 ( .A1(n12215), .A2(n12766), .ZN(n9521) );
  NAND2_X1 U12041 ( .A1(n12753), .A2(n9521), .ZN(n12741) );
  AND2_X2 U12042 ( .A1(n12741), .A2(n12740), .ZN(n12743) );
  NOR2_X1 U12043 ( .A1(n12731), .A2(n12744), .ZN(n12355) );
  NAND2_X1 U12044 ( .A1(n12731), .A2(n12744), .ZN(n12353) );
  INV_X1 U12045 ( .A(n12708), .ZN(n12679) );
  NOR2_X1 U12046 ( .A1(n9664), .A2(n12679), .ZN(n9522) );
  NAND2_X1 U12047 ( .A1(n9044), .A2(n12529), .ZN(n9526) );
  NAND2_X1 U12048 ( .A1(n12398), .A2(n9582), .ZN(n9525) );
  OAI211_X1 U12049 ( .C1(n9527), .C2(n12511), .A(n9558), .B(n12832), .ZN(n9537) );
  INV_X1 U12050 ( .A(n9528), .ZN(n12632) );
  NAND2_X1 U12051 ( .A1(n6486), .A2(n12632), .ZN(n12345) );
  NAND2_X1 U12052 ( .A1(n6483), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U12053 ( .A1(n9529), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9531) );
  NAND2_X1 U12054 ( .A1(n12341), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9530) );
  NAND4_X1 U12055 ( .A1(n12345), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(
        n12534) );
  INV_X1 U12056 ( .A(n11956), .ZN(n12527) );
  NAND2_X1 U12057 ( .A1(n12527), .A2(n6475), .ZN(n10057) );
  NAND2_X1 U12058 ( .A1(n12534), .A2(n12797), .ZN(n9535) );
  NAND2_X1 U12059 ( .A1(n12535), .A2(n12827), .ZN(n9534) );
  NAND2_X1 U12060 ( .A1(n9535), .A2(n9534), .ZN(n12181) );
  INV_X1 U12061 ( .A(n12181), .ZN(n9536) );
  OAI21_X1 U12062 ( .B1(n14372), .B2(n12648), .A(n12652), .ZN(n9552) );
  XNOR2_X1 U12063 ( .A(n12956), .B(n12954), .ZN(n9542) );
  NAND2_X1 U12064 ( .A1(n10043), .A2(n9540), .ZN(n9541) );
  OAI22_X1 U12065 ( .A1(n9044), .A2(n9543), .B1(n9582), .B2(n15068), .ZN(n9544) );
  NAND2_X1 U12066 ( .A1(n9544), .A2(n9547), .ZN(n9545) );
  NAND2_X1 U12067 ( .A1(n9545), .A2(n12514), .ZN(n9546) );
  NAND2_X1 U12068 ( .A1(n9546), .A2(n10803), .ZN(n9550) );
  NAND2_X1 U12069 ( .A1(n9547), .A2(n12504), .ZN(n9690) );
  NAND2_X1 U12070 ( .A1(n9548), .A2(n12514), .ZN(n10805) );
  NAND2_X1 U12071 ( .A1(n9690), .A2(n10805), .ZN(n10804) );
  NAND2_X1 U12072 ( .A1(n10804), .A2(n12954), .ZN(n9549) );
  NAND2_X1 U12073 ( .A1(n9552), .A2(n15085), .ZN(n9556) );
  INV_X1 U12074 ( .A(n15085), .ZN(n9553) );
  AOI22_X1 U12075 ( .A1(n12647), .A2(n9554), .B1(P3_REG1_REG_28__SCAN_IN), 
        .B2(n9553), .ZN(n9555) );
  NAND2_X1 U12076 ( .A1(n9556), .A2(n9555), .ZN(P3_U3487) );
  NOR2_X1 U12077 ( .A1(n9559), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U12078 ( .A1(n9559), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9560) );
  OAI21_X2 U12079 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n12187) );
  XNOR2_X1 U12080 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12186) );
  XNOR2_X1 U12081 ( .A(n12187), .B(n12186), .ZN(n12964) );
  NAND2_X1 U12082 ( .A1(n12964), .A2(n12338), .ZN(n9564) );
  NAND2_X1 U12083 ( .A1(n12340), .A2(SI_29_), .ZN(n9563) );
  NAND2_X1 U12084 ( .A1(n9564), .A2(n9563), .ZN(n9578) );
  INV_X1 U12085 ( .A(n12534), .ZN(n9565) );
  NAND2_X1 U12086 ( .A1(n9578), .A2(n9565), .ZN(n12519) );
  XNOR2_X1 U12087 ( .A(n9566), .B(n12379), .ZN(n9572) );
  NAND2_X1 U12088 ( .A1(n6482), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U12089 ( .A1(n9529), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U12090 ( .A1(n12341), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U12091 ( .A1(n12527), .A2(P3_B_REG_SCAN_IN), .ZN(n9570) );
  NAND2_X1 U12092 ( .A1(n12797), .A2(n9570), .ZN(n12629) );
  OAI22_X1 U12093 ( .A1(n12348), .A2(n12629), .B1(n12655), .B2(n15042), .ZN(
        n9571) );
  NAND2_X1 U12094 ( .A1(n9574), .A2(n9573), .ZN(n12394) );
  INV_X1 U12095 ( .A(n12379), .ZN(n9576) );
  XNOR2_X1 U12096 ( .A(n12346), .B(n9576), .ZN(n12640) );
  NAND2_X1 U12097 ( .A1(n12640), .A2(n15054), .ZN(n9577) );
  INV_X1 U12098 ( .A(n9578), .ZN(n12637) );
  NAND2_X1 U12099 ( .A1(n9579), .A2(n7442), .ZN(P3_U3488) );
  NAND2_X1 U12100 ( .A1(n9581), .A2(n7443), .ZN(P3_U3456) );
  XNOR2_X1 U12102 ( .A(n6484), .B(n10821), .ZN(n9603) );
  INV_X1 U12103 ( .A(n9603), .ZN(n9604) );
  XNOR2_X1 U12104 ( .A(n9587), .B(n6484), .ZN(n9601) );
  INV_X1 U12105 ( .A(n9588), .ZN(n9589) );
  NAND2_X1 U12106 ( .A1(n9589), .A2(n10737), .ZN(n9597) );
  INV_X1 U12107 ( .A(n15031), .ZN(n10742) );
  AND2_X1 U12108 ( .A1(n6484), .A2(n10742), .ZN(n9593) );
  AOI21_X1 U12109 ( .B1(n9592), .B2(n9590), .A(n9591), .ZN(n9594) );
  NOR2_X1 U12110 ( .A1(n9594), .A2(n9593), .ZN(n9598) );
  NAND3_X1 U12111 ( .A1(n9597), .A2(n10741), .A3(n9596), .ZN(n10740) );
  INV_X1 U12112 ( .A(n9598), .ZN(n9599) );
  XNOR2_X1 U12113 ( .A(n9590), .B(n10905), .ZN(n9600) );
  XNOR2_X1 U12114 ( .A(n9600), .B(n12553), .ZN(n10612) );
  XOR2_X1 U12115 ( .A(n12551), .B(n9603), .Z(n10832) );
  XNOR2_X1 U12116 ( .A(n9675), .B(n10971), .ZN(n9605) );
  XNOR2_X1 U12117 ( .A(n9605), .B(n12550), .ZN(n10970) );
  XNOR2_X1 U12118 ( .A(n9675), .B(n10947), .ZN(n9606) );
  XOR2_X1 U12119 ( .A(n12549), .B(n9606), .Z(n11026) );
  NAND2_X1 U12120 ( .A1(n9606), .A2(n12549), .ZN(n9607) );
  NAND2_X1 U12121 ( .A1(n11025), .A2(n9607), .ZN(n14845) );
  XNOR2_X1 U12122 ( .A(n12436), .B(n9675), .ZN(n14844) );
  INV_X1 U12123 ( .A(n14844), .ZN(n9608) );
  NAND2_X1 U12124 ( .A1(n9608), .A2(n12548), .ZN(n9609) );
  NAND2_X1 U12125 ( .A1(n14843), .A2(n9609), .ZN(n11231) );
  XNOR2_X1 U12126 ( .A(n9675), .B(n11236), .ZN(n9610) );
  XOR2_X1 U12127 ( .A(n12547), .B(n9610), .Z(n11230) );
  NAND2_X1 U12128 ( .A1(n9610), .A2(n12547), .ZN(n9611) );
  NAND2_X1 U12129 ( .A1(n11229), .A2(n9611), .ZN(n11366) );
  INV_X1 U12130 ( .A(n11366), .ZN(n9613) );
  XNOR2_X1 U12131 ( .A(n9675), .B(n15069), .ZN(n9614) );
  XOR2_X1 U12132 ( .A(n12546), .B(n9614), .Z(n11367) );
  INV_X1 U12133 ( .A(n11367), .ZN(n9612) );
  NAND2_X1 U12134 ( .A1(n9614), .A2(n11233), .ZN(n9615) );
  XNOR2_X1 U12135 ( .A(n9675), .B(n11572), .ZN(n9617) );
  XOR2_X1 U12136 ( .A(n12545), .B(n9617), .Z(n11576) );
  INV_X1 U12137 ( .A(n9617), .ZN(n9618) );
  NAND2_X1 U12138 ( .A1(n9618), .A2(n12545), .ZN(n9619) );
  XNOR2_X1 U12139 ( .A(n9675), .B(n12294), .ZN(n9620) );
  XNOR2_X1 U12140 ( .A(n9675), .B(n11497), .ZN(n12231) );
  NAND2_X1 U12141 ( .A1(n12231), .A2(n12543), .ZN(n9622) );
  OAI21_X1 U12142 ( .B1(n9620), .B2(n12290), .A(n9622), .ZN(n9625) );
  INV_X1 U12143 ( .A(n9620), .ZN(n12229) );
  NOR2_X1 U12144 ( .A1(n12229), .A2(n12544), .ZN(n9623) );
  INV_X1 U12145 ( .A(n12231), .ZN(n9621) );
  AOI22_X1 U12146 ( .A1(n9623), .A2(n9622), .B1(n11504), .B2(n9621), .ZN(n9624) );
  XNOR2_X1 U12147 ( .A(n14376), .B(n9675), .ZN(n12022) );
  NOR2_X1 U12148 ( .A1(n12022), .A2(n12828), .ZN(n12193) );
  XNOR2_X1 U12149 ( .A(n14369), .B(n9675), .ZN(n9628) );
  NAND2_X1 U12150 ( .A1(n9628), .A2(n12325), .ZN(n9627) );
  INV_X1 U12151 ( .A(n9627), .ZN(n9630) );
  OR2_X1 U12152 ( .A1(n12193), .A2(n9630), .ZN(n9626) );
  NOR2_X1 U12153 ( .A1(n12021), .A2(n9626), .ZN(n9633) );
  OAI21_X1 U12154 ( .B1(n9628), .B2(n12325), .A(n9627), .ZN(n12199) );
  INV_X1 U12155 ( .A(n12199), .ZN(n9629) );
  NAND2_X1 U12156 ( .A1(n12022), .A2(n12828), .ZN(n12194) );
  AND2_X1 U12157 ( .A1(n9629), .A2(n12194), .ZN(n12195) );
  NOR2_X1 U12158 ( .A1(n9630), .A2(n12195), .ZN(n9631) );
  XNOR2_X1 U12159 ( .A(n14364), .B(n9675), .ZN(n12321) );
  OR2_X1 U12160 ( .A1(n9631), .A2(n12830), .ZN(n9632) );
  OR2_X1 U12161 ( .A1(n9633), .A2(n9632), .ZN(n9634) );
  NAND2_X1 U12162 ( .A1(n9635), .A2(n9634), .ZN(n12250) );
  XNOR2_X1 U12163 ( .A(n12470), .B(n9675), .ZN(n9637) );
  XNOR2_X1 U12164 ( .A(n9637), .B(n12541), .ZN(n12249) );
  INV_X1 U12165 ( .A(n12249), .ZN(n9636) );
  NAND2_X1 U12166 ( .A1(n9637), .A2(n12541), .ZN(n9638) );
  XNOR2_X1 U12167 ( .A(n12948), .B(n9675), .ZN(n9642) );
  XNOR2_X1 U12168 ( .A(n9642), .B(n12796), .ZN(n12258) );
  XNOR2_X1 U12169 ( .A(n12885), .B(n10737), .ZN(n9641) );
  NAND2_X1 U12170 ( .A1(n9641), .A2(n9640), .ZN(n9639) );
  AND2_X1 U12171 ( .A1(n12258), .A2(n9639), .ZN(n9646) );
  INV_X1 U12172 ( .A(n9639), .ZN(n12301) );
  NOR2_X1 U12173 ( .A1(n9641), .A2(n9640), .ZN(n12302) );
  INV_X1 U12174 ( .A(n12302), .ZN(n9644) );
  INV_X1 U12175 ( .A(n9642), .ZN(n9643) );
  NAND2_X1 U12176 ( .A1(n9643), .A2(n12796), .ZN(n12299) );
  AND2_X1 U12177 ( .A1(n9644), .A2(n12299), .ZN(n9645) );
  XNOR2_X1 U12178 ( .A(n12215), .B(n9675), .ZN(n9647) );
  XNOR2_X1 U12179 ( .A(n9647), .B(n12766), .ZN(n12213) );
  NAND2_X1 U12180 ( .A1(n9647), .A2(n12766), .ZN(n9648) );
  XNOR2_X1 U12181 ( .A(n12486), .B(n9675), .ZN(n9649) );
  XOR2_X1 U12182 ( .A(n12539), .B(n9649), .Z(n12274) );
  INV_X1 U12183 ( .A(n9649), .ZN(n9650) );
  XNOR2_X1 U12184 ( .A(n12731), .B(n10737), .ZN(n9651) );
  NAND2_X1 U12185 ( .A1(n9651), .A2(n12277), .ZN(n9652) );
  OAI21_X1 U12186 ( .B1(n9651), .B2(n12277), .A(n9652), .ZN(n12223) );
  NAND2_X1 U12187 ( .A1(n12220), .A2(n9652), .ZN(n9657) );
  INV_X1 U12188 ( .A(n9657), .ZN(n9655) );
  XOR2_X1 U12189 ( .A(n9675), .B(n9653), .Z(n9656) );
  INV_X1 U12190 ( .A(n9656), .ZN(n9654) );
  INV_X1 U12191 ( .A(n9663), .ZN(n9661) );
  XOR2_X1 U12192 ( .A(n9675), .B(n12395), .Z(n9662) );
  INV_X1 U12193 ( .A(n9662), .ZN(n9660) );
  XNOR2_X1 U12194 ( .A(n9664), .B(n10737), .ZN(n9665) );
  NAND2_X1 U12195 ( .A1(n9665), .A2(n12708), .ZN(n12242) );
  INV_X1 U12196 ( .A(n9665), .ZN(n9666) );
  NAND2_X1 U12197 ( .A1(n9666), .A2(n12679), .ZN(n9667) );
  XNOR2_X1 U12198 ( .A(n12501), .B(n10737), .ZN(n9669) );
  NAND2_X1 U12199 ( .A1(n9669), .A2(n12669), .ZN(n9672) );
  INV_X1 U12200 ( .A(n9669), .ZN(n9670) );
  NAND2_X1 U12201 ( .A1(n9670), .A2(n12536), .ZN(n9671) );
  NAND2_X1 U12202 ( .A1(n9672), .A2(n9671), .ZN(n12241) );
  XNOR2_X1 U12203 ( .A(n12506), .B(n9675), .ZN(n9673) );
  NOR2_X1 U12204 ( .A1(n9673), .A2(n12678), .ZN(n9674) );
  AOI21_X1 U12205 ( .B1(n9673), .B2(n12678), .A(n9674), .ZN(n12313) );
  INV_X1 U12206 ( .A(n9674), .ZN(n12174) );
  XNOR2_X1 U12207 ( .A(n9676), .B(n9675), .ZN(n9677) );
  NOR2_X1 U12208 ( .A1(n9677), .A2(n12535), .ZN(n12173) );
  XNOR2_X1 U12209 ( .A(n9678), .B(n12176), .ZN(n9682) );
  NAND2_X1 U12210 ( .A1(n9687), .A2(n15068), .ZN(n9680) );
  INV_X1 U12211 ( .A(n9689), .ZN(n9679) );
  OAI22_X1 U12212 ( .A1(n9680), .A2(n9688), .B1(n9694), .B2(n9679), .ZN(n9681)
         );
  NAND2_X1 U12213 ( .A1(n9682), .A2(n14857), .ZN(n9705) );
  INV_X1 U12214 ( .A(n10043), .ZN(n9683) );
  NAND2_X1 U12215 ( .A1(n9684), .A2(n9685), .ZN(n9686) );
  NAND2_X1 U12216 ( .A1(n9688), .A2(n9687), .ZN(n9692) );
  NAND2_X1 U12217 ( .A1(n9694), .A2(n9689), .ZN(n9691) );
  NAND4_X1 U12218 ( .A1(n9692), .A2(n9709), .A3(n9691), .A4(n9690), .ZN(n9693)
         );
  NAND2_X1 U12219 ( .A1(n9693), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9696) );
  NAND3_X1 U12220 ( .A1(n10606), .A2(n10043), .A3(n9694), .ZN(n9695) );
  AND2_X1 U12221 ( .A1(n9696), .A2(n9695), .ZN(n10613) );
  INV_X1 U12222 ( .A(n10040), .ZN(n9697) );
  NAND2_X1 U12223 ( .A1(n9697), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12531) );
  AND2_X1 U12224 ( .A1(n12524), .A2(n10043), .ZN(n12526) );
  NAND2_X1 U12225 ( .A1(n14865), .A2(n12827), .ZN(n12317) );
  NOR2_X1 U12226 ( .A1(n12505), .A2(n12317), .ZN(n9701) );
  NAND2_X1 U12227 ( .A1(n14865), .A2(n12797), .ZN(n12276) );
  INV_X1 U12228 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9699) );
  OAI22_X1 U12229 ( .A1(n12655), .A2(n12276), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9699), .ZN(n9700) );
  AOI211_X1 U12230 ( .C1(n12660), .C2(n12326), .A(n9701), .B(n9700), .ZN(n9702) );
  INV_X1 U12231 ( .A(n9703), .ZN(n9704) );
  NAND2_X1 U12232 ( .A1(n9705), .A2(n9704), .ZN(P3_U3154) );
  INV_X1 U12233 ( .A(n9706), .ZN(n9707) );
  INV_X1 U12234 ( .A(n9730), .ZN(n9708) );
  INV_X1 U12235 ( .A(n9709), .ZN(n9710) );
  NOR2_X1 U12236 ( .A1(n9735), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13543) );
  NAND2_X1 U12237 ( .A1(n9735), .A2(P2_U3088), .ZN(n13559) );
  OAI222_X1 U12238 ( .A1(n13550), .A2(n9711), .B1(n13559), .B2(n9760), .C1(
        n14660), .C2(P2_U3088), .ZN(P2_U3326) );
  NAND2_X1 U12239 ( .A1(n7495), .A2(P3_U3151), .ZN(n12191) );
  NAND2_X1 U12240 ( .A1(n9735), .A2(P3_U3151), .ZN(n12968) );
  OAI222_X1 U12241 ( .A1(n12191), .A2(n9713), .B1(n12968), .B2(n9712), .C1(
        P3_U3151), .C2(n10182), .ZN(P3_U3294) );
  INV_X1 U12242 ( .A(SI_8_), .ZN(n9714) );
  OAI222_X1 U12243 ( .A1(n12191), .A2(n9715), .B1(n12968), .B2(n9714), .C1(
        P3_U3151), .C2(n11203), .ZN(P3_U3287) );
  OAI222_X1 U12244 ( .A1(P3_U3151), .A2(n10754), .B1(n12968), .B2(n9717), .C1(
        n12191), .C2(n9716), .ZN(P3_U3288) );
  INV_X1 U12245 ( .A(SI_9_), .ZN(n9718) );
  OAI222_X1 U12246 ( .A1(n11195), .A2(P3_U3151), .B1(n12191), .B2(n9719), .C1(
        n9718), .C2(n12968), .ZN(P3_U3286) );
  INV_X1 U12247 ( .A(n13559), .ZN(n11389) );
  INV_X1 U12248 ( .A(n11389), .ZN(n13552) );
  INV_X1 U12249 ( .A(n9720), .ZN(n9742) );
  OAI222_X1 U12250 ( .A1(n13550), .A2(n9721), .B1(n13552), .B2(n9742), .C1(
        P2_U3088), .C2(n10004), .ZN(P2_U3325) );
  INV_X1 U12251 ( .A(n9722), .ZN(n9737) );
  INV_X1 U12252 ( .A(n9881), .ZN(n10106) );
  OAI222_X1 U12253 ( .A1(n13550), .A2(n9723), .B1(n13552), .B2(n9737), .C1(
        P2_U3088), .C2(n10106), .ZN(P2_U3323) );
  INV_X1 U12254 ( .A(n9724), .ZN(n9762) );
  INV_X1 U12255 ( .A(n9880), .ZN(n14679) );
  OAI222_X1 U12256 ( .A1(n13550), .A2(n9725), .B1(n13552), .B2(n9762), .C1(
        P2_U3088), .C2(n14679), .ZN(P2_U3324) );
  INV_X1 U12257 ( .A(n9726), .ZN(n9740) );
  OAI222_X1 U12258 ( .A1(n13550), .A2(n9727), .B1(n13552), .B2(n9740), .C1(
        P2_U3088), .C2(n10093), .ZN(P2_U3322) );
  NAND2_X1 U12259 ( .A1(n9943), .A2(n10125), .ZN(n14581) );
  INV_X1 U12260 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9729) );
  INV_X1 U12261 ( .A(n10123), .ZN(n9728) );
  AOI22_X1 U12262 ( .A1(n14581), .A2(n9729), .B1(n9730), .B2(n9728), .ZN(
        P1_U3446) );
  INV_X1 U12263 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9732) );
  AND2_X1 U12264 ( .A1(n9730), .A2(n14160), .ZN(n9731) );
  AOI22_X1 U12265 ( .A1(n14581), .A2(n9732), .B1(n9731), .B2(n14167), .ZN(
        P1_U3445) );
  INV_X1 U12266 ( .A(n12191), .ZN(n10931) );
  INV_X1 U12267 ( .A(n12968), .ZN(n12961) );
  AOI222_X1 U12268 ( .A1(n9733), .A2(n10931), .B1(n10456), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n12961), .C2(SI_3_), .ZN(n9734) );
  INV_X1 U12269 ( .A(n9734), .ZN(P3_U3292) );
  INV_X1 U12270 ( .A(n13762), .ZN(n9738) );
  OAI222_X1 U12271 ( .A1(n9738), .A2(P1_U3086), .B1(n14166), .B2(n9737), .C1(
        n9736), .C2(n14163), .ZN(P1_U3351) );
  OAI222_X1 U12272 ( .A1(n9816), .A2(P1_U3086), .B1(n14166), .B2(n9740), .C1(
        n9739), .C2(n14163), .ZN(P1_U3350) );
  OAI222_X1 U12273 ( .A1(n9795), .A2(P1_U3086), .B1(n14166), .B2(n9742), .C1(
        n9741), .C2(n14163), .ZN(P1_U3353) );
  INV_X1 U12274 ( .A(n9943), .ZN(n9744) );
  INV_X1 U12275 ( .A(n9743), .ZN(n9745) );
  NAND2_X1 U12276 ( .A1(n9745), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11934) );
  NAND2_X1 U12277 ( .A1(n9744), .A2(n11934), .ZN(n9789) );
  OR2_X1 U12278 ( .A1(n11872), .A2(n9745), .ZN(n9747) );
  AND2_X1 U12279 ( .A1(n9747), .A2(n9746), .ZN(n9788) );
  INV_X1 U12280 ( .A(n9788), .ZN(n9748) );
  AND2_X1 U12281 ( .A1(n9789), .A2(n9748), .ZN(n14570) );
  NOR2_X1 U12282 ( .A1(n14570), .A2(n13728), .ZN(P1_U3085) );
  INV_X1 U12283 ( .A(n13778), .ZN(n13772) );
  INV_X1 U12284 ( .A(n9749), .ZN(n9751) );
  OAI222_X1 U12285 ( .A1(n13772), .A2(P1_U3086), .B1(n14166), .B2(n9751), .C1(
        n9750), .C2(n14163), .ZN(P1_U3349) );
  INV_X1 U12286 ( .A(n9883), .ZN(n9928) );
  OAI222_X1 U12287 ( .A1(n13550), .A2(n9752), .B1(n13552), .B2(n9751), .C1(
        P2_U3088), .C2(n9928), .ZN(P2_U3321) );
  INV_X1 U12288 ( .A(n12961), .ZN(n11489) );
  OAI222_X1 U12289 ( .A1(P3_U3151), .A2(n12557), .B1(n11489), .B2(n9754), .C1(
        n12191), .C2(n9753), .ZN(P3_U3285) );
  OAI222_X1 U12290 ( .A1(P3_U3151), .A2(n14962), .B1(n11489), .B2(n15213), 
        .C1(n12191), .C2(n9755), .ZN(P3_U3284) );
  INV_X1 U12291 ( .A(n12596), .ZN(n14981) );
  OAI222_X1 U12292 ( .A1(P3_U3151), .A2(n14981), .B1(n11489), .B2(n15176), 
        .C1(n12191), .C2(n9756), .ZN(P3_U3283) );
  INV_X1 U12293 ( .A(n9757), .ZN(n9759) );
  OAI222_X1 U12294 ( .A1(P3_U3151), .A2(n6746), .B1(n12191), .B2(n9759), .C1(
        n9758), .C2(n11489), .ZN(P3_U3295) );
  OAI222_X1 U12295 ( .A1(P1_U3086), .A2(n9856), .B1(n14166), .B2(n9760), .C1(
        n7211), .C2(n14163), .ZN(P1_U3354) );
  INV_X1 U12296 ( .A(n13750), .ZN(n9796) );
  OAI222_X1 U12297 ( .A1(n9796), .A2(P1_U3086), .B1(n14166), .B2(n9762), .C1(
        n9761), .C2(n14163), .ZN(P1_U3352) );
  INV_X1 U12298 ( .A(n10624), .ZN(n10628) );
  OAI222_X1 U12299 ( .A1(P3_U3151), .A2(n10628), .B1(n12967), .B2(n9763), .C1(
        n9176), .C2(n11489), .ZN(P3_U3289) );
  INV_X1 U12300 ( .A(n9818), .ZN(n9835) );
  INV_X1 U12301 ( .A(n9764), .ZN(n9767) );
  OAI222_X1 U12302 ( .A1(n9835), .A2(P1_U3086), .B1(n14166), .B2(n9767), .C1(
        n9765), .C2(n14163), .ZN(P1_U3348) );
  INV_X1 U12303 ( .A(n9971), .ZN(n9766) );
  OAI222_X1 U12304 ( .A1(n13550), .A2(n9768), .B1(n13552), .B2(n9767), .C1(
        P2_U3088), .C2(n9766), .ZN(P2_U3320) );
  INV_X1 U12305 ( .A(SI_5_), .ZN(n9770) );
  OAI222_X1 U12306 ( .A1(P3_U3151), .A2(n14924), .B1(n12968), .B2(n9770), .C1(
        n12967), .C2(n9769), .ZN(P3_U3290) );
  INV_X1 U12307 ( .A(SI_2_), .ZN(n15165) );
  OAI222_X1 U12308 ( .A1(P3_U3151), .A2(n10444), .B1(n12968), .B2(n15165), 
        .C1(n12967), .C2(n9771), .ZN(P3_U3293) );
  INV_X1 U12309 ( .A(SI_4_), .ZN(n9773) );
  OAI222_X1 U12310 ( .A1(P3_U3151), .A2(n14902), .B1(n12968), .B2(n9773), .C1(
        n12967), .C2(n9772), .ZN(P3_U3291) );
  OAI222_X1 U12311 ( .A1(P3_U3151), .A2(n14997), .B1(n11489), .B2(n15175), 
        .C1(n12191), .C2(n9774), .ZN(P3_U3282) );
  INV_X1 U12312 ( .A(n9901), .ZN(n9826) );
  INV_X1 U12313 ( .A(n9775), .ZN(n9777) );
  OAI222_X1 U12314 ( .A1(n9826), .A2(P1_U3086), .B1(n14166), .B2(n9777), .C1(
        n9776), .C2(n14163), .ZN(P1_U3347) );
  INV_X1 U12315 ( .A(n9972), .ZN(n10019) );
  OAI222_X1 U12316 ( .A1(n13550), .A2(n9778), .B1(n13552), .B2(n9777), .C1(
        P2_U3088), .C2(n10019), .ZN(P2_U3319) );
  AND2_X1 U12317 ( .A1(n9968), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12318 ( .A1(n9968), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12319 ( .A1(n9968), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12320 ( .A1(n9968), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12321 ( .A1(n9968), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12322 ( .A1(n9968), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12323 ( .A1(n9968), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12324 ( .A1(n9968), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12325 ( .A1(n9968), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12326 ( .A1(n9968), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12327 ( .A1(n9968), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12328 ( .A1(n9968), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12329 ( .A1(n9968), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12330 ( .A1(n9968), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12331 ( .A1(n9968), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12332 ( .A1(n9968), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  INV_X1 U12333 ( .A(n12578), .ZN(n15017) );
  OAI222_X1 U12334 ( .A1(P3_U3151), .A2(n15017), .B1(n11489), .B2(n15127), 
        .C1(n12191), .C2(n9779), .ZN(P3_U3281) );
  MUX2_X1 U12335 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9805), .S(n9816), .Z(n9787)
         );
  INV_X1 U12336 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10142) );
  MUX2_X1 U12337 ( .A(n10142), .B(P1_REG1_REG_2__SCAN_IN), .S(n9795), .Z(
        n13738) );
  INV_X1 U12338 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14644) );
  MUX2_X1 U12339 ( .A(n14644), .B(P1_REG1_REG_1__SCAN_IN), .S(n9856), .Z(n9847) );
  NAND2_X1 U12340 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9851) );
  INV_X1 U12341 ( .A(n9851), .ZN(n9780) );
  NAND2_X1 U12342 ( .A1(n9847), .A2(n9780), .ZN(n9848) );
  INV_X1 U12343 ( .A(n9856), .ZN(n9794) );
  NAND2_X1 U12344 ( .A1(n9794), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U12345 ( .A1(n9848), .A2(n9781), .ZN(n13737) );
  NAND2_X1 U12346 ( .A1(n13738), .A2(n13737), .ZN(n13736) );
  OR2_X1 U12347 ( .A1(n9795), .A2(n10142), .ZN(n9782) );
  NAND2_X1 U12348 ( .A1(n13736), .A2(n9782), .ZN(n13748) );
  MUX2_X1 U12349 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7518), .S(n13750), .Z(
        n13749) );
  NAND2_X1 U12350 ( .A1(n13748), .A2(n13749), .ZN(n13747) );
  NAND2_X1 U12351 ( .A1(n13750), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9783) );
  NAND2_X1 U12352 ( .A1(n13747), .A2(n9783), .ZN(n13759) );
  MUX2_X1 U12353 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7541), .S(n13762), .Z(
        n13760) );
  NAND2_X1 U12354 ( .A1(n13759), .A2(n13760), .ZN(n13758) );
  NAND2_X1 U12355 ( .A1(n13762), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U12356 ( .A1(n13758), .A2(n9784), .ZN(n9786) );
  OR2_X1 U12357 ( .A1(n9786), .A2(n9787), .ZN(n9807) );
  INV_X1 U12358 ( .A(n9807), .ZN(n9785) );
  AOI21_X1 U12359 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9804) );
  NAND2_X1 U12360 ( .A1(n9789), .A2(n9788), .ZN(n14550) );
  INV_X1 U12361 ( .A(n14157), .ZN(n14546) );
  AND2_X1 U12362 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9791) );
  OR2_X1 U12363 ( .A1(n14550), .A2(n13726), .ZN(n13838) );
  NOR2_X1 U12364 ( .A1(n13838), .A2(n9816), .ZN(n9790) );
  AOI211_X1 U12365 ( .C1(n14570), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9791), .B(
        n9790), .ZN(n9803) );
  NAND2_X1 U12366 ( .A1(n13726), .A2(n14546), .ZN(n9792) );
  OR2_X1 U12367 ( .A1(n14550), .A2(n9792), .ZN(n14579) );
  INV_X1 U12368 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10558) );
  MUX2_X1 U12369 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10558), .S(n9856), .Z(n9845) );
  INV_X1 U12370 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9793) );
  NOR3_X1 U12371 ( .A1(n9845), .A2(n14547), .A3(n9793), .ZN(n9844) );
  AOI21_X1 U12372 ( .B1(n9794), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9844), .ZN(
        n13734) );
  INV_X1 U12373 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U12374 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10424), .S(n9795), .Z(
        n13733) );
  OR2_X1 U12375 ( .A1(n13734), .A2(n13733), .ZN(n13744) );
  INV_X1 U12376 ( .A(n9795), .ZN(n13732) );
  NAND2_X1 U12377 ( .A1(n13732), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13743) );
  MUX2_X1 U12378 ( .A(n7519), .B(P1_REG2_REG_3__SCAN_IN), .S(n13750), .Z(
        n13742) );
  AOI21_X1 U12379 ( .B1(n13744), .B2(n13743), .A(n13742), .ZN(n13767) );
  NOR2_X1 U12380 ( .A1(n9796), .A2(n7519), .ZN(n13761) );
  INV_X1 U12381 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10402) );
  MUX2_X1 U12382 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10402), .S(n13762), .Z(
        n9797) );
  OAI21_X1 U12383 ( .B1(n13767), .B2(n13761), .A(n9797), .ZN(n13765) );
  NAND2_X1 U12384 ( .A1(n13762), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9799) );
  INV_X1 U12385 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U12386 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9815), .S(n9816), .Z(n9798)
         );
  AOI21_X1 U12387 ( .B1(n13765), .B2(n9799), .A(n9798), .ZN(n13784) );
  INV_X1 U12388 ( .A(n13784), .ZN(n9801) );
  NAND3_X1 U12389 ( .A1(n13765), .A2(n9799), .A3(n9798), .ZN(n9800) );
  NAND3_X1 U12390 ( .A1(n14560), .A2(n9801), .A3(n9800), .ZN(n9802) );
  OAI211_X1 U12391 ( .C1(n9804), .C2(n11539), .A(n9803), .B(n9802), .ZN(
        P1_U3248) );
  MUX2_X1 U12392 ( .A(n7624), .B(P1_REG1_REG_8__SCAN_IN), .S(n9901), .Z(n9814)
         );
  NAND2_X1 U12393 ( .A1(n9816), .A2(n9805), .ZN(n9806) );
  AND2_X1 U12394 ( .A1(n9807), .A2(n9806), .ZN(n13776) );
  INV_X1 U12395 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9808) );
  XNOR2_X1 U12396 ( .A(n13778), .B(n9808), .ZN(n13777) );
  NAND2_X1 U12397 ( .A1(n13776), .A2(n13777), .ZN(n13775) );
  NAND2_X1 U12398 ( .A1(n13778), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9809) );
  NAND2_X1 U12399 ( .A1(n13775), .A2(n9809), .ZN(n9838) );
  INV_X1 U12400 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9810) );
  XNOR2_X1 U12401 ( .A(n9818), .B(n9810), .ZN(n9839) );
  NAND2_X1 U12402 ( .A1(n9838), .A2(n9839), .ZN(n9837) );
  NAND2_X1 U12403 ( .A1(n9818), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U12404 ( .A1(n9837), .A2(n9811), .ZN(n9813) );
  OR2_X1 U12405 ( .A1(n9813), .A2(n9814), .ZN(n9903) );
  INV_X1 U12406 ( .A(n9903), .ZN(n9812) );
  AOI21_X1 U12407 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9831) );
  NOR2_X1 U12408 ( .A1(n9816), .A2(n9815), .ZN(n13779) );
  INV_X1 U12409 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10652) );
  MUX2_X1 U12410 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10652), .S(n13778), .Z(
        n9817) );
  OAI21_X1 U12411 ( .B1(n13784), .B2(n13779), .A(n9817), .ZN(n13782) );
  NAND2_X1 U12412 ( .A1(n13778), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9833) );
  INV_X1 U12413 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9819) );
  MUX2_X1 U12414 ( .A(n9819), .B(P1_REG2_REG_7__SCAN_IN), .S(n9818), .Z(n9832)
         );
  AOI21_X1 U12415 ( .B1(n13782), .B2(n9833), .A(n9832), .ZN(n9843) );
  NOR2_X1 U12416 ( .A1(n9835), .A2(n9819), .ZN(n9824) );
  INV_X1 U12417 ( .A(n9824), .ZN(n9822) );
  INV_X1 U12418 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9820) );
  MUX2_X1 U12419 ( .A(n9820), .B(P1_REG2_REG_8__SCAN_IN), .S(n9901), .Z(n9821)
         );
  NAND2_X1 U12420 ( .A1(n9822), .A2(n9821), .ZN(n9825) );
  MUX2_X1 U12421 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9820), .S(n9901), .Z(n9823)
         );
  OAI21_X1 U12422 ( .B1(n9843), .B2(n9824), .A(n9823), .ZN(n9896) );
  OAI211_X1 U12423 ( .C1(n9843), .C2(n9825), .A(n9896), .B(n14560), .ZN(n9830)
         );
  AND2_X1 U12424 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U12425 ( .A1(n13838), .A2(n9826), .ZN(n9827) );
  AOI211_X1 U12426 ( .C1(n14570), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9828), .B(
        n9827), .ZN(n9829) );
  OAI211_X1 U12427 ( .C1(n9831), .C2(n11539), .A(n9830), .B(n9829), .ZN(
        P1_U3251) );
  NAND3_X1 U12428 ( .A1(n13782), .A2(n9833), .A3(n9832), .ZN(n9834) );
  NAND2_X1 U12429 ( .A1(n9834), .A2(n14560), .ZN(n9842) );
  NOR2_X1 U12430 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7620), .ZN(n11060) );
  NOR2_X1 U12431 ( .A1(n13838), .A2(n9835), .ZN(n9836) );
  AOI211_X1 U12432 ( .C1(n14570), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n11060), .B(
        n9836), .ZN(n9841) );
  OAI211_X1 U12433 ( .C1(n9839), .C2(n9838), .A(n14575), .B(n9837), .ZN(n9840)
         );
  OAI211_X1 U12434 ( .C1(n9843), .C2(n9842), .A(n9841), .B(n9840), .ZN(
        P1_U3250) );
  NOR2_X1 U12435 ( .A1(n14547), .A2(n9793), .ZN(n13725) );
  INV_X1 U12436 ( .A(n13725), .ZN(n9846) );
  AOI211_X1 U12437 ( .C1(n9846), .C2(n9845), .A(n9844), .B(n14579), .ZN(n9853)
         );
  INV_X1 U12438 ( .A(n9847), .ZN(n9850) );
  INV_X1 U12439 ( .A(n9848), .ZN(n9849) );
  AOI211_X1 U12440 ( .C1(n9851), .C2(n9850), .A(n9849), .B(n11539), .ZN(n9852)
         );
  NOR2_X1 U12441 ( .A1(n9853), .A2(n9852), .ZN(n9855) );
  AOI22_X1 U12442 ( .A1(n14570), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9854) );
  OAI211_X1 U12443 ( .C1(n9856), .C2(n13838), .A(n9855), .B(n9854), .ZN(
        P1_U3244) );
  INV_X1 U12444 ( .A(n10183), .ZN(n10190) );
  INV_X1 U12445 ( .A(n9857), .ZN(n9859) );
  OAI222_X1 U12446 ( .A1(n10190), .A2(P1_U3086), .B1(n14166), .B2(n9859), .C1(
        n9858), .C2(n14163), .ZN(P1_U3346) );
  INV_X1 U12447 ( .A(n10221), .ZN(n9988) );
  OAI222_X1 U12448 ( .A1(n13550), .A2(n9860), .B1(n13552), .B2(n9859), .C1(
        P2_U3088), .C2(n9988), .ZN(P2_U3318) );
  INV_X1 U12449 ( .A(n10004), .ZN(n9863) );
  INV_X1 U12450 ( .A(n14660), .ZN(n9862) );
  NAND2_X1 U12451 ( .A1(n9862), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9991) );
  MUX2_X1 U12452 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8180), .S(n10004), .Z(n9992) );
  AOI21_X1 U12453 ( .B1(n14665), .B2(n9991), .A(n9992), .ZN(n9994) );
  MUX2_X1 U12454 ( .A(n8194), .B(P2_REG2_REG_3__SCAN_IN), .S(n9880), .Z(n14682) );
  MUX2_X1 U12455 ( .A(n10479), .B(P2_REG2_REG_4__SCAN_IN), .S(n9881), .Z(
        n10095) );
  AOI21_X1 U12456 ( .B1(n9881), .B2(P2_REG2_REG_4__SCAN_IN), .A(n10094), .ZN(
        n10086) );
  MUX2_X1 U12457 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10522), .S(n10093), .Z(
        n10085) );
  NOR2_X1 U12458 ( .A1(n10093), .A2(n10522), .ZN(n9917) );
  MUX2_X1 U12459 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10676), .S(n9883), .Z(n9916) );
  NAND2_X1 U12460 ( .A1(n9883), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9865) );
  MUX2_X1 U12461 ( .A(n8252), .B(P2_REG2_REG_7__SCAN_IN), .S(n9971), .Z(n9864)
         );
  NAND3_X1 U12462 ( .A1(n9919), .A2(n9865), .A3(n9864), .ZN(n9872) );
  INV_X1 U12463 ( .A(n9866), .ZN(n9871) );
  INV_X1 U12464 ( .A(n9867), .ZN(n9869) );
  OAI21_X1 U12465 ( .B1(n9869), .B2(n9958), .A(n9868), .ZN(n9870) );
  NAND2_X1 U12466 ( .A1(n9871), .A2(n9870), .ZN(n9874) );
  NOR2_X1 U12467 ( .A1(n9873), .A2(P2_U3088), .ZN(n13542) );
  NAND2_X1 U12468 ( .A1(n9874), .A2(n13542), .ZN(n9886) );
  NOR2_X2 U12469 ( .A1(n9886), .A2(n13547), .ZN(n14727) );
  NAND2_X1 U12470 ( .A1(n9872), .A2(n14727), .ZN(n9892) );
  AND2_X1 U12471 ( .A1(n9874), .A2(n9873), .ZN(n14659) );
  AND2_X1 U12472 ( .A1(n14659), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14741) );
  INV_X1 U12473 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U12474 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10719) );
  OAI21_X1 U12475 ( .B1(n14752), .B2(n9875), .A(n10719), .ZN(n9876) );
  AOI21_X1 U12476 ( .B1(n9971), .B2(n14741), .A(n9876), .ZN(n9891) );
  MUX2_X1 U12477 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8169), .S(n14660), .Z(
        n14671) );
  NAND2_X1 U12478 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n14663), .ZN(n14670) );
  NOR2_X1 U12479 ( .A1(n14671), .A2(n14670), .ZN(n14669) );
  NOR2_X1 U12480 ( .A1(n14660), .A2(n8169), .ZN(n9997) );
  MUX2_X1 U12481 ( .A(n9877), .B(P2_REG1_REG_2__SCAN_IN), .S(n10004), .Z(n9878) );
  OAI21_X1 U12482 ( .B1(n14669), .B2(n9997), .A(n9878), .ZN(n10000) );
  OAI21_X1 U12483 ( .B1(n9877), .B2(n10004), .A(n10000), .ZN(n14687) );
  MUX2_X1 U12484 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9879), .S(n9880), .Z(n14686) );
  NAND2_X1 U12485 ( .A1(n14687), .A2(n14686), .ZN(n14685) );
  NAND2_X1 U12486 ( .A1(n9880), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10100) );
  MUX2_X1 U12487 ( .A(n8213), .B(P2_REG1_REG_4__SCAN_IN), .S(n9881), .Z(n10099) );
  AOI21_X1 U12488 ( .B1(n14685), .B2(n10100), .A(n10099), .ZN(n10102) );
  AOI21_X1 U12489 ( .B1(n9881), .B2(P2_REG1_REG_4__SCAN_IN), .A(n10102), .ZN(
        n10082) );
  MUX2_X1 U12490 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n8229), .S(n10093), .Z(
        n10081) );
  NOR2_X1 U12491 ( .A1(n10082), .A2(n10081), .ZN(n10080) );
  AOI21_X1 U12492 ( .B1(n9882), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10080), .ZN(
        n9922) );
  MUX2_X1 U12493 ( .A(n8242), .B(P2_REG1_REG_6__SCAN_IN), .S(n9883), .Z(n9921)
         );
  NOR2_X1 U12494 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  NOR2_X1 U12495 ( .A1(n9928), .A2(n8242), .ZN(n9888) );
  MUX2_X1 U12496 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9884), .S(n9971), .Z(n9887)
         );
  OAI21_X1 U12497 ( .B1(n9920), .B2(n9888), .A(n9887), .ZN(n10008) );
  OR3_X1 U12498 ( .A1(n9920), .A2(n9888), .A3(n9887), .ZN(n9889) );
  NAND3_X1 U12499 ( .A1(n10008), .A2(n14743), .A3(n9889), .ZN(n9890) );
  OAI211_X1 U12500 ( .C1(n9969), .C2(n9892), .A(n9891), .B(n9890), .ZN(
        P2_U3221) );
  NAND2_X1 U12501 ( .A1(n9901), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9895) );
  INV_X1 U12502 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9893) );
  MUX2_X1 U12503 ( .A(n9893), .B(P1_REG2_REG_9__SCAN_IN), .S(n10183), .Z(n9894) );
  AOI21_X1 U12504 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n13794) );
  NAND3_X1 U12505 ( .A1(n9896), .A2(n9895), .A3(n9894), .ZN(n9897) );
  NAND2_X1 U12506 ( .A1(n9897), .A2(n14560), .ZN(n9909) );
  NOR2_X1 U12507 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11354), .ZN(n9899) );
  NOR2_X1 U12508 ( .A1(n13838), .A2(n10190), .ZN(n9898) );
  AOI211_X1 U12509 ( .C1(n14570), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9899), .B(
        n9898), .ZN(n9908) );
  MUX2_X1 U12510 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9900), .S(n10183), .Z(n9905) );
  OR2_X1 U12511 ( .A1(n9901), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U12512 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  NAND2_X1 U12513 ( .A1(n9904), .A2(n9905), .ZN(n10185) );
  OAI21_X1 U12514 ( .B1(n9905), .B2(n9904), .A(n10185), .ZN(n9906) );
  NAND2_X1 U12515 ( .A1(n9906), .A2(n14575), .ZN(n9907) );
  OAI211_X1 U12516 ( .C1(n13794), .C2(n9909), .A(n9908), .B(n9907), .ZN(
        P1_U3252) );
  INV_X1 U12517 ( .A(n9910), .ZN(n9913) );
  INV_X1 U12518 ( .A(n10293), .ZN(n10226) );
  OAI222_X1 U12519 ( .A1(n13550), .A2(n9911), .B1(n13552), .B2(n9913), .C1(
        P2_U3088), .C2(n10226), .ZN(P2_U3317) );
  INV_X1 U12520 ( .A(n13788), .ZN(n13796) );
  OAI222_X1 U12521 ( .A1(n13796), .A2(P1_U3086), .B1(n14166), .B2(n9913), .C1(
        n9912), .C2(n14163), .ZN(P1_U3345) );
  OAI222_X1 U12522 ( .A1(P3_U3151), .A2(n12604), .B1(n11489), .B2(n9915), .C1(
        n12191), .C2(n9914), .ZN(P3_U3280) );
  OR3_X1 U12523 ( .A1(n10084), .A2(n9917), .A3(n9916), .ZN(n9918) );
  NAND3_X1 U12524 ( .A1(n9919), .A2(n14727), .A3(n9918), .ZN(n9927) );
  INV_X1 U12525 ( .A(n14752), .ZN(n14724) );
  NAND2_X1 U12526 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10549) );
  AOI211_X1 U12527 ( .C1(n9922), .C2(n9921), .A(n9920), .B(n14668), .ZN(n9923)
         );
  INV_X1 U12528 ( .A(n9923), .ZN(n9924) );
  NAND2_X1 U12529 ( .A1(n10549), .A2(n9924), .ZN(n9925) );
  AOI21_X1 U12530 ( .B1(n14724), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9925), .ZN(
        n9926) );
  OAI211_X1 U12531 ( .C1(n14694), .C2(n9928), .A(n9927), .B(n9926), .ZN(
        P2_U3220) );
  INV_X1 U12532 ( .A(n9930), .ZN(n9929) );
  INV_X1 U12533 ( .A(n9931), .ZN(n9932) );
  INV_X1 U12534 ( .A(n12148), .ZN(n12109) );
  OAI22_X1 U12535 ( .A1(n12109), .A2(n11694), .B1(n9931), .B2(n14547), .ZN(
        n9933) );
  NOR2_X1 U12536 ( .A1(n9935), .A2(n10107), .ZN(n10108) );
  AOI21_X1 U12537 ( .B1(n10107), .B2(n9935), .A(n10108), .ZN(n13724) );
  NAND2_X1 U12538 ( .A1(n10130), .A2(n9936), .ZN(n9941) );
  INV_X1 U12539 ( .A(n9941), .ZN(n9940) );
  NAND2_X1 U12540 ( .A1(n9943), .A2(n11872), .ZN(n9938) );
  NOR2_X1 U12541 ( .A1(n14124), .A2(n9938), .ZN(n9939) );
  AND2_X1 U12542 ( .A1(n13658), .A2(n14008), .ZN(n13681) );
  NAND2_X1 U12543 ( .A1(n9941), .A2(n10127), .ZN(n10343) );
  NAND2_X1 U12544 ( .A1(n10343), .A2(n9942), .ZN(n10239) );
  AOI22_X1 U12545 ( .A1(n13681), .A2(n13722), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10239), .ZN(n9945) );
  AND2_X1 U12546 ( .A1(n10343), .A2(n9943), .ZN(n13580) );
  NAND2_X1 U12547 ( .A1(n14490), .A2(n7408), .ZN(n9944) );
  OAI211_X1 U12548 ( .C1(n13724), .C2(n14467), .A(n9945), .B(n9944), .ZN(
        P1_U3232) );
  NAND2_X1 U12549 ( .A1(n13129), .A2(n13065), .ZN(n10035) );
  NAND3_X1 U12550 ( .A1(n10276), .A2(n9947), .A3(n9946), .ZN(n9949) );
  INV_X1 U12551 ( .A(n9949), .ZN(n9952) );
  OAI211_X1 U12552 ( .C1(n9952), .C2(n9953), .A(n9951), .B(n9950), .ZN(n10206)
         );
  OR2_X1 U12553 ( .A1(n10206), .A2(P2_U3088), .ZN(n10162) );
  NOR2_X1 U12554 ( .A1(n10033), .A2(n11023), .ZN(n10481) );
  NAND2_X1 U12555 ( .A1(n9960), .A2(n10481), .ZN(n9954) );
  AOI22_X1 U12556 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n10162), .B1(n13095), 
        .B2(n8554), .ZN(n9963) );
  NOR2_X1 U12557 ( .A1(n9955), .A2(n12001), .ZN(n9961) );
  NAND2_X1 U12558 ( .A1(n10263), .A2(n8554), .ZN(n9957) );
  NAND2_X1 U12559 ( .A1(n10249), .A2(n9957), .ZN(n10025) );
  AND2_X1 U12560 ( .A1(n14828), .A2(n9958), .ZN(n9959) );
  OAI21_X1 U12561 ( .B1(n9961), .B2(n10025), .A(n13060), .ZN(n9962) );
  OAI211_X1 U12562 ( .C1(n10035), .C2(n13066), .A(n9963), .B(n9962), .ZN(
        P2_U3204) );
  INV_X1 U12563 ( .A(n9964), .ZN(n9966) );
  INV_X1 U12564 ( .A(n13143), .ZN(n13133) );
  OAI222_X1 U12565 ( .A1(n13550), .A2(n9965), .B1(n13552), .B2(n9966), .C1(
        P2_U3088), .C2(n13133), .ZN(P2_U3316) );
  INV_X1 U12566 ( .A(n10324), .ZN(n10198) );
  OAI222_X1 U12567 ( .A1(n14163), .A2(n9967), .B1(n14166), .B2(n9966), .C1(
        P1_U3086), .C2(n10198), .ZN(P1_U3344) );
  AND2_X1 U12568 ( .A1(n9968), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12569 ( .A1(n9968), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12570 ( .A1(n9968), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12571 ( .A1(n9968), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12572 ( .A1(n9968), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12573 ( .A1(n9968), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12574 ( .A1(n9968), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12575 ( .A1(n9968), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12576 ( .A1(n9968), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12577 ( .A1(n9968), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12578 ( .A1(n9968), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12579 ( .A1(n9968), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12580 ( .A1(n9968), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12581 ( .A1(n9968), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AOI21_X1 U12582 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n9971), .A(n9969), .ZN(
        n10013) );
  INV_X1 U12583 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U12584 ( .A(n9970), .B(P2_REG2_REG_8__SCAN_IN), .S(n9972), .Z(n10012) );
  NOR2_X1 U12585 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  INV_X1 U12586 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9982) );
  INV_X1 U12587 ( .A(n14727), .ZN(n14747) );
  NOR3_X1 U12588 ( .A1(n9984), .A2(n9982), .A3(n14747), .ZN(n9974) );
  NAND2_X1 U12589 ( .A1(n9971), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10007) );
  MUX2_X1 U12590 ( .A(n8274), .B(P2_REG1_REG_8__SCAN_IN), .S(n9972), .Z(n10006) );
  AOI21_X1 U12591 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(n10005) );
  AOI21_X1 U12592 ( .B1(n9972), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10005), .ZN(
        n9978) );
  NOR3_X1 U12593 ( .A1(n9978), .A2(n9975), .A3(n14668), .ZN(n9973) );
  NOR3_X1 U12594 ( .A1(n9974), .A2(n14741), .A3(n9973), .ZN(n9989) );
  NAND2_X1 U12595 ( .A1(n9988), .A2(n9975), .ZN(n9977) );
  MUX2_X1 U12596 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9975), .S(n10221), .Z(n9976) );
  NAND2_X1 U12597 ( .A1(n9978), .A2(n9976), .ZN(n10220) );
  OAI21_X1 U12598 ( .B1(n9978), .B2(n9977), .A(n10220), .ZN(n9981) );
  INV_X1 U12599 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U12600 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n9979) );
  OAI21_X1 U12601 ( .B1(n14752), .B2(n14243), .A(n9979), .ZN(n9980) );
  AOI21_X1 U12602 ( .B1(n9981), .B2(n14743), .A(n9980), .ZN(n9987) );
  OR2_X1 U12603 ( .A1(n10221), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10216) );
  MUX2_X1 U12604 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9982), .S(n10221), .Z(n9983) );
  NAND2_X1 U12605 ( .A1(n9984), .A2(n9983), .ZN(n10217) );
  OAI21_X1 U12606 ( .B1(n9984), .B2(n10216), .A(n10217), .ZN(n9985) );
  NAND2_X1 U12607 ( .A1(n9985), .A2(n14727), .ZN(n9986) );
  OAI211_X1 U12608 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(
        P2_U3223) );
  OAI222_X1 U12609 ( .A1(n12968), .A2(n15194), .B1(n12967), .B2(n9990), .C1(
        n12610), .C2(P3_U3151), .ZN(P3_U3279) );
  NOR2_X1 U12610 ( .A1(n10690), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9996) );
  AND3_X1 U12611 ( .A1(n14665), .A2(n9992), .A3(n9991), .ZN(n9993) );
  NOR3_X1 U12612 ( .A1(n14747), .A2(n9994), .A3(n9993), .ZN(n9995) );
  AOI211_X1 U12613 ( .C1(n14724), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9996), .B(
        n9995), .ZN(n10003) );
  MUX2_X1 U12614 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9877), .S(n10004), .Z(n9999) );
  INV_X1 U12615 ( .A(n9997), .ZN(n9998) );
  NAND2_X1 U12616 ( .A1(n9999), .A2(n9998), .ZN(n10001) );
  OAI211_X1 U12617 ( .C1(n14669), .C2(n10001), .A(n14743), .B(n10000), .ZN(
        n10002) );
  OAI211_X1 U12618 ( .C1(n14694), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        P2_U3216) );
  INV_X1 U12619 ( .A(n10005), .ZN(n10010) );
  NAND3_X1 U12620 ( .A1(n10008), .A2(n10007), .A3(n10006), .ZN(n10009) );
  NAND3_X1 U12621 ( .A1(n10010), .A2(n14743), .A3(n10009), .ZN(n10018) );
  NAND2_X1 U12622 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10927) );
  AOI211_X1 U12623 ( .C1(n10013), .C2(n10012), .A(n10011), .B(n14747), .ZN(
        n10014) );
  INV_X1 U12624 ( .A(n10014), .ZN(n10015) );
  NAND2_X1 U12625 ( .A1(n10927), .A2(n10015), .ZN(n10016) );
  AOI21_X1 U12626 ( .B1(n14724), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10016), .ZN(
        n10017) );
  OAI211_X1 U12627 ( .C1(n14694), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        P2_U3222) );
  INV_X1 U12628 ( .A(n10020), .ZN(n10038) );
  INV_X1 U12629 ( .A(n14163), .ZN(n14149) );
  AOI22_X1 U12630 ( .A1(n14562), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14149), .ZN(n10021) );
  OAI21_X1 U12631 ( .B1(n10038), .B2(n14166), .A(n10021), .ZN(P1_U3343) );
  INV_X1 U12632 ( .A(n13095), .ZN(n13071) );
  NAND2_X1 U12633 ( .A1(n13129), .A2(n9956), .ZN(n10154) );
  INV_X1 U12634 ( .A(n10025), .ZN(n10026) );
  NAND2_X1 U12635 ( .A1(n10026), .A2(n6588), .ZN(n10027) );
  OAI21_X1 U12636 ( .B1(n10028), .B2(n10027), .A(n10157), .ZN(n10029) );
  NAND2_X1 U12637 ( .A1(n10029), .A2(n13060), .ZN(n10032) );
  AOI22_X1 U12638 ( .A1(n13064), .A2(n13131), .B1(n13128), .B2(n13065), .ZN(
        n10250) );
  INV_X1 U12639 ( .A(n10250), .ZN(n10030) );
  AOI22_X1 U12640 ( .A1(n10162), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n13085), 
        .B2(n10030), .ZN(n10031) );
  OAI211_X1 U12641 ( .C1(n10683), .C2(n13071), .A(n10032), .B(n10031), .ZN(
        P2_U3194) );
  INV_X1 U12642 ( .A(n14805), .ZN(n14835) );
  NOR2_X1 U12643 ( .A1(n10034), .A2(n10033), .ZN(n10281) );
  INV_X1 U12644 ( .A(n10023), .ZN(n14810) );
  OAI21_X1 U12645 ( .B1(n14810), .B2(n14399), .A(n10285), .ZN(n10036) );
  NAND2_X1 U12646 ( .A1(n10036), .A2(n10035), .ZN(n10279) );
  AOI211_X1 U12647 ( .C1(n14835), .C2(n10285), .A(n10281), .B(n10279), .ZN(
        n14793) );
  NAND2_X1 U12648 ( .A1(n8665), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10037) );
  OAI21_X1 U12649 ( .B1(n14793), .B2(n8665), .A(n10037), .ZN(P2_U3499) );
  INV_X1 U12650 ( .A(n13144), .ZN(n13167) );
  OAI222_X1 U12651 ( .A1(n13550), .A2(n10039), .B1(n13552), .B2(n10038), .C1(
        n13167), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U12652 ( .A1(n12504), .A2(n10040), .ZN(n10041) );
  NAND2_X1 U12653 ( .A1(n9102), .A2(n10041), .ZN(n10073) );
  INV_X1 U12654 ( .A(n10073), .ZN(n10044) );
  INV_X1 U12655 ( .A(n12531), .ZN(n10042) );
  OR2_X1 U12656 ( .A1(n10043), .A2(n10042), .ZN(n10072) );
  INV_X1 U12657 ( .A(n10066), .ZN(n10045) );
  INV_X2 U12658 ( .A(P3_U3897), .ZN(n12554) );
  MUX2_X1 U12659 ( .A(n10045), .B(n12554), .S(n12527), .Z(n15018) );
  INV_X1 U12660 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10046) );
  INV_X1 U12661 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10168) );
  INV_X1 U12662 ( .A(n10182), .ZN(n10047) );
  INV_X1 U12663 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10059) );
  INV_X1 U12664 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U12665 ( .A(n10059), .B(n10048), .S(n9533), .Z(n14869) );
  NAND2_X1 U12666 ( .A1(n14869), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14868) );
  NOR2_X1 U12667 ( .A1(n10176), .A2(n14868), .ZN(n10175) );
  INV_X1 U12668 ( .A(n10049), .ZN(n10054) );
  INV_X1 U12669 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10909) );
  INV_X1 U12670 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U12671 ( .A(n10909), .B(n10067), .S(n9533), .Z(n10050) );
  INV_X1 U12672 ( .A(n10444), .ZN(n10455) );
  NAND2_X1 U12673 ( .A1(n10050), .A2(n10455), .ZN(n14881) );
  INV_X1 U12674 ( .A(n10050), .ZN(n10051) );
  NAND2_X1 U12675 ( .A1(n10051), .A2(n10444), .ZN(n10052) );
  AND2_X1 U12676 ( .A1(n14881), .A2(n10052), .ZN(n10053) );
  INV_X1 U12677 ( .A(n14882), .ZN(n10056) );
  NOR3_X1 U12678 ( .A1(n10175), .A2(n10054), .A3(n10053), .ZN(n10055) );
  NAND2_X1 U12679 ( .A1(P3_U3897), .A2(n11956), .ZN(n15003) );
  OAI21_X1 U12680 ( .B1(n10056), .B2(n10055), .A(n15022), .ZN(n10078) );
  INV_X1 U12681 ( .A(n10057), .ZN(n10058) );
  MUX2_X1 U12682 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n10909), .S(n10444), .Z(
        n10064) );
  NOR2_X1 U12683 ( .A1(n10059), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U12684 ( .A1(n10060), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U12685 ( .A1(n10167), .A2(n10062), .ZN(n10063) );
  OAI21_X1 U12686 ( .B1(n10064), .B2(n10063), .A(n10446), .ZN(n10065) );
  NAND2_X1 U12687 ( .A1(n14355), .A2(n10065), .ZN(n10076) );
  MUX2_X1 U12688 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10067), .S(n10444), .Z(
        n10070) );
  AND2_X1 U12689 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n6746), .ZN(n10068) );
  OAI21_X1 U12690 ( .B1(n10182), .B2(n10068), .A(n7435), .ZN(n10169) );
  OR2_X1 U12691 ( .A1(n10169), .A2(n10168), .ZN(n10171) );
  NAND2_X1 U12692 ( .A1(n10171), .A2(n7435), .ZN(n10069) );
  NAND2_X1 U12693 ( .A1(n10070), .A2(n10069), .ZN(n10454) );
  OAI21_X1 U12694 ( .B1(n10070), .B2(n10069), .A(n10454), .ZN(n10071) );
  NAND2_X1 U12695 ( .A1(n15014), .A2(n10071), .ZN(n10075) );
  AOI22_X1 U12696 ( .A1(n15021), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10074) );
  AND3_X1 U12697 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(n10077) );
  OAI211_X1 U12698 ( .C1(n15018), .C2(n10444), .A(n10078), .B(n10077), .ZN(
        P3_U3184) );
  INV_X1 U12699 ( .A(SI_17_), .ZN(n15253) );
  OAI222_X1 U12700 ( .A1(P3_U3151), .A2(n12612), .B1(n11489), .B2(n15253), 
        .C1(n12191), .C2(n10079), .ZN(P3_U3278) );
  AOI211_X1 U12701 ( .C1(n10082), .C2(n10081), .A(n10080), .B(n14668), .ZN(
        n10083) );
  INV_X1 U12702 ( .A(n10083), .ZN(n10089) );
  AOI211_X1 U12703 ( .C1(n10086), .C2(n10085), .A(n10084), .B(n14747), .ZN(
        n10087) );
  INV_X1 U12704 ( .A(n10087), .ZN(n10088) );
  NAND2_X1 U12705 ( .A1(n10089), .A2(n10088), .ZN(n10091) );
  NAND2_X1 U12706 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10507) );
  INV_X1 U12707 ( .A(n10507), .ZN(n10090) );
  AOI211_X1 U12708 ( .C1(n14724), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10091), .B(
        n10090), .ZN(n10092) );
  OAI21_X1 U12709 ( .B1(n14694), .B2(n10093), .A(n10092), .ZN(P2_U3219) );
  NAND2_X1 U12710 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10378) );
  AOI211_X1 U12711 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n14747), .ZN(
        n10097) );
  INV_X1 U12712 ( .A(n10097), .ZN(n10098) );
  NAND2_X1 U12713 ( .A1(n10378), .A2(n10098), .ZN(n10104) );
  AND3_X1 U12714 ( .A1(n14685), .A2(n10100), .A3(n10099), .ZN(n10101) );
  NOR3_X1 U12715 ( .A1(n14668), .A2(n10102), .A3(n10101), .ZN(n10103) );
  AOI211_X1 U12716 ( .C1(n14724), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10104), .B(
        n10103), .ZN(n10105) );
  OAI21_X1 U12717 ( .B1(n10106), .B2(n14694), .A(n10105), .ZN(P2_U3218) );
  NAND2_X1 U12718 ( .A1(n13722), .A2(n12148), .ZN(n10110) );
  NAND2_X1 U12719 ( .A1(n11700), .A2(n12147), .ZN(n10109) );
  NAND2_X1 U12720 ( .A1(n10110), .A2(n10109), .ZN(n10111) );
  XNOR2_X1 U12721 ( .A(n10111), .B(n12129), .ZN(n10114) );
  NAND2_X1 U12722 ( .A1(n10114), .A2(n10113), .ZN(n10234) );
  INV_X1 U12723 ( .A(n10235), .ZN(n10116) );
  AOI21_X1 U12724 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10122) );
  AND2_X1 U12725 ( .A1(n13658), .A2(n14006), .ZN(n13673) );
  AOI22_X1 U12726 ( .A1(n13681), .A2(n13721), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10239), .ZN(n10119) );
  OAI21_X1 U12727 ( .B1(n10565), .B2(n14477), .A(n10119), .ZN(n10120) );
  AOI21_X1 U12728 ( .B1(n14490), .B2(n11700), .A(n10120), .ZN(n10121) );
  OAI21_X1 U12729 ( .B1(n10122), .B2(n14467), .A(n10121), .ZN(P1_U3222) );
  OAI21_X1 U12730 ( .B1(n10125), .B2(P1_D_REG_1__SCAN_IN), .A(n10123), .ZN(
        n10128) );
  OR2_X1 U12731 ( .A1(n10125), .A2(n10124), .ZN(n10126) );
  NAND3_X1 U12732 ( .A1(n10128), .A2(n10127), .A3(n10126), .ZN(n10129) );
  NOR2_X1 U12733 ( .A1(n10129), .A2(n11931), .ZN(n10144) );
  OAI21_X1 U12734 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(n10429) );
  INV_X1 U12735 ( .A(n10429), .ZN(n10140) );
  OR2_X1 U12736 ( .A1(n13843), .A2(n11871), .ZN(n14130) );
  XNOR2_X1 U12737 ( .A(n10135), .B(n11891), .ZN(n10136) );
  OAI22_X1 U12738 ( .A1(n14046), .A2(n14021), .B1(n10579), .B2(n14045), .ZN(
        n10240) );
  AOI21_X1 U12739 ( .B1(n10136), .B2(n14028), .A(n10240), .ZN(n10432) );
  NAND2_X1 U12740 ( .A1(n10560), .A2(n7516), .ZN(n10137) );
  NAND2_X1 U12741 ( .A1(n10137), .A2(n14126), .ZN(n10138) );
  NOR2_X1 U12742 ( .A1(n10353), .A2(n10138), .ZN(n10428) );
  AOI21_X1 U12743 ( .B1(n7516), .B2(n14124), .A(n10428), .ZN(n10139) );
  OAI211_X1 U12744 ( .C1(n10140), .C2(n14583), .A(n10432), .B(n10139), .ZN(
        n10145) );
  NAND2_X1 U12745 ( .A1(n10145), .A2(n14654), .ZN(n10141) );
  OAI21_X1 U12746 ( .B1(n14654), .B2(n10142), .A(n10141), .ZN(P1_U3530) );
  INV_X1 U12747 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10147) );
  NAND2_X1 U12748 ( .A1(n10145), .A2(n14641), .ZN(n10146) );
  OAI21_X1 U12749 ( .B1(n14641), .B2(n10147), .A(n10146), .ZN(P1_U3465) );
  NAND2_X1 U12750 ( .A1(n13128), .A2(n9956), .ZN(n10149) );
  NAND2_X1 U12751 ( .A1(n10148), .A2(n10149), .ZN(n10204) );
  INV_X1 U12752 ( .A(n10148), .ZN(n10151) );
  INV_X1 U12753 ( .A(n10149), .ZN(n10150) );
  NAND2_X1 U12754 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  AND2_X1 U12755 ( .A1(n10204), .A2(n10152), .ZN(n10159) );
  INV_X1 U12756 ( .A(n10153), .ZN(n10155) );
  NAND2_X1 U12757 ( .A1(n10155), .A2(n10154), .ZN(n10156) );
  OAI21_X1 U12758 ( .B1(n10159), .B2(n10158), .A(n10205), .ZN(n10160) );
  NAND2_X1 U12759 ( .A1(n10160), .A2(n13060), .ZN(n10164) );
  AOI22_X1 U12760 ( .A1(n13064), .A2(n13129), .B1(n13127), .B2(n13065), .ZN(
        n10268) );
  INV_X1 U12761 ( .A(n10268), .ZN(n10161) );
  AOI22_X1 U12762 ( .A1(n10162), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n13085), 
        .B2(n10161), .ZN(n10163) );
  OAI211_X1 U12763 ( .C1(n10689), .C2(n13071), .A(n10164), .B(n10163), .ZN(
        P2_U3209) );
  NAND2_X1 U12764 ( .A1(n10165), .A2(n10046), .ZN(n10166) );
  NAND2_X1 U12765 ( .A1(n10167), .A2(n10166), .ZN(n10180) );
  INV_X1 U12766 ( .A(n15021), .ZN(n14953) );
  NAND2_X1 U12767 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  NAND2_X1 U12768 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  NAND2_X1 U12769 ( .A1(n15014), .A2(n10172), .ZN(n10174) );
  NAND2_X1 U12770 ( .A1(P3_U3151), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n10173) );
  OAI211_X1 U12771 ( .C1(n14173), .C2(n14953), .A(n10174), .B(n10173), .ZN(
        n10179) );
  AOI21_X1 U12772 ( .B1(n14868), .B2(n10176), .A(n10175), .ZN(n10177) );
  NOR2_X1 U12773 ( .A1(n10177), .A2(n15003), .ZN(n10178) );
  AOI211_X1 U12774 ( .C1(n14355), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10181) );
  OAI21_X1 U12775 ( .B1(n10182), .B2(n15018), .A(n10181), .ZN(P3_U3183) );
  MUX2_X1 U12776 ( .A(n7682), .B(P1_REG1_REG_11__SCAN_IN), .S(n10324), .Z(
        n10189) );
  OR2_X1 U12777 ( .A1(n10183), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10184) );
  AND2_X1 U12778 ( .A1(n10185), .A2(n10184), .ZN(n13801) );
  INV_X1 U12779 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14652) );
  MUX2_X1 U12780 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n14652), .S(n13788), .Z(
        n13800) );
  NAND2_X1 U12781 ( .A1(n13801), .A2(n13800), .ZN(n13799) );
  NAND2_X1 U12782 ( .A1(n13788), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U12783 ( .A1(n13799), .A2(n10186), .ZN(n10188) );
  INV_X1 U12784 ( .A(n14554), .ZN(n10187) );
  AOI21_X1 U12785 ( .B1(n10189), .B2(n10188), .A(n10187), .ZN(n10203) );
  NOR2_X1 U12786 ( .A1(n10190), .A2(n9893), .ZN(n13789) );
  INV_X1 U12787 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10191) );
  MUX2_X1 U12788 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10191), .S(n13788), .Z(
        n10192) );
  OAI21_X1 U12789 ( .B1(n13794), .B2(n13789), .A(n10192), .ZN(n13792) );
  NAND2_X1 U12790 ( .A1(n13788), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10195) );
  INV_X1 U12791 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10193) );
  MUX2_X1 U12792 ( .A(n10193), .B(P1_REG2_REG_11__SCAN_IN), .S(n10324), .Z(
        n10194) );
  AOI21_X1 U12793 ( .B1(n13792), .B2(n10195), .A(n10194), .ZN(n10316) );
  INV_X1 U12794 ( .A(n10316), .ZN(n10197) );
  NAND3_X1 U12795 ( .A1(n13792), .A2(n10195), .A3(n10194), .ZN(n10196) );
  NAND3_X1 U12796 ( .A1(n10197), .A2(n14560), .A3(n10196), .ZN(n10202) );
  NAND2_X1 U12797 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14491)
         );
  INV_X1 U12798 ( .A(n14491), .ZN(n10200) );
  NOR2_X1 U12799 ( .A1(n13838), .A2(n10198), .ZN(n10199) );
  AOI211_X1 U12800 ( .C1(n14570), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10200), 
        .B(n10199), .ZN(n10201) );
  OAI211_X1 U12801 ( .C1(n10203), .C2(n11539), .A(n10202), .B(n10201), .ZN(
        P1_U3254) );
  XNOR2_X1 U12802 ( .A(n12009), .B(n10305), .ZN(n10366) );
  XNOR2_X1 U12803 ( .A(n10365), .B(n10366), .ZN(n10368) );
  XNOR2_X1 U12804 ( .A(n10369), .B(n10368), .ZN(n10211) );
  INV_X1 U12805 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U12806 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10208), .ZN(n14677) );
  AOI22_X1 U12807 ( .A1(n13064), .A2(n13128), .B1(n13126), .B2(n13065), .ZN(
        n10308) );
  NOR2_X1 U12808 ( .A1(n13066), .A2(n10308), .ZN(n10207) );
  AOI211_X1 U12809 ( .C1(n13068), .C2(n10208), .A(n14677), .B(n10207), .ZN(
        n10210) );
  NAND2_X1 U12810 ( .A1(n13095), .A2(n10305), .ZN(n10209) );
  OAI211_X1 U12811 ( .C1(n10211), .C2(n13091), .A(n10210), .B(n10209), .ZN(
        P2_U3190) );
  INV_X1 U12812 ( .A(n10587), .ZN(n10594) );
  INV_X1 U12813 ( .A(n10212), .ZN(n10215) );
  OAI222_X1 U12814 ( .A1(P1_U3086), .A2(n10594), .B1(n14166), .B2(n10215), 
        .C1(n10213), .C2(n14163), .ZN(P1_U3342) );
  OAI222_X1 U12815 ( .A1(P2_U3088), .A2(n14693), .B1(n13559), .B2(n10215), 
        .C1(n10214), .C2(n13550), .ZN(P2_U3314) );
  NAND2_X1 U12816 ( .A1(n10217), .A2(n10216), .ZN(n10219) );
  MUX2_X1 U12817 ( .A(n11016), .B(P2_REG2_REG_10__SCAN_IN), .S(n10293), .Z(
        n10218) );
  NOR2_X1 U12818 ( .A1(n10219), .A2(n10218), .ZN(n10292) );
  AOI211_X1 U12819 ( .C1(n10219), .C2(n10218), .A(n14747), .B(n10292), .ZN(
        n10229) );
  OAI21_X1 U12820 ( .B1(n10221), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10220), .ZN(
        n10224) );
  MUX2_X1 U12821 ( .A(n8302), .B(P2_REG1_REG_10__SCAN_IN), .S(n10293), .Z(
        n10223) );
  INV_X1 U12822 ( .A(n10290), .ZN(n10222) );
  AOI211_X1 U12823 ( .C1(n10224), .C2(n10223), .A(n14668), .B(n10222), .ZN(
        n10228) );
  NAND2_X1 U12824 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11145)
         );
  NAND2_X1 U12825 ( .A1(n14724), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10225) );
  OAI211_X1 U12826 ( .C1(n14694), .C2(n10226), .A(n11145), .B(n10225), .ZN(
        n10227) );
  OR3_X1 U12827 ( .A1(n10229), .A2(n10228), .A3(n10227), .ZN(P2_U3224) );
  NAND2_X1 U12828 ( .A1(n13721), .A2(n12148), .ZN(n10231) );
  NAND2_X1 U12829 ( .A1(n7516), .A2(n12147), .ZN(n10230) );
  NAND2_X1 U12830 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  XNOR2_X1 U12831 ( .A(n10232), .B(n12158), .ZN(n10336) );
  OAI22_X1 U12832 ( .A1(n10566), .A2(n10334), .B1(n10425), .B2(n12062), .ZN(
        n10335) );
  NAND2_X1 U12833 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  OAI21_X1 U12834 ( .B1(n10237), .B2(n10236), .A(n10339), .ZN(n10238) );
  NAND2_X1 U12835 ( .A1(n10238), .A2(n14483), .ZN(n10242) );
  AOI22_X1 U12836 ( .A1(n10240), .A2(n13658), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10239), .ZN(n10241) );
  OAI211_X1 U12837 ( .C1(n10425), .C2(n13699), .A(n10242), .B(n10241), .ZN(
        P1_U3237) );
  OAI21_X1 U12838 ( .B1(n10248), .B2(n10244), .A(n10243), .ZN(n10685) );
  INV_X1 U12839 ( .A(n10264), .ZN(n10245) );
  AOI211_X1 U12840 ( .C1(n8554), .C2(n10246), .A(n13295), .B(n10245), .ZN(
        n10680) );
  XOR2_X1 U12841 ( .A(n10249), .B(n10248), .Z(n10251) );
  OAI21_X1 U12842 ( .B1(n10251), .B2(n13393), .A(n10250), .ZN(n10679) );
  AOI211_X1 U12843 ( .C1(n14816), .C2(n10685), .A(n10680), .B(n10679), .ZN(
        n10257) );
  INV_X1 U12844 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10252) );
  OAI22_X1 U12845 ( .A1(n13531), .A2(n10683), .B1(n14836), .B2(n10252), .ZN(
        n10253) );
  INV_X1 U12846 ( .A(n10253), .ZN(n10254) );
  OAI21_X1 U12847 ( .B1(n10257), .B2(n7143), .A(n10254), .ZN(P2_U3433) );
  OAI22_X1 U12848 ( .A1(n13474), .A2(n10683), .B1(n14842), .B2(n8169), .ZN(
        n10255) );
  INV_X1 U12849 ( .A(n10255), .ZN(n10256) );
  OAI21_X1 U12850 ( .B1(n10257), .B2(n8665), .A(n10256), .ZN(P2_U3500) );
  INV_X1 U12851 ( .A(n10258), .ZN(n10260) );
  OAI222_X1 U12852 ( .A1(n12614), .A2(P3_U3151), .B1(n12967), .B2(n10260), 
        .C1(n10259), .C2(n11489), .ZN(P3_U3277) );
  OAI21_X1 U12853 ( .B1(n10262), .B2(n10266), .A(n10261), .ZN(n10694) );
  AOI211_X1 U12854 ( .C1(n10265), .C2(n10264), .A(n14410), .B(n10303), .ZN(
        n10693) );
  XNOR2_X1 U12855 ( .A(n10266), .B(n10267), .ZN(n10269) );
  OAI21_X1 U12856 ( .B1(n10269), .B2(n13393), .A(n10268), .ZN(n10688) );
  AOI211_X1 U12857 ( .C1(n14816), .C2(n10694), .A(n10693), .B(n10688), .ZN(
        n10275) );
  INV_X1 U12858 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10270) );
  OAI22_X1 U12859 ( .A1(n13531), .A2(n10689), .B1(n14836), .B2(n10270), .ZN(
        n10271) );
  INV_X1 U12860 ( .A(n10271), .ZN(n10272) );
  OAI21_X1 U12861 ( .B1(n10275), .B2(n7143), .A(n10272), .ZN(P2_U3436) );
  OAI22_X1 U12862 ( .A1(n13474), .A2(n10689), .B1(n14842), .B2(n9877), .ZN(
        n10273) );
  INV_X1 U12863 ( .A(n10273), .ZN(n10274) );
  OAI21_X1 U12864 ( .B1(n10275), .B2(n8665), .A(n10274), .ZN(P2_U3501) );
  NAND2_X1 U12865 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  AOI21_X1 U12866 ( .B1(n10281), .B2(n10280), .A(n10279), .ZN(n10287) );
  NAND2_X1 U12867 ( .A1(n8670), .A2(n10282), .ZN(n10475) );
  OR2_X1 U12868 ( .A1(n14420), .A2(n10475), .ZN(n13389) );
  INV_X1 U12869 ( .A(n13389), .ZN(n11226) );
  OAI22_X1 U12870 ( .A1(n13336), .A2(n8158), .B1(n10283), .B2(n13300), .ZN(
        n10284) );
  AOI21_X1 U12871 ( .B1(n11226), .B2(n10285), .A(n10284), .ZN(n10286) );
  OAI21_X1 U12872 ( .B1(n13411), .B2(n10287), .A(n10286), .ZN(P2_U3265) );
  NAND2_X1 U12873 ( .A1(n10293), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10289) );
  MUX2_X1 U12874 ( .A(n8316), .B(P2_REG1_REG_11__SCAN_IN), .S(n13143), .Z(
        n10288) );
  AOI21_X1 U12875 ( .B1(n10290), .B2(n10289), .A(n10288), .ZN(n13142) );
  NAND3_X1 U12876 ( .A1(n10290), .A2(n10289), .A3(n10288), .ZN(n10291) );
  NAND2_X1 U12877 ( .A1(n10291), .A2(n14743), .ZN(n10300) );
  INV_X1 U12878 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13132) );
  MUX2_X1 U12879 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13132), .S(n13143), .Z(
        n10294) );
  NAND2_X1 U12880 ( .A1(n10295), .A2(n10294), .ZN(n13137) );
  OAI21_X1 U12881 ( .B1(n10295), .B2(n10294), .A(n13137), .ZN(n10296) );
  NAND2_X1 U12882 ( .A1(n10296), .A2(n14727), .ZN(n10299) );
  AND2_X1 U12883 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11269) );
  NOR2_X1 U12884 ( .A1(n14694), .A2(n13133), .ZN(n10297) );
  AOI211_X1 U12885 ( .C1(n14724), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11269), 
        .B(n10297), .ZN(n10298) );
  OAI211_X1 U12886 ( .C1(n13142), .C2(n10300), .A(n10299), .B(n10298), .ZN(
        P2_U3225) );
  OAI21_X1 U12887 ( .B1(n10302), .B2(n10306), .A(n10301), .ZN(n10489) );
  INV_X1 U12888 ( .A(n10303), .ZN(n10304) );
  AOI211_X1 U12889 ( .C1(n10305), .C2(n10304), .A(n13295), .B(n6932), .ZN(
        n10492) );
  XNOR2_X1 U12890 ( .A(n10306), .B(n10307), .ZN(n10309) );
  OAI21_X1 U12891 ( .B1(n10309), .B2(n13393), .A(n10308), .ZN(n10493) );
  AOI211_X1 U12892 ( .C1(n14816), .C2(n10489), .A(n10492), .B(n10493), .ZN(
        n10315) );
  INV_X1 U12893 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10310) );
  OAI22_X1 U12894 ( .A1(n13531), .A2(n8204), .B1(n14836), .B2(n10310), .ZN(
        n10311) );
  INV_X1 U12895 ( .A(n10311), .ZN(n10312) );
  OAI21_X1 U12896 ( .B1(n10315), .B2(n7143), .A(n10312), .ZN(P2_U3439) );
  OAI22_X1 U12897 ( .A1(n13474), .A2(n8204), .B1(n14842), .B2(n9879), .ZN(
        n10313) );
  INV_X1 U12898 ( .A(n10313), .ZN(n10314) );
  OAI21_X1 U12899 ( .B1(n10315), .B2(n8665), .A(n10314), .ZN(P2_U3502) );
  AOI21_X1 U12900 ( .B1(n10324), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10316), 
        .ZN(n14559) );
  INV_X1 U12901 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U12902 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10317), .S(n14562), .Z(
        n14558) );
  NAND2_X1 U12903 ( .A1(n14559), .A2(n14558), .ZN(n14557) );
  OAI21_X1 U12904 ( .B1(n14562), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14557), 
        .ZN(n10319) );
  INV_X1 U12905 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10593) );
  MUX2_X1 U12906 ( .A(n10593), .B(P1_REG2_REG_13__SCAN_IN), .S(n10587), .Z(
        n10318) );
  NOR2_X1 U12907 ( .A1(n10319), .A2(n10318), .ZN(n10600) );
  AOI211_X1 U12908 ( .C1(n10319), .C2(n10318), .A(n14579), .B(n10600), .ZN(
        n10323) );
  NOR2_X1 U12909 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13649), .ZN(n10320) );
  AOI21_X1 U12910 ( .B1(n14570), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10320), 
        .ZN(n10321) );
  OAI21_X1 U12911 ( .B1(n13838), .B2(n10594), .A(n10321), .ZN(n10322) );
  NOR2_X1 U12912 ( .A1(n10323), .A2(n10322), .ZN(n10332) );
  OR2_X1 U12913 ( .A1(n10324), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n14553) );
  NAND2_X1 U12914 ( .A1(n14554), .A2(n14553), .ZN(n10327) );
  INV_X1 U12915 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10325) );
  MUX2_X1 U12916 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10325), .S(n14562), .Z(
        n10326) );
  NAND2_X1 U12917 ( .A1(n10327), .A2(n10326), .ZN(n14556) );
  OR2_X1 U12918 ( .A1(n14562), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10328) );
  INV_X1 U12919 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11484) );
  MUX2_X1 U12920 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11484), .S(n10587), .Z(
        n10329) );
  NAND2_X1 U12921 ( .A1(n10330), .A2(n10329), .ZN(n10589) );
  OAI211_X1 U12922 ( .C1(n10330), .C2(n10329), .A(n10589), .B(n14575), .ZN(
        n10331) );
  NAND2_X1 U12923 ( .A1(n10332), .A2(n10331), .ZN(P1_U3256) );
  OR2_X1 U12924 ( .A1(n10354), .A2(n12161), .ZN(n10333) );
  OAI22_X1 U12925 ( .A1(n10579), .A2(n10334), .B1(n10354), .B2(n12062), .ZN(
        n10575) );
  AOI211_X1 U12926 ( .C1(n10341), .C2(n10340), .A(n14467), .B(n10573), .ZN(
        n10349) );
  NAND3_X1 U12927 ( .A1(n10343), .A2(n10342), .A3(n9931), .ZN(n10344) );
  NAND2_X1 U12928 ( .A1(n10344), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10345) );
  MUX2_X1 U12929 ( .A(n14494), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n10347) );
  AOI22_X1 U12930 ( .A1(n13673), .A2(n13721), .B1(n13681), .B2(n13720), .ZN(
        n10346) );
  OAI211_X1 U12931 ( .C1(n10354), .C2(n13699), .A(n10347), .B(n10346), .ZN(
        n10348) );
  OR2_X1 U12932 ( .A1(n10349), .A2(n10348), .ZN(P1_U3218) );
  INV_X1 U12933 ( .A(n14130), .ZN(n14618) );
  OR2_X1 U12934 ( .A1(n10350), .A2(n10356), .ZN(n10351) );
  NAND2_X1 U12935 ( .A1(n10352), .A2(n10351), .ZN(n10704) );
  OAI211_X1 U12936 ( .C1(n10353), .C2(n10354), .A(n10394), .B(n14126), .ZN(
        n10700) );
  OAI21_X1 U12937 ( .B1(n10354), .B2(n14634), .A(n10700), .ZN(n10360) );
  INV_X1 U12938 ( .A(n14028), .ZN(n14584) );
  XNOR2_X1 U12939 ( .A(n10355), .B(n10356), .ZN(n10359) );
  INV_X1 U12940 ( .A(n14025), .ZN(n13924) );
  NAND2_X1 U12941 ( .A1(n10704), .A2(n13924), .ZN(n10358) );
  AOI22_X1 U12942 ( .A1(n13720), .A2(n14008), .B1(n14006), .B2(n13721), .ZN(
        n10357) );
  OAI211_X1 U12943 ( .C1(n14584), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10701) );
  AOI211_X1 U12944 ( .C1(n14618), .C2(n10704), .A(n10360), .B(n10701), .ZN(
        n10362) );
  OR2_X1 U12945 ( .A1(n10362), .A2(n14651), .ZN(n10361) );
  OAI21_X1 U12946 ( .B1(n14654), .B2(n7518), .A(n10361), .ZN(P1_U3531) );
  INV_X1 U12947 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10364) );
  OR2_X1 U12948 ( .A1(n10362), .A2(n14639), .ZN(n10363) );
  OAI21_X1 U12949 ( .B1(n14641), .B2(n10364), .A(n10363), .ZN(P1_U3468) );
  NAND2_X1 U12950 ( .A1(n10366), .A2(n10365), .ZN(n10367) );
  XNOR2_X1 U12951 ( .A(n10413), .B(n11975), .ZN(n10370) );
  INV_X2 U12952 ( .A(n12001), .ZN(n13295) );
  NAND2_X1 U12953 ( .A1(n13126), .A2(n14410), .ZN(n10371) );
  NAND2_X1 U12954 ( .A1(n10370), .A2(n10371), .ZN(n10502) );
  INV_X1 U12955 ( .A(n10370), .ZN(n10373) );
  INV_X1 U12956 ( .A(n10371), .ZN(n10372) );
  NAND2_X1 U12957 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  NAND2_X1 U12958 ( .A1(n10502), .A2(n10374), .ZN(n10376) );
  INV_X1 U12959 ( .A(n10503), .ZN(n10375) );
  AOI21_X1 U12960 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n10382) );
  NOR2_X1 U12961 ( .A1(n13087), .A2(n10483), .ZN(n10380) );
  AOI22_X1 U12962 ( .A1(n13064), .A2(n13127), .B1(n13125), .B2(n13065), .ZN(
        n10411) );
  OAI21_X1 U12963 ( .B1(n13066), .B2(n10411), .A(n10378), .ZN(n10379) );
  AOI211_X1 U12964 ( .C1(n10413), .C2(n13095), .A(n10380), .B(n10379), .ZN(
        n10381) );
  OAI21_X1 U12965 ( .B1(n10382), .B2(n13091), .A(n10381), .ZN(P2_U3202) );
  INV_X1 U12966 ( .A(n11534), .ZN(n13809) );
  INV_X1 U12967 ( .A(n10383), .ZN(n10386) );
  OAI222_X1 U12968 ( .A1(P1_U3086), .A2(n13809), .B1(n14166), .B2(n10386), 
        .C1(n10384), .C2(n14163), .ZN(P1_U3339) );
  INV_X1 U12969 ( .A(n14725), .ZN(n13174) );
  OAI222_X1 U12970 ( .A1(P2_U3088), .A2(n13174), .B1(n13559), .B2(n10386), 
        .C1(n10385), .C2(n13550), .ZN(P2_U3311) );
  INV_X1 U12971 ( .A(n11526), .ZN(n11547) );
  INV_X1 U12972 ( .A(n10387), .ZN(n10390) );
  OAI222_X1 U12973 ( .A1(P1_U3086), .A2(n11547), .B1(n14166), .B2(n10390), 
        .C1(n10388), .C2(n14163), .ZN(P1_U3341) );
  INV_X1 U12974 ( .A(n14710), .ZN(n13170) );
  OAI222_X1 U12975 ( .A1(P2_U3088), .A2(n13170), .B1(n13559), .B2(n10390), 
        .C1(n10389), .C2(n13550), .ZN(P2_U3313) );
  AND2_X1 U12976 ( .A1(n10392), .A2(n10391), .ZN(n11894) );
  XOR2_X1 U12977 ( .A(n10393), .B(n11894), .Z(n14595) );
  AOI21_X1 U12978 ( .B1(n10394), .B2(n11715), .A(n14509), .ZN(n10395) );
  AND2_X1 U12979 ( .A1(n10395), .A2(n10539), .ZN(n14597) );
  OAI22_X1 U12980 ( .A1(n14035), .A2(n11713), .B1(n14011), .B2(n10583), .ZN(
        n10396) );
  AOI21_X1 U12981 ( .B1(n14597), .B2(n13999), .A(n10396), .ZN(n10404) );
  INV_X1 U12982 ( .A(n11894), .ZN(n10397) );
  XNOR2_X1 U12983 ( .A(n10398), .B(n10397), .ZN(n10400) );
  NOR2_X1 U12984 ( .A1(n10579), .A2(n14021), .ZN(n10399) );
  AOI21_X1 U12985 ( .B1(n10400), .B2(n14028), .A(n10399), .ZN(n14601) );
  NAND2_X1 U12986 ( .A1(n13719), .A2(n14008), .ZN(n14599) );
  AND2_X1 U12987 ( .A1(n14601), .A2(n14599), .ZN(n10401) );
  MUX2_X1 U12988 ( .A(n10402), .B(n10401), .S(n14047), .Z(n10403) );
  OAI211_X1 U12989 ( .C1(n14595), .C2(n14019), .A(n10404), .B(n10403), .ZN(
        P1_U3289) );
  OAI21_X1 U12990 ( .B1(n10406), .B2(n10410), .A(n10405), .ZN(n10474) );
  INV_X1 U12991 ( .A(n10523), .ZN(n10407) );
  AOI211_X1 U12992 ( .C1(n10413), .C2(n10408), .A(n13295), .B(n10407), .ZN(
        n10485) );
  XNOR2_X1 U12993 ( .A(n10409), .B(n10410), .ZN(n10412) );
  OAI21_X1 U12994 ( .B1(n10412), .B2(n13393), .A(n10411), .ZN(n10477) );
  AOI211_X1 U12995 ( .C1(n14816), .C2(n10474), .A(n10485), .B(n10477), .ZN(
        n10419) );
  OAI22_X1 U12996 ( .A1(n13474), .A2(n6931), .B1(n14842), .B2(n8213), .ZN(
        n10414) );
  INV_X1 U12997 ( .A(n10414), .ZN(n10415) );
  OAI21_X1 U12998 ( .B1(n10419), .B2(n8665), .A(n10415), .ZN(P2_U3503) );
  INV_X1 U12999 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10416) );
  OAI22_X1 U13000 ( .A1(n13531), .A2(n6931), .B1(n14836), .B2(n10416), .ZN(
        n10417) );
  INV_X1 U13001 ( .A(n10417), .ZN(n10418) );
  OAI21_X1 U13002 ( .B1(n10419), .B2(n7143), .A(n10418), .ZN(P2_U3442) );
  INV_X1 U13003 ( .A(n11545), .ZN(n13821) );
  INV_X1 U13004 ( .A(n10420), .ZN(n10422) );
  OAI222_X1 U13005 ( .A1(P1_U3086), .A2(n13821), .B1(n14166), .B2(n10422), 
        .C1(n10421), .C2(n14163), .ZN(P1_U3338) );
  INV_X1 U13006 ( .A(n13177), .ZN(n13189) );
  OAI222_X1 U13007 ( .A1(n13550), .A2(n10423), .B1(n13559), .B2(n10422), .C1(
        n13189), .C2(P2_U3088), .ZN(P2_U3310) );
  OAI22_X1 U13008 ( .A1(n14047), .A2(n10424), .B1(n13730), .B2(n14011), .ZN(
        n10427) );
  NOR2_X1 U13009 ( .A1(n14035), .A2(n10425), .ZN(n10426) );
  AOI211_X1 U13010 ( .C1(n10428), .C2(n13999), .A(n10427), .B(n10426), .ZN(
        n10431) );
  INV_X1 U13011 ( .A(n14019), .ZN(n13951) );
  NAND2_X1 U13012 ( .A1(n10429), .A2(n13951), .ZN(n10430) );
  OAI211_X1 U13013 ( .C1(n10432), .C2(n14041), .A(n10431), .B(n10430), .ZN(
        P1_U3291) );
  MUX2_X1 U13014 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12586), .Z(n10619) );
  XNOR2_X1 U13015 ( .A(n10619), .B(n10624), .ZN(n10621) );
  INV_X1 U13016 ( .A(n14902), .ZN(n10459) );
  MUX2_X1 U13017 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12586), .Z(n10440) );
  INV_X1 U13018 ( .A(n10440), .ZN(n10441) );
  INV_X1 U13019 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10434) );
  INV_X1 U13020 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U13021 ( .A(n10434), .B(n10433), .S(n9533), .Z(n10435) );
  NAND2_X1 U13022 ( .A1(n10435), .A2(n10456), .ZN(n10438) );
  INV_X1 U13023 ( .A(n10435), .ZN(n10436) );
  INV_X1 U13024 ( .A(n10456), .ZN(n14889) );
  NAND2_X1 U13025 ( .A1(n10436), .A2(n14889), .ZN(n10437) );
  NAND2_X1 U13026 ( .A1(n10438), .A2(n10437), .ZN(n14880) );
  AOI21_X1 U13027 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14884) );
  INV_X1 U13028 ( .A(n10438), .ZN(n10439) );
  XNOR2_X1 U13029 ( .A(n10440), .B(n14902), .ZN(n14900) );
  MUX2_X1 U13030 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12586), .Z(n10442) );
  AND2_X1 U13031 ( .A1(n10442), .A2(n14924), .ZN(n14920) );
  NOR2_X1 U13032 ( .A1(n10442), .A2(n14924), .ZN(n14921) );
  INV_X1 U13033 ( .A(n14921), .ZN(n10443) );
  XOR2_X1 U13034 ( .A(n10621), .B(n10622), .Z(n10468) );
  NAND2_X1 U13035 ( .A1(n10444), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10445) );
  MUX2_X1 U13036 ( .A(n10812), .B(P3_REG2_REG_4__SCAN_IN), .S(n14902), .Z(
        n14897) );
  NOR2_X1 U13037 ( .A1(n14898), .A2(n14897), .ZN(n14896) );
  INV_X1 U13038 ( .A(n14924), .ZN(n10447) );
  NOR2_X1 U13039 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  INV_X1 U13040 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14919) );
  INV_X1 U13041 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10450) );
  MUX2_X1 U13042 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10450), .S(n10624), .Z(
        n10451) );
  AOI21_X1 U13043 ( .B1(n10452), .B2(n10451), .A(n10627), .ZN(n10453) );
  NOR2_X1 U13044 ( .A1(n15028), .A2(n10453), .ZN(n10466) );
  INV_X1 U13045 ( .A(n15014), .ZN(n14913) );
  INV_X1 U13046 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15079) );
  MUX2_X1 U13047 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15079), .S(n10624), .Z(
        n10462) );
  INV_X1 U13048 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10458) );
  OAI21_X1 U13049 ( .B1(n10455), .B2(n10067), .A(n10454), .ZN(n10457) );
  XNOR2_X1 U13050 ( .A(n10457), .B(n10456), .ZN(n14891) );
  AOI22_X1 U13051 ( .A1(n14891), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n14889), 
        .B2(n10457), .ZN(n14911) );
  MUX2_X1 U13052 ( .A(n10458), .B(P3_REG1_REG_4__SCAN_IN), .S(n14902), .Z(
        n14910) );
  NAND2_X1 U13053 ( .A1(n14924), .A2(n10460), .ZN(n10461) );
  AOI21_X1 U13054 ( .B1(n10462), .B2(n6514), .A(n10623), .ZN(n10464) );
  NAND2_X1 U13055 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13056 ( .A1(n15021), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10463) );
  OAI211_X1 U13057 ( .C1(n14913), .C2(n10464), .A(n11028), .B(n10463), .ZN(
        n10465) );
  AOI211_X1 U13058 ( .C1(n14944), .C2(n10624), .A(n10466), .B(n10465), .ZN(
        n10467) );
  OAI21_X1 U13059 ( .B1(n10468), .B2(n15003), .A(n10467), .ZN(P3_U3188) );
  INV_X1 U13060 ( .A(n10469), .ZN(n10472) );
  OAI222_X1 U13061 ( .A1(P1_U3086), .A2(n11530), .B1(n14166), .B2(n10472), 
        .C1(n10470), .C2(n14163), .ZN(P1_U3340) );
  INV_X1 U13062 ( .A(n14715), .ZN(n13171) );
  OAI222_X1 U13063 ( .A1(P2_U3088), .A2(n13171), .B1(n13559), .B2(n10472), 
        .C1(n10471), .C2(n13550), .ZN(P2_U3312) );
  NAND2_X1 U13064 ( .A1(n12554), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10473) );
  OAI21_X1 U13065 ( .B1(n12655), .B2(n12554), .A(n10473), .ZN(P3_U3519) );
  INV_X1 U13066 ( .A(n10474), .ZN(n10488) );
  AND2_X1 U13067 ( .A1(n10023), .A2(n10475), .ZN(n10476) );
  INV_X1 U13068 ( .A(n10477), .ZN(n10478) );
  MUX2_X1 U13069 ( .A(n10479), .B(n10478), .S(n13336), .Z(n10487) );
  INV_X1 U13070 ( .A(n10481), .ZN(n10482) );
  OAI22_X1 U13071 ( .A1(n13406), .A2(n6931), .B1(n13300), .B2(n10483), .ZN(
        n10484) );
  AOI21_X1 U13072 ( .B1(n10485), .B2(n13402), .A(n10484), .ZN(n10486) );
  OAI211_X1 U13073 ( .C1(n10488), .C2(n13372), .A(n10487), .B(n10486), .ZN(
        P2_U3261) );
  INV_X1 U13074 ( .A(n10489), .ZN(n10496) );
  NOR2_X1 U13075 ( .A1(n13406), .A2(n8204), .ZN(n10491) );
  OAI22_X1 U13076 ( .A1(n13336), .A2(n8194), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n13300), .ZN(n10490) );
  AOI211_X1 U13077 ( .C1(n10492), .C2(n13402), .A(n10491), .B(n10490), .ZN(
        n10495) );
  NAND2_X1 U13078 ( .A1(n10493), .A2(n13336), .ZN(n10494) );
  OAI211_X1 U13079 ( .C1(n13372), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        P2_U3262) );
  INV_X1 U13080 ( .A(n14796), .ZN(n10525) );
  XNOR2_X1 U13081 ( .A(n14796), .B(n11975), .ZN(n10497) );
  NAND2_X1 U13082 ( .A1(n13125), .A2(n14410), .ZN(n10498) );
  NAND2_X1 U13083 ( .A1(n10497), .A2(n10498), .ZN(n10545) );
  INV_X1 U13084 ( .A(n10497), .ZN(n10500) );
  INV_X1 U13085 ( .A(n10498), .ZN(n10499) );
  NAND2_X1 U13086 ( .A1(n10500), .A2(n10499), .ZN(n10501) );
  AND2_X1 U13087 ( .A1(n10545), .A2(n10501), .ZN(n10505) );
  OAI21_X1 U13088 ( .B1(n10505), .B2(n10504), .A(n10546), .ZN(n10506) );
  NAND2_X1 U13089 ( .A1(n10506), .A2(n13060), .ZN(n10511) );
  INV_X1 U13090 ( .A(n10524), .ZN(n10509) );
  AOI22_X1 U13091 ( .A1(n13064), .A2(n13126), .B1(n13124), .B2(n13065), .ZN(
        n10519) );
  OAI21_X1 U13092 ( .B1(n13066), .B2(n10519), .A(n10507), .ZN(n10508) );
  AOI21_X1 U13093 ( .B1(n10509), .B2(n13068), .A(n10508), .ZN(n10510) );
  OAI211_X1 U13094 ( .C1(n10525), .C2(n13071), .A(n10511), .B(n10510), .ZN(
        P2_U3199) );
  INV_X1 U13095 ( .A(n10512), .ZN(n10514) );
  OAI222_X1 U13096 ( .A1(P3_U3151), .A2(n10515), .B1(n12967), .B2(n10514), 
        .C1(n10513), .C2(n12968), .ZN(P3_U3275) );
  XNOR2_X1 U13097 ( .A(n10516), .B(n10517), .ZN(n14798) );
  XOR2_X1 U13098 ( .A(n10518), .B(n10517), .Z(n10520) );
  OAI21_X1 U13099 ( .B1(n10520), .B2(n13393), .A(n10519), .ZN(n14794) );
  INV_X1 U13100 ( .A(n14794), .ZN(n10521) );
  MUX2_X1 U13101 ( .A(n10522), .B(n10521), .S(n13336), .Z(n10528) );
  AOI211_X1 U13102 ( .C1(n14796), .C2(n10523), .A(n13295), .B(n10666), .ZN(
        n14795) );
  OAI22_X1 U13103 ( .A1(n13406), .A2(n10525), .B1(n13300), .B2(n10524), .ZN(
        n10526) );
  AOI21_X1 U13104 ( .B1(n14795), .B2(n13402), .A(n10526), .ZN(n10527) );
  OAI211_X1 U13105 ( .C1(n13372), .C2(n14798), .A(n10528), .B(n10527), .ZN(
        P2_U3260) );
  INV_X1 U13106 ( .A(n10529), .ZN(n10531) );
  OAI21_X1 U13107 ( .B1(n10531), .B2(n11895), .A(n10530), .ZN(n14607) );
  INV_X1 U13108 ( .A(n14607), .ZN(n10544) );
  OR2_X1 U13109 ( .A1(n9930), .A2(n13843), .ZN(n11874) );
  INV_X1 U13110 ( .A(n11874), .ZN(n10532) );
  NAND2_X1 U13111 ( .A1(n14047), .A2(n10532), .ZN(n14037) );
  NAND2_X1 U13112 ( .A1(n10533), .A2(n11895), .ZN(n10534) );
  AOI21_X1 U13113 ( .B1(n10535), .B2(n10534), .A(n14584), .ZN(n10537) );
  OAI22_X1 U13114 ( .A1(n11062), .A2(n14045), .B1(n11714), .B2(n14021), .ZN(
        n10536) );
  AOI211_X1 U13115 ( .C1(n14607), .C2(n13924), .A(n10537), .B(n10536), .ZN(
        n14609) );
  MUX2_X1 U13116 ( .A(n9815), .B(n14609), .S(n14047), .Z(n10543) );
  INV_X1 U13117 ( .A(n10642), .ZN(n10538) );
  AOI211_X1 U13118 ( .C1(n11721), .C2(n10539), .A(n14509), .B(n10538), .ZN(
        n14605) );
  INV_X1 U13119 ( .A(n11721), .ZN(n10540) );
  OAI22_X1 U13120 ( .A1(n10540), .A2(n14035), .B1(n10796), .B2(n14011), .ZN(
        n10541) );
  AOI21_X1 U13121 ( .B1(n14605), .B2(n13999), .A(n10541), .ZN(n10542) );
  OAI211_X1 U13122 ( .C1(n10544), .C2(n14037), .A(n10543), .B(n10542), .ZN(
        P1_U3288) );
  XNOR2_X1 U13123 ( .A(n14803), .B(n11975), .ZN(n10710) );
  NAND2_X1 U13124 ( .A1(n13124), .A2(n14410), .ZN(n10711) );
  XNOR2_X1 U13125 ( .A(n10710), .B(n10711), .ZN(n10715) );
  XNOR2_X1 U13126 ( .A(n10716), .B(n10715), .ZN(n10553) );
  NOR2_X1 U13127 ( .A1(n13087), .A2(n10668), .ZN(n10551) );
  NAND2_X1 U13128 ( .A1(n13123), .A2(n13065), .ZN(n10548) );
  NAND2_X1 U13129 ( .A1(n13125), .A2(n13064), .ZN(n10547) );
  AND2_X1 U13130 ( .A1(n10548), .A2(n10547), .ZN(n10673) );
  OAI21_X1 U13131 ( .B1(n13066), .B2(n10673), .A(n10549), .ZN(n10550) );
  AOI211_X1 U13132 ( .C1(n14803), .C2(n13095), .A(n10551), .B(n10550), .ZN(
        n10552) );
  OAI21_X1 U13133 ( .B1(n10553), .B2(n13091), .A(n10552), .ZN(P2_U3211) );
  OAI21_X1 U13134 ( .B1(n10556), .B2(n10555), .A(n10554), .ZN(n14593) );
  INV_X1 U13135 ( .A(n14593), .ZN(n10572) );
  OAI22_X1 U13136 ( .A1(n14047), .A2(n10558), .B1(n10557), .B2(n14011), .ZN(
        n10562) );
  INV_X1 U13137 ( .A(n13999), .ZN(n13948) );
  NAND2_X1 U13138 ( .A1(n7408), .A2(n11700), .ZN(n10559) );
  NAND2_X1 U13139 ( .A1(n10560), .A2(n10559), .ZN(n10563) );
  OR2_X1 U13140 ( .A1(n10563), .A2(n14509), .ZN(n14589) );
  NOR2_X1 U13141 ( .A1(n13948), .A2(n14589), .ZN(n10561) );
  AOI211_X1 U13142 ( .C1(n14049), .C2(n11700), .A(n10562), .B(n10561), .ZN(
        n10571) );
  XNOR2_X1 U13143 ( .A(n10563), .B(n14046), .ZN(n10564) );
  MUX2_X1 U13144 ( .A(n11893), .B(n10564), .S(n10565), .Z(n10569) );
  OAI22_X1 U13145 ( .A1(n10566), .A2(n14045), .B1(n10565), .B2(n14021), .ZN(
        n10567) );
  AOI21_X1 U13146 ( .B1(n14593), .B2(n13924), .A(n10567), .ZN(n10568) );
  OAI21_X1 U13147 ( .B1(n14584), .B2(n10569), .A(n10568), .ZN(n14591) );
  NAND2_X1 U13148 ( .A1(n14591), .A2(n14047), .ZN(n10570) );
  OAI211_X1 U13149 ( .C1(n10572), .C2(n14037), .A(n10571), .B(n10570), .ZN(
        P1_U3292) );
  OR2_X1 U13150 ( .A1(n11713), .A2(n12062), .ZN(n10577) );
  NAND2_X1 U13151 ( .A1(n13720), .A2(n12152), .ZN(n10576) );
  NAND2_X1 U13152 ( .A1(n10577), .A2(n10576), .ZN(n10782) );
  OAI22_X1 U13153 ( .A1(n11713), .A2(n12161), .B1(n11714), .B2(n12062), .ZN(
        n10578) );
  XNOR2_X1 U13154 ( .A(n10578), .B(n12158), .ZN(n10784) );
  XNOR2_X1 U13155 ( .A(n10785), .B(n10784), .ZN(n10586) );
  NOR2_X1 U13156 ( .A1(n11713), .A2(n14634), .ZN(n14596) );
  INV_X1 U13157 ( .A(n13681), .ZN(n14478) );
  NAND2_X1 U13158 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13755) );
  OAI21_X1 U13159 ( .B1(n14478), .B2(n10580), .A(n13755), .ZN(n10581) );
  AOI21_X1 U13160 ( .B1(n13673), .B2(n6478), .A(n10581), .ZN(n10582) );
  OAI21_X1 U13161 ( .B1(n14494), .B2(n10583), .A(n10582), .ZN(n10584) );
  AOI21_X1 U13162 ( .B1(n13580), .B2(n14596), .A(n10584), .ZN(n10585) );
  OAI21_X1 U13163 ( .B1(n10586), .B2(n14467), .A(n10585), .ZN(P1_U3230) );
  MUX2_X1 U13164 ( .A(n7733), .B(P1_REG1_REG_14__SCAN_IN), .S(n11526), .Z(
        n10592) );
  NAND2_X1 U13165 ( .A1(n10587), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13166 ( .A1(n10589), .A2(n10588), .ZN(n10591) );
  INV_X1 U13167 ( .A(n11528), .ZN(n10590) );
  AOI21_X1 U13168 ( .B1(n10592), .B2(n10591), .A(n10590), .ZN(n10605) );
  MUX2_X1 U13169 ( .A(n11548), .B(P1_REG2_REG_14__SCAN_IN), .S(n11526), .Z(
        n10596) );
  NOR2_X1 U13170 ( .A1(n10594), .A2(n10593), .ZN(n10598) );
  INV_X1 U13171 ( .A(n10598), .ZN(n10595) );
  NAND2_X1 U13172 ( .A1(n10596), .A2(n10595), .ZN(n10599) );
  MUX2_X1 U13173 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11548), .S(n11526), .Z(
        n10597) );
  OAI21_X1 U13174 ( .B1(n10600), .B2(n10598), .A(n10597), .ZN(n11546) );
  OAI211_X1 U13175 ( .C1(n10600), .C2(n10599), .A(n11546), .B(n14560), .ZN(
        n10604) );
  NAND2_X1 U13176 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14459)
         );
  INV_X1 U13177 ( .A(n14459), .ZN(n10602) );
  NOR2_X1 U13178 ( .A1(n13838), .A2(n11547), .ZN(n10601) );
  AOI211_X1 U13179 ( .C1(n14570), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n10602), 
        .B(n10601), .ZN(n10603) );
  OAI211_X1 U13180 ( .C1(n10605), .C2(n11539), .A(n10604), .B(n10603), .ZN(
        P1_U3257) );
  NOR2_X1 U13181 ( .A1(n15030), .A2(n12400), .ZN(n12360) );
  OR3_X1 U13182 ( .A1(n12360), .A2(n14383), .A3(n10606), .ZN(n10608) );
  NAND2_X1 U13183 ( .A1(n9495), .A2(n12797), .ZN(n10607) );
  NAND2_X1 U13184 ( .A1(n10608), .A2(n10607), .ZN(n11677) );
  INV_X1 U13185 ( .A(n11677), .ZN(n10610) );
  AOI22_X1 U13186 ( .A1(n9554), .A2(n10636), .B1(n9553), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n10609) );
  OAI21_X1 U13187 ( .B1(n10610), .B2(n9553), .A(n10609), .ZN(P3_U3459) );
  XOR2_X1 U13188 ( .A(n10612), .B(n10611), .Z(n10618) );
  NAND2_X1 U13189 ( .A1(n10613), .A2(n12955), .ZN(n10743) );
  NAND2_X1 U13190 ( .A1(n9495), .A2(n12827), .ZN(n10615) );
  NAND2_X1 U13191 ( .A1(n12552), .A2(n12797), .ZN(n10614) );
  AND2_X1 U13192 ( .A1(n10615), .A2(n10614), .ZN(n10660) );
  INV_X1 U13193 ( .A(n14865), .ZN(n14851) );
  OAI22_X1 U13194 ( .A1(n10660), .A2(n14851), .B1(n14856), .B2(n10905), .ZN(
        n10616) );
  AOI21_X1 U13195 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10743), .A(n10616), .ZN(
        n10617) );
  OAI21_X1 U13196 ( .B1(n10618), .B2(n12310), .A(n10617), .ZN(P3_U3177) );
  MUX2_X1 U13197 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12586), .Z(n10755) );
  XNOR2_X1 U13198 ( .A(n10755), .B(n10754), .ZN(n10756) );
  INV_X1 U13199 ( .A(n10619), .ZN(n10620) );
  XOR2_X1 U13200 ( .A(n10756), .B(n10757), .Z(n10635) );
  INV_X1 U13201 ( .A(n10754), .ZN(n10762) );
  NAND2_X1 U13202 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10625), .ZN(n10750) );
  OAI21_X1 U13203 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10625), .A(n10750), .ZN(
        n10633) );
  AND2_X1 U13204 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n14846) );
  AOI21_X1 U13205 ( .B1(n15021), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n14846), .ZN(
        n10626) );
  OAI21_X1 U13206 ( .B1(n15018), .B2(n10754), .A(n10626), .ZN(n10632) );
  NOR2_X1 U13207 ( .A1(n9185), .A2(n10629), .ZN(n10763) );
  AOI21_X1 U13208 ( .B1(n10629), .B2(n9185), .A(n10763), .ZN(n10630) );
  NOR2_X1 U13209 ( .A1(n10630), .A2(n15028), .ZN(n10631) );
  AOI211_X1 U13210 ( .C1(n15014), .C2(n10633), .A(n10632), .B(n10631), .ZN(
        n10634) );
  OAI21_X1 U13211 ( .B1(n10635), .B2(n15003), .A(n10634), .ZN(P3_U3189) );
  AOI22_X1 U13212 ( .A1(n12315), .A2(n9495), .B1(n10636), .B2(n14847), .ZN(
        n10638) );
  NAND2_X1 U13213 ( .A1(n10743), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10637) );
  OAI211_X1 U13214 ( .C1(n12360), .C2(n12310), .A(n10638), .B(n10637), .ZN(
        P3_U3172) );
  OAI21_X1 U13215 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(n14617) );
  NAND2_X1 U13216 ( .A1(n10642), .A2(n11725), .ZN(n10643) );
  NAND2_X1 U13217 ( .A1(n10643), .A2(n14126), .ZN(n10644) );
  OR2_X1 U13218 ( .A1(n10644), .A2(n11038), .ZN(n14614) );
  NOR2_X1 U13219 ( .A1(n14614), .A2(n13948), .ZN(n10647) );
  INV_X1 U13220 ( .A(n11725), .ZN(n10645) );
  OAI22_X1 U13221 ( .A1(n10645), .A2(n14035), .B1(n14011), .B2(n10899), .ZN(
        n10646) );
  AOI211_X1 U13222 ( .C1(n14617), .C2(n13951), .A(n10647), .B(n10646), .ZN(
        n10655) );
  XNOR2_X1 U13223 ( .A(n10648), .B(n11897), .ZN(n10649) );
  AND2_X1 U13224 ( .A1(n10649), .A2(n14028), .ZN(n14615) );
  NAND2_X1 U13225 ( .A1(n13719), .A2(n14006), .ZN(n10651) );
  NAND2_X1 U13226 ( .A1(n13717), .A2(n14008), .ZN(n10650) );
  NAND2_X1 U13227 ( .A1(n10651), .A2(n10650), .ZN(n14611) );
  NOR2_X1 U13228 ( .A1(n14615), .A2(n14611), .ZN(n10653) );
  MUX2_X1 U13229 ( .A(n10653), .B(n10652), .S(n14041), .Z(n10654) );
  NAND2_X1 U13230 ( .A1(n10655), .A2(n10654), .ZN(P1_U3287) );
  OAI21_X1 U13231 ( .B1(n10656), .B2(n10657), .A(n10658), .ZN(n10903) );
  XNOR2_X1 U13232 ( .A(n10659), .B(n10657), .ZN(n10661) );
  OAI21_X1 U13233 ( .B1(n10661), .B2(n15038), .A(n10660), .ZN(n10907) );
  AOI21_X1 U13234 ( .B1(n15054), .B2(n10903), .A(n10907), .ZN(n10828) );
  AOI22_X1 U13235 ( .A1(n9554), .A2(n12405), .B1(n9553), .B2(
        P3_REG1_REG_2__SCAN_IN), .ZN(n10662) );
  OAI21_X1 U13236 ( .B1(n10828), .B2(n9553), .A(n10662), .ZN(P3_U3461) );
  INV_X1 U13237 ( .A(n10663), .ZN(n10664) );
  AOI21_X1 U13238 ( .B1(n7128), .B2(n10665), .A(n10664), .ZN(n14809) );
  INV_X1 U13239 ( .A(n14809), .ZN(n14806) );
  INV_X1 U13240 ( .A(n10666), .ZN(n10667) );
  AOI211_X1 U13241 ( .C1(n14803), .C2(n10667), .A(n13295), .B(n10849), .ZN(
        n14802) );
  OAI22_X1 U13242 ( .A1(n13406), .A2(n10669), .B1(n13300), .B2(n10668), .ZN(
        n10670) );
  AOI21_X1 U13243 ( .B1(n14802), .B2(n13402), .A(n10670), .ZN(n10678) );
  XNOR2_X1 U13244 ( .A(n10671), .B(n10672), .ZN(n10674) );
  OAI21_X1 U13245 ( .B1(n10674), .B2(n13393), .A(n10673), .ZN(n14808) );
  INV_X1 U13246 ( .A(n14808), .ZN(n10675) );
  MUX2_X1 U13247 ( .A(n10676), .B(n10675), .S(n13336), .Z(n10677) );
  OAI211_X1 U13248 ( .C1(n14806), .C2(n13372), .A(n10678), .B(n10677), .ZN(
        P2_U3259) );
  INV_X1 U13249 ( .A(n10679), .ZN(n10687) );
  NAND2_X1 U13250 ( .A1(n13402), .A2(n10680), .ZN(n10682) );
  INV_X1 U13251 ( .A(n13300), .ZN(n14402) );
  AOI22_X1 U13252 ( .A1(n13411), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14402), .ZN(n10681) );
  OAI211_X1 U13253 ( .C1(n10683), .C2(n13406), .A(n10682), .B(n10681), .ZN(
        n10684) );
  AOI21_X1 U13254 ( .B1(n14417), .B2(n10685), .A(n10684), .ZN(n10686) );
  OAI21_X1 U13255 ( .B1(n13411), .B2(n10687), .A(n10686), .ZN(P2_U3264) );
  INV_X1 U13256 ( .A(n10688), .ZN(n10697) );
  NOR2_X1 U13257 ( .A1(n13406), .A2(n10689), .ZN(n10692) );
  OAI22_X1 U13258 ( .A1(n13336), .A2(n8180), .B1(n10690), .B2(n13300), .ZN(
        n10691) );
  AOI211_X1 U13259 ( .C1(n10693), .C2(n13402), .A(n10692), .B(n10691), .ZN(
        n10696) );
  NAND2_X1 U13260 ( .A1(n14417), .A2(n10694), .ZN(n10695) );
  OAI211_X1 U13261 ( .C1(n13411), .C2(n10697), .A(n10696), .B(n10695), .ZN(
        P2_U3263) );
  INV_X1 U13262 ( .A(n14037), .ZN(n13932) );
  INV_X1 U13263 ( .A(n14011), .ZN(n14051) );
  INV_X1 U13264 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13265 ( .A1(n14049), .A2(n6646), .B1(n14051), .B2(n10698), .ZN(
        n10699) );
  OAI21_X1 U13266 ( .B1(n13948), .B2(n10700), .A(n10699), .ZN(n10703) );
  MUX2_X1 U13267 ( .A(n10701), .B(P1_REG2_REG_3__SCAN_IN), .S(n14041), .Z(
        n10702) );
  AOI211_X1 U13268 ( .C1(n13932), .C2(n10704), .A(n10703), .B(n10702), .ZN(
        n10705) );
  INV_X1 U13269 ( .A(n10705), .ZN(P1_U3290) );
  INV_X1 U13270 ( .A(n10706), .ZN(n10708) );
  INV_X1 U13271 ( .A(SI_21_), .ZN(n10707) );
  OAI222_X1 U13272 ( .A1(P3_U3151), .A2(n10709), .B1(n12967), .B2(n10708), 
        .C1(n10707), .C2(n12968), .ZN(P3_U3274) );
  INV_X1 U13273 ( .A(n10710), .ZN(n10713) );
  INV_X1 U13274 ( .A(n10711), .ZN(n10712) );
  NAND2_X1 U13275 ( .A1(n10713), .A2(n10712), .ZN(n10714) );
  XNOR2_X1 U13276 ( .A(n10852), .B(n6637), .ZN(n10920) );
  NAND2_X1 U13277 ( .A1(n13123), .A2(n13295), .ZN(n10918) );
  XNOR2_X1 U13278 ( .A(n10920), .B(n10918), .ZN(n10916) );
  XNOR2_X1 U13279 ( .A(n10917), .B(n10916), .ZN(n10723) );
  NOR2_X1 U13280 ( .A1(n13087), .A2(n10850), .ZN(n10721) );
  NAND2_X1 U13281 ( .A1(n13122), .A2(n13065), .ZN(n10718) );
  NAND2_X1 U13282 ( .A1(n13124), .A2(n13064), .ZN(n10717) );
  AND2_X1 U13283 ( .A1(n10718), .A2(n10717), .ZN(n10858) );
  OAI21_X1 U13284 ( .B1(n13066), .B2(n10858), .A(n10719), .ZN(n10720) );
  AOI211_X1 U13285 ( .C1(n10852), .C2(n13095), .A(n10721), .B(n10720), .ZN(
        n10722) );
  OAI21_X1 U13286 ( .B1(n10723), .B2(n13091), .A(n10722), .ZN(P2_U3185) );
  XNOR2_X1 U13287 ( .A(n6721), .B(n10724), .ZN(n10725) );
  NAND2_X1 U13288 ( .A1(n10725), .A2(n14028), .ZN(n10727) );
  AOI22_X1 U13289 ( .A1(n14006), .A2(n13717), .B1(n13715), .B2(n14008), .ZN(
        n10726) );
  NAND2_X1 U13290 ( .A1(n10727), .A2(n10726), .ZN(n14628) );
  INV_X1 U13291 ( .A(n14628), .ZN(n10735) );
  OAI21_X1 U13292 ( .B1(n10729), .B2(n6721), .A(n10728), .ZN(n14630) );
  NAND2_X1 U13293 ( .A1(n14630), .A2(n13951), .ZN(n10734) );
  INV_X1 U13294 ( .A(n10963), .ZN(n10730) );
  AOI211_X1 U13295 ( .C1(n11739), .C2(n11037), .A(n14509), .B(n10730), .ZN(
        n14627) );
  INV_X1 U13296 ( .A(n11739), .ZN(n11165) );
  NOR2_X1 U13297 ( .A1(n11165), .A2(n14035), .ZN(n10732) );
  OAI22_X1 U13298 ( .A1(n14047), .A2(n9820), .B1(n11168), .B2(n14011), .ZN(
        n10731) );
  AOI211_X1 U13299 ( .C1(n14627), .C2(n13999), .A(n10732), .B(n10731), .ZN(
        n10733) );
  OAI211_X1 U13300 ( .C1(n10735), .C2(n14041), .A(n10734), .B(n10733), .ZN(
        P1_U3285) );
  INV_X1 U13301 ( .A(n10736), .ZN(n15036) );
  INV_X1 U13302 ( .A(n15030), .ZN(n10738) );
  NAND3_X1 U13303 ( .A1(n10736), .A2(n10738), .A3(n10737), .ZN(n10739) );
  OAI211_X1 U13304 ( .C1(n10741), .C2(n9596), .A(n10740), .B(n10739), .ZN(
        n10747) );
  INV_X1 U13305 ( .A(n12555), .ZN(n15041) );
  AOI22_X1 U13306 ( .A1(n12315), .A2(n12553), .B1(n10742), .B2(n14847), .ZN(
        n10745) );
  NAND2_X1 U13307 ( .A1(n10743), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n10744) );
  OAI211_X1 U13308 ( .C1(n15041), .C2(n12317), .A(n10745), .B(n10744), .ZN(
        n10746) );
  AOI21_X1 U13309 ( .B1(n10747), .B2(n14857), .A(n10746), .ZN(n10748) );
  INV_X1 U13310 ( .A(n10748), .ZN(P3_U3162) );
  INV_X1 U13311 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15081) );
  MUX2_X1 U13312 ( .A(n15081), .B(P3_REG1_REG_8__SCAN_IN), .S(n11203), .Z(
        n10753) );
  NAND2_X1 U13313 ( .A1(n10754), .A2(n10749), .ZN(n10751) );
  AOI21_X1 U13314 ( .B1(n10753), .B2(n10752), .A(n11185), .ZN(n10773) );
  OAI22_X1 U13315 ( .A1(n10757), .A2(n10756), .B1(n10755), .B2(n10754), .ZN(
        n10759) );
  MUX2_X1 U13316 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12586), .Z(n11192) );
  XNOR2_X1 U13317 ( .A(n11192), .B(n11186), .ZN(n10758) );
  NAND2_X1 U13318 ( .A1(n10759), .A2(n10758), .ZN(n11193) );
  OAI21_X1 U13319 ( .B1(n10759), .B2(n10758), .A(n11193), .ZN(n10760) );
  NAND2_X1 U13320 ( .A1(n10760), .A2(n15022), .ZN(n10772) );
  NOR2_X1 U13321 ( .A1(n10762), .A2(n10761), .ZN(n10764) );
  NOR2_X1 U13322 ( .A1(n10764), .A2(n10763), .ZN(n10767) );
  INV_X1 U13323 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10765) );
  MUX2_X1 U13324 ( .A(n10765), .B(P3_REG2_REG_8__SCAN_IN), .S(n11203), .Z(
        n10766) );
  AOI21_X1 U13325 ( .B1(n10767), .B2(n10766), .A(n11202), .ZN(n10769) );
  AND2_X1 U13326 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11235) );
  AOI21_X1 U13327 ( .B1(n15021), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11235), .ZN(
        n10768) );
  OAI21_X1 U13328 ( .B1(n15028), .B2(n10769), .A(n10768), .ZN(n10770) );
  AOI21_X1 U13329 ( .B1(n11186), .B2(n14944), .A(n10770), .ZN(n10771) );
  OAI211_X1 U13330 ( .C1(n10773), .C2(n14913), .A(n10772), .B(n10771), .ZN(
        P3_U3190) );
  OAI21_X1 U13331 ( .B1(n10774), .B2(n12359), .A(n10775), .ZN(n10814) );
  NAND2_X1 U13332 ( .A1(n10937), .A2(n12414), .ZN(n10869) );
  OAI211_X1 U13333 ( .C1(n10937), .C2(n12414), .A(n10869), .B(n12832), .ZN(
        n10779) );
  NAND2_X1 U13334 ( .A1(n12552), .A2(n12827), .ZN(n10778) );
  NAND2_X1 U13335 ( .A1(n12550), .A2(n12829), .ZN(n10777) );
  AND2_X1 U13336 ( .A1(n10778), .A2(n10777), .ZN(n10835) );
  NAND2_X1 U13337 ( .A1(n10779), .A2(n10835), .ZN(n10802) );
  AOI21_X1 U13338 ( .B1(n15054), .B2(n10814), .A(n10802), .ZN(n10824) );
  AOI22_X1 U13339 ( .A1(n9554), .A2(n10833), .B1(n9553), .B2(
        P3_REG1_REG_4__SCAN_IN), .ZN(n10780) );
  OAI21_X1 U13340 ( .B1(n10824), .B2(n9553), .A(n10780), .ZN(P3_U3463) );
  INV_X1 U13341 ( .A(n13580), .ZN(n13636) );
  NAND2_X1 U13342 ( .A1(n11721), .A2(n14124), .ZN(n14604) );
  INV_X1 U13343 ( .A(n10781), .ZN(n10783) );
  NAND2_X1 U13344 ( .A1(n11721), .A2(n12147), .ZN(n10787) );
  NAND2_X1 U13345 ( .A1(n13719), .A2(n12148), .ZN(n10786) );
  NAND2_X1 U13346 ( .A1(n10787), .A2(n10786), .ZN(n10788) );
  XNOR2_X1 U13347 ( .A(n10788), .B(n12158), .ZN(n10792) );
  NAND2_X1 U13348 ( .A1(n11721), .A2(n12148), .ZN(n10790) );
  NAND2_X1 U13349 ( .A1(n13719), .A2(n12152), .ZN(n10789) );
  NAND2_X1 U13350 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  NOR2_X1 U13351 ( .A1(n10792), .A2(n10791), .ZN(n10893) );
  NAND2_X1 U13352 ( .A1(n10792), .A2(n10791), .ZN(n10892) );
  INV_X1 U13353 ( .A(n10892), .ZN(n10793) );
  NOR2_X1 U13354 ( .A1(n10893), .A2(n10793), .ZN(n10794) );
  XNOR2_X1 U13355 ( .A(n10894), .B(n10794), .ZN(n10795) );
  NAND2_X1 U13356 ( .A1(n10795), .A2(n14483), .ZN(n10801) );
  NOR2_X1 U13357 ( .A1(n14494), .A2(n10796), .ZN(n10799) );
  OAI22_X1 U13358 ( .A1(n14478), .A2(n11062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10797), .ZN(n10798) );
  AOI211_X1 U13359 ( .C1(n13673), .C2(n13720), .A(n10799), .B(n10798), .ZN(
        n10800) );
  OAI211_X1 U13360 ( .C1(n13636), .C2(n14604), .A(n10801), .B(n10800), .ZN(
        P1_U3227) );
  INV_X1 U13361 ( .A(n10802), .ZN(n10816) );
  NAND2_X1 U13362 ( .A1(n10804), .A2(n10803), .ZN(n10807) );
  NAND2_X1 U13363 ( .A1(n10805), .A2(n12954), .ZN(n10806) );
  AND2_X1 U13364 ( .A1(n10807), .A2(n10806), .ZN(n10808) );
  NAND2_X1 U13365 ( .A1(n10809), .A2(n10808), .ZN(n10810) );
  AND2_X1 U13366 ( .A1(n15034), .A2(n12398), .ZN(n10946) );
  OR2_X1 U13367 ( .A1(n12683), .A2(n10946), .ZN(n15044) );
  INV_X1 U13368 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10812) );
  OR2_X1 U13369 ( .A1(n15034), .A2(n15068), .ZN(n10904) );
  INV_X1 U13370 ( .A(n12807), .ZN(n12837) );
  AOI22_X1 U13371 ( .A1(n12837), .A2(n10833), .B1(n12805), .B2(n10837), .ZN(
        n10811) );
  OAI21_X1 U13372 ( .B1(n10812), .B2(n15045), .A(n10811), .ZN(n10813) );
  AOI21_X1 U13373 ( .B1(n10814), .B2(n12841), .A(n10813), .ZN(n10815) );
  OAI21_X1 U13374 ( .B1(n10816), .B2(n12844), .A(n10815), .ZN(P3_U3229) );
  INV_X1 U13375 ( .A(n10817), .ZN(n10819) );
  OAI22_X1 U13376 ( .A1(n12529), .A2(P3_U3151), .B1(SI_22_), .B2(n11489), .ZN(
        n10818) );
  AOI21_X1 U13377 ( .B1(n10819), .B2(n10931), .A(n10818), .ZN(P3_U3273) );
  INV_X1 U13378 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10820) );
  OAI22_X1 U13379 ( .A1(n12952), .A2(n10821), .B1(n15076), .B2(n10820), .ZN(
        n10822) );
  INV_X1 U13380 ( .A(n10822), .ZN(n10823) );
  OAI21_X1 U13381 ( .B1(n10824), .B2(n15074), .A(n10823), .ZN(P3_U3402) );
  INV_X1 U13382 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n10825) );
  OAI22_X1 U13383 ( .A1(n12952), .A2(n10905), .B1(n15076), .B2(n10825), .ZN(
        n10826) );
  INV_X1 U13384 ( .A(n10826), .ZN(n10827) );
  OAI21_X1 U13385 ( .B1(n10828), .B2(n15074), .A(n10827), .ZN(P3_U3396) );
  INV_X1 U13386 ( .A(n10829), .ZN(n10830) );
  AOI21_X1 U13387 ( .B1(n10832), .B2(n10831), .A(n10830), .ZN(n10839) );
  AOI22_X1 U13388 ( .A1(n10833), .A2(n14847), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10834) );
  OAI21_X1 U13389 ( .B1(n10835), .B2(n14851), .A(n10834), .ZN(n10836) );
  AOI21_X1 U13390 ( .B1(n10837), .B2(n12326), .A(n10836), .ZN(n10838) );
  OAI21_X1 U13391 ( .B1(n10839), .B2(n12310), .A(n10838), .ZN(P3_U3170) );
  INV_X1 U13392 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10840) );
  OAI22_X1 U13393 ( .A1(n12952), .A2(n11678), .B1(n15076), .B2(n10840), .ZN(
        n10841) );
  AOI21_X1 U13394 ( .B1(n11677), .B2(n15076), .A(n10841), .ZN(n10842) );
  INV_X1 U13395 ( .A(n10842), .ZN(P3_U3390) );
  INV_X1 U13396 ( .A(n10843), .ZN(n10846) );
  OAI222_X1 U13397 ( .A1(n11554), .A2(P1_U3086), .B1(n14166), .B2(n10846), 
        .C1(n10844), .C2(n14163), .ZN(P1_U3337) );
  INV_X1 U13398 ( .A(n14740), .ZN(n10845) );
  OAI222_X1 U13399 ( .A1(n13550), .A2(n10847), .B1(n13559), .B2(n10846), .C1(
        P2_U3088), .C2(n10845), .ZN(P2_U3309) );
  XOR2_X1 U13400 ( .A(n10848), .B(n10854), .Z(n14817) );
  OAI211_X1 U13401 ( .C1(n14813), .C2(n10849), .A(n12001), .B(n10985), .ZN(
        n14812) );
  INV_X1 U13402 ( .A(n10850), .ZN(n10851) );
  AOI22_X1 U13403 ( .A1(n14403), .A2(n10852), .B1(n14402), .B2(n10851), .ZN(
        n10853) );
  OAI21_X1 U13404 ( .B1(n14812), .B2(n14415), .A(n10853), .ZN(n10861) );
  INV_X1 U13405 ( .A(n10854), .ZN(n10855) );
  XNOR2_X1 U13406 ( .A(n10856), .B(n10855), .ZN(n10857) );
  NAND2_X1 U13407 ( .A1(n10857), .A2(n14399), .ZN(n10859) );
  NAND2_X1 U13408 ( .A1(n10859), .A2(n10858), .ZN(n14814) );
  MUX2_X1 U13409 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n14814), .S(n13336), .Z(
        n10860) );
  AOI211_X1 U13410 ( .C1(n14417), .C2(n14817), .A(n10861), .B(n10860), .ZN(
        n10862) );
  INV_X1 U13411 ( .A(n10862), .ZN(P2_U3258) );
  OAI21_X1 U13412 ( .B1(n10864), .B2(n12423), .A(n10863), .ZN(n10865) );
  INV_X1 U13413 ( .A(n10865), .ZN(n11156) );
  AND2_X1 U13414 ( .A1(n10869), .A2(n10866), .ZN(n10871) );
  NAND2_X1 U13415 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  OAI21_X1 U13416 ( .B1(n10871), .B2(n12364), .A(n10870), .ZN(n10873) );
  OAI22_X1 U13417 ( .A1(n11093), .A2(n15042), .B1(n10872), .B2(n15040), .ZN(
        n10973) );
  AOI21_X1 U13418 ( .B1(n10873), .B2(n12832), .A(n10973), .ZN(n11152) );
  OAI21_X1 U13419 ( .B1(n14372), .B2(n11156), .A(n11152), .ZN(n10879) );
  INV_X1 U13420 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10874) );
  OAI22_X1 U13421 ( .A1(n12898), .A2(n10971), .B1(n15085), .B2(n10874), .ZN(
        n10875) );
  AOI21_X1 U13422 ( .B1(n10879), .B2(n15085), .A(n10875), .ZN(n10876) );
  INV_X1 U13423 ( .A(n10876), .ZN(P3_U3464) );
  INV_X1 U13424 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10877) );
  OAI22_X1 U13425 ( .A1(n12952), .A2(n10971), .B1(n15076), .B2(n10877), .ZN(
        n10878) );
  AOI21_X1 U13426 ( .B1(n10879), .B2(n15076), .A(n10878), .ZN(n10880) );
  INV_X1 U13427 ( .A(n10880), .ZN(P3_U3405) );
  XNOR2_X1 U13428 ( .A(n10883), .B(n10882), .ZN(n11069) );
  INV_X1 U13429 ( .A(n11069), .ZN(n10891) );
  XNOR2_X1 U13430 ( .A(n10885), .B(n10884), .ZN(n10886) );
  AOI22_X1 U13431 ( .A1(n13064), .A2(n13122), .B1(n13119), .B2(n13065), .ZN(
        n11109) );
  OAI21_X1 U13432 ( .B1(n10886), .B2(n13393), .A(n11109), .ZN(n11067) );
  NAND2_X1 U13433 ( .A1(n11067), .A2(n13336), .ZN(n10890) );
  AOI211_X1 U13434 ( .C1(n11112), .C2(n10986), .A(n13295), .B(n11013), .ZN(
        n11068) );
  NOR2_X1 U13435 ( .A1(n7297), .A2(n13406), .ZN(n10888) );
  OAI22_X1 U13436 ( .A1(n13336), .A2(n9982), .B1(n11107), .B2(n13300), .ZN(
        n10887) );
  AOI211_X1 U13437 ( .C1(n11068), .C2(n13402), .A(n10888), .B(n10887), .ZN(
        n10889) );
  OAI211_X1 U13438 ( .C1(n10891), .C2(n13372), .A(n10890), .B(n10889), .ZN(
        P2_U3256) );
  NAND2_X1 U13439 ( .A1(n11725), .A2(n14124), .ZN(n14612) );
  AND2_X1 U13440 ( .A1(n13718), .A2(n12152), .ZN(n10895) );
  AOI21_X1 U13441 ( .B1(n11725), .B2(n12132), .A(n10895), .ZN(n11050) );
  AOI22_X1 U13442 ( .A1(n11725), .A2(n12147), .B1(n12148), .B2(n13718), .ZN(
        n10896) );
  XNOR2_X1 U13443 ( .A(n10896), .B(n12158), .ZN(n11049) );
  XOR2_X1 U13444 ( .A(n11050), .B(n11049), .Z(n10897) );
  NAND2_X1 U13445 ( .A1(n10898), .A2(n10897), .ZN(n11054) );
  OAI211_X1 U13446 ( .C1(n10898), .C2(n10897), .A(n11054), .B(n14483), .ZN(
        n10902) );
  AND2_X1 U13447 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13774) );
  NOR2_X1 U13448 ( .A1(n14494), .A2(n10899), .ZN(n10900) );
  AOI211_X1 U13449 ( .C1(n13658), .C2(n14611), .A(n13774), .B(n10900), .ZN(
        n10901) );
  OAI211_X1 U13450 ( .C1(n13636), .C2(n14612), .A(n10902), .B(n10901), .ZN(
        P1_U3239) );
  INV_X1 U13451 ( .A(n12841), .ZN(n12791) );
  INV_X1 U13452 ( .A(n10903), .ZN(n10911) );
  INV_X1 U13453 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15199) );
  OAI22_X1 U13454 ( .A1(n10905), .A2(n10904), .B1(n15199), .B2(n15032), .ZN(
        n10906) );
  NOR2_X1 U13455 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  MUX2_X1 U13456 ( .A(n10909), .B(n10908), .S(n15045), .Z(n10910) );
  OAI21_X1 U13457 ( .B1(n12791), .B2(n10911), .A(n10910), .ZN(P3_U3231) );
  XNOR2_X1 U13458 ( .A(n14820), .B(n11975), .ZN(n10912) );
  NAND2_X1 U13459 ( .A1(n13122), .A2(n13295), .ZN(n10913) );
  NAND2_X1 U13460 ( .A1(n10912), .A2(n10913), .ZN(n11100) );
  INV_X1 U13461 ( .A(n10912), .ZN(n10915) );
  INV_X1 U13462 ( .A(n10913), .ZN(n10914) );
  NAND2_X1 U13463 ( .A1(n10915), .A2(n10914), .ZN(n11102) );
  NAND2_X1 U13464 ( .A1(n11100), .A2(n11102), .ZN(n10923) );
  NAND2_X1 U13465 ( .A1(n10917), .A2(n10916), .ZN(n10922) );
  INV_X1 U13466 ( .A(n10918), .ZN(n10919) );
  NAND2_X1 U13467 ( .A1(n10920), .A2(n10919), .ZN(n10921) );
  NAND2_X1 U13468 ( .A1(n10922), .A2(n10921), .ZN(n11101) );
  XOR2_X1 U13469 ( .A(n10923), .B(n11101), .Z(n10930) );
  NAND2_X1 U13470 ( .A1(n13120), .A2(n13065), .ZN(n10925) );
  NAND2_X1 U13471 ( .A1(n13123), .A2(n13064), .ZN(n10924) );
  NAND2_X1 U13472 ( .A1(n10925), .A2(n10924), .ZN(n10981) );
  NAND2_X1 U13473 ( .A1(n13085), .A2(n10981), .ZN(n10926) );
  OAI211_X1 U13474 ( .C1(n13087), .C2(n10988), .A(n10927), .B(n10926), .ZN(
        n10928) );
  AOI21_X1 U13475 ( .B1(n14820), .B2(n13095), .A(n10928), .ZN(n10929) );
  OAI21_X1 U13476 ( .B1(n10930), .B2(n13091), .A(n10929), .ZN(P2_U3193) );
  INV_X1 U13477 ( .A(SI_23_), .ZN(n10934) );
  NAND2_X1 U13478 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  OAI211_X1 U13479 ( .C1(n10934), .C2(n11489), .A(n10933), .B(n12531), .ZN(
        P3_U3272) );
  XNOR2_X1 U13480 ( .A(n10935), .B(n6476), .ZN(n10945) );
  INV_X1 U13481 ( .A(n12683), .ZN(n11282) );
  NAND2_X1 U13482 ( .A1(n10937), .A2(n10936), .ZN(n10938) );
  AND2_X1 U13483 ( .A1(n10940), .A2(n10941), .ZN(n10942) );
  OAI211_X1 U13484 ( .C1(n7434), .C2(n6476), .A(n12832), .B(n10942), .ZN(
        n10944) );
  AOI22_X1 U13485 ( .A1(n12548), .A2(n12797), .B1(n12827), .B2(n12550), .ZN(
        n10943) );
  OAI211_X1 U13486 ( .C1(n10945), .C2(n11282), .A(n10944), .B(n10943), .ZN(
        n15058) );
  INV_X1 U13487 ( .A(n15058), .ZN(n10951) );
  INV_X1 U13488 ( .A(n10945), .ZN(n15060) );
  AND2_X1 U13489 ( .A1(n15045), .A2(n10946), .ZN(n12690) );
  AOI22_X1 U13490 ( .A1(n12837), .A2(n10947), .B1(n12805), .B2(n11031), .ZN(
        n10948) );
  OAI21_X1 U13491 ( .B1(n10450), .B2(n15045), .A(n10948), .ZN(n10949) );
  AOI21_X1 U13492 ( .B1(n15060), .B2(n12690), .A(n10949), .ZN(n10950) );
  OAI21_X1 U13493 ( .B1(n10951), .B2(n12844), .A(n10950), .ZN(P3_U3227) );
  INV_X1 U13494 ( .A(n10952), .ZN(n10955) );
  OAI222_X1 U13495 ( .A1(n13550), .A2(n10953), .B1(n13559), .B2(n10955), .C1(
        n8653), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13496 ( .A1(P1_U3086), .A2(n13843), .B1(n14166), .B2(n10955), 
        .C1(n10954), .C2(n14163), .ZN(P1_U3336) );
  OAI21_X1 U13497 ( .B1(n10957), .B2(n11902), .A(n10956), .ZN(n11115) );
  INV_X1 U13498 ( .A(n10958), .ZN(n10959) );
  AOI21_X1 U13499 ( .B1(n11902), .B2(n10960), .A(n10959), .ZN(n10961) );
  AOI22_X1 U13500 ( .A1(n14006), .A2(n13716), .B1(n13714), .B2(n14008), .ZN(
        n11355) );
  OAI21_X1 U13501 ( .B1(n10961), .B2(n14584), .A(n11355), .ZN(n10962) );
  AOI21_X1 U13502 ( .B1(n13924), .B2(n11115), .A(n10962), .ZN(n11118) );
  INV_X1 U13503 ( .A(n11748), .ZN(n11360) );
  AOI211_X1 U13504 ( .C1(n11748), .C2(n10963), .A(n14509), .B(n11082), .ZN(
        n11116) );
  NAND2_X1 U13505 ( .A1(n11116), .A2(n13999), .ZN(n10966) );
  INV_X1 U13506 ( .A(n10964), .ZN(n11357) );
  AOI22_X1 U13507 ( .A1(n14041), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11357), 
        .B2(n14051), .ZN(n10965) );
  OAI211_X1 U13508 ( .C1(n11360), .C2(n14035), .A(n10966), .B(n10965), .ZN(
        n10967) );
  AOI21_X1 U13509 ( .B1(n11115), .B2(n13932), .A(n10967), .ZN(n10968) );
  OAI21_X1 U13510 ( .B1(n11118), .B2(n14041), .A(n10968), .ZN(P1_U3284) );
  XOR2_X1 U13511 ( .A(n10970), .B(n10969), .Z(n10976) );
  OAI22_X1 U13512 ( .A1(n14856), .A2(n10971), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15191), .ZN(n10972) );
  AOI21_X1 U13513 ( .B1(n10973), .B2(n14865), .A(n10972), .ZN(n10975) );
  NAND2_X1 U13514 ( .A1(n12326), .A2(n11153), .ZN(n10974) );
  OAI211_X1 U13515 ( .C1(n10976), .C2(n12310), .A(n10975), .B(n10974), .ZN(
        P3_U3167) );
  XNOR2_X1 U13516 ( .A(n10977), .B(n10980), .ZN(n14824) );
  INV_X1 U13517 ( .A(n14824), .ZN(n10993) );
  NAND2_X1 U13518 ( .A1(n14824), .A2(n14810), .ZN(n10984) );
  OAI21_X1 U13519 ( .B1(n10980), .B2(n10978), .A(n10979), .ZN(n10982) );
  AOI21_X1 U13520 ( .B1(n10982), .B2(n14399), .A(n10981), .ZN(n10983) );
  AND2_X1 U13521 ( .A1(n10984), .A2(n10983), .ZN(n14826) );
  MUX2_X1 U13522 ( .A(n9970), .B(n14826), .S(n13336), .Z(n10992) );
  AOI21_X1 U13523 ( .B1(n10985), .B2(n14820), .A(n13295), .ZN(n10987) );
  AND2_X1 U13524 ( .A1(n10987), .A2(n10986), .ZN(n14822) );
  INV_X1 U13525 ( .A(n14820), .ZN(n10989) );
  OAI22_X1 U13526 ( .A1(n10989), .A2(n13406), .B1(n13300), .B2(n10988), .ZN(
        n10990) );
  AOI21_X1 U13527 ( .B1(n14822), .B2(n13402), .A(n10990), .ZN(n10991) );
  OAI211_X1 U13528 ( .C1(n10993), .C2(n13389), .A(n10992), .B(n10991), .ZN(
        P2_U3257) );
  OAI21_X1 U13529 ( .B1(n10995), .B2(n12358), .A(n10994), .ZN(n11308) );
  NAND2_X1 U13530 ( .A1(n12549), .A2(n12827), .ZN(n10998) );
  NAND2_X1 U13531 ( .A1(n12547), .A2(n12797), .ZN(n10997) );
  AND2_X1 U13532 ( .A1(n10998), .A2(n10997), .ZN(n14852) );
  NAND2_X1 U13533 ( .A1(n10999), .A2(n14852), .ZN(n11305) );
  AOI21_X1 U13534 ( .B1(n15054), .B2(n11308), .A(n11305), .ZN(n11005) );
  INV_X1 U13535 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11000) );
  OAI22_X1 U13536 ( .A1(n12898), .A2(n11304), .B1(n15085), .B2(n11000), .ZN(
        n11001) );
  INV_X1 U13537 ( .A(n11001), .ZN(n11002) );
  OAI21_X1 U13538 ( .B1(n11005), .B2(n9553), .A(n11002), .ZN(P3_U3466) );
  OAI22_X1 U13539 ( .A1(n12952), .A2(n11304), .B1(n15076), .B2(n9186), .ZN(
        n11003) );
  INV_X1 U13540 ( .A(n11003), .ZN(n11004) );
  OAI21_X1 U13541 ( .B1(n11005), .B2(n15074), .A(n11004), .ZN(P3_U3411) );
  XNOR2_X1 U13542 ( .A(n11007), .B(n11006), .ZN(n11124) );
  INV_X1 U13543 ( .A(n11124), .ZN(n11021) );
  XNOR2_X1 U13544 ( .A(n11009), .B(n11008), .ZN(n11012) );
  NAND2_X1 U13545 ( .A1(n13118), .A2(n13065), .ZN(n11011) );
  NAND2_X1 U13546 ( .A1(n13120), .A2(n13064), .ZN(n11010) );
  AND2_X1 U13547 ( .A1(n11011), .A2(n11010), .ZN(n11146) );
  OAI21_X1 U13548 ( .B1(n11012), .B2(n13393), .A(n11146), .ZN(n11122) );
  NAND2_X1 U13549 ( .A1(n11122), .A2(n13336), .ZN(n11020) );
  INV_X1 U13550 ( .A(n11013), .ZN(n11015) );
  INV_X1 U13551 ( .A(n11014), .ZN(n11247) );
  AOI211_X1 U13552 ( .C1(n11133), .C2(n11015), .A(n13295), .B(n11247), .ZN(
        n11123) );
  NOR2_X1 U13553 ( .A1(n11151), .A2(n13406), .ZN(n11018) );
  OAI22_X1 U13554 ( .A1(n13336), .A2(n11016), .B1(n11144), .B2(n13300), .ZN(
        n11017) );
  AOI211_X1 U13555 ( .C1(n11123), .C2(n13402), .A(n11018), .B(n11017), .ZN(
        n11019) );
  OAI211_X1 U13556 ( .C1(n11021), .C2(n13372), .A(n11020), .B(n11019), .ZN(
        P2_U3255) );
  INV_X1 U13557 ( .A(n11022), .ZN(n11937) );
  OAI222_X1 U13558 ( .A1(n13550), .A2(n11024), .B1(P2_U3088), .B2(n11023), 
        .C1(n13552), .C2(n11937), .ZN(P2_U3307) );
  OAI211_X1 U13559 ( .C1(n11027), .C2(n11026), .A(n11025), .B(n14857), .ZN(
        n11033) );
  INV_X1 U13560 ( .A(n12317), .ZN(n12025) );
  AOI22_X1 U13561 ( .A1(n12548), .A2(n12315), .B1(n12025), .B2(n12550), .ZN(
        n11029) );
  OAI211_X1 U13562 ( .C1(n15057), .C2(n14856), .A(n11029), .B(n11028), .ZN(
        n11030) );
  AOI21_X1 U13563 ( .B1(n11031), .B2(n12326), .A(n11030), .ZN(n11032) );
  NAND2_X1 U13564 ( .A1(n11033), .A2(n11032), .ZN(P3_U3179) );
  OR2_X1 U13565 ( .A1(n11034), .A2(n11041), .ZN(n11035) );
  NAND2_X1 U13566 ( .A1(n11036), .A2(n11035), .ZN(n14619) );
  OAI211_X1 U13567 ( .C1(n11038), .C2(n14622), .A(n11037), .B(n14126), .ZN(
        n14620) );
  INV_X1 U13568 ( .A(n11039), .ZN(n11064) );
  AOI22_X1 U13569 ( .A1(n11734), .A2(n14049), .B1(n11064), .B2(n14051), .ZN(
        n11040) );
  OAI21_X1 U13570 ( .B1(n14620), .B2(n13948), .A(n11040), .ZN(n11047) );
  XNOR2_X1 U13571 ( .A(n11042), .B(n11041), .ZN(n11045) );
  NAND2_X1 U13572 ( .A1(n14619), .A2(n13924), .ZN(n11044) );
  AOI22_X1 U13573 ( .A1(n14006), .A2(n13718), .B1(n13716), .B2(n14008), .ZN(
        n11043) );
  OAI211_X1 U13574 ( .C1(n14584), .C2(n11045), .A(n11044), .B(n11043), .ZN(
        n14624) );
  MUX2_X1 U13575 ( .A(n14624), .B(P1_REG2_REG_7__SCAN_IN), .S(n14041), .Z(
        n11046) );
  AOI211_X1 U13576 ( .C1(n13932), .C2(n14619), .A(n11047), .B(n11046), .ZN(
        n11048) );
  INV_X1 U13577 ( .A(n11048), .ZN(P1_U3286) );
  INV_X1 U13578 ( .A(n11049), .ZN(n11052) );
  INV_X1 U13579 ( .A(n11050), .ZN(n11051) );
  NAND2_X1 U13580 ( .A1(n11054), .A2(n11053), .ZN(n11059) );
  OAI22_X1 U13581 ( .A1(n14622), .A2(n12161), .B1(n11055), .B2(n12062), .ZN(
        n11056) );
  XNOR2_X1 U13582 ( .A(n11056), .B(n12158), .ZN(n11158) );
  AND2_X1 U13583 ( .A1(n13717), .A2(n12152), .ZN(n11057) );
  AOI21_X1 U13584 ( .B1(n11734), .B2(n12132), .A(n11057), .ZN(n11159) );
  XNOR2_X1 U13585 ( .A(n11158), .B(n11159), .ZN(n11058) );
  NAND2_X2 U13586 ( .A1(n11059), .A2(n11058), .ZN(n11162) );
  OAI211_X1 U13587 ( .C1(n11059), .C2(n11058), .A(n11162), .B(n14483), .ZN(
        n11066) );
  INV_X1 U13588 ( .A(n14494), .ZN(n13695) );
  AOI21_X1 U13589 ( .B1(n13681), .B2(n13716), .A(n11060), .ZN(n11061) );
  OAI21_X1 U13590 ( .B1(n14477), .B2(n11062), .A(n11061), .ZN(n11063) );
  AOI21_X1 U13591 ( .B1(n11064), .B2(n13695), .A(n11063), .ZN(n11065) );
  OAI211_X1 U13592 ( .C1(n14622), .C2(n13699), .A(n11066), .B(n11065), .ZN(
        P1_U3213) );
  AOI211_X1 U13593 ( .C1(n14816), .C2(n11069), .A(n11068), .B(n11067), .ZN(
        n11073) );
  NOR2_X1 U13594 ( .A1(n14836), .A2(n8286), .ZN(n11070) );
  AOI21_X1 U13595 ( .B1(n11112), .B2(n8940), .A(n11070), .ZN(n11071) );
  OAI21_X1 U13596 ( .B1(n11073), .B2(n7143), .A(n11071), .ZN(P2_U3457) );
  INV_X1 U13597 ( .A(n13474), .ZN(n11125) );
  AOI22_X1 U13598 ( .A1(n11112), .A2(n11125), .B1(n8665), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11072) );
  OAI21_X1 U13599 ( .B1(n11073), .B2(n8665), .A(n11072), .ZN(P2_U3508) );
  INV_X1 U13600 ( .A(n11074), .ZN(n11078) );
  OAI222_X1 U13601 ( .A1(n13550), .A2(n11076), .B1(n13559), .B2(n11078), .C1(
        n11075), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13602 ( .A1(P1_U3086), .A2(n11691), .B1(n14166), .B2(n11078), 
        .C1(n11077), .C2(n14163), .ZN(P1_U3334) );
  OAI21_X1 U13603 ( .B1(n6703), .B2(n11903), .A(n11079), .ZN(n14637) );
  INV_X1 U13604 ( .A(n14637), .ZN(n11091) );
  OAI22_X1 U13605 ( .A1(n14047), .A2(n10191), .B1(n11472), .B2(n14011), .ZN(
        n11081) );
  AOI21_X1 U13606 ( .B1(n11757), .B2(n14049), .A(n11081), .ZN(n11090) );
  INV_X1 U13607 ( .A(n11082), .ZN(n11083) );
  AOI21_X1 U13608 ( .B1(n11083), .B2(n11757), .A(n14509), .ZN(n11084) );
  AOI22_X1 U13609 ( .A1(n11084), .A2(n11294), .B1(n14008), .B2(n13713), .ZN(
        n14632) );
  AOI21_X1 U13610 ( .B1(n11085), .B2(n11903), .A(n14584), .ZN(n11087) );
  AOI22_X1 U13611 ( .A1(n11087), .A2(n11086), .B1(n14006), .B2(n13715), .ZN(
        n14633) );
  OAI21_X1 U13612 ( .B1(n11688), .B2(n14632), .A(n14633), .ZN(n11088) );
  NAND2_X1 U13613 ( .A1(n11088), .A2(n14047), .ZN(n11089) );
  OAI211_X1 U13614 ( .C1(n11091), .C2(n14019), .A(n11090), .B(n11089), .ZN(
        P1_U3283) );
  AOI21_X1 U13615 ( .B1(n11092), .B2(n12357), .A(n15038), .ZN(n11095) );
  OAI22_X1 U13616 ( .A1(n15039), .A2(n15042), .B1(n11093), .B2(n15040), .ZN(
        n14864) );
  AOI21_X1 U13617 ( .B1(n11095), .B2(n11094), .A(n14864), .ZN(n15051) );
  OAI22_X1 U13618 ( .A1(n12807), .A2(n15052), .B1(n15032), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n11096) );
  AOI21_X1 U13619 ( .B1(n12844), .B2(P3_REG2_REG_3__SCAN_IN), .A(n11096), .ZN(
        n11099) );
  XNOR2_X1 U13620 ( .A(n12357), .B(n11097), .ZN(n15055) );
  NAND2_X1 U13621 ( .A1(n15055), .A2(n12841), .ZN(n11098) );
  OAI211_X1 U13622 ( .C1(n15051), .C2(n12844), .A(n11099), .B(n11098), .ZN(
        P3_U3230) );
  XNOR2_X1 U13623 ( .A(n11112), .B(n11975), .ZN(n11132) );
  NAND2_X1 U13624 ( .A1(n13120), .A2(n13295), .ZN(n11131) );
  XNOR2_X1 U13625 ( .A(n11132), .B(n11131), .ZN(n11106) );
  INV_X1 U13626 ( .A(n11141), .ZN(n11104) );
  AOI21_X1 U13627 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n11114) );
  NOR2_X1 U13628 ( .A1(n13087), .A2(n11107), .ZN(n11111) );
  OAI22_X1 U13629 ( .A1(n13066), .A2(n11109), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11108), .ZN(n11110) );
  AOI211_X1 U13630 ( .C1(n11112), .C2(n13095), .A(n11111), .B(n11110), .ZN(
        n11113) );
  OAI21_X1 U13631 ( .B1(n11114), .B2(n13091), .A(n11113), .ZN(P2_U3203) );
  INV_X1 U13632 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11121) );
  INV_X1 U13633 ( .A(n11115), .ZN(n11119) );
  AOI21_X1 U13634 ( .B1(n11748), .B2(n14124), .A(n11116), .ZN(n11117) );
  OAI211_X1 U13635 ( .C1(n11119), .C2(n14130), .A(n11118), .B(n11117), .ZN(
        n14132) );
  NAND2_X1 U13636 ( .A1(n14132), .A2(n14641), .ZN(n11120) );
  OAI21_X1 U13637 ( .B1(n14641), .B2(n11121), .A(n11120), .ZN(P1_U3486) );
  AOI211_X1 U13638 ( .C1(n14816), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        n11130) );
  AOI22_X1 U13639 ( .A1(n11133), .A2(n11125), .B1(n8665), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11126) );
  OAI21_X1 U13640 ( .B1(n11130), .B2(n8665), .A(n11126), .ZN(P2_U3509) );
  INV_X1 U13641 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11127) );
  OAI22_X1 U13642 ( .A1(n11151), .A2(n13531), .B1(n14836), .B2(n11127), .ZN(
        n11128) );
  INV_X1 U13643 ( .A(n11128), .ZN(n11129) );
  OAI21_X1 U13644 ( .B1(n11130), .B2(n7143), .A(n11129), .ZN(P2_U3460) );
  NAND2_X1 U13645 ( .A1(n11132), .A2(n11131), .ZN(n11139) );
  AND2_X1 U13646 ( .A1(n11141), .A2(n11139), .ZN(n11143) );
  XNOR2_X1 U13647 ( .A(n11133), .B(n6637), .ZN(n11134) );
  AND2_X1 U13648 ( .A1(n13119), .A2(n13295), .ZN(n11135) );
  NAND2_X1 U13649 ( .A1(n11134), .A2(n11135), .ZN(n11261) );
  INV_X1 U13650 ( .A(n11134), .ZN(n11137) );
  INV_X1 U13651 ( .A(n11135), .ZN(n11136) );
  NAND2_X1 U13652 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  AND2_X1 U13653 ( .A1(n11261), .A2(n11138), .ZN(n11142) );
  AND2_X1 U13654 ( .A1(n11142), .A2(n11139), .ZN(n11140) );
  OAI211_X1 U13655 ( .C1(n11143), .C2(n11142), .A(n6650), .B(n13060), .ZN(
        n11150) );
  INV_X1 U13656 ( .A(n11144), .ZN(n11148) );
  OAI21_X1 U13657 ( .B1(n13066), .B2(n11146), .A(n11145), .ZN(n11147) );
  AOI21_X1 U13658 ( .B1(n11148), .B2(n13068), .A(n11147), .ZN(n11149) );
  OAI211_X1 U13659 ( .C1(n11151), .C2(n13071), .A(n11150), .B(n11149), .ZN(
        P2_U3189) );
  MUX2_X1 U13660 ( .A(n11152), .B(n14919), .S(n12844), .Z(n11155) );
  AOI22_X1 U13661 ( .A1(n12837), .A2(n12418), .B1(n12805), .B2(n11153), .ZN(
        n11154) );
  OAI211_X1 U13662 ( .C1(n11156), .C2(n12791), .A(n11155), .B(n11154), .ZN(
        P3_U3228) );
  AOI22_X1 U13663 ( .A1(n11739), .A2(n12147), .B1(n12148), .B2(n13716), .ZN(
        n11157) );
  XNOR2_X1 U13664 ( .A(n11157), .B(n12158), .ZN(n11346) );
  AOI22_X1 U13665 ( .A1(n11739), .A2(n12132), .B1(n12152), .B2(n13716), .ZN(
        n11345) );
  XNOR2_X1 U13666 ( .A(n11346), .B(n11345), .ZN(n11164) );
  INV_X1 U13667 ( .A(n11159), .ZN(n11160) );
  NAND2_X1 U13668 ( .A1(n11158), .A2(n11160), .ZN(n11161) );
  AOI21_X1 U13669 ( .B1(n11164), .B2(n11163), .A(n11347), .ZN(n11171) );
  NOR2_X1 U13670 ( .A1(n11165), .A2(n14634), .ZN(n14626) );
  AOI22_X1 U13671 ( .A1(n13681), .A2(n13715), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11167) );
  NAND2_X1 U13672 ( .A1(n13673), .A2(n13717), .ZN(n11166) );
  OAI211_X1 U13673 ( .C1(n14494), .C2(n11168), .A(n11167), .B(n11166), .ZN(
        n11169) );
  AOI21_X1 U13674 ( .B1(n14626), .B2(n13580), .A(n11169), .ZN(n11170) );
  OAI21_X1 U13675 ( .B1(n11171), .B2(n14467), .A(n11170), .ZN(P1_U3221) );
  INV_X1 U13676 ( .A(n11172), .ZN(n11173) );
  OAI222_X1 U13677 ( .A1(n13550), .A2(n11174), .B1(n13559), .B2(n11173), .C1(
        n8148), .C2(P2_U3088), .ZN(P2_U3305) );
  XOR2_X1 U13678 ( .A(n12435), .B(n11175), .Z(n11180) );
  XNOR2_X1 U13679 ( .A(n11176), .B(n12435), .ZN(n11178) );
  OAI22_X1 U13680 ( .A1(n11233), .A2(n15040), .B1(n11232), .B2(n15042), .ZN(
        n11177) );
  AOI21_X1 U13681 ( .B1(n11178), .B2(n12832), .A(n11177), .ZN(n11179) );
  OAI21_X1 U13682 ( .B1(n11180), .B2(n11282), .A(n11179), .ZN(n15063) );
  INV_X1 U13683 ( .A(n15063), .ZN(n11184) );
  INV_X1 U13684 ( .A(n11180), .ZN(n15065) );
  AOI22_X1 U13685 ( .A1(n12837), .A2(n11236), .B1(n12805), .B2(n11228), .ZN(
        n11181) );
  OAI21_X1 U13686 ( .B1(n10765), .B2(n15045), .A(n11181), .ZN(n11182) );
  AOI21_X1 U13687 ( .B1(n15065), .B2(n12690), .A(n11182), .ZN(n11183) );
  OAI21_X1 U13688 ( .B1(n11184), .B2(n12844), .A(n11183), .ZN(P3_U3225) );
  NAND2_X1 U13689 ( .A1(n11195), .A2(n11187), .ZN(n11188) );
  XOR2_X1 U13690 ( .A(n11195), .B(n11187), .Z(n14943) );
  NAND2_X1 U13691 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14943), .ZN(n14942) );
  INV_X1 U13692 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11189) );
  MUX2_X1 U13693 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11189), .S(n12557), .Z(
        n11190) );
  OAI21_X1 U13694 ( .B1(n11191), .B2(n11190), .A(n12571), .ZN(n11211) );
  OR2_X1 U13695 ( .A1(n11192), .A2(n11203), .ZN(n11194) );
  NAND2_X1 U13696 ( .A1(n11194), .A2(n11193), .ZN(n14937) );
  INV_X1 U13697 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14940) );
  INV_X1 U13698 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15083) );
  MUX2_X1 U13699 ( .A(n14940), .B(n15083), .S(n12586), .Z(n11196) );
  INV_X1 U13700 ( .A(n11195), .ZN(n14945) );
  OR2_X1 U13701 ( .A1(n11196), .A2(n14945), .ZN(n14934) );
  NAND2_X1 U13702 ( .A1(n11196), .A2(n14945), .ZN(n14935) );
  INV_X1 U13703 ( .A(n14935), .ZN(n11197) );
  MUX2_X1 U13704 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12586), .Z(n12587) );
  XNOR2_X1 U13705 ( .A(n12587), .B(n12557), .ZN(n11198) );
  NOR2_X1 U13706 ( .A1(n11199), .A2(n11198), .ZN(n12588) );
  AOI21_X1 U13707 ( .B1(n11199), .B2(n11198), .A(n12588), .ZN(n11201) );
  INV_X1 U13708 ( .A(n12557), .ZN(n12590) );
  AOI22_X1 U13709 ( .A1(n14944), .A2(n12590), .B1(n15021), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n11200) );
  OAI21_X1 U13710 ( .B1(n11201), .B2(n15003), .A(n11200), .ZN(n11210) );
  NOR2_X1 U13711 ( .A1(n14945), .A2(n11204), .ZN(n11205) );
  INV_X1 U13712 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11206) );
  MUX2_X1 U13713 ( .A(n11206), .B(P3_REG2_REG_10__SCAN_IN), .S(n12557), .Z(
        n11207) );
  AOI21_X1 U13714 ( .B1(n6618), .B2(n11207), .A(n12556), .ZN(n11208) );
  NAND2_X1 U13715 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n11570)
         );
  OAI21_X1 U13716 ( .B1(n11208), .B2(n15028), .A(n11570), .ZN(n11209) );
  AOI211_X1 U13717 ( .C1(n15014), .C2(n11211), .A(n11210), .B(n11209), .ZN(
        n11212) );
  INV_X1 U13718 ( .A(n11212), .ZN(P3_U3192) );
  XNOR2_X1 U13719 ( .A(n11213), .B(n11214), .ZN(n14442) );
  NAND2_X1 U13720 ( .A1(n14442), .A2(n14810), .ZN(n11221) );
  INV_X1 U13721 ( .A(n11214), .ZN(n11215) );
  XNOR2_X1 U13722 ( .A(n11216), .B(n11215), .ZN(n11219) );
  NAND2_X1 U13723 ( .A1(n13116), .A2(n13065), .ZN(n11218) );
  NAND2_X1 U13724 ( .A1(n13118), .A2(n13064), .ZN(n11217) );
  NAND2_X1 U13725 ( .A1(n11218), .A2(n11217), .ZN(n11404) );
  AOI21_X1 U13726 ( .B1(n11219), .B2(n14399), .A(n11404), .ZN(n11220) );
  AND2_X1 U13727 ( .A1(n11221), .A2(n11220), .ZN(n14444) );
  AOI21_X1 U13728 ( .B1(n14439), .B2(n11246), .A(n14410), .ZN(n11222) );
  NAND2_X1 U13729 ( .A1(n11222), .A2(n11382), .ZN(n14440) );
  OAI22_X1 U13730 ( .A1(n13336), .A2(n13134), .B1(n11406), .B2(n13300), .ZN(
        n11223) );
  AOI21_X1 U13731 ( .B1(n14439), .B2(n14403), .A(n11223), .ZN(n11224) );
  OAI21_X1 U13732 ( .B1(n14440), .B2(n14415), .A(n11224), .ZN(n11225) );
  AOI21_X1 U13733 ( .B1(n14442), .B2(n11226), .A(n11225), .ZN(n11227) );
  OAI21_X1 U13734 ( .B1(n14444), .B2(n14420), .A(n11227), .ZN(P2_U3253) );
  INV_X1 U13735 ( .A(n11228), .ZN(n11239) );
  OAI211_X1 U13736 ( .C1(n11231), .C2(n11230), .A(n11229), .B(n14857), .ZN(
        n11238) );
  OAI22_X1 U13737 ( .A1(n11233), .A2(n12276), .B1(n11232), .B2(n12317), .ZN(
        n11234) );
  AOI211_X1 U13738 ( .C1(n11236), .C2(n14847), .A(n11235), .B(n11234), .ZN(
        n11237) );
  OAI211_X1 U13739 ( .C1(n11239), .C2(n14867), .A(n11238), .B(n11237), .ZN(
        P3_U3161) );
  XNOR2_X1 U13740 ( .A(n11240), .B(n11245), .ZN(n11243) );
  NAND2_X1 U13741 ( .A1(n13117), .A2(n13065), .ZN(n11242) );
  NAND2_X1 U13742 ( .A1(n13119), .A2(n13064), .ZN(n11241) );
  NAND2_X1 U13743 ( .A1(n11242), .A2(n11241), .ZN(n11270) );
  AOI21_X1 U13744 ( .B1(n11243), .B2(n14399), .A(n11270), .ZN(n14830) );
  XOR2_X1 U13745 ( .A(n11245), .B(n11244), .Z(n14831) );
  INV_X1 U13746 ( .A(n14831), .ZN(n14834) );
  INV_X1 U13747 ( .A(n11263), .ZN(n14829) );
  OAI211_X1 U13748 ( .C1(n11247), .C2(n14829), .A(n12001), .B(n11246), .ZN(
        n14827) );
  OAI22_X1 U13749 ( .A1(n13336), .A2(n13132), .B1(n11267), .B2(n13300), .ZN(
        n11248) );
  AOI21_X1 U13750 ( .B1(n11263), .B2(n14403), .A(n11248), .ZN(n11249) );
  OAI21_X1 U13751 ( .B1(n14827), .B2(n14415), .A(n11249), .ZN(n11250) );
  AOI21_X1 U13752 ( .B1(n14834), .B2(n14417), .A(n11250), .ZN(n11251) );
  OAI21_X1 U13753 ( .B1(n13411), .B2(n14830), .A(n11251), .ZN(P2_U3254) );
  XNOR2_X1 U13754 ( .A(n11252), .B(n7000), .ZN(n11253) );
  AOI222_X1 U13755 ( .A1(n12832), .A2(n11253), .B1(n12546), .B2(n12827), .C1(
        n12544), .C2(n12797), .ZN(n11312) );
  INV_X1 U13756 ( .A(n11579), .ZN(n11254) );
  OAI22_X1 U13757 ( .A1(n12807), .A2(n11572), .B1(n11254), .B2(n15032), .ZN(
        n11255) );
  AOI21_X1 U13758 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12844), .A(n11255), 
        .ZN(n11260) );
  NAND2_X1 U13759 ( .A1(n11258), .A2(n11257), .ZN(n11310) );
  NAND3_X1 U13760 ( .A1(n11256), .A2(n11310), .A3(n12841), .ZN(n11259) );
  OAI211_X1 U13761 ( .C1(n11312), .C2(n12844), .A(n11260), .B(n11259), .ZN(
        P3_U3223) );
  NAND2_X1 U13762 ( .A1(n13118), .A2(n13295), .ZN(n11408) );
  XNOR2_X1 U13763 ( .A(n11407), .B(n11408), .ZN(n11264) );
  OAI21_X1 U13764 ( .B1(n11265), .B2(n11264), .A(n11410), .ZN(n11266) );
  NAND2_X1 U13765 ( .A1(n11266), .A2(n13060), .ZN(n11272) );
  NOR2_X1 U13766 ( .A1(n13087), .A2(n11267), .ZN(n11268) );
  AOI211_X1 U13767 ( .C1(n13085), .C2(n11270), .A(n11269), .B(n11268), .ZN(
        n11271) );
  OAI211_X1 U13768 ( .C1(n14829), .C2(n13071), .A(n11272), .B(n11271), .ZN(
        P2_U3208) );
  XNOR2_X1 U13769 ( .A(n11273), .B(n11276), .ZN(n15067) );
  INV_X1 U13770 ( .A(n12690), .ZN(n11287) );
  XNOR2_X1 U13771 ( .A(n11275), .B(n7001), .ZN(n11280) );
  OAI22_X1 U13772 ( .A1(n11278), .A2(n15042), .B1(n11277), .B2(n15040), .ZN(
        n11279) );
  AOI21_X1 U13773 ( .B1(n11280), .B2(n12832), .A(n11279), .ZN(n11281) );
  OAI21_X1 U13774 ( .B1(n11282), .B2(n15067), .A(n11281), .ZN(n15070) );
  NAND2_X1 U13775 ( .A1(n15070), .A2(n15045), .ZN(n11286) );
  INV_X1 U13776 ( .A(n11370), .ZN(n11283) );
  OAI22_X1 U13777 ( .A1(n12807), .A2(n15069), .B1(n11283), .B2(n15032), .ZN(
        n11284) );
  AOI21_X1 U13778 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n12844), .A(n11284), .ZN(
        n11285) );
  OAI211_X1 U13779 ( .C1(n15067), .C2(n11287), .A(n11286), .B(n11285), .ZN(
        P3_U3224) );
  INV_X1 U13780 ( .A(n11288), .ZN(n11290) );
  INV_X1 U13781 ( .A(SI_24_), .ZN(n11289) );
  OAI222_X1 U13782 ( .A1(P3_U3151), .A2(n11291), .B1(n12967), .B2(n11290), 
        .C1(n11289), .C2(n11489), .ZN(P3_U3271) );
  XNOR2_X1 U13783 ( .A(n11292), .B(n11904), .ZN(n11293) );
  AOI222_X1 U13784 ( .A1(n13712), .A2(n14008), .B1(n13714), .B2(n14006), .C1(
        n14028), .C2(n11293), .ZN(n11420) );
  AOI21_X1 U13785 ( .B1(n11294), .B2(n14489), .A(n14509), .ZN(n11295) );
  AND2_X1 U13786 ( .A1(n11295), .A2(n11326), .ZN(n11418) );
  NAND2_X1 U13787 ( .A1(n14489), .A2(n14049), .ZN(n11297) );
  NAND2_X1 U13788 ( .A1(n14041), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11296) );
  OAI211_X1 U13789 ( .C1(n14011), .C2(n14493), .A(n11297), .B(n11296), .ZN(
        n11302) );
  OAI21_X1 U13790 ( .B1(n11299), .B2(n11904), .A(n11298), .ZN(n11300) );
  INV_X1 U13791 ( .A(n11300), .ZN(n11421) );
  NOR2_X1 U13792 ( .A1(n11421), .A2(n14019), .ZN(n11301) );
  AOI211_X1 U13793 ( .C1(n11418), .C2(n13999), .A(n11302), .B(n11301), .ZN(
        n11303) );
  OAI21_X1 U13794 ( .B1(n14041), .B2(n11420), .A(n11303), .ZN(P1_U3282) );
  OAI22_X1 U13795 ( .A1(n12807), .A2(n11304), .B1(n14855), .B2(n15032), .ZN(
        n11307) );
  MUX2_X1 U13796 ( .A(n11305), .B(P3_REG2_REG_7__SCAN_IN), .S(n12844), .Z(
        n11306) );
  AOI211_X1 U13797 ( .C1(n12841), .C2(n11308), .A(n11307), .B(n11306), .ZN(
        n11309) );
  INV_X1 U13798 ( .A(n11309), .ZN(P3_U3226) );
  NAND3_X1 U13799 ( .A1(n11256), .A2(n11310), .A3(n15054), .ZN(n11311) );
  AND2_X1 U13800 ( .A1(n11312), .A2(n11311), .ZN(n11318) );
  INV_X1 U13801 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11313) );
  OAI22_X1 U13802 ( .A1(n12952), .A2(n11572), .B1(n15076), .B2(n11313), .ZN(
        n11314) );
  INV_X1 U13803 ( .A(n11314), .ZN(n11315) );
  OAI21_X1 U13804 ( .B1(n11318), .B2(n15074), .A(n11315), .ZN(P3_U3420) );
  AOI22_X1 U13805 ( .A1(n9554), .A2(n11316), .B1(n9553), .B2(
        P3_REG1_REG_10__SCAN_IN), .ZN(n11317) );
  OAI21_X1 U13806 ( .B1(n11318), .B2(n9553), .A(n11317), .ZN(P3_U3469) );
  XNOR2_X1 U13807 ( .A(n11319), .B(n11905), .ZN(n11325) );
  OAI21_X1 U13808 ( .B1(n11322), .B2(n11321), .A(n11320), .ZN(n14292) );
  NAND2_X1 U13809 ( .A1(n14292), .A2(n13924), .ZN(n11324) );
  AOI22_X1 U13810 ( .A1(n14006), .A2(n13713), .B1(n13711), .B2(n14008), .ZN(
        n11323) );
  OAI211_X1 U13811 ( .C1(n14584), .C2(n11325), .A(n11324), .B(n11323), .ZN(
        n14290) );
  INV_X1 U13812 ( .A(n14290), .ZN(n11333) );
  INV_X1 U13813 ( .A(n11326), .ZN(n11327) );
  OAI211_X1 U13814 ( .C1(n6896), .C2(n11327), .A(n6898), .B(n14126), .ZN(
        n14289) );
  INV_X1 U13815 ( .A(n11328), .ZN(n11645) );
  AOI22_X1 U13816 ( .A1(n14041), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11645), 
        .B2(n14051), .ZN(n11330) );
  NAND2_X1 U13817 ( .A1(n11768), .A2(n14049), .ZN(n11329) );
  OAI211_X1 U13818 ( .C1(n14289), .C2(n13948), .A(n11330), .B(n11329), .ZN(
        n11331) );
  AOI21_X1 U13819 ( .B1(n14292), .B2(n13932), .A(n11331), .ZN(n11332) );
  OAI21_X1 U13820 ( .B1(n11333), .B2(n14041), .A(n11332), .ZN(P1_U3281) );
  XNOR2_X1 U13821 ( .A(n11334), .B(n11906), .ZN(n11335) );
  AOI22_X1 U13822 ( .A1(n13710), .A2(n14008), .B1(n14006), .B2(n13712), .ZN(
        n13650) );
  OAI21_X1 U13823 ( .B1(n11335), .B2(n14584), .A(n13650), .ZN(n11480) );
  INV_X1 U13824 ( .A(n11480), .ZN(n11344) );
  OAI21_X1 U13825 ( .B1(n11338), .B2(n11337), .A(n11336), .ZN(n11482) );
  OAI211_X1 U13826 ( .C1(n13655), .C2(n11339), .A(n14126), .B(n11457), .ZN(
        n11479) );
  OAI22_X1 U13827 ( .A1(n14047), .A2(n10593), .B1(n13648), .B2(n14011), .ZN(
        n11340) );
  AOI21_X1 U13828 ( .B1(n12040), .B2(n14049), .A(n11340), .ZN(n11341) );
  OAI21_X1 U13829 ( .B1(n11479), .B2(n13948), .A(n11341), .ZN(n11342) );
  AOI21_X1 U13830 ( .B1(n11482), .B2(n13951), .A(n11342), .ZN(n11343) );
  OAI21_X1 U13831 ( .B1(n14041), .B2(n11344), .A(n11343), .ZN(P1_U3280) );
  NAND2_X1 U13832 ( .A1(n11748), .A2(n12147), .ZN(n11349) );
  NAND2_X1 U13833 ( .A1(n13715), .A2(n12148), .ZN(n11348) );
  NAND2_X1 U13834 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  XNOR2_X1 U13835 ( .A(n11350), .B(n12158), .ZN(n11463) );
  AND2_X1 U13836 ( .A1(n13715), .A2(n12152), .ZN(n11351) );
  AOI21_X1 U13837 ( .B1(n11748), .B2(n12132), .A(n11351), .ZN(n11464) );
  XNOR2_X1 U13838 ( .A(n11463), .B(n11464), .ZN(n11352) );
  OAI211_X1 U13839 ( .C1(n11353), .C2(n11352), .A(n11467), .B(n14483), .ZN(
        n11359) );
  INV_X1 U13840 ( .A(n13658), .ZN(n13692) );
  OAI22_X1 U13841 ( .A1(n11355), .A2(n13692), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11354), .ZN(n11356) );
  AOI21_X1 U13842 ( .B1(n11357), .B2(n13695), .A(n11356), .ZN(n11358) );
  OAI211_X1 U13843 ( .C1(n11360), .C2(n13699), .A(n11359), .B(n11358), .ZN(
        P1_U3231) );
  INV_X1 U13844 ( .A(n11361), .ZN(n11363) );
  OAI222_X1 U13845 ( .A1(n12191), .A2(n11363), .B1(n12968), .B2(n15186), .C1(
        P3_U3151), .C2(n11362), .ZN(P3_U3269) );
  INV_X1 U13846 ( .A(n11364), .ZN(n11365) );
  AOI21_X1 U13847 ( .B1(n11367), .B2(n11366), .A(n11365), .ZN(n11372) );
  AOI22_X1 U13848 ( .A1(n12025), .A2(n12547), .B1(n12315), .B2(n12545), .ZN(
        n11368) );
  NAND2_X1 U13849 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n14951) );
  OAI211_X1 U13850 ( .C1(n14856), .C2(n15069), .A(n11368), .B(n14951), .ZN(
        n11369) );
  AOI21_X1 U13851 ( .B1(n11370), .B2(n12326), .A(n11369), .ZN(n11371) );
  OAI21_X1 U13852 ( .B1(n11372), .B2(n12310), .A(n11371), .ZN(P3_U3171) );
  INV_X1 U13853 ( .A(n11390), .ZN(n11374) );
  NAND2_X1 U13854 ( .A1(n14149), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11373) );
  OAI211_X1 U13855 ( .C1(n11374), .C2(n14166), .A(n11373), .B(n11934), .ZN(
        P1_U3332) );
  XOR2_X1 U13856 ( .A(n11375), .B(n11381), .Z(n11379) );
  NAND2_X1 U13857 ( .A1(n13115), .A2(n13065), .ZN(n11377) );
  NAND2_X1 U13858 ( .A1(n13117), .A2(n13064), .ZN(n11376) );
  NAND2_X1 U13859 ( .A1(n11377), .A2(n11376), .ZN(n11445) );
  INV_X1 U13860 ( .A(n11445), .ZN(n11378) );
  OAI21_X1 U13861 ( .B1(n11379), .B2(n13393), .A(n11378), .ZN(n14436) );
  INV_X1 U13862 ( .A(n14436), .ZN(n11388) );
  XOR2_X1 U13863 ( .A(n11381), .B(n11380), .Z(n14438) );
  INV_X1 U13864 ( .A(n11431), .ZN(n14435) );
  INV_X1 U13865 ( .A(n11382), .ZN(n11383) );
  OAI211_X1 U13866 ( .C1(n14435), .C2(n11383), .A(n12001), .B(n14411), .ZN(
        n14434) );
  OAI22_X1 U13867 ( .A1(n13336), .A2(n13152), .B1(n11443), .B2(n13300), .ZN(
        n11384) );
  AOI21_X1 U13868 ( .B1(n11431), .B2(n14403), .A(n11384), .ZN(n11385) );
  OAI21_X1 U13869 ( .B1(n14434), .B2(n14415), .A(n11385), .ZN(n11386) );
  AOI21_X1 U13870 ( .B1(n14438), .B2(n14417), .A(n11386), .ZN(n11387) );
  OAI21_X1 U13871 ( .B1(n11388), .B2(n14420), .A(n11387), .ZN(P2_U3252) );
  NAND2_X1 U13872 ( .A1(n11390), .A2(n11389), .ZN(n11392) );
  OAI211_X1 U13873 ( .C1(n11393), .C2(n13550), .A(n11392), .B(n11391), .ZN(
        P2_U3304) );
  XNOR2_X1 U13874 ( .A(n11394), .B(n9266), .ZN(n11397) );
  NAND2_X1 U13875 ( .A1(n12545), .A2(n12827), .ZN(n11396) );
  NAND2_X1 U13876 ( .A1(n12543), .A2(n12797), .ZN(n11395) );
  NAND2_X1 U13877 ( .A1(n11396), .A2(n11395), .ZN(n12292) );
  AOI21_X1 U13878 ( .B1(n11397), .B2(n12832), .A(n12292), .ZN(n14387) );
  NAND2_X1 U13879 ( .A1(n11398), .A2(n12447), .ZN(n11399) );
  NAND2_X1 U13880 ( .A1(n11400), .A2(n11399), .ZN(n14385) );
  AOI22_X1 U13881 ( .A1(n12844), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n12805), 
        .B2(n12296), .ZN(n11401) );
  OAI21_X1 U13882 ( .B1(n12294), .B2(n12807), .A(n11401), .ZN(n11402) );
  AOI21_X1 U13883 ( .B1(n14385), .B2(n12841), .A(n11402), .ZN(n11403) );
  OAI21_X1 U13884 ( .B1(n14387), .B2(n12844), .A(n11403), .ZN(P3_U3222) );
  NAND2_X1 U13885 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n13139)
         );
  NAND2_X1 U13886 ( .A1(n13085), .A2(n11404), .ZN(n11405) );
  OAI211_X1 U13887 ( .C1(n13087), .C2(n11406), .A(n13139), .B(n11405), .ZN(
        n11416) );
  INV_X1 U13888 ( .A(n11407), .ZN(n11409) );
  NAND2_X1 U13889 ( .A1(n11409), .A2(n11408), .ZN(n11412) );
  XNOR2_X1 U13890 ( .A(n14439), .B(n6637), .ZN(n11426) );
  NAND2_X1 U13891 ( .A1(n13117), .A2(n13295), .ZN(n11427) );
  XNOR2_X1 U13892 ( .A(n11426), .B(n11427), .ZN(n11411) );
  INV_X1 U13893 ( .A(n11411), .ZN(n11413) );
  NAND3_X1 U13894 ( .A1(n11410), .A2(n11413), .A3(n11412), .ZN(n11414) );
  AOI21_X1 U13895 ( .B1(n11430), .B2(n11414), .A(n13091), .ZN(n11415) );
  AOI211_X1 U13896 ( .C1(n14439), .C2(n13095), .A(n11416), .B(n11415), .ZN(
        n11417) );
  INV_X1 U13897 ( .A(n11417), .ZN(P2_U3196) );
  AOI21_X1 U13898 ( .B1(n14489), .B2(n14124), .A(n11418), .ZN(n11419) );
  OAI211_X1 U13899 ( .C1(n14583), .C2(n11421), .A(n11420), .B(n11419), .ZN(
        n11423) );
  NAND2_X1 U13900 ( .A1(n11423), .A2(n14654), .ZN(n11422) );
  OAI21_X1 U13901 ( .B1(n14654), .B2(n7682), .A(n11422), .ZN(P1_U3539) );
  INV_X1 U13902 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11425) );
  NAND2_X1 U13903 ( .A1(n11423), .A2(n14641), .ZN(n11424) );
  OAI21_X1 U13904 ( .B1(n14641), .B2(n11425), .A(n11424), .ZN(P1_U3492) );
  INV_X1 U13905 ( .A(n11426), .ZN(n11428) );
  NAND2_X1 U13906 ( .A1(n11428), .A2(n11427), .ZN(n11429) );
  XNOR2_X1 U13907 ( .A(n11431), .B(n6637), .ZN(n11432) );
  AND2_X1 U13908 ( .A1(n13116), .A2(n13295), .ZN(n11433) );
  NAND2_X1 U13909 ( .A1(n11432), .A2(n11433), .ZN(n11558) );
  INV_X1 U13910 ( .A(n11432), .ZN(n11435) );
  INV_X1 U13911 ( .A(n11433), .ZN(n11434) );
  NAND2_X1 U13912 ( .A1(n11435), .A2(n11434), .ZN(n11436) );
  NAND2_X1 U13913 ( .A1(n11558), .A2(n11436), .ZN(n11438) );
  AOI21_X1 U13914 ( .B1(n11437), .B2(n11438), .A(n13091), .ZN(n11441) );
  INV_X1 U13915 ( .A(n11437), .ZN(n11440) );
  NAND2_X1 U13916 ( .A1(n11441), .A2(n11559), .ZN(n11447) );
  NOR2_X1 U13917 ( .A1(n11442), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14691) );
  NOR2_X1 U13918 ( .A1(n13087), .A2(n11443), .ZN(n11444) );
  AOI211_X1 U13919 ( .C1(n13085), .C2(n11445), .A(n14691), .B(n11444), .ZN(
        n11446) );
  OAI211_X1 U13920 ( .C1(n14435), .C2(n13071), .A(n11447), .B(n11446), .ZN(
        P2_U3206) );
  INV_X1 U13921 ( .A(n11448), .ZN(n11449) );
  AOI21_X1 U13922 ( .B1(n11451), .B2(n11450), .A(n11449), .ZN(n14513) );
  INV_X1 U13923 ( .A(n14513), .ZN(n11462) );
  AOI22_X1 U13924 ( .A1(n14507), .A2(n14049), .B1(n14041), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n11461) );
  XNOR2_X1 U13925 ( .A(n11452), .B(n7738), .ZN(n11453) );
  NAND2_X1 U13926 ( .A1(n11453), .A2(n14028), .ZN(n11455) );
  AOI22_X1 U13927 ( .A1(n13709), .A2(n14008), .B1(n14006), .B2(n13711), .ZN(
        n11454) );
  NAND2_X1 U13928 ( .A1(n11455), .A2(n11454), .ZN(n14512) );
  INV_X1 U13929 ( .A(n11456), .ZN(n11514) );
  NAND2_X1 U13930 ( .A1(n14507), .A2(n11457), .ZN(n11458) );
  NAND2_X1 U13931 ( .A1(n11514), .A2(n11458), .ZN(n14510) );
  OAI22_X1 U13932 ( .A1(n14510), .A2(n14013), .B1(n14461), .B2(n14011), .ZN(
        n11459) );
  OAI21_X1 U13933 ( .B1(n14512), .B2(n11459), .A(n14047), .ZN(n11460) );
  OAI211_X1 U13934 ( .C1(n11462), .C2(n14019), .A(n11461), .B(n11460), .ZN(
        P1_U3279) );
  INV_X1 U13935 ( .A(n11464), .ZN(n11465) );
  NAND2_X1 U13936 ( .A1(n11463), .A2(n11465), .ZN(n11466) );
  OAI22_X1 U13937 ( .A1(n14635), .A2(n12161), .B1(n14476), .B2(n12062), .ZN(
        n11468) );
  XNOR2_X1 U13938 ( .A(n11468), .B(n12158), .ZN(n11632) );
  AND2_X1 U13939 ( .A1(n13714), .A2(n12152), .ZN(n11469) );
  AOI21_X1 U13940 ( .B1(n11757), .B2(n12132), .A(n11469), .ZN(n11630) );
  XNOR2_X1 U13941 ( .A(n11632), .B(n11630), .ZN(n11470) );
  OAI211_X1 U13942 ( .C1(n6682), .C2(n11470), .A(n14482), .B(n14483), .ZN(
        n11478) );
  INV_X1 U13943 ( .A(n11472), .ZN(n11476) );
  NAND2_X1 U13944 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n13795)
         );
  NAND2_X1 U13945 ( .A1(n13681), .A2(n13713), .ZN(n11473) );
  OAI211_X1 U13946 ( .C1(n14477), .C2(n11474), .A(n13795), .B(n11473), .ZN(
        n11475) );
  AOI21_X1 U13947 ( .B1(n11476), .B2(n13695), .A(n11475), .ZN(n11477) );
  OAI211_X1 U13948 ( .C1(n14635), .C2(n13699), .A(n11478), .B(n11477), .ZN(
        P1_U3217) );
  OAI21_X1 U13949 ( .B1(n13655), .B2(n14634), .A(n11479), .ZN(n11481) );
  AOI211_X1 U13950 ( .C1(n14638), .C2(n11482), .A(n11481), .B(n11480), .ZN(
        n11485) );
  OR2_X1 U13951 ( .A1(n11485), .A2(n14651), .ZN(n11483) );
  OAI21_X1 U13952 ( .B1(n14654), .B2(n11484), .A(n11483), .ZN(P1_U3541) );
  INV_X1 U13953 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11487) );
  OR2_X1 U13954 ( .A1(n11485), .A2(n14639), .ZN(n11486) );
  OAI21_X1 U13955 ( .B1(n14641), .B2(n11487), .A(n11486), .ZN(P1_U3498) );
  INV_X1 U13956 ( .A(n11488), .ZN(n11490) );
  INV_X1 U13957 ( .A(SI_27_), .ZN(n15218) );
  OAI222_X1 U13958 ( .A1(P3_U3151), .A2(n12586), .B1(n12967), .B2(n11490), 
        .C1(n15218), .C2(n11489), .ZN(P3_U3268) );
  XNOR2_X1 U13959 ( .A(n11492), .B(n6982), .ZN(n11494) );
  AOI22_X1 U13960 ( .A1(n12544), .A2(n12827), .B1(n12829), .B2(n12828), .ZN(
        n12234) );
  INV_X1 U13961 ( .A(n12234), .ZN(n11493) );
  AOI21_X1 U13962 ( .B1(n11494), .B2(n12832), .A(n11493), .ZN(n14378) );
  INV_X1 U13963 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12559) );
  INV_X1 U13964 ( .A(n12237), .ZN(n11495) );
  OAI22_X1 U13965 ( .A1(n15045), .A2(n12559), .B1(n11495), .B2(n15032), .ZN(
        n11496) );
  AOI21_X1 U13966 ( .B1(n12837), .B2(n11497), .A(n11496), .ZN(n11500) );
  XNOR2_X1 U13967 ( .A(n11498), .B(n6982), .ZN(n14381) );
  NAND2_X1 U13968 ( .A1(n14381), .A2(n12841), .ZN(n11499) );
  OAI211_X1 U13969 ( .C1(n14378), .C2(n12844), .A(n11500), .B(n11499), .ZN(
        P3_U3221) );
  XNOR2_X1 U13970 ( .A(n11501), .B(n12454), .ZN(n14373) );
  XNOR2_X1 U13971 ( .A(n11502), .B(n12454), .ZN(n11503) );
  OAI222_X1 U13972 ( .A1(n15040), .A2(n12325), .B1(n15042), .B2(n11504), .C1(
        n11503), .C2(n15038), .ZN(n14374) );
  INV_X1 U13973 ( .A(n14376), .ZN(n11506) );
  AOI22_X1 U13974 ( .A1(n12844), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12805), 
        .B2(n12024), .ZN(n11505) );
  OAI21_X1 U13975 ( .B1(n11506), .B2(n12807), .A(n11505), .ZN(n11507) );
  AOI21_X1 U13976 ( .B1(n14374), .B2(n15045), .A(n11507), .ZN(n11508) );
  OAI21_X1 U13977 ( .B1(n12791), .B2(n14373), .A(n11508), .ZN(P3_U3220) );
  INV_X1 U13978 ( .A(n11509), .ZN(n11510) );
  AOI21_X1 U13979 ( .B1(n11512), .B2(n11511), .A(n11510), .ZN(n11585) );
  INV_X1 U13980 ( .A(n11513), .ZN(n11591) );
  AOI211_X1 U13981 ( .C1(n12047), .C2(n11514), .A(n14509), .B(n11591), .ZN(
        n11581) );
  INV_X1 U13982 ( .A(n12047), .ZN(n13700) );
  INV_X1 U13983 ( .A(n11515), .ZN(n13696) );
  AOI22_X1 U13984 ( .A1(n14041), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13696), 
        .B2(n14051), .ZN(n11516) );
  OAI21_X1 U13985 ( .B1(n13700), .B2(n14035), .A(n11516), .ZN(n11517) );
  AOI21_X1 U13986 ( .B1(n11581), .B2(n13999), .A(n11517), .ZN(n11524) );
  XNOR2_X1 U13987 ( .A(n11518), .B(n11910), .ZN(n11519) );
  NAND2_X1 U13988 ( .A1(n11519), .A2(n14028), .ZN(n11583) );
  INV_X1 U13989 ( .A(n11583), .ZN(n11522) );
  NAND2_X1 U13990 ( .A1(n13710), .A2(n14006), .ZN(n11521) );
  NAND2_X1 U13991 ( .A1(n13708), .A2(n14008), .ZN(n11520) );
  AND2_X1 U13992 ( .A1(n11521), .A2(n11520), .ZN(n13693) );
  INV_X1 U13993 ( .A(n13693), .ZN(n11582) );
  OAI21_X1 U13994 ( .B1(n11522), .B2(n11582), .A(n14047), .ZN(n11523) );
  OAI211_X1 U13995 ( .C1(n11585), .C2(n14019), .A(n11524), .B(n11523), .ZN(
        P1_U3278) );
  INV_X1 U13996 ( .A(n13838), .ZN(n14573) );
  INV_X1 U13997 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U13998 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13670)
         );
  OAI21_X1 U13999 ( .B1(n14566), .B2(n11525), .A(n13670), .ZN(n11543) );
  INV_X1 U14000 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11541) );
  OR2_X1 U14001 ( .A1(n11526), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14002 ( .A1(n11528), .A2(n11527), .ZN(n11531) );
  XNOR2_X1 U14003 ( .A(n11531), .B(n14574), .ZN(n14572) );
  NAND2_X1 U14004 ( .A1(n14572), .A2(n7758), .ZN(n14571) );
  INV_X1 U14005 ( .A(n14571), .ZN(n11529) );
  AOI21_X1 U14006 ( .B1(n11531), .B2(n11530), .A(n11529), .ZN(n13814) );
  INV_X1 U14007 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14008 ( .A1(n11534), .A2(n11533), .ZN(n11532) );
  OAI21_X1 U14009 ( .B1(n11534), .B2(n11533), .A(n11532), .ZN(n13813) );
  NAND2_X1 U14010 ( .A1(n13814), .A2(n13813), .ZN(n13812) );
  NAND2_X1 U14011 ( .A1(n11534), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14012 ( .A1(n13812), .A2(n11535), .ZN(n13826) );
  INV_X1 U14013 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14500) );
  MUX2_X1 U14014 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14500), .S(n11545), .Z(
        n13825) );
  NAND2_X1 U14015 ( .A1(n13826), .A2(n13825), .ZN(n13824) );
  NAND2_X1 U14016 ( .A1(n11545), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U14017 ( .A1(n13824), .A2(n11536), .ZN(n11537) );
  AND2_X1 U14018 ( .A1(n11537), .A2(n13833), .ZN(n13830) );
  NOR2_X1 U14019 ( .A1(n11537), .A2(n13833), .ZN(n11538) );
  NOR2_X1 U14020 ( .A1(n11540), .A2(n11541), .ZN(n13831) );
  AOI211_X1 U14021 ( .C1(n11541), .C2(n11540), .A(n11539), .B(n13831), .ZN(
        n11542) );
  AOI211_X1 U14022 ( .C1(n14573), .C2(n13833), .A(n11543), .B(n11542), .ZN(
        n11557) );
  NAND2_X1 U14023 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n11545), .ZN(n11553) );
  INV_X1 U14024 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14025 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n11545), .B1(n13821), 
        .B2(n11544), .ZN(n13819) );
  INV_X1 U14026 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U14027 ( .B1(n11548), .B2(n11547), .A(n11546), .ZN(n11549) );
  NOR2_X1 U14028 ( .A1(n14574), .A2(n11549), .ZN(n11550) );
  XNOR2_X1 U14029 ( .A(n11549), .B(n14574), .ZN(n14569) );
  NOR2_X1 U14030 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14569), .ZN(n14568) );
  NOR2_X1 U14031 ( .A1(n11550), .A2(n14568), .ZN(n13808) );
  NAND2_X1 U14032 ( .A1(n13809), .A2(n11552), .ZN(n11551) );
  OAI211_X1 U14033 ( .C1(n13809), .C2(n11552), .A(n13808), .B(n11551), .ZN(
        n13806) );
  OAI21_X1 U14034 ( .B1(n11552), .B2(n13809), .A(n13806), .ZN(n13820) );
  NAND2_X1 U14035 ( .A1(n13819), .A2(n13820), .ZN(n13818) );
  NAND2_X1 U14036 ( .A1(n11553), .A2(n13818), .ZN(n13834) );
  XNOR2_X1 U14037 ( .A(n13834), .B(n11554), .ZN(n11555) );
  NAND2_X1 U14038 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11555), .ZN(n13836) );
  OAI211_X1 U14039 ( .C1(n11555), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14560), 
        .B(n13836), .ZN(n11556) );
  NAND2_X1 U14040 ( .A1(n11557), .A2(n11556), .ZN(P1_U3261) );
  INV_X1 U14041 ( .A(n14412), .ZN(n14429) );
  XNOR2_X1 U14042 ( .A(n14412), .B(n6637), .ZN(n11957) );
  NAND2_X1 U14043 ( .A1(n13115), .A2(n13295), .ZN(n11958) );
  XNOR2_X1 U14044 ( .A(n11957), .B(n11958), .ZN(n11560) );
  OAI21_X1 U14045 ( .B1(n11561), .B2(n11560), .A(n11961), .ZN(n11562) );
  NAND2_X1 U14046 ( .A1(n11562), .A2(n13060), .ZN(n11569) );
  INV_X1 U14047 ( .A(n11563), .ZN(n14401) );
  NAND2_X1 U14048 ( .A1(n13114), .A2(n13065), .ZN(n11565) );
  NAND2_X1 U14049 ( .A1(n13116), .A2(n13064), .ZN(n11564) );
  AND2_X1 U14050 ( .A1(n11565), .A2(n11564), .ZN(n14397) );
  OAI22_X1 U14051 ( .A1(n13066), .A2(n14397), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11566), .ZN(n11567) );
  AOI21_X1 U14052 ( .B1(n14401), .B2(n13068), .A(n11567), .ZN(n11568) );
  OAI211_X1 U14053 ( .C1(n14429), .C2(n13071), .A(n11569), .B(n11568), .ZN(
        P2_U3187) );
  AOI22_X1 U14054 ( .A1(n12544), .A2(n12315), .B1(n12025), .B2(n12546), .ZN(
        n11571) );
  OAI211_X1 U14055 ( .C1(n14856), .C2(n11572), .A(n11571), .B(n11570), .ZN(
        n11578) );
  INV_X1 U14056 ( .A(n11573), .ZN(n11574) );
  AOI211_X1 U14057 ( .C1(n11576), .C2(n11575), .A(n12310), .B(n11574), .ZN(
        n11577) );
  AOI211_X1 U14058 ( .C1(n11579), .C2(n12326), .A(n11578), .B(n11577), .ZN(
        n11580) );
  INV_X1 U14059 ( .A(n11580), .ZN(P3_U3157) );
  AOI211_X1 U14060 ( .C1(n12047), .C2(n14124), .A(n11582), .B(n11581), .ZN(
        n11584) );
  OAI211_X1 U14061 ( .C1(n11585), .C2(n14583), .A(n11584), .B(n11583), .ZN(
        n11587) );
  NAND2_X1 U14062 ( .A1(n11587), .A2(n14654), .ZN(n11586) );
  OAI21_X1 U14063 ( .B1(n14654), .B2(n7758), .A(n11586), .ZN(P1_U3543) );
  INV_X1 U14064 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U14065 ( .A1(n11587), .A2(n14641), .ZN(n11588) );
  OAI21_X1 U14066 ( .B1(n14641), .B2(n11589), .A(n11588), .ZN(P1_U3504) );
  XNOR2_X1 U14067 ( .A(n11590), .B(n11594), .ZN(n14506) );
  INV_X1 U14068 ( .A(n14506), .ZN(n11603) );
  OAI22_X1 U14069 ( .A1(n14047), .A2(n11552), .B1(n14475), .B2(n14011), .ZN(
        n11593) );
  INV_X1 U14070 ( .A(n14472), .ZN(n14503) );
  OAI211_X1 U14071 ( .C1(n11591), .C2(n14503), .A(n14126), .B(n11655), .ZN(
        n14502) );
  NOR2_X1 U14072 ( .A1(n14502), .A2(n13948), .ZN(n11592) );
  AOI211_X1 U14073 ( .C1(n14049), .C2(n14472), .A(n11593), .B(n11592), .ZN(
        n11602) );
  NAND2_X1 U14074 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  AOI21_X1 U14075 ( .B1(n11597), .B2(n11596), .A(n14584), .ZN(n14505) );
  NAND2_X1 U14076 ( .A1(n13707), .A2(n14008), .ZN(n11599) );
  NAND2_X1 U14077 ( .A1(n13709), .A2(n14006), .ZN(n11598) );
  AND2_X1 U14078 ( .A1(n11599), .A2(n11598), .ZN(n14501) );
  INV_X1 U14079 ( .A(n14501), .ZN(n11600) );
  OAI21_X1 U14080 ( .B1(n14505), .B2(n11600), .A(n14047), .ZN(n11601) );
  OAI211_X1 U14081 ( .C1(n11603), .C2(n14019), .A(n11602), .B(n11601), .ZN(
        P1_U3277) );
  INV_X1 U14082 ( .A(n11604), .ZN(n13019) );
  OAI211_X1 U14083 ( .C1(n6616), .C2(n8585), .A(n14399), .B(n11665), .ZN(
        n11605) );
  AOI22_X1 U14084 ( .A1(n13112), .A2(n13065), .B1(n13064), .B2(n13114), .ZN(
        n13017) );
  NAND2_X1 U14085 ( .A1(n11605), .A2(n13017), .ZN(n13486) );
  AOI21_X1 U14086 ( .B1(n13019), .B2(n14402), .A(n13486), .ZN(n11610) );
  AOI211_X1 U14087 ( .C1(n13488), .C2(n11620), .A(n13295), .B(n11670), .ZN(
        n13487) );
  INV_X1 U14088 ( .A(n13488), .ZN(n13022) );
  OAI22_X1 U14089 ( .A1(n13022), .A2(n13406), .B1(n8394), .B2(n13336), .ZN(
        n11606) );
  AOI21_X1 U14090 ( .B1(n13487), .B2(n13402), .A(n11606), .ZN(n11609) );
  NAND2_X1 U14091 ( .A1(n11607), .A2(n8585), .ZN(n13489) );
  NAND3_X1 U14092 ( .A1(n13490), .A2(n13489), .A3(n14417), .ZN(n11608) );
  OAI211_X1 U14093 ( .C1(n11610), .C2(n14420), .A(n11609), .B(n11608), .ZN(
        P2_U3249) );
  OAI21_X1 U14094 ( .B1(n11612), .B2(n8384), .A(n11611), .ZN(n14427) );
  INV_X1 U14095 ( .A(n14427), .ZN(n11625) );
  XNOR2_X1 U14096 ( .A(n11614), .B(n11613), .ZN(n11615) );
  NOR2_X1 U14097 ( .A1(n11615), .A2(n13393), .ZN(n14425) );
  NAND2_X1 U14098 ( .A1(n13113), .A2(n13065), .ZN(n11617) );
  NAND2_X1 U14099 ( .A1(n13115), .A2(n13064), .ZN(n11616) );
  NAND2_X1 U14100 ( .A1(n11617), .A2(n11616), .ZN(n14421) );
  OAI21_X1 U14101 ( .B1(n14425), .B2(n14421), .A(n13336), .ZN(n11624) );
  OAI22_X1 U14102 ( .A1(n13336), .A2(n11618), .B1(n13088), .B2(n13300), .ZN(
        n11622) );
  INV_X1 U14103 ( .A(n13096), .ZN(n14424) );
  OAI211_X1 U14104 ( .C1(n14424), .C2(n11619), .A(n12001), .B(n11620), .ZN(
        n14423) );
  NOR2_X1 U14105 ( .A1(n14423), .A2(n14415), .ZN(n11621) );
  AOI211_X1 U14106 ( .C1(n14403), .C2(n13096), .A(n11622), .B(n11621), .ZN(
        n11623) );
  OAI211_X1 U14107 ( .C1(n11625), .C2(n13372), .A(n11624), .B(n11623), .ZN(
        P2_U3250) );
  NAND2_X1 U14108 ( .A1(n14489), .A2(n12147), .ZN(n11627) );
  NAND2_X1 U14109 ( .A1(n13713), .A2(n12132), .ZN(n11626) );
  NAND2_X1 U14110 ( .A1(n11627), .A2(n11626), .ZN(n11628) );
  XNOR2_X1 U14111 ( .A(n11628), .B(n12158), .ZN(n11634) );
  AND2_X1 U14112 ( .A1(n13713), .A2(n12152), .ZN(n11629) );
  AOI21_X1 U14113 ( .B1(n14489), .B2(n12132), .A(n11629), .ZN(n11635) );
  XNOR2_X1 U14114 ( .A(n11634), .B(n11635), .ZN(n14480) );
  INV_X1 U14115 ( .A(n11630), .ZN(n11631) );
  NAND2_X1 U14116 ( .A1(n11632), .A2(n11631), .ZN(n14481) );
  AND2_X1 U14117 ( .A1(n14480), .A2(n14481), .ZN(n11633) );
  INV_X1 U14118 ( .A(n11634), .ZN(n11636) );
  NAND2_X1 U14119 ( .A1(n11768), .A2(n12147), .ZN(n11638) );
  NAND2_X1 U14120 ( .A1(n13712), .A2(n12132), .ZN(n11637) );
  NAND2_X1 U14121 ( .A1(n11638), .A2(n11637), .ZN(n11639) );
  XNOR2_X1 U14122 ( .A(n11639), .B(n12158), .ZN(n12033) );
  AND2_X1 U14123 ( .A1(n13712), .A2(n12152), .ZN(n11640) );
  AOI21_X1 U14124 ( .B1(n11768), .B2(n12132), .A(n11640), .ZN(n12034) );
  XNOR2_X1 U14125 ( .A(n12033), .B(n12034), .ZN(n11641) );
  OAI211_X1 U14126 ( .C1(n11642), .C2(n11641), .A(n12037), .B(n14483), .ZN(
        n11647) );
  NAND2_X1 U14127 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14564)
         );
  NAND2_X1 U14128 ( .A1(n13673), .A2(n13713), .ZN(n11643) );
  OAI211_X1 U14129 ( .C1(n14478), .C2(n14452), .A(n14564), .B(n11643), .ZN(
        n11644) );
  AOI21_X1 U14130 ( .B1(n11645), .B2(n13695), .A(n11644), .ZN(n11646) );
  OAI211_X1 U14131 ( .C1(n6896), .C2(n13699), .A(n11647), .B(n11646), .ZN(
        P1_U3224) );
  NAND2_X1 U14132 ( .A1(n11648), .A2(n7236), .ZN(n11649) );
  NAND3_X1 U14133 ( .A1(n11650), .A2(n14028), .A3(n11649), .ZN(n11652) );
  AOI22_X1 U14134 ( .A1(n14007), .A2(n14008), .B1(n14006), .B2(n13708), .ZN(
        n11651) );
  NAND2_X1 U14135 ( .A1(n11652), .A2(n11651), .ZN(n14498) );
  INV_X1 U14136 ( .A(n14498), .ZN(n11660) );
  NAND2_X1 U14137 ( .A1(n11654), .A2(n11911), .ZN(n14495) );
  NAND3_X1 U14138 ( .A1(n11653), .A2(n14495), .A3(n13951), .ZN(n11659) );
  OAI22_X1 U14139 ( .A1(n14047), .A2(n11544), .B1(n13621), .B2(n14011), .ZN(
        n11657) );
  OAI211_X1 U14140 ( .C1(n6891), .C2(n6890), .A(n14126), .B(n14031), .ZN(
        n14496) );
  NOR2_X1 U14141 ( .A1(n14496), .A2(n13948), .ZN(n11656) );
  AOI211_X1 U14142 ( .C1(n14049), .C2(n13623), .A(n11657), .B(n11656), .ZN(
        n11658) );
  OAI211_X1 U14143 ( .C1(n14041), .C2(n11660), .A(n11659), .B(n11658), .ZN(
        P1_U3276) );
  OAI21_X1 U14144 ( .B1(n11662), .B2(n11664), .A(n11661), .ZN(n13484) );
  NAND3_X1 U14145 ( .A1(n11665), .A2(n11664), .A3(n11663), .ZN(n11666) );
  NAND3_X1 U14146 ( .A1(n11667), .A2(n14399), .A3(n11666), .ZN(n11669) );
  AND2_X1 U14147 ( .A1(n13113), .A2(n13064), .ZN(n11668) );
  AOI21_X1 U14148 ( .B1(n13111), .B2(n13065), .A(n11668), .ZN(n13028) );
  NAND2_X1 U14149 ( .A1(n11669), .A2(n13028), .ZN(n13480) );
  INV_X1 U14150 ( .A(n13399), .ZN(n11671) );
  AOI211_X1 U14151 ( .C1(n13482), .C2(n6938), .A(n13295), .B(n11671), .ZN(
        n13481) );
  NAND2_X1 U14152 ( .A1(n13481), .A2(n13402), .ZN(n11674) );
  INV_X1 U14153 ( .A(n11672), .ZN(n13030) );
  AOI22_X1 U14154 ( .A1(n13411), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13030), 
        .B2(n14402), .ZN(n11673) );
  OAI211_X1 U14155 ( .C1(n13033), .C2(n13406), .A(n11674), .B(n11673), .ZN(
        n11675) );
  AOI21_X1 U14156 ( .B1(n13336), .B2(n13480), .A(n11675), .ZN(n11676) );
  OAI21_X1 U14157 ( .B1(n13372), .B2(n13484), .A(n11676), .ZN(P2_U3248) );
  MUX2_X1 U14158 ( .A(n11677), .B(P3_REG2_REG_0__SCAN_IN), .S(n12844), .Z(
        n11680) );
  INV_X1 U14159 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14872) );
  OAI22_X1 U14160 ( .A1(n12807), .A2(n11678), .B1(n15032), .B2(n14872), .ZN(
        n11679) );
  OR2_X1 U14161 ( .A1(n11680), .A2(n11679), .ZN(P3_U3233) );
  INV_X1 U14162 ( .A(n11681), .ZN(n11683) );
  OAI222_X1 U14163 ( .A1(n12967), .A2(n11683), .B1(n12968), .B2(n15221), .C1(
        P3_U3151), .C2(n11682), .ZN(P3_U3270) );
  INV_X1 U14164 ( .A(n11684), .ZN(n13545) );
  INV_X1 U14165 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11685) );
  OAI222_X1 U14166 ( .A1(n8098), .A2(P1_U3086), .B1(n14166), .B2(n13545), .C1(
        n11685), .C2(n14163), .ZN(P1_U3327) );
  INV_X1 U14167 ( .A(n11686), .ZN(n11712) );
  NAND2_X1 U14168 ( .A1(n11688), .A2(n11687), .ZN(n11690) );
  NAND2_X1 U14169 ( .A1(n11690), .A2(n11689), .ZN(n11692) );
  NAND2_X1 U14170 ( .A1(n11692), .A2(n11691), .ZN(n11858) );
  NAND2_X1 U14171 ( .A1(n11858), .A2(n11693), .ZN(n11738) );
  INV_X2 U14172 ( .A(n11839), .ZN(n11842) );
  MUX2_X1 U14173 ( .A(n6478), .B(n6646), .S(n11842), .Z(n11711) );
  NAND2_X1 U14174 ( .A1(n11890), .A2(n9930), .ZN(n11695) );
  NAND2_X1 U14175 ( .A1(n13723), .A2(n11694), .ZN(n11889) );
  NAND2_X1 U14176 ( .A1(n11695), .A2(n11889), .ZN(n11697) );
  INV_X4 U14177 ( .A(n11839), .ZN(n11878) );
  OAI211_X1 U14178 ( .C1(n11697), .C2(n11878), .A(n11893), .B(n11696), .ZN(
        n11703) );
  NAND2_X1 U14179 ( .A1(n13722), .A2(n11860), .ZN(n11698) );
  NOR2_X1 U14180 ( .A1(n11698), .A2(n11700), .ZN(n11699) );
  AOI21_X1 U14181 ( .B1(n11701), .B2(n11700), .A(n11699), .ZN(n11702) );
  NAND2_X1 U14182 ( .A1(n11703), .A2(n11702), .ZN(n11707) );
  MUX2_X1 U14183 ( .A(n13721), .B(n7516), .S(n11839), .Z(n11704) );
  INV_X1 U14184 ( .A(n11704), .ZN(n11705) );
  NAND3_X1 U14185 ( .A1(n11707), .A2(n13721), .A3(n7516), .ZN(n11708) );
  NAND3_X1 U14186 ( .A1(n11709), .A2(n11708), .A3(n11892), .ZN(n11710) );
  OAI21_X1 U14187 ( .B1(n11712), .B2(n11711), .A(n11710), .ZN(n11718) );
  MUX2_X1 U14188 ( .A(n11714), .B(n11713), .S(n11842), .Z(n11717) );
  MUX2_X1 U14189 ( .A(n13720), .B(n11715), .S(n11839), .Z(n11716) );
  NAND2_X1 U14190 ( .A1(n11718), .A2(n11717), .ZN(n11719) );
  MUX2_X1 U14191 ( .A(n13719), .B(n11721), .S(n11839), .Z(n11723) );
  MUX2_X1 U14192 ( .A(n13719), .B(n11721), .S(n11842), .Z(n11722) );
  INV_X1 U14193 ( .A(n11723), .ZN(n11724) );
  MUX2_X1 U14194 ( .A(n13718), .B(n11725), .S(n11878), .Z(n11729) );
  NAND2_X1 U14195 ( .A1(n11728), .A2(n11729), .ZN(n11727) );
  MUX2_X1 U14196 ( .A(n13718), .B(n11725), .S(n11839), .Z(n11726) );
  NAND2_X1 U14197 ( .A1(n11727), .A2(n11726), .ZN(n11733) );
  INV_X1 U14198 ( .A(n11728), .ZN(n11731) );
  INV_X1 U14199 ( .A(n11729), .ZN(n11730) );
  NAND2_X1 U14200 ( .A1(n11731), .A2(n11730), .ZN(n11732) );
  MUX2_X1 U14201 ( .A(n13717), .B(n11734), .S(n11839), .Z(n11736) );
  MUX2_X1 U14202 ( .A(n13717), .B(n11734), .S(n11842), .Z(n11735) );
  INV_X1 U14203 ( .A(n11736), .ZN(n11737) );
  MUX2_X1 U14204 ( .A(n13716), .B(n11739), .S(n11842), .Z(n11743) );
  NAND2_X1 U14205 ( .A1(n11742), .A2(n11743), .ZN(n11741) );
  MUX2_X1 U14206 ( .A(n13716), .B(n11739), .S(n11860), .Z(n11740) );
  NAND2_X1 U14207 ( .A1(n11741), .A2(n11740), .ZN(n11747) );
  INV_X1 U14208 ( .A(n11742), .ZN(n11745) );
  INV_X1 U14209 ( .A(n11743), .ZN(n11744) );
  NAND2_X1 U14210 ( .A1(n11745), .A2(n11744), .ZN(n11746) );
  NAND2_X1 U14211 ( .A1(n11747), .A2(n11746), .ZN(n11751) );
  MUX2_X1 U14212 ( .A(n13715), .B(n11748), .S(n11860), .Z(n11752) );
  NAND2_X1 U14213 ( .A1(n11751), .A2(n11752), .ZN(n11750) );
  MUX2_X1 U14214 ( .A(n13715), .B(n11748), .S(n11878), .Z(n11749) );
  NAND2_X1 U14215 ( .A1(n11750), .A2(n11749), .ZN(n11756) );
  INV_X1 U14216 ( .A(n11751), .ZN(n11754) );
  INV_X1 U14217 ( .A(n11752), .ZN(n11753) );
  NAND2_X1 U14218 ( .A1(n11754), .A2(n11753), .ZN(n11755) );
  MUX2_X1 U14219 ( .A(n13714), .B(n11757), .S(n11842), .Z(n11759) );
  MUX2_X1 U14220 ( .A(n13714), .B(n11757), .S(n11860), .Z(n11758) );
  MUX2_X1 U14221 ( .A(n13713), .B(n14489), .S(n11860), .Z(n11763) );
  NAND2_X1 U14222 ( .A1(n11762), .A2(n11763), .ZN(n11761) );
  MUX2_X1 U14223 ( .A(n13713), .B(n14489), .S(n11842), .Z(n11760) );
  NAND2_X1 U14224 ( .A1(n11761), .A2(n11760), .ZN(n11767) );
  INV_X1 U14225 ( .A(n11762), .ZN(n11765) );
  INV_X1 U14226 ( .A(n11763), .ZN(n11764) );
  NAND2_X1 U14227 ( .A1(n11765), .A2(n11764), .ZN(n11766) );
  NAND2_X1 U14228 ( .A1(n11767), .A2(n11766), .ZN(n11772) );
  MUX2_X1 U14229 ( .A(n13712), .B(n11768), .S(n11878), .Z(n11771) );
  NAND2_X1 U14230 ( .A1(n11772), .A2(n11771), .ZN(n11770) );
  MUX2_X1 U14231 ( .A(n13712), .B(n11768), .S(n11860), .Z(n11769) );
  MUX2_X1 U14233 ( .A(n13711), .B(n12040), .S(n11860), .Z(n11779) );
  NOR2_X1 U14234 ( .A1(n12040), .A2(n11860), .ZN(n11777) );
  NOR2_X1 U14235 ( .A1(n13711), .A2(n11878), .ZN(n11780) );
  OR3_X1 U14236 ( .A1(n11779), .A2(n11777), .A3(n11780), .ZN(n11776) );
  AND2_X1 U14237 ( .A1(n11785), .A2(n11775), .ZN(n11778) );
  AOI22_X1 U14238 ( .A1(n7738), .A2(n11878), .B1(n11777), .B2(n11779), .ZN(
        n11788) );
  INV_X1 U14239 ( .A(n11778), .ZN(n11787) );
  INV_X1 U14240 ( .A(n11781), .ZN(n11782) );
  MUX2_X1 U14241 ( .A(n11785), .B(n11784), .S(n11878), .Z(n11786) );
  MUX2_X1 U14242 ( .A(n13708), .B(n14472), .S(n11860), .Z(n11790) );
  MUX2_X1 U14243 ( .A(n14007), .B(n14125), .S(n11842), .Z(n11795) );
  NAND2_X1 U14244 ( .A1(n11795), .A2(n11789), .ZN(n11794) );
  NAND2_X1 U14245 ( .A1(n11791), .A2(n11790), .ZN(n11793) );
  MUX2_X1 U14246 ( .A(n13708), .B(n14472), .S(n11842), .Z(n11792) );
  INV_X1 U14247 ( .A(n11795), .ZN(n11802) );
  AND2_X1 U14248 ( .A1(n13707), .A2(n11842), .ZN(n11797) );
  NOR2_X1 U14249 ( .A1(n13707), .A2(n11878), .ZN(n11796) );
  MUX2_X1 U14250 ( .A(n11797), .B(n11796), .S(n13623), .Z(n11799) );
  OR2_X1 U14251 ( .A1(n11798), .A2(n11799), .ZN(n11801) );
  AOI22_X1 U14252 ( .A1(n11802), .A2(n11801), .B1(n11800), .B2(n11799), .ZN(
        n11803) );
  MUX2_X1 U14253 ( .A(n13984), .B(n14119), .S(n11860), .Z(n11804) );
  OR2_X1 U14254 ( .A1(n13994), .A2(n11804), .ZN(n11805) );
  MUX2_X1 U14255 ( .A(n13598), .B(n13991), .S(n11860), .Z(n11807) );
  MUX2_X1 U14256 ( .A(n14009), .B(n14115), .S(n11878), .Z(n11806) );
  OAI21_X1 U14257 ( .B1(n11808), .B2(n11807), .A(n11806), .ZN(n11810) );
  NAND2_X1 U14258 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  MUX2_X1 U14259 ( .A(n13656), .B(n13971), .S(n11839), .Z(n11812) );
  MUX2_X1 U14260 ( .A(n13983), .B(n14109), .S(n11842), .Z(n11811) );
  MUX2_X1 U14261 ( .A(n14104), .B(n13706), .S(n11842), .Z(n11814) );
  MUX2_X1 U14262 ( .A(n13597), .B(n13957), .S(n11878), .Z(n11813) );
  MUX2_X1 U14263 ( .A(n13657), .B(n13943), .S(n11860), .Z(n11815) );
  MUX2_X1 U14264 ( .A(n13657), .B(n13943), .S(n11842), .Z(n11816) );
  MUX2_X1 U14265 ( .A(n13704), .B(n13928), .S(n11860), .Z(n11820) );
  NAND2_X1 U14266 ( .A1(n11819), .A2(n11820), .ZN(n11818) );
  MUX2_X1 U14267 ( .A(n13704), .B(n13928), .S(n11878), .Z(n11817) );
  NAND2_X1 U14268 ( .A1(n11818), .A2(n11817), .ZN(n11824) );
  INV_X1 U14269 ( .A(n11819), .ZN(n11822) );
  INV_X1 U14270 ( .A(n11820), .ZN(n11821) );
  NAND2_X1 U14271 ( .A1(n11822), .A2(n11821), .ZN(n11823) );
  NAND2_X1 U14272 ( .A1(n11824), .A2(n11823), .ZN(n11826) );
  MUX2_X1 U14273 ( .A(n13886), .B(n14084), .S(n11842), .Z(n11827) );
  MUX2_X1 U14274 ( .A(n13886), .B(n14084), .S(n11860), .Z(n11825) );
  MUX2_X1 U14275 ( .A(n13703), .B(n14079), .S(n11839), .Z(n11829) );
  MUX2_X1 U14276 ( .A(n13703), .B(n14079), .S(n11842), .Z(n11828) );
  INV_X1 U14277 ( .A(n11829), .ZN(n11830) );
  MUX2_X1 U14278 ( .A(n13887), .B(n14075), .S(n11878), .Z(n11834) );
  NAND2_X1 U14279 ( .A1(n11833), .A2(n11834), .ZN(n11832) );
  MUX2_X1 U14280 ( .A(n13887), .B(n14075), .S(n11839), .Z(n11831) );
  NAND2_X1 U14281 ( .A1(n11832), .A2(n11831), .ZN(n11838) );
  INV_X1 U14282 ( .A(n11833), .ZN(n11836) );
  INV_X1 U14283 ( .A(n11834), .ZN(n11835) );
  NAND2_X1 U14284 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  MUX2_X1 U14285 ( .A(n13702), .B(n14070), .S(n11878), .Z(n11840) );
  MUX2_X1 U14286 ( .A(n13862), .B(n14065), .S(n11842), .Z(n11844) );
  NAND2_X1 U14287 ( .A1(n11843), .A2(n11844), .ZN(n11848) );
  MUX2_X1 U14288 ( .A(n14065), .B(n13862), .S(n11878), .Z(n11847) );
  INV_X1 U14289 ( .A(n11843), .ZN(n11846) );
  INV_X1 U14290 ( .A(n11844), .ZN(n11845) );
  NAND2_X1 U14291 ( .A1(n11953), .A2(n7965), .ZN(n11850) );
  NAND2_X1 U14292 ( .A1(n8000), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11849) );
  INV_X1 U14293 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11851) );
  OR2_X1 U14294 ( .A1(n7561), .A2(n11851), .ZN(n11857) );
  INV_X1 U14295 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13849) );
  OR2_X1 U14296 ( .A1(n11852), .A2(n13849), .ZN(n11856) );
  INV_X1 U14297 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11853) );
  OR2_X1 U14298 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  OAI21_X1 U14299 ( .B1(n11877), .B2(n11860), .A(n11858), .ZN(n11859) );
  AOI22_X1 U14300 ( .A1(n11919), .A2(n11860), .B1(n13701), .B2(n11859), .ZN(
        n11864) );
  NAND2_X1 U14301 ( .A1(n11863), .A2(n11864), .ZN(n11868) );
  INV_X1 U14302 ( .A(n11877), .ZN(n13851) );
  OAI21_X1 U14303 ( .B1(n11861), .B2(n13851), .A(n13701), .ZN(n11862) );
  MUX2_X1 U14304 ( .A(n11862), .B(n14060), .S(n11878), .Z(n11867) );
  INV_X1 U14305 ( .A(n11863), .ZN(n11866) );
  INV_X1 U14306 ( .A(n11864), .ZN(n11865) );
  AOI22_X1 U14307 ( .A1(n11868), .A2(n11867), .B1(n11866), .B2(n11865), .ZN(
        n11887) );
  INV_X1 U14308 ( .A(n11887), .ZN(n11876) );
  NAND2_X1 U14309 ( .A1(n13536), .A2(n7965), .ZN(n11870) );
  NAND2_X1 U14310 ( .A1(n8000), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11869) );
  XNOR2_X1 U14311 ( .A(n14055), .B(n11877), .ZN(n11888) );
  NAND2_X1 U14312 ( .A1(n11872), .A2(n11871), .ZN(n11873) );
  AND2_X1 U14313 ( .A1(n11874), .A2(n11873), .ZN(n11883) );
  INV_X1 U14314 ( .A(n11883), .ZN(n11875) );
  NAND2_X1 U14315 ( .A1(n11876), .A2(n7440), .ZN(n11930) );
  NOR2_X1 U14316 ( .A1(n14055), .A2(n11877), .ZN(n11880) );
  AND2_X1 U14317 ( .A1(n14055), .A2(n11877), .ZN(n11879) );
  MUX2_X1 U14318 ( .A(n11880), .B(n11879), .S(n11878), .Z(n11881) );
  INV_X1 U14319 ( .A(n11881), .ZN(n11884) );
  NAND3_X1 U14320 ( .A1(n11884), .A2(n11883), .A3(n11888), .ZN(n11882) );
  OAI211_X1 U14321 ( .C1(n11884), .C2(n11883), .A(n11882), .B(n11925), .ZN(
        n11885) );
  AOI21_X1 U14322 ( .B1(n11887), .B2(n11886), .A(n11885), .ZN(n11929) );
  INV_X1 U14323 ( .A(n11888), .ZN(n11923) );
  AND2_X1 U14324 ( .A1(n11890), .A2(n11889), .ZN(n14582) );
  NAND4_X1 U14325 ( .A1(n14582), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11896) );
  NOR3_X1 U14326 ( .A1(n11896), .A2(n11895), .A3(n11894), .ZN(n11899) );
  NAND4_X1 U14327 ( .A1(n11898), .A2(n11899), .A3(n11900), .A4(n11897), .ZN(
        n11901) );
  NOR4_X1 U14328 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11907) );
  NAND4_X1 U14329 ( .A1(n11908), .A2(n11907), .A3(n11906), .A4(n11905), .ZN(
        n11909) );
  NOR3_X1 U14330 ( .A1(n11910), .A2(n7738), .A3(n11909), .ZN(n11912) );
  NAND4_X1 U14331 ( .A1(n14024), .A2(n11912), .A3(n14005), .A4(n11911), .ZN(
        n11913) );
  NOR4_X1 U14332 ( .A1(n13959), .A2(n13976), .A3(n11914), .A4(n11913), .ZN(
        n11915) );
  NAND4_X1 U14333 ( .A1(n13898), .A2(n11915), .A3(n13914), .A4(n13938), .ZN(
        n11916) );
  NOR4_X1 U14334 ( .A1(n13873), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11922) );
  XOR2_X1 U14335 ( .A(n14062), .B(n11919), .Z(n11921) );
  NAND4_X1 U14336 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n11924) );
  XOR2_X1 U14337 ( .A(n13843), .B(n11924), .Z(n11927) );
  INV_X1 U14338 ( .A(n11925), .ZN(n11926) );
  AOI21_X1 U14339 ( .B1(n11930), .B2(n11929), .A(n11928), .ZN(n11935) );
  NOR3_X1 U14340 ( .A1(n11931), .A2(n14157), .A3(n14021), .ZN(n11933) );
  OAI21_X1 U14341 ( .B1(n11934), .B2(n14168), .A(P1_B_REG_SCAN_IN), .ZN(n11932) );
  OAI22_X1 U14342 ( .A1(n11935), .A2(n11934), .B1(n11933), .B2(n11932), .ZN(
        P1_U3242) );
  OAI222_X1 U14343 ( .A1(n8056), .A2(P1_U3086), .B1(n14166), .B2(n11937), .C1(
        n11936), .C2(n14163), .ZN(P1_U3335) );
  AOI21_X1 U14344 ( .B1(n11942), .B2(n11939), .A(n11938), .ZN(n14078) );
  OAI21_X1 U14345 ( .B1(n11942), .B2(n11941), .A(n11940), .ZN(n11944) );
  OAI22_X1 U14346 ( .A1(n13603), .A2(n14021), .B1(n12160), .B2(n14045), .ZN(
        n11943) );
  INV_X1 U14347 ( .A(n13867), .ZN(n11947) );
  AOI211_X1 U14348 ( .C1(n14075), .C2(n13880), .A(n14509), .B(n11947), .ZN(
        n14074) );
  INV_X1 U14349 ( .A(n11948), .ZN(n13567) );
  AOI22_X1 U14350 ( .A1(n14041), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13567), 
        .B2(n14051), .ZN(n11949) );
  OAI21_X1 U14351 ( .B1(n13569), .B2(n14035), .A(n11949), .ZN(n11951) );
  NOR2_X1 U14352 ( .A1(n14078), .A2(n14037), .ZN(n11950) );
  AOI211_X1 U14353 ( .C1(n14074), .C2(n13999), .A(n11951), .B(n11950), .ZN(
        n11952) );
  OAI21_X1 U14354 ( .B1(n14077), .B2(n14041), .A(n11952), .ZN(P1_U3266) );
  INV_X1 U14355 ( .A(n11953), .ZN(n12172) );
  INV_X1 U14356 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12332) );
  OAI222_X1 U14357 ( .A1(P1_U3086), .A2(n7468), .B1(n14166), .B2(n12172), .C1(
        n12332), .C2(n14163), .ZN(P1_U3325) );
  INV_X1 U14358 ( .A(n11954), .ZN(n11955) );
  OAI222_X1 U14359 ( .A1(n12968), .A2(n15184), .B1(P3_U3151), .B2(n11956), 
        .C1(n12191), .C2(n11955), .ZN(P3_U3267) );
  XNOR2_X1 U14360 ( .A(n13477), .B(n6637), .ZN(n11973) );
  NAND2_X1 U14361 ( .A1(n13111), .A2(n13295), .ZN(n11974) );
  XNOR2_X1 U14362 ( .A(n13482), .B(n11975), .ZN(n11972) );
  NAND2_X1 U14363 ( .A1(n13112), .A2(n13295), .ZN(n11971) );
  INV_X1 U14364 ( .A(n11957), .ZN(n11959) );
  NAND2_X1 U14365 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  XOR2_X1 U14366 ( .A(n6637), .B(n13096), .Z(n11963) );
  NAND2_X1 U14367 ( .A1(n13114), .A2(n13295), .ZN(n13092) );
  INV_X1 U14368 ( .A(n11962), .ZN(n11965) );
  INV_X1 U14369 ( .A(n11963), .ZN(n11964) );
  NOR2_X1 U14370 ( .A1(n11966), .A2(n10263), .ZN(n11968) );
  XNOR2_X1 U14371 ( .A(n13488), .B(n6637), .ZN(n11967) );
  XOR2_X1 U14372 ( .A(n11968), .B(n11967), .Z(n13013) );
  INV_X1 U14373 ( .A(n11967), .ZN(n11970) );
  INV_X1 U14374 ( .A(n11968), .ZN(n11969) );
  NAND2_X1 U14375 ( .A1(n11970), .A2(n11969), .ZN(n13023) );
  XNOR2_X1 U14376 ( .A(n11972), .B(n11971), .ZN(n13024) );
  XNOR2_X1 U14377 ( .A(n11973), .B(n11974), .ZN(n13062) );
  XNOR2_X1 U14378 ( .A(n13383), .B(n11975), .ZN(n11977) );
  NAND2_X1 U14379 ( .A1(n13110), .A2(n13295), .ZN(n11976) );
  NAND2_X1 U14380 ( .A1(n11977), .A2(n11976), .ZN(n12986) );
  NOR2_X1 U14381 ( .A1(n11977), .A2(n11976), .ZN(n12988) );
  AND2_X1 U14382 ( .A1(n13109), .A2(n13295), .ZN(n11979) );
  XNOR2_X1 U14383 ( .A(n13465), .B(n6637), .ZN(n11978) );
  NOR2_X1 U14384 ( .A1(n11978), .A2(n11979), .ZN(n11980) );
  AOI21_X1 U14385 ( .B1(n11979), .B2(n11978), .A(n11980), .ZN(n13044) );
  INV_X1 U14386 ( .A(n11980), .ZN(n11981) );
  NAND2_X1 U14387 ( .A1(n13108), .A2(n13295), .ZN(n11983) );
  XNOR2_X1 U14388 ( .A(n13348), .B(n6637), .ZN(n11982) );
  XOR2_X1 U14389 ( .A(n11983), .B(n11982), .Z(n12995) );
  XNOR2_X1 U14390 ( .A(n13332), .B(n6637), .ZN(n11985) );
  INV_X1 U14391 ( .A(n11985), .ZN(n11984) );
  NOR2_X1 U14392 ( .A1(n12981), .A2(n12001), .ZN(n13053) );
  XNOR2_X1 U14393 ( .A(n13313), .B(n6637), .ZN(n11990) );
  XNOR2_X1 U14394 ( .A(n11989), .B(n11990), .ZN(n12978) );
  NOR2_X1 U14395 ( .A1(n11988), .A2(n12001), .ZN(n12979) );
  NAND2_X1 U14396 ( .A1(n12978), .A2(n12979), .ZN(n11993) );
  INV_X1 U14397 ( .A(n11989), .ZN(n11991) );
  XNOR2_X1 U14398 ( .A(n13441), .B(n6637), .ZN(n11995) );
  NAND2_X1 U14399 ( .A1(n13105), .A2(n13295), .ZN(n11994) );
  XNOR2_X1 U14400 ( .A(n11995), .B(n11994), .ZN(n13034) );
  INV_X1 U14401 ( .A(n11994), .ZN(n11996) );
  XNOR2_X1 U14402 ( .A(n13010), .B(n6637), .ZN(n11997) );
  NOR2_X1 U14403 ( .A1(n13079), .A2(n12001), .ZN(n11998) );
  XNOR2_X1 U14404 ( .A(n11997), .B(n11998), .ZN(n13003) );
  INV_X1 U14405 ( .A(n11997), .ZN(n12000) );
  INV_X1 U14406 ( .A(n11998), .ZN(n11999) );
  XNOR2_X1 U14407 ( .A(n13507), .B(n6637), .ZN(n12003) );
  OR2_X1 U14408 ( .A1(n13005), .A2(n12001), .ZN(n12002) );
  NAND2_X1 U14409 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  OAI21_X1 U14410 ( .B1(n12003), .B2(n12002), .A(n12004), .ZN(n13074) );
  XNOR2_X1 U14411 ( .A(n13424), .B(n6637), .ZN(n12005) );
  NOR2_X1 U14412 ( .A1(n13077), .A2(n12001), .ZN(n12006) );
  XNOR2_X1 U14413 ( .A(n12005), .B(n12006), .ZN(n12969) );
  INV_X1 U14414 ( .A(n12005), .ZN(n12008) );
  INV_X1 U14415 ( .A(n12006), .ZN(n12007) );
  NOR2_X1 U14416 ( .A1(n12971), .A2(n12001), .ZN(n12010) );
  XNOR2_X1 U14417 ( .A(n12010), .B(n6637), .ZN(n12011) );
  XNOR2_X1 U14418 ( .A(n13502), .B(n12011), .ZN(n12012) );
  OR2_X1 U14419 ( .A1(n12013), .A2(n13076), .ZN(n12015) );
  OR2_X1 U14420 ( .A1(n13077), .A2(n13078), .ZN(n12014) );
  NAND2_X1 U14421 ( .A1(n12015), .A2(n12014), .ZN(n13237) );
  AOI22_X1 U14422 ( .A1(n13085), .A2(n13237), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12016) );
  OAI21_X1 U14423 ( .B1(n13240), .B2(n13087), .A(n12016), .ZN(n12017) );
  AOI21_X1 U14424 ( .B1(n12018), .B2(n13095), .A(n12017), .ZN(n12019) );
  OAI21_X1 U14425 ( .B1(n12020), .B2(n13091), .A(n12019), .ZN(P2_U3192) );
  XNOR2_X1 U14426 ( .A(n12022), .B(n12828), .ZN(n12023) );
  XNOR2_X1 U14427 ( .A(n12021), .B(n12023), .ZN(n12030) );
  NAND2_X1 U14428 ( .A1(n12326), .A2(n12024), .ZN(n12027) );
  AOI22_X1 U14429 ( .A1(n12025), .A2(n12543), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12026) );
  OAI211_X1 U14430 ( .C1(n12325), .C2(n12276), .A(n12027), .B(n12026), .ZN(
        n12028) );
  AOI21_X1 U14431 ( .B1(n14376), .B2(n14847), .A(n12028), .ZN(n12029) );
  OAI21_X1 U14432 ( .B1(n12030), .B2(n12310), .A(n12029), .ZN(P3_U3174) );
  OAI222_X1 U14433 ( .A1(n12967), .A2(n12031), .B1(n12968), .B2(n15160), .C1(
        P3_U3151), .C2(n6490), .ZN(P3_U3276) );
  AOI22_X1 U14434 ( .A1(n14507), .A2(n12147), .B1(n12148), .B2(n13710), .ZN(
        n12032) );
  XNOR2_X1 U14435 ( .A(n12032), .B(n12158), .ZN(n12046) );
  AOI22_X1 U14436 ( .A1(n14507), .A2(n12132), .B1(n12152), .B2(n13710), .ZN(
        n12045) );
  NAND2_X1 U14437 ( .A1(n12033), .A2(n12035), .ZN(n12036) );
  NAND2_X1 U14438 ( .A1(n12037), .A2(n12036), .ZN(n13647) );
  OAI22_X1 U14439 ( .A1(n13655), .A2(n12161), .B1(n14452), .B2(n12062), .ZN(
        n12038) );
  XNOR2_X1 U14440 ( .A(n12038), .B(n12158), .ZN(n12041) );
  AND2_X1 U14441 ( .A1(n13711), .A2(n12152), .ZN(n12039) );
  AOI21_X1 U14442 ( .B1(n12040), .B2(n12132), .A(n12039), .ZN(n12042) );
  XNOR2_X1 U14443 ( .A(n12041), .B(n12042), .ZN(n13646) );
  INV_X1 U14444 ( .A(n12042), .ZN(n12043) );
  NAND2_X1 U14445 ( .A1(n12041), .A2(n12043), .ZN(n12044) );
  XNOR2_X1 U14446 ( .A(n12046), .B(n12045), .ZN(n14453) );
  NAND2_X1 U14447 ( .A1(n12047), .A2(n12147), .ZN(n12049) );
  NAND2_X1 U14448 ( .A1(n13709), .A2(n12148), .ZN(n12048) );
  NAND2_X1 U14449 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  XNOR2_X1 U14450 ( .A(n12050), .B(n12158), .ZN(n12051) );
  OAI22_X1 U14451 ( .A1(n13700), .A2(n12062), .B1(n14462), .B2(n10334), .ZN(
        n13689) );
  NAND2_X1 U14452 ( .A1(n13690), .A2(n13689), .ZN(n13687) );
  INV_X1 U14453 ( .A(n12051), .ZN(n12052) );
  NOR2_X1 U14454 ( .A1(n12053), .A2(n12052), .ZN(n14465) );
  NAND2_X1 U14455 ( .A1(n14472), .A2(n12147), .ZN(n12055) );
  NAND2_X1 U14456 ( .A1(n13708), .A2(n12148), .ZN(n12054) );
  NAND2_X1 U14457 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  XNOR2_X1 U14458 ( .A(n12056), .B(n6648), .ZN(n12060) );
  AND2_X1 U14459 ( .A1(n13708), .A2(n12152), .ZN(n12057) );
  AOI21_X1 U14460 ( .B1(n14472), .B2(n12132), .A(n12057), .ZN(n12059) );
  XNOR2_X1 U14461 ( .A(n12060), .B(n12059), .ZN(n14464) );
  NOR2_X1 U14462 ( .A1(n14465), .A2(n14464), .ZN(n12058) );
  NAND2_X1 U14463 ( .A1(n12060), .A2(n12059), .ZN(n12061) );
  NAND2_X1 U14464 ( .A1(n13623), .A2(n12147), .ZN(n12064) );
  NAND2_X1 U14465 ( .A1(n13707), .A2(n12132), .ZN(n12063) );
  NAND2_X1 U14466 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  XNOR2_X1 U14467 ( .A(n12065), .B(n12158), .ZN(n12068) );
  NAND2_X1 U14468 ( .A1(n13623), .A2(n12132), .ZN(n12067) );
  NAND2_X1 U14469 ( .A1(n13707), .A2(n12152), .ZN(n12066) );
  NAND2_X1 U14470 ( .A1(n12067), .A2(n12066), .ZN(n12069) );
  NAND2_X1 U14471 ( .A1(n12068), .A2(n12069), .ZN(n13616) );
  INV_X1 U14472 ( .A(n12068), .ZN(n12071) );
  INV_X1 U14473 ( .A(n12069), .ZN(n12070) );
  NAND2_X1 U14474 ( .A1(n12071), .A2(n12070), .ZN(n13617) );
  NAND2_X1 U14475 ( .A1(n14125), .A2(n12147), .ZN(n12073) );
  NAND2_X1 U14476 ( .A1(n14007), .A2(n12132), .ZN(n12072) );
  NAND2_X1 U14477 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  XNOR2_X1 U14478 ( .A(n12074), .B(n12158), .ZN(n12081) );
  AOI22_X1 U14479 ( .A1(n14125), .A2(n12132), .B1(n12152), .B2(n14007), .ZN(
        n12079) );
  XNOR2_X1 U14480 ( .A(n12081), .B(n12079), .ZN(n13668) );
  NAND2_X1 U14481 ( .A1(n14119), .A2(n12147), .ZN(n12076) );
  NAND2_X1 U14482 ( .A1(n13984), .A2(n12132), .ZN(n12075) );
  NAND2_X1 U14483 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  XNOR2_X1 U14484 ( .A(n12077), .B(n6648), .ZN(n12083) );
  AND2_X1 U14485 ( .A1(n13984), .A2(n12152), .ZN(n12078) );
  AOI21_X1 U14486 ( .B1(n14119), .B2(n12132), .A(n12078), .ZN(n12084) );
  XNOR2_X1 U14487 ( .A(n12083), .B(n12084), .ZN(n13584) );
  INV_X1 U14488 ( .A(n12079), .ZN(n12080) );
  NOR2_X1 U14489 ( .A1(n12081), .A2(n12080), .ZN(n13585) );
  NOR2_X1 U14490 ( .A1(n13584), .A2(n13585), .ZN(n12082) );
  NAND2_X1 U14491 ( .A1(n13583), .A2(n12082), .ZN(n13587) );
  INV_X1 U14492 ( .A(n12083), .ZN(n12086) );
  INV_X1 U14493 ( .A(n12084), .ZN(n12085) );
  NAND2_X1 U14494 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  NAND2_X1 U14495 ( .A1(n13587), .A2(n12087), .ZN(n13637) );
  OAI22_X1 U14496 ( .A1(n13991), .A2(n12062), .B1(n13598), .B2(n10334), .ZN(
        n12089) );
  OAI22_X1 U14497 ( .A1(n13991), .A2(n12161), .B1(n13598), .B2(n12062), .ZN(
        n12088) );
  XNOR2_X1 U14498 ( .A(n12088), .B(n12158), .ZN(n12090) );
  XOR2_X1 U14499 ( .A(n12089), .B(n12090), .Z(n13638) );
  NAND2_X1 U14500 ( .A1(n12090), .A2(n12089), .ZN(n12091) );
  OAI22_X1 U14501 ( .A1(n13971), .A2(n12161), .B1(n13656), .B2(n12062), .ZN(
        n12092) );
  XNOR2_X1 U14502 ( .A(n12092), .B(n6648), .ZN(n12096) );
  OR2_X1 U14503 ( .A1(n13971), .A2(n12109), .ZN(n12094) );
  NAND2_X1 U14504 ( .A1(n13983), .A2(n12152), .ZN(n12093) );
  AND2_X1 U14505 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  NAND2_X1 U14506 ( .A1(n12096), .A2(n12095), .ZN(n13662) );
  OAI21_X1 U14507 ( .B1(n12096), .B2(n12095), .A(n13662), .ZN(n13595) );
  NAND2_X1 U14508 ( .A1(n13593), .A2(n13662), .ZN(n12107) );
  NAND2_X1 U14509 ( .A1(n14104), .A2(n12147), .ZN(n12099) );
  NAND2_X1 U14510 ( .A1(n13706), .A2(n12132), .ZN(n12098) );
  NAND2_X1 U14511 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  XNOR2_X1 U14512 ( .A(n12100), .B(n6648), .ZN(n12102) );
  AND2_X1 U14513 ( .A1(n13706), .A2(n12152), .ZN(n12101) );
  AOI21_X1 U14514 ( .B1(n14104), .B2(n12132), .A(n12101), .ZN(n12103) );
  NAND2_X1 U14515 ( .A1(n12102), .A2(n12103), .ZN(n13570) );
  INV_X1 U14516 ( .A(n12102), .ZN(n12105) );
  INV_X1 U14517 ( .A(n12103), .ZN(n12104) );
  NAND2_X1 U14518 ( .A1(n12105), .A2(n12104), .ZN(n12106) );
  AND2_X1 U14519 ( .A1(n13570), .A2(n12106), .ZN(n13660) );
  NAND2_X1 U14520 ( .A1(n12107), .A2(n13660), .ZN(n13573) );
  NAND2_X1 U14521 ( .A1(n13573), .A2(n13570), .ZN(n12117) );
  OAI22_X1 U14522 ( .A1(n13943), .A2(n12161), .B1(n13657), .B2(n12062), .ZN(
        n12108) );
  XNOR2_X1 U14523 ( .A(n12108), .B(n6648), .ZN(n12112) );
  OR2_X1 U14524 ( .A1(n13943), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U14525 ( .A1(n13705), .A2(n12152), .ZN(n12110) );
  AND2_X1 U14526 ( .A1(n12111), .A2(n12110), .ZN(n12113) );
  NAND2_X1 U14527 ( .A1(n12112), .A2(n12113), .ZN(n13626) );
  INV_X1 U14528 ( .A(n12112), .ZN(n12115) );
  INV_X1 U14529 ( .A(n12113), .ZN(n12114) );
  NAND2_X1 U14530 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  NAND2_X1 U14531 ( .A1(n13928), .A2(n12147), .ZN(n12119) );
  NAND2_X1 U14532 ( .A1(n13704), .A2(n12132), .ZN(n12118) );
  NAND2_X1 U14533 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  XNOR2_X1 U14534 ( .A(n12120), .B(n6648), .ZN(n12122) );
  AND2_X1 U14535 ( .A1(n13704), .A2(n12152), .ZN(n12121) );
  AOI21_X1 U14536 ( .B1(n13928), .B2(n12132), .A(n12121), .ZN(n12123) );
  NAND2_X1 U14537 ( .A1(n12122), .A2(n12123), .ZN(n13609) );
  INV_X1 U14538 ( .A(n12122), .ZN(n12125) );
  INV_X1 U14539 ( .A(n12123), .ZN(n12124) );
  NAND2_X1 U14540 ( .A1(n12125), .A2(n12124), .ZN(n12126) );
  NAND2_X1 U14541 ( .A1(n14084), .A2(n12147), .ZN(n12128) );
  NAND2_X1 U14542 ( .A1(n13886), .A2(n12148), .ZN(n12127) );
  NAND2_X1 U14543 ( .A1(n12128), .A2(n12127), .ZN(n12130) );
  XNOR2_X1 U14544 ( .A(n12130), .B(n6648), .ZN(n12133) );
  AND2_X1 U14545 ( .A1(n13886), .A2(n12152), .ZN(n12131) );
  AOI21_X1 U14546 ( .B1(n14084), .B2(n12132), .A(n12131), .ZN(n12134) );
  NAND2_X1 U14547 ( .A1(n12133), .A2(n12134), .ZN(n12138) );
  INV_X1 U14548 ( .A(n12133), .ZN(n12136) );
  INV_X1 U14549 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U14550 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  AND2_X1 U14551 ( .A1(n12138), .A2(n12137), .ZN(n13607) );
  NAND2_X1 U14552 ( .A1(n14079), .A2(n12147), .ZN(n12140) );
  NAND2_X1 U14553 ( .A1(n13703), .A2(n12132), .ZN(n12139) );
  NAND2_X1 U14554 ( .A1(n12140), .A2(n12139), .ZN(n12141) );
  XNOR2_X1 U14555 ( .A(n12141), .B(n12158), .ZN(n12145) );
  NAND2_X1 U14556 ( .A1(n14079), .A2(n12148), .ZN(n12143) );
  NAND2_X1 U14557 ( .A1(n13703), .A2(n12152), .ZN(n12142) );
  NAND2_X1 U14558 ( .A1(n12143), .A2(n12142), .ZN(n12144) );
  NOR2_X1 U14559 ( .A1(n12145), .A2(n12144), .ZN(n12146) );
  AOI21_X1 U14560 ( .B1(n12145), .B2(n12144), .A(n12146), .ZN(n13678) );
  NAND2_X1 U14561 ( .A1(n14075), .A2(n12147), .ZN(n12150) );
  NAND2_X1 U14562 ( .A1(n13887), .A2(n12148), .ZN(n12149) );
  NAND2_X1 U14563 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  XNOR2_X1 U14564 ( .A(n12151), .B(n12158), .ZN(n12156) );
  NAND2_X1 U14565 ( .A1(n14075), .A2(n12148), .ZN(n12154) );
  NAND2_X1 U14566 ( .A1(n13887), .A2(n12152), .ZN(n12153) );
  NAND2_X1 U14567 ( .A1(n12154), .A2(n12153), .ZN(n12155) );
  NOR2_X1 U14568 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  AOI21_X1 U14569 ( .B1(n12156), .B2(n12155), .A(n12157), .ZN(n13563) );
  OAI22_X1 U14570 ( .A1(n12162), .A2(n12062), .B1(n12160), .B2(n10334), .ZN(
        n12159) );
  XNOR2_X1 U14571 ( .A(n12159), .B(n12158), .ZN(n12164) );
  OAI22_X1 U14572 ( .A1(n12162), .A2(n12161), .B1(n12160), .B2(n12062), .ZN(
        n12163) );
  XNOR2_X1 U14573 ( .A(n12164), .B(n12163), .ZN(n12165) );
  XNOR2_X1 U14574 ( .A(n12166), .B(n12165), .ZN(n12171) );
  AOI22_X1 U14575 ( .A1(n13673), .A2(n13887), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12168) );
  NAND2_X1 U14576 ( .A1(n13681), .A2(n13862), .ZN(n12167) );
  OAI211_X1 U14577 ( .C1(n14494), .C2(n13871), .A(n12168), .B(n12167), .ZN(
        n12169) );
  AOI21_X1 U14578 ( .B1(n14070), .B2(n14490), .A(n12169), .ZN(n12170) );
  OAI21_X1 U14579 ( .B1(n12171), .B2(n14467), .A(n12170), .ZN(P1_U3220) );
  OAI222_X1 U14580 ( .A1(n13552), .A2(n12172), .B1(P2_U3088), .B2(n8159), .C1(
        n12189), .C2(n13550), .ZN(P2_U3297) );
  INV_X1 U14581 ( .A(n12173), .ZN(n12175) );
  AND2_X1 U14582 ( .A1(n12174), .A2(n12175), .ZN(n12177) );
  XOR2_X1 U14583 ( .A(n9675), .B(n12511), .Z(n12178) );
  XNOR2_X1 U14584 ( .A(n12179), .B(n12178), .ZN(n12185) );
  INV_X1 U14585 ( .A(n12180), .ZN(n12644) );
  AOI22_X1 U14586 ( .A1(n12181), .A2(n14865), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12182) );
  OAI21_X1 U14587 ( .B1(n12644), .B2(n14867), .A(n12182), .ZN(n12183) );
  AOI21_X1 U14588 ( .B1(n12647), .B2(n14847), .A(n12183), .ZN(n12184) );
  OAI21_X1 U14589 ( .B1(n12185), .B2(n12310), .A(n12184), .ZN(P3_U3160) );
  NAND2_X1 U14590 ( .A1(n14152), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12188) );
  XNOR2_X1 U14591 ( .A(n12189), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12333) );
  XNOR2_X1 U14592 ( .A(n12334), .B(n12333), .ZN(n12339) );
  INV_X1 U14593 ( .A(n12339), .ZN(n12190) );
  OAI222_X1 U14594 ( .A1(n12192), .A2(P3_U3151), .B1(n12968), .B2(n15215), 
        .C1(n12191), .C2(n12190), .ZN(P3_U3265) );
  OR2_X1 U14595 ( .A1(n12021), .A2(n12193), .ZN(n12196) );
  NAND2_X1 U14596 ( .A1(n12196), .A2(n12194), .ZN(n12198) );
  AND2_X1 U14597 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  AOI21_X1 U14598 ( .B1(n12199), .B2(n12198), .A(n12197), .ZN(n12205) );
  NAND2_X1 U14599 ( .A1(n12830), .A2(n12315), .ZN(n12200) );
  NAND2_X1 U14600 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15016)
         );
  OAI211_X1 U14601 ( .C1(n12201), .C2(n12317), .A(n12200), .B(n15016), .ZN(
        n12203) );
  NOR2_X1 U14602 ( .A1(n14369), .A2(n14856), .ZN(n12202) );
  AOI211_X1 U14603 ( .C1(n12833), .C2(n12326), .A(n12203), .B(n12202), .ZN(
        n12204) );
  OAI21_X1 U14604 ( .B1(n12205), .B2(n12310), .A(n12204), .ZN(P3_U3155) );
  AOI21_X1 U14605 ( .B1(n12537), .B2(n12206), .A(n6518), .ZN(n12212) );
  NOR2_X1 U14606 ( .A1(n12729), .A2(n12317), .ZN(n12209) );
  INV_X1 U14607 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12207) );
  OAI22_X1 U14608 ( .A1(n12708), .A2(n12276), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12207), .ZN(n12208) );
  AOI211_X1 U14609 ( .C1(n12709), .C2(n12326), .A(n12209), .B(n12208), .ZN(
        n12211) );
  NAND2_X1 U14610 ( .A1(n12395), .A2(n14847), .ZN(n12210) );
  OAI211_X1 U14611 ( .C1(n12212), .C2(n12310), .A(n12211), .B(n12210), .ZN(
        P3_U3156) );
  XNOR2_X1 U14612 ( .A(n12214), .B(n12213), .ZN(n12219) );
  AOI22_X1 U14613 ( .A1(n12540), .A2(n12827), .B1(n12829), .B2(n12539), .ZN(
        n12756) );
  OAI22_X1 U14614 ( .A1(n12756), .A2(n14851), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15251), .ZN(n12217) );
  INV_X1 U14615 ( .A(n12215), .ZN(n12943) );
  NOR2_X1 U14616 ( .A1(n12943), .A2(n14856), .ZN(n12216) );
  AOI211_X1 U14617 ( .C1(n12759), .C2(n12326), .A(n12217), .B(n12216), .ZN(
        n12218) );
  OAI21_X1 U14618 ( .B1(n12219), .B2(n12310), .A(n12218), .ZN(P3_U3159) );
  INV_X1 U14619 ( .A(n12220), .ZN(n12221) );
  AOI21_X1 U14620 ( .B1(n12223), .B2(n12222), .A(n12221), .ZN(n12228) );
  NAND2_X1 U14621 ( .A1(n12326), .A2(n12732), .ZN(n12225) );
  AOI22_X1 U14622 ( .A1(n12315), .A2(n12538), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12224) );
  OAI211_X1 U14623 ( .C1(n12730), .C2(n12317), .A(n12225), .B(n12224), .ZN(
        n12226) );
  AOI21_X1 U14624 ( .B1(n12731), .B2(n14847), .A(n12226), .ZN(n12227) );
  OAI21_X1 U14625 ( .B1(n12228), .B2(n12310), .A(n12227), .ZN(P3_U3163) );
  XNOR2_X1 U14626 ( .A(n12230), .B(n12229), .ZN(n12291) );
  OAI22_X1 U14627 ( .A1(n12291), .A2(n12544), .B1(n12230), .B2(n12229), .ZN(
        n12233) );
  XNOR2_X1 U14628 ( .A(n12231), .B(n12543), .ZN(n12232) );
  XNOR2_X1 U14629 ( .A(n12233), .B(n12232), .ZN(n12239) );
  NOR2_X1 U14630 ( .A1(n14379), .A2(n14856), .ZN(n12236) );
  INV_X1 U14631 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n14978) );
  OAI22_X1 U14632 ( .A1(n12234), .A2(n14851), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14978), .ZN(n12235) );
  AOI211_X1 U14633 ( .C1(n12237), .C2(n12326), .A(n12236), .B(n12235), .ZN(
        n12238) );
  OAI21_X1 U14634 ( .B1(n12239), .B2(n12310), .A(n12238), .ZN(P3_U3164) );
  AND3_X1 U14635 ( .A1(n12240), .A2(n12242), .A3(n12241), .ZN(n12243) );
  OAI21_X1 U14636 ( .B1(n12244), .B2(n12243), .A(n14857), .ZN(n12248) );
  AOI22_X1 U14637 ( .A1(n12315), .A2(n12678), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12245) );
  OAI21_X1 U14638 ( .B1(n12708), .B2(n12317), .A(n12245), .ZN(n12246) );
  AOI21_X1 U14639 ( .B1(n12687), .B2(n12326), .A(n12246), .ZN(n12247) );
  OAI211_X1 U14640 ( .C1(n12919), .C2(n14856), .A(n12248), .B(n12247), .ZN(
        P3_U3165) );
  AOI21_X1 U14641 ( .B1(n12250), .B2(n12249), .A(n12310), .ZN(n12252) );
  NAND2_X1 U14642 ( .A1(n12252), .A2(n12251), .ZN(n12257) );
  AOI22_X1 U14643 ( .A1(n12315), .A2(n12796), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12253) );
  OAI21_X1 U14644 ( .B1(n12254), .B2(n12317), .A(n12253), .ZN(n12255) );
  AOI21_X1 U14645 ( .B1(n12804), .B2(n12326), .A(n12255), .ZN(n12256) );
  OAI211_X1 U14646 ( .C1(n12953), .C2(n14856), .A(n12257), .B(n12256), .ZN(
        P3_U3166) );
  NAND2_X1 U14647 ( .A1(n12259), .A2(n12258), .ZN(n12300) );
  OAI211_X1 U14648 ( .C1(n12259), .C2(n12258), .A(n12300), .B(n14857), .ZN(
        n12263) );
  AOI22_X1 U14649 ( .A1(n12540), .A2(n12797), .B1(n12827), .B2(n12541), .ZN(
        n12785) );
  OAI22_X1 U14650 ( .A1(n12785), .A2(n14851), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12260), .ZN(n12261) );
  AOI21_X1 U14651 ( .B1(n12787), .B2(n12326), .A(n12261), .ZN(n12262) );
  OAI211_X1 U14652 ( .C1(n14856), .C2(n12948), .A(n12263), .B(n12262), .ZN(
        P3_U3168) );
  INV_X1 U14653 ( .A(n12264), .ZN(n12266) );
  NOR3_X1 U14654 ( .A1(n6518), .A2(n12266), .A3(n12265), .ZN(n12268) );
  INV_X1 U14655 ( .A(n12240), .ZN(n12267) );
  OAI21_X1 U14656 ( .B1(n12268), .B2(n12267), .A(n14857), .ZN(n12272) );
  AOI22_X1 U14657 ( .A1(n12536), .A2(n12829), .B1(n12827), .B2(n12537), .ZN(
        n12694) );
  INV_X1 U14658 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12269) );
  OAI22_X1 U14659 ( .A1(n12694), .A2(n14851), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12269), .ZN(n12270) );
  AOI21_X1 U14660 ( .B1(n12699), .B2(n12326), .A(n12270), .ZN(n12271) );
  OAI211_X1 U14661 ( .C1(n12923), .C2(n14856), .A(n12272), .B(n12271), .ZN(
        P3_U3169) );
  XNOR2_X1 U14662 ( .A(n12273), .B(n12274), .ZN(n12282) );
  NOR2_X1 U14663 ( .A1(n12275), .A2(n12317), .ZN(n12279) );
  OAI22_X1 U14664 ( .A1(n12277), .A2(n12276), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15270), .ZN(n12278) );
  AOI211_X1 U14665 ( .C1(n12747), .C2(n12326), .A(n12279), .B(n12278), .ZN(
        n12281) );
  NAND2_X1 U14666 ( .A1(n12486), .A2(n14847), .ZN(n12280) );
  OAI211_X1 U14667 ( .C1(n12282), .C2(n12310), .A(n12281), .B(n12280), .ZN(
        P3_U3173) );
  INV_X1 U14668 ( .A(n12284), .ZN(n12285) );
  AOI21_X1 U14669 ( .B1(n12538), .B2(n12283), .A(n12285), .ZN(n12289) );
  AOI22_X1 U14670 ( .A1(n12744), .A2(n12827), .B1(n12829), .B2(n12537), .ZN(
        n12718) );
  OAI22_X1 U14671 ( .A1(n12718), .A2(n14851), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15219), .ZN(n12287) );
  NOR2_X1 U14672 ( .A1(n12931), .A2(n14856), .ZN(n12286) );
  AOI211_X1 U14673 ( .C1(n12720), .C2(n12326), .A(n12287), .B(n12286), .ZN(
        n12288) );
  OAI21_X1 U14674 ( .B1(n12289), .B2(n12310), .A(n12288), .ZN(P3_U3175) );
  XNOR2_X1 U14675 ( .A(n12291), .B(n12290), .ZN(n12298) );
  AOI22_X1 U14676 ( .A1(n12292), .A2(n14865), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12293) );
  OAI21_X1 U14677 ( .B1(n14856), .B2(n12294), .A(n12293), .ZN(n12295) );
  AOI21_X1 U14678 ( .B1(n12296), .B2(n12326), .A(n12295), .ZN(n12297) );
  OAI21_X1 U14679 ( .B1(n12298), .B2(n12310), .A(n12297), .ZN(P3_U3176) );
  NAND2_X1 U14680 ( .A1(n12300), .A2(n12299), .ZN(n12304) );
  NOR2_X1 U14681 ( .A1(n12302), .A2(n12301), .ZN(n12303) );
  XNOR2_X1 U14682 ( .A(n12304), .B(n12303), .ZN(n12311) );
  NAND2_X1 U14683 ( .A1(n12326), .A2(n12768), .ZN(n12306) );
  AOI22_X1 U14684 ( .A1(n12315), .A2(n12766), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12305) );
  OAI211_X1 U14685 ( .C1(n12307), .C2(n12317), .A(n12306), .B(n12305), .ZN(
        n12308) );
  AOI21_X1 U14686 ( .B1(n12885), .B2(n14847), .A(n12308), .ZN(n12309) );
  OAI21_X1 U14687 ( .B1(n12311), .B2(n12310), .A(n12309), .ZN(P3_U3178) );
  NAND2_X1 U14688 ( .A1(n12314), .A2(n14857), .ZN(n12320) );
  AOI22_X1 U14689 ( .A1(n12315), .A2(n12535), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12316) );
  OAI21_X1 U14690 ( .B1(n12669), .B2(n12317), .A(n12316), .ZN(n12318) );
  AOI21_X1 U14691 ( .B1(n12671), .B2(n12326), .A(n12318), .ZN(n12319) );
  OAI211_X1 U14692 ( .C1(n12915), .C2(n14856), .A(n12320), .B(n12319), .ZN(
        P3_U3180) );
  XNOR2_X1 U14693 ( .A(n12321), .B(n12830), .ZN(n12322) );
  XNOR2_X1 U14694 ( .A(n12323), .B(n12322), .ZN(n12330) );
  NAND2_X1 U14695 ( .A1(n12541), .A2(n12829), .ZN(n12324) );
  OAI21_X1 U14696 ( .B1(n12325), .B2(n15042), .A(n12324), .ZN(n12812) );
  AOI22_X1 U14697 ( .A1(n12812), .A2(n14865), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12328) );
  NAND2_X1 U14698 ( .A1(n12326), .A2(n12814), .ZN(n12327) );
  OAI211_X1 U14699 ( .C1(n14364), .C2(n14856), .A(n12328), .B(n12327), .ZN(
        n12329) );
  AOI21_X1 U14700 ( .B1(n12330), .B2(n14857), .A(n12329), .ZN(n12331) );
  INV_X1 U14701 ( .A(n12331), .ZN(P3_U3181) );
  XNOR2_X1 U14702 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12335) );
  NAND2_X1 U14703 ( .A1(n12957), .A2(n12338), .ZN(n12337) );
  NAND2_X1 U14704 ( .A1(n12340), .A2(SI_31_), .ZN(n12336) );
  INV_X1 U14705 ( .A(n12348), .ZN(n12533) );
  NAND2_X1 U14706 ( .A1(n12907), .A2(n12533), .ZN(n12383) );
  NAND2_X1 U14707 ( .A1(n6482), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12344) );
  NAND2_X1 U14708 ( .A1(n9529), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U14709 ( .A1(n12341), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12342) );
  NAND4_X1 U14710 ( .A1(n12345), .A2(n12344), .A3(n12343), .A4(n12342), .ZN(
        n12631) );
  NAND2_X1 U14711 ( .A1(n12383), .A2(n12631), .ZN(n12381) );
  NAND2_X1 U14712 ( .A1(n6490), .A2(n12398), .ZN(n12385) );
  INV_X1 U14713 ( .A(n12346), .ZN(n12347) );
  INV_X1 U14714 ( .A(n12631), .ZN(n12351) );
  OR2_X1 U14715 ( .A1(n12900), .A2(n12351), .ZN(n12350) );
  INV_X1 U14716 ( .A(n12907), .ZN(n12352) );
  NAND2_X1 U14717 ( .A1(n12352), .A2(n12348), .ZN(n12349) );
  NAND2_X1 U14718 ( .A1(n12350), .A2(n12349), .ZN(n12522) );
  NAND2_X1 U14719 ( .A1(n12352), .A2(n12351), .ZN(n12387) );
  NOR2_X1 U14720 ( .A1(n12846), .A2(n12631), .ZN(n12520) );
  INV_X1 U14721 ( .A(n12383), .ZN(n12517) );
  INV_X1 U14722 ( .A(n12697), .ZN(n12376) );
  INV_X1 U14723 ( .A(n12353), .ZN(n12354) );
  INV_X1 U14724 ( .A(n12754), .ZN(n12373) );
  NAND4_X1 U14725 ( .A1(n15036), .A2(n12357), .A3(n12356), .A4(n7000), .ZN(
        n12362) );
  NAND4_X1 U14726 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12435), .ZN(
        n12361) );
  NOR2_X1 U14727 ( .A1(n12362), .A2(n12361), .ZN(n12366) );
  NOR2_X1 U14728 ( .A1(n12364), .A2(n12363), .ZN(n12365) );
  NAND4_X1 U14729 ( .A1(n12366), .A2(n9266), .A3(n7001), .A4(n12365), .ZN(
        n12368) );
  NOR3_X1 U14730 ( .A1(n12368), .A2(n12367), .A3(n12454), .ZN(n12369) );
  AND2_X1 U14731 ( .A1(n12466), .A2(n12800), .ZN(n12821) );
  INV_X1 U14732 ( .A(n12839), .ZN(n12826) );
  NAND4_X1 U14733 ( .A1(n12802), .A2(n12369), .A3(n12821), .A4(n12826), .ZN(
        n12370) );
  NOR2_X1 U14734 ( .A1(n12472), .A2(n12370), .ZN(n12371) );
  NAND4_X1 U14735 ( .A1(n12726), .A2(n12373), .A3(n12372), .A4(n12371), .ZN(
        n12374) );
  OR4_X1 U14736 ( .A1(n12705), .A2(n12716), .A3(n12740), .A4(n12374), .ZN(
        n12375) );
  XNOR2_X1 U14737 ( .A(n12506), .B(n12678), .ZN(n12666) );
  NAND4_X1 U14738 ( .A1(n12379), .A2(n12378), .A3(n12377), .A4(n12666), .ZN(
        n12380) );
  NOR4_X1 U14739 ( .A1(n12520), .A2(n12522), .A3(n12517), .A4(n12380), .ZN(
        n12392) );
  INV_X1 U14740 ( .A(n12381), .ZN(n12382) );
  NOR3_X1 U14741 ( .A1(n12382), .A2(n12846), .A3(n6490), .ZN(n12390) );
  NAND3_X1 U14742 ( .A1(n12383), .A2(n6490), .A3(n12631), .ZN(n12384) );
  OAI211_X1 U14743 ( .C1(n12900), .C2(n9044), .A(n12384), .B(n12398), .ZN(
        n12389) );
  INV_X1 U14744 ( .A(n12385), .ZN(n12386) );
  NAND3_X1 U14745 ( .A1(n12387), .A2(n12386), .A3(n12519), .ZN(n12388) );
  OAI22_X1 U14746 ( .A1(n12390), .A2(n12389), .B1(n12522), .B2(n12388), .ZN(
        n12391) );
  OAI21_X1 U14747 ( .B1(n12394), .B2(n12514), .A(n12393), .ZN(n12515) );
  INV_X1 U14748 ( .A(n12395), .ZN(n12927) );
  MUX2_X1 U14749 ( .A(n12396), .B(n6495), .S(n12504), .Z(n12494) );
  AND2_X1 U14750 ( .A1(n12397), .A2(n12450), .ZN(n12453) );
  NOR2_X1 U14751 ( .A1(n12400), .A2(n12529), .ZN(n12399) );
  MUX2_X1 U14752 ( .A(n15030), .B(n12399), .S(n12398), .Z(n12403) );
  INV_X1 U14753 ( .A(n12400), .ZN(n12401) );
  AOI21_X1 U14754 ( .B1(n6526), .B2(n12401), .A(n12514), .ZN(n12402) );
  NOR3_X1 U14755 ( .A1(n12403), .A2(n12404), .A3(n12402), .ZN(n12409) );
  NAND2_X1 U14756 ( .A1(n10657), .A2(n6526), .ZN(n12408) );
  OAI211_X1 U14757 ( .C1(n12409), .C2(n12408), .A(n12407), .B(n12406), .ZN(
        n12411) );
  NAND2_X1 U14758 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  MUX2_X1 U14759 ( .A(n12413), .B(n12412), .S(n12514), .Z(n12415) );
  OR2_X1 U14760 ( .A1(n12415), .A2(n12414), .ZN(n12421) );
  NAND3_X1 U14761 ( .A1(n12421), .A2(n12423), .A3(n12416), .ZN(n12417) );
  OAI211_X1 U14762 ( .C1(n12419), .C2(n12418), .A(n12417), .B(n12428), .ZN(
        n12420) );
  NAND2_X1 U14763 ( .A1(n12420), .A2(n12425), .ZN(n12431) );
  INV_X1 U14764 ( .A(n12421), .ZN(n12427) );
  NAND2_X1 U14765 ( .A1(n12423), .A2(n12422), .ZN(n12426) );
  OAI211_X1 U14766 ( .C1(n12427), .C2(n12426), .A(n12425), .B(n12424), .ZN(
        n12429) );
  NAND2_X1 U14767 ( .A1(n12429), .A2(n12428), .ZN(n12430) );
  MUX2_X1 U14768 ( .A(n12431), .B(n12430), .S(n12504), .Z(n12437) );
  MUX2_X1 U14769 ( .A(n12433), .B(n12432), .S(n12504), .Z(n12434) );
  OAI211_X1 U14770 ( .C1(n12437), .C2(n12436), .A(n12435), .B(n12434), .ZN(
        n12441) );
  MUX2_X1 U14771 ( .A(n12439), .B(n12438), .S(n12514), .Z(n12440) );
  MUX2_X1 U14772 ( .A(n12504), .B(n15069), .S(n12546), .Z(n12442) );
  OAI21_X1 U14773 ( .B1(n12443), .B2(n12514), .A(n12442), .ZN(n12444) );
  MUX2_X1 U14774 ( .A(n12446), .B(n12445), .S(n12514), .Z(n12448) );
  AOI21_X1 U14775 ( .B1(n12457), .B2(n12449), .A(n12504), .ZN(n12451) );
  OAI21_X1 U14776 ( .B1(n12453), .B2(n12514), .A(n12452), .ZN(n12456) );
  INV_X1 U14777 ( .A(n12454), .ZN(n12455) );
  OAI211_X1 U14778 ( .C1(n12457), .C2(n12514), .A(n12456), .B(n12455), .ZN(
        n12461) );
  MUX2_X1 U14779 ( .A(n12459), .B(n12458), .S(n12504), .Z(n12460) );
  MUX2_X1 U14780 ( .A(n12462), .B(n12819), .S(n12504), .Z(n12463) );
  AOI21_X1 U14781 ( .B1(n12464), .B2(n12800), .A(n12504), .ZN(n12465) );
  INV_X1 U14782 ( .A(n12779), .ZN(n12468) );
  INV_X1 U14783 ( .A(n12466), .ZN(n12467) );
  OAI21_X1 U14784 ( .B1(n12468), .B2(n12467), .A(n12504), .ZN(n12471) );
  NOR3_X1 U14785 ( .A1(n12473), .A2(n12472), .A3(n12773), .ZN(n12485) );
  INV_X1 U14786 ( .A(n12477), .ZN(n12476) );
  OAI211_X1 U14787 ( .C1(n12476), .C2(n12475), .A(n12481), .B(n12474), .ZN(
        n12480) );
  OAI211_X1 U14788 ( .C1(n12773), .C2(n12478), .A(n12482), .B(n12477), .ZN(
        n12479) );
  MUX2_X1 U14789 ( .A(n12480), .B(n12479), .S(n12514), .Z(n12484) );
  MUX2_X1 U14790 ( .A(n12482), .B(n12481), .S(n12514), .Z(n12483) );
  OAI211_X1 U14791 ( .C1(n12485), .C2(n12484), .A(n7083), .B(n12483), .ZN(
        n12490) );
  NAND2_X1 U14792 ( .A1(n12486), .A2(n12730), .ZN(n12488) );
  MUX2_X1 U14793 ( .A(n12488), .B(n12487), .S(n12504), .Z(n12489) );
  NAND3_X1 U14794 ( .A1(n12490), .A2(n12726), .A3(n12489), .ZN(n12493) );
  INV_X1 U14795 ( .A(n12716), .ZN(n12714) );
  MUX2_X1 U14796 ( .A(n12491), .B(n6577), .S(n12514), .Z(n12492) );
  INV_X1 U14797 ( .A(n12495), .ZN(n12499) );
  AOI21_X1 U14798 ( .B1(n12497), .B2(n12496), .A(n12499), .ZN(n12498) );
  MUX2_X1 U14799 ( .A(n12499), .B(n12498), .S(n12514), .Z(n12500) );
  MUX2_X1 U14800 ( .A(n12504), .B(n12501), .S(n12536), .Z(n12502) );
  AOI21_X1 U14801 ( .B1(n12919), .B2(n12514), .A(n12502), .ZN(n12503) );
  NOR2_X1 U14802 ( .A1(n12505), .A2(n12504), .ZN(n12508) );
  NOR2_X1 U14803 ( .A1(n12678), .A2(n12514), .ZN(n12507) );
  MUX2_X1 U14804 ( .A(n12508), .B(n12507), .S(n12506), .Z(n12509) );
  OAI21_X1 U14805 ( .B1(n12510), .B2(n12509), .A(n6991), .ZN(n12513) );
  NAND3_X1 U14806 ( .A1(n12911), .A2(n12535), .A3(n12514), .ZN(n12512) );
  INV_X1 U14807 ( .A(n12516), .ZN(n12518) );
  INV_X1 U14808 ( .A(n12520), .ZN(n12521) );
  NAND3_X1 U14809 ( .A1(n12827), .A2(n12527), .A3(n12526), .ZN(n12528) );
  OAI211_X1 U14810 ( .C1(n12529), .C2(n12531), .A(n12528), .B(P3_B_REG_SCAN_IN), .ZN(n12530) );
  OAI21_X1 U14811 ( .B1(n12532), .B2(n12531), .A(n12530), .ZN(P3_U3296) );
  MUX2_X1 U14812 ( .A(n12631), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12554), .Z(
        P3_U3522) );
  MUX2_X1 U14813 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12533), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14814 ( .A(n12534), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12554), .Z(
        P3_U3520) );
  MUX2_X1 U14815 ( .A(n12535), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12554), .Z(
        P3_U3518) );
  MUX2_X1 U14816 ( .A(n12678), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12554), .Z(
        P3_U3517) );
  MUX2_X1 U14817 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12536), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14818 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12679), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14819 ( .A(n12537), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12554), .Z(
        P3_U3514) );
  MUX2_X1 U14820 ( .A(n12538), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12554), .Z(
        P3_U3513) );
  MUX2_X1 U14821 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12744), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14822 ( .A(n12539), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12554), .Z(
        P3_U3511) );
  MUX2_X1 U14823 ( .A(n12766), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12554), .Z(
        P3_U3510) );
  MUX2_X1 U14824 ( .A(n12540), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12554), .Z(
        P3_U3509) );
  MUX2_X1 U14825 ( .A(n12796), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12554), .Z(
        P3_U3508) );
  MUX2_X1 U14826 ( .A(n12541), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12554), .Z(
        P3_U3507) );
  MUX2_X1 U14827 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12830), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14828 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12542), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14829 ( .A(n12828), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12554), .Z(
        P3_U3504) );
  MUX2_X1 U14830 ( .A(n12543), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12554), .Z(
        P3_U3503) );
  MUX2_X1 U14831 ( .A(n12544), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12554), .Z(
        P3_U3502) );
  MUX2_X1 U14832 ( .A(n12545), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12554), .Z(
        P3_U3501) );
  MUX2_X1 U14833 ( .A(n12546), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12554), .Z(
        P3_U3500) );
  MUX2_X1 U14834 ( .A(n12547), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12554), .Z(
        P3_U3499) );
  MUX2_X1 U14835 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12548), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14836 ( .A(n12549), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12554), .Z(
        P3_U3497) );
  MUX2_X1 U14837 ( .A(n12550), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12554), .Z(
        P3_U3496) );
  MUX2_X1 U14838 ( .A(n12551), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12554), .Z(
        P3_U3495) );
  MUX2_X1 U14839 ( .A(n12552), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12554), .Z(
        P3_U3494) );
  MUX2_X1 U14840 ( .A(n12553), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12554), .Z(
        P3_U3493) );
  MUX2_X1 U14841 ( .A(n9495), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12554), .Z(
        P3_U3492) );
  MUX2_X1 U14842 ( .A(n12555), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12554), .Z(
        P3_U3491) );
  INV_X1 U14843 ( .A(n14962), .ZN(n12593) );
  XNOR2_X1 U14844 ( .A(n12593), .B(n12558), .ZN(n14956) );
  MUX2_X1 U14845 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n12559), .S(n12596), .Z(
        n14973) );
  NOR2_X1 U14846 ( .A1(n12599), .A2(n12560), .ZN(n12561) );
  INV_X1 U14847 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14992) );
  NOR2_X1 U14848 ( .A1(n14992), .A2(n14991), .ZN(n14990) );
  OR2_X1 U14849 ( .A1(n12578), .A2(n12835), .ZN(n12602) );
  NAND2_X1 U14850 ( .A1(n12578), .A2(n12835), .ZN(n12562) );
  NAND2_X1 U14851 ( .A1(n12602), .A2(n12562), .ZN(n15009) );
  AND2_X1 U14852 ( .A1(n12604), .A2(n12563), .ZN(n12564) );
  NAND2_X1 U14853 ( .A1(n12610), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12565) );
  OAI21_X1 U14854 ( .B1(n12610), .B2(P3_REG2_REG_16__SCAN_IN), .A(n12565), 
        .ZN(n14324) );
  INV_X1 U14855 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14340) );
  OR2_X1 U14856 ( .A1(n12614), .A2(n12770), .ZN(n12568) );
  NAND2_X1 U14857 ( .A1(n12614), .A2(n12770), .ZN(n12567) );
  AND2_X1 U14858 ( .A1(n12568), .A2(n12567), .ZN(n14356) );
  INV_X1 U14859 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12569) );
  MUX2_X1 U14860 ( .A(n12569), .B(P3_REG2_REG_19__SCAN_IN), .S(n9044), .Z(
        n12617) );
  XNOR2_X1 U14861 ( .A(n12570), .B(n12617), .ZN(n12628) );
  NAND2_X1 U14862 ( .A1(n15017), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12601) );
  INV_X1 U14863 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U14864 ( .A1(n14962), .A2(n12572), .ZN(n12573) );
  NAND2_X1 U14865 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n14958), .ZN(n14957) );
  MUX2_X1 U14866 ( .A(n14382), .B(P3_REG1_REG_12__SCAN_IN), .S(n12596), .Z(
        n14976) );
  NAND2_X1 U14867 ( .A1(n14997), .A2(n12574), .ZN(n12575) );
  NAND2_X1 U14868 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n14994), .ZN(n14993) );
  NAND2_X1 U14869 ( .A1(n12575), .A2(n14993), .ZN(n15012) );
  INV_X1 U14870 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12577) );
  INV_X1 U14871 ( .A(n12601), .ZN(n12576) );
  AOI21_X1 U14872 ( .B1(n12578), .B2(n12577), .A(n12576), .ZN(n15013) );
  NAND2_X1 U14873 ( .A1(n15012), .A2(n15013), .ZN(n15011) );
  NAND2_X1 U14874 ( .A1(n12604), .A2(n12579), .ZN(n12580) );
  XOR2_X1 U14875 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12610), .Z(n14319) );
  AOI22_X1 U14876 ( .A1(n14320), .A2(n14319), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n12610), .ZN(n12581) );
  NAND2_X1 U14877 ( .A1(n12612), .A2(n12582), .ZN(n12583) );
  XOR2_X1 U14878 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12614), .Z(n14347) );
  AOI22_X1 U14879 ( .A1(n14348), .A2(n14347), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12614), .ZN(n12584) );
  XNOR2_X1 U14880 ( .A(n6490), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12616) );
  XNOR2_X1 U14881 ( .A(n12584), .B(n12616), .ZN(n12626) );
  MUX2_X1 U14882 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12586), .Z(n12613) );
  MUX2_X1 U14883 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12586), .Z(n12585) );
  MUX2_X1 U14884 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12586), .Z(n12597) );
  INV_X1 U14885 ( .A(n12597), .ZN(n12598) );
  MUX2_X1 U14886 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12586), .Z(n12594) );
  INV_X1 U14887 ( .A(n12594), .ZN(n12595) );
  MUX2_X1 U14888 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12586), .Z(n12591) );
  INV_X1 U14889 ( .A(n12591), .ZN(n12592) );
  INV_X1 U14890 ( .A(n12587), .ZN(n12589) );
  AOI21_X1 U14891 ( .B1(n12590), .B2(n12589), .A(n12588), .ZN(n14967) );
  XNOR2_X1 U14892 ( .A(n12591), .B(n14962), .ZN(n14966) );
  XNOR2_X1 U14893 ( .A(n12594), .B(n12596), .ZN(n14985) );
  XNOR2_X1 U14894 ( .A(n12597), .B(n14997), .ZN(n15002) );
  NOR2_X1 U14895 ( .A1(n15001), .A2(n15002), .ZN(n15000) );
  INV_X1 U14896 ( .A(n15009), .ZN(n12600) );
  MUX2_X1 U14897 ( .A(n12600), .B(n15013), .S(n12586), .Z(n15024) );
  MUX2_X1 U14898 ( .A(n12602), .B(n12601), .S(n12586), .Z(n12603) );
  INV_X1 U14899 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14367) );
  MUX2_X1 U14900 ( .A(n12816), .B(n14367), .S(n12586), .Z(n14308) );
  INV_X1 U14901 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12609) );
  INV_X1 U14902 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12896) );
  MUX2_X1 U14903 ( .A(n12609), .B(n12896), .S(n12586), .Z(n12611) );
  INV_X1 U14904 ( .A(n12610), .ZN(n14315) );
  NAND2_X1 U14905 ( .A1(n12611), .A2(n14315), .ZN(n14316) );
  XNOR2_X1 U14906 ( .A(n12613), .B(n12612), .ZN(n14335) );
  INV_X1 U14907 ( .A(n12614), .ZN(n14346) );
  XOR2_X1 U14908 ( .A(n12614), .B(n12615), .Z(n14350) );
  MUX2_X1 U14909 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12586), .Z(n14351) );
  NOR2_X1 U14910 ( .A1(n14350), .A2(n14351), .ZN(n14349) );
  AOI21_X1 U14911 ( .B1(n12615), .B2(n14346), .A(n14349), .ZN(n12620) );
  INV_X1 U14912 ( .A(n12616), .ZN(n12618) );
  MUX2_X1 U14913 ( .A(n12618), .B(n12617), .S(n6475), .Z(n12619) );
  NOR2_X1 U14914 ( .A1(n7449), .A2(n15003), .ZN(n12625) );
  NAND2_X1 U14915 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n12622)
         );
  NAND2_X1 U14916 ( .A1(n15021), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12621) );
  OAI211_X1 U14917 ( .C1(n15018), .C2(n6490), .A(n12622), .B(n12621), .ZN(
        n12624) );
  AOI211_X1 U14918 ( .C1(n12626), .C2(n15014), .A(n12625), .B(n12624), .ZN(
        n12627) );
  OAI21_X1 U14919 ( .B1(n12628), .B2(n15028), .A(n12627), .ZN(P3_U3201) );
  INV_X1 U14920 ( .A(n12629), .ZN(n12630) );
  NAND2_X1 U14921 ( .A1(n12631), .A2(n12630), .ZN(n12901) );
  NAND2_X1 U14922 ( .A1(n12805), .A2(n12632), .ZN(n12636) );
  OAI21_X1 U14923 ( .B1(n12844), .B2(n12901), .A(n12636), .ZN(n12634) );
  AOI21_X1 U14924 ( .B1(n12844), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12634), 
        .ZN(n12633) );
  OAI21_X1 U14925 ( .B1(n12846), .B2(n12807), .A(n12633), .ZN(P3_U3202) );
  AOI21_X1 U14926 ( .B1(n12844), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12634), 
        .ZN(n12635) );
  OAI21_X1 U14927 ( .B1(n12907), .B2(n12807), .A(n12635), .ZN(P3_U3203) );
  INV_X1 U14928 ( .A(n12636), .ZN(n12639) );
  NOR2_X1 U14929 ( .A1(n12637), .A2(n12807), .ZN(n12638) );
  AOI211_X1 U14930 ( .C1(n12844), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12639), 
        .B(n12638), .ZN(n12642) );
  NAND2_X1 U14931 ( .A1(n12640), .A2(n12841), .ZN(n12641) );
  OAI211_X1 U14932 ( .C1(n12643), .C2(n12844), .A(n12642), .B(n12641), .ZN(
        P3_U3204) );
  OAI22_X1 U14933 ( .A1(n15045), .A2(n12645), .B1(n12644), .B2(n15032), .ZN(
        n12646) );
  AOI21_X1 U14934 ( .B1(n12647), .B2(n12837), .A(n12646), .ZN(n12651) );
  INV_X1 U14935 ( .A(n12648), .ZN(n12649) );
  NAND2_X1 U14936 ( .A1(n12649), .A2(n12841), .ZN(n12650) );
  OAI211_X1 U14937 ( .C1(n12652), .C2(n12844), .A(n12651), .B(n12650), .ZN(
        P3_U3205) );
  XNOR2_X1 U14938 ( .A(n12653), .B(n12658), .ZN(n12657) );
  NAND2_X1 U14939 ( .A1(n12678), .A2(n12827), .ZN(n12654) );
  OAI21_X1 U14940 ( .B1(n12655), .B2(n15040), .A(n12654), .ZN(n12656) );
  AOI21_X1 U14941 ( .B1(n12659), .B2(n12658), .A(n9575), .ZN(n12850) );
  INV_X1 U14942 ( .A(n12850), .ZN(n12663) );
  AOI22_X1 U14943 ( .A1(n12844), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n12805), 
        .B2(n12660), .ZN(n12661) );
  OAI21_X1 U14944 ( .B1(n12911), .B2(n12807), .A(n12661), .ZN(n12662) );
  AOI21_X1 U14945 ( .B1(n12663), .B2(n12841), .A(n12662), .ZN(n12664) );
  OAI21_X1 U14946 ( .B1(n12849), .B2(n12844), .A(n12664), .ZN(P3_U3206) );
  XNOR2_X1 U14947 ( .A(n12665), .B(n12666), .ZN(n12854) );
  INV_X1 U14948 ( .A(n12854), .ZN(n12675) );
  XNOR2_X1 U14949 ( .A(n12667), .B(n12666), .ZN(n12668) );
  OAI222_X1 U14950 ( .A1(n15040), .A2(n12670), .B1(n15042), .B2(n12669), .C1(
        n15038), .C2(n12668), .ZN(n12853) );
  AOI22_X1 U14951 ( .A1(n12844), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n12805), 
        .B2(n12671), .ZN(n12672) );
  OAI21_X1 U14952 ( .B1(n12915), .B2(n12807), .A(n12672), .ZN(n12673) );
  AOI21_X1 U14953 ( .B1(n12853), .B2(n15045), .A(n12673), .ZN(n12674) );
  OAI21_X1 U14954 ( .B1(n12675), .B2(n12791), .A(n12674), .ZN(P3_U3207) );
  XNOR2_X1 U14955 ( .A(n12677), .B(n12676), .ZN(n12686) );
  AOI22_X1 U14956 ( .A1(n12679), .A2(n12827), .B1(n12829), .B2(n12678), .ZN(
        n12685) );
  OAI21_X1 U14957 ( .B1(n12682), .B2(n12681), .A(n12680), .ZN(n12858) );
  NAND2_X1 U14958 ( .A1(n12858), .A2(n12683), .ZN(n12684) );
  OAI211_X1 U14959 ( .C1(n12686), .C2(n15038), .A(n12685), .B(n12684), .ZN(
        n12857) );
  INV_X1 U14960 ( .A(n12857), .ZN(n12692) );
  AOI22_X1 U14961 ( .A1(n12844), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12805), 
        .B2(n12687), .ZN(n12688) );
  OAI21_X1 U14962 ( .B1(n12919), .B2(n12807), .A(n12688), .ZN(n12689) );
  AOI21_X1 U14963 ( .B1(n12858), .B2(n12690), .A(n12689), .ZN(n12691) );
  OAI21_X1 U14964 ( .B1(n12692), .B2(n12844), .A(n12691), .ZN(P3_U3208) );
  XNOR2_X1 U14965 ( .A(n12693), .B(n12697), .ZN(n12695) );
  OAI21_X1 U14966 ( .B1(n12695), .B2(n15038), .A(n12694), .ZN(n12861) );
  INV_X1 U14967 ( .A(n12861), .ZN(n12703) );
  OAI21_X1 U14968 ( .B1(n12698), .B2(n12697), .A(n12696), .ZN(n12862) );
  AOI22_X1 U14969 ( .A1(n12844), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12805), 
        .B2(n12699), .ZN(n12700) );
  OAI21_X1 U14970 ( .B1(n12923), .B2(n12807), .A(n12700), .ZN(n12701) );
  AOI21_X1 U14971 ( .B1(n12862), .B2(n12841), .A(n12701), .ZN(n12702) );
  OAI21_X1 U14972 ( .B1(n12703), .B2(n12844), .A(n12702), .ZN(P3_U3209) );
  XNOR2_X1 U14973 ( .A(n12704), .B(n12705), .ZN(n12866) );
  INV_X1 U14974 ( .A(n12866), .ZN(n12713) );
  XNOR2_X1 U14975 ( .A(n12706), .B(n12705), .ZN(n12707) );
  OAI222_X1 U14976 ( .A1(n15040), .A2(n12708), .B1(n15042), .B2(n12729), .C1(
        n15038), .C2(n12707), .ZN(n12865) );
  AOI22_X1 U14977 ( .A1(n12844), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12805), 
        .B2(n12709), .ZN(n12710) );
  OAI21_X1 U14978 ( .B1(n12927), .B2(n12807), .A(n12710), .ZN(n12711) );
  AOI21_X1 U14979 ( .B1(n12865), .B2(n15045), .A(n12711), .ZN(n12712) );
  OAI21_X1 U14980 ( .B1(n12713), .B2(n12791), .A(n12712), .ZN(P3_U3210) );
  XNOR2_X1 U14981 ( .A(n12715), .B(n12714), .ZN(n12870) );
  INV_X1 U14982 ( .A(n12870), .ZN(n12724) );
  XNOR2_X1 U14983 ( .A(n12717), .B(n12716), .ZN(n12719) );
  OAI21_X1 U14984 ( .B1(n12719), .B2(n15038), .A(n12718), .ZN(n12869) );
  AOI22_X1 U14985 ( .A1(n12844), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12805), 
        .B2(n12720), .ZN(n12721) );
  OAI21_X1 U14986 ( .B1(n12931), .B2(n12807), .A(n12721), .ZN(n12722) );
  AOI21_X1 U14987 ( .B1(n12869), .B2(n15045), .A(n12722), .ZN(n12723) );
  OAI21_X1 U14988 ( .B1(n12791), .B2(n12724), .A(n12723), .ZN(P3_U3211) );
  XOR2_X1 U14989 ( .A(n12726), .B(n12725), .Z(n12874) );
  INV_X1 U14990 ( .A(n12874), .ZN(n12736) );
  XNOR2_X1 U14991 ( .A(n12727), .B(n12726), .ZN(n12728) );
  OAI222_X1 U14992 ( .A1(n15042), .A2(n12730), .B1(n15040), .B2(n12729), .C1(
        n15038), .C2(n12728), .ZN(n12873) );
  INV_X1 U14993 ( .A(n12731), .ZN(n12935) );
  AOI22_X1 U14994 ( .A1(n12844), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12805), 
        .B2(n12732), .ZN(n12733) );
  OAI21_X1 U14995 ( .B1(n12935), .B2(n12807), .A(n12733), .ZN(n12734) );
  AOI21_X1 U14996 ( .B1(n12873), .B2(n15045), .A(n12734), .ZN(n12735) );
  OAI21_X1 U14997 ( .B1(n12791), .B2(n12736), .A(n12735), .ZN(P3_U3212) );
  NAND2_X1 U14998 ( .A1(n12738), .A2(n12740), .ZN(n12739) );
  NAND2_X1 U14999 ( .A1(n12737), .A2(n12739), .ZN(n12878) );
  OAI21_X1 U15000 ( .B1(n12741), .B2(n12740), .A(n12832), .ZN(n12742) );
  OR2_X1 U15001 ( .A1(n12743), .A2(n12742), .ZN(n12746) );
  AOI22_X1 U15002 ( .A1(n12744), .A2(n12829), .B1(n12827), .B2(n12766), .ZN(
        n12745) );
  INV_X1 U15003 ( .A(n12877), .ZN(n12750) );
  AOI22_X1 U15004 ( .A1(n12844), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12805), 
        .B2(n12747), .ZN(n12748) );
  OAI21_X1 U15005 ( .B1(n12939), .B2(n12807), .A(n12748), .ZN(n12749) );
  AOI21_X1 U15006 ( .B1(n12750), .B2(n15045), .A(n12749), .ZN(n12751) );
  OAI21_X1 U15007 ( .B1(n12791), .B2(n12878), .A(n12751), .ZN(P3_U3213) );
  XNOR2_X1 U15008 ( .A(n12752), .B(n12754), .ZN(n12882) );
  INV_X1 U15009 ( .A(n12882), .ZN(n12763) );
  NAND2_X1 U15010 ( .A1(n12753), .A2(n12832), .ZN(n12758) );
  AOI21_X1 U15011 ( .B1(n12764), .B2(n12755), .A(n12754), .ZN(n12757) );
  OAI21_X1 U15012 ( .B1(n12758), .B2(n12757), .A(n12756), .ZN(n12881) );
  AOI22_X1 U15013 ( .A1(n12844), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12759), 
        .B2(n12805), .ZN(n12760) );
  OAI21_X1 U15014 ( .B1(n12943), .B2(n12807), .A(n12760), .ZN(n12761) );
  AOI21_X1 U15015 ( .B1(n12881), .B2(n15045), .A(n12761), .ZN(n12762) );
  OAI21_X1 U15016 ( .B1(n12763), .B2(n12791), .A(n12762), .ZN(P3_U3214) );
  OAI21_X1 U15017 ( .B1(n12765), .B2(n12773), .A(n12764), .ZN(n12767) );
  AOI222_X1 U15018 ( .A1(n12832), .A2(n12767), .B1(n12766), .B2(n12797), .C1(
        n12796), .C2(n12827), .ZN(n12888) );
  INV_X1 U15019 ( .A(n12768), .ZN(n12769) );
  OAI22_X1 U15020 ( .A1(n15045), .A2(n12770), .B1(n12769), .B2(n15032), .ZN(
        n12771) );
  AOI21_X1 U15021 ( .B1(n12885), .B2(n12837), .A(n12771), .ZN(n12776) );
  NAND2_X1 U15022 ( .A1(n12774), .A2(n12773), .ZN(n12886) );
  NAND3_X1 U15023 ( .A1(n12772), .A2(n12886), .A3(n12841), .ZN(n12775) );
  OAI211_X1 U15024 ( .C1(n12888), .C2(n12844), .A(n12776), .B(n12775), .ZN(
        P3_U3215) );
  NAND2_X1 U15025 ( .A1(n12777), .A2(n12778), .ZN(n12801) );
  NAND2_X1 U15026 ( .A1(n12801), .A2(n12779), .ZN(n12780) );
  XNOR2_X1 U15027 ( .A(n12780), .B(n12783), .ZN(n12891) );
  INV_X1 U15028 ( .A(n12891), .ZN(n12792) );
  NAND3_X1 U15029 ( .A1(n7450), .A2(n12783), .A3(n12782), .ZN(n12784) );
  NAND3_X1 U15030 ( .A1(n12781), .A2(n12832), .A3(n12784), .ZN(n12786) );
  NAND2_X1 U15031 ( .A1(n12786), .A2(n12785), .ZN(n12890) );
  AOI22_X1 U15032 ( .A1(n12844), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12805), 
        .B2(n12787), .ZN(n12788) );
  OAI21_X1 U15033 ( .B1(n12948), .B2(n12807), .A(n12788), .ZN(n12789) );
  AOI21_X1 U15034 ( .B1(n12890), .B2(n15045), .A(n12789), .ZN(n12790) );
  OAI21_X1 U15035 ( .B1(n12792), .B2(n12791), .A(n12790), .ZN(P3_U3216) );
  INV_X1 U15036 ( .A(n12793), .ZN(n12795) );
  INV_X1 U15037 ( .A(n12802), .ZN(n12794) );
  OAI211_X1 U15038 ( .C1(n12795), .C2(n12794), .A(n12832), .B(n7450), .ZN(
        n12799) );
  AOI22_X1 U15039 ( .A1(n12830), .A2(n12827), .B1(n12797), .B2(n12796), .ZN(
        n12798) );
  NAND2_X1 U15040 ( .A1(n12799), .A2(n12798), .ZN(n12894) );
  INV_X1 U15041 ( .A(n12894), .ZN(n12810) );
  AND2_X1 U15042 ( .A1(n12777), .A2(n12800), .ZN(n12803) );
  OAI21_X1 U15043 ( .B1(n12803), .B2(n12802), .A(n12801), .ZN(n12895) );
  AOI22_X1 U15044 ( .A1(n12844), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12805), 
        .B2(n12804), .ZN(n12806) );
  OAI21_X1 U15045 ( .B1(n12953), .B2(n12807), .A(n12806), .ZN(n12808) );
  AOI21_X1 U15046 ( .B1(n12895), .B2(n12841), .A(n12808), .ZN(n12809) );
  OAI21_X1 U15047 ( .B1(n12810), .B2(n12844), .A(n12809), .ZN(P3_U3217) );
  XNOR2_X1 U15048 ( .A(n12811), .B(n12821), .ZN(n12813) );
  AOI21_X1 U15049 ( .B1(n12813), .B2(n12832), .A(n12812), .ZN(n14363) );
  INV_X1 U15050 ( .A(n14364), .ZN(n12818) );
  INV_X1 U15051 ( .A(n12814), .ZN(n12815) );
  OAI22_X1 U15052 ( .A1(n15045), .A2(n12816), .B1(n12815), .B2(n15032), .ZN(
        n12817) );
  AOI21_X1 U15053 ( .B1(n12818), .B2(n12837), .A(n12817), .ZN(n12824) );
  NAND2_X1 U15054 ( .A1(n12820), .A2(n12819), .ZN(n12822) );
  XNOR2_X1 U15055 ( .A(n12822), .B(n12821), .ZN(n14366) );
  NAND2_X1 U15056 ( .A1(n14366), .A2(n12841), .ZN(n12823) );
  OAI211_X1 U15057 ( .C1(n14363), .C2(n12844), .A(n12824), .B(n12823), .ZN(
        P3_U3218) );
  XNOR2_X1 U15058 ( .A(n12825), .B(n12826), .ZN(n12831) );
  AOI222_X1 U15059 ( .A1(n12832), .A2(n12831), .B1(n12830), .B2(n12829), .C1(
        n12828), .C2(n12827), .ZN(n14368) );
  INV_X1 U15060 ( .A(n14369), .ZN(n12838) );
  INV_X1 U15061 ( .A(n12833), .ZN(n12834) );
  OAI22_X1 U15062 ( .A1(n15045), .A2(n12835), .B1(n12834), .B2(n15032), .ZN(
        n12836) );
  AOI21_X1 U15063 ( .B1(n12838), .B2(n12837), .A(n12836), .ZN(n12843) );
  XNOR2_X1 U15064 ( .A(n12840), .B(n12839), .ZN(n14371) );
  NAND2_X1 U15065 ( .A1(n14371), .A2(n12841), .ZN(n12842) );
  OAI211_X1 U15066 ( .C1(n14368), .C2(n12844), .A(n12843), .B(n12842), .ZN(
        P3_U3219) );
  NOR2_X1 U15067 ( .A1(n12901), .A2(n9553), .ZN(n12847) );
  AOI21_X1 U15068 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n9553), .A(n12847), .ZN(
        n12845) );
  OAI21_X1 U15069 ( .B1(n12846), .B2(n12898), .A(n12845), .ZN(P3_U3490) );
  AOI21_X1 U15070 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n9553), .A(n12847), .ZN(
        n12848) );
  OAI21_X1 U15071 ( .B1(n12907), .B2(n12898), .A(n12848), .ZN(P3_U3489) );
  OAI21_X1 U15072 ( .B1(n14372), .B2(n12850), .A(n12849), .ZN(n12908) );
  INV_X1 U15073 ( .A(n12851), .ZN(n12852) );
  OAI21_X1 U15074 ( .B1(n12911), .B2(n12898), .A(n12852), .ZN(P3_U3486) );
  INV_X1 U15075 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12855) );
  AOI21_X1 U15076 ( .B1(n15054), .B2(n12854), .A(n12853), .ZN(n12912) );
  MUX2_X1 U15077 ( .A(n12855), .B(n12912), .S(n15085), .Z(n12856) );
  OAI21_X1 U15078 ( .B1(n12915), .B2(n12898), .A(n12856), .ZN(P3_U3485) );
  INV_X1 U15079 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12859) );
  AOI21_X1 U15080 ( .B1(n15072), .B2(n12858), .A(n12857), .ZN(n12916) );
  MUX2_X1 U15081 ( .A(n12859), .B(n12916), .S(n15085), .Z(n12860) );
  OAI21_X1 U15082 ( .B1(n12919), .B2(n12898), .A(n12860), .ZN(P3_U3484) );
  INV_X1 U15083 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12863) );
  AOI21_X1 U15084 ( .B1(n15054), .B2(n12862), .A(n12861), .ZN(n12920) );
  MUX2_X1 U15085 ( .A(n12863), .B(n12920), .S(n15085), .Z(n12864) );
  OAI21_X1 U15086 ( .B1(n12923), .B2(n12898), .A(n12864), .ZN(P3_U3483) );
  INV_X1 U15087 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12867) );
  AOI21_X1 U15088 ( .B1(n15054), .B2(n12866), .A(n12865), .ZN(n12924) );
  MUX2_X1 U15089 ( .A(n12867), .B(n12924), .S(n15085), .Z(n12868) );
  OAI21_X1 U15090 ( .B1(n12927), .B2(n12898), .A(n12868), .ZN(P3_U3482) );
  INV_X1 U15091 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12871) );
  AOI21_X1 U15092 ( .B1(n12870), .B2(n15054), .A(n12869), .ZN(n12928) );
  MUX2_X1 U15093 ( .A(n12871), .B(n12928), .S(n15085), .Z(n12872) );
  OAI21_X1 U15094 ( .B1(n12931), .B2(n12898), .A(n12872), .ZN(P3_U3481) );
  INV_X1 U15095 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12875) );
  AOI21_X1 U15096 ( .B1(n12874), .B2(n15054), .A(n12873), .ZN(n12932) );
  MUX2_X1 U15097 ( .A(n12875), .B(n12932), .S(n15085), .Z(n12876) );
  OAI21_X1 U15098 ( .B1(n12935), .B2(n12898), .A(n12876), .ZN(P3_U3480) );
  OAI21_X1 U15099 ( .B1(n12878), .B2(n14372), .A(n12877), .ZN(n12936) );
  MUX2_X1 U15100 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12936), .S(n15085), .Z(
        n12879) );
  INV_X1 U15101 ( .A(n12879), .ZN(n12880) );
  OAI21_X1 U15102 ( .B1(n12939), .B2(n12898), .A(n12880), .ZN(P3_U3479) );
  INV_X1 U15103 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12883) );
  AOI21_X1 U15104 ( .B1(n15054), .B2(n12882), .A(n12881), .ZN(n12940) );
  MUX2_X1 U15105 ( .A(n12883), .B(n12940), .S(n15085), .Z(n12884) );
  OAI21_X1 U15106 ( .B1(n12943), .B2(n12898), .A(n12884), .ZN(P3_U3478) );
  INV_X1 U15107 ( .A(n12885), .ZN(n12889) );
  NAND3_X1 U15108 ( .A1(n12772), .A2(n15054), .A3(n12886), .ZN(n12887) );
  OAI211_X1 U15109 ( .C1(n12889), .C2(n15068), .A(n12888), .B(n12887), .ZN(
        n12944) );
  MUX2_X1 U15110 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12944), .S(n15085), .Z(
        P3_U3477) );
  INV_X1 U15111 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12892) );
  AOI21_X1 U15112 ( .B1(n12891), .B2(n15054), .A(n12890), .ZN(n12945) );
  MUX2_X1 U15113 ( .A(n12892), .B(n12945), .S(n15085), .Z(n12893) );
  OAI21_X1 U15114 ( .B1(n12898), .B2(n12948), .A(n12893), .ZN(P3_U3476) );
  AOI21_X1 U15115 ( .B1(n15054), .B2(n12895), .A(n12894), .ZN(n12949) );
  MUX2_X1 U15116 ( .A(n12896), .B(n12949), .S(n15085), .Z(n12897) );
  OAI21_X1 U15117 ( .B1(n12953), .B2(n12898), .A(n12897), .ZN(P3_U3475) );
  INV_X1 U15118 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12904) );
  INV_X1 U15119 ( .A(n12952), .ZN(n12899) );
  NAND2_X1 U15120 ( .A1(n12900), .A2(n12899), .ZN(n12903) );
  INV_X1 U15121 ( .A(n12901), .ZN(n12902) );
  NAND2_X1 U15122 ( .A1(n12902), .A2(n15076), .ZN(n12906) );
  OAI211_X1 U15123 ( .C1(n15076), .C2(n12904), .A(n12903), .B(n12906), .ZN(
        P3_U3458) );
  NAND2_X1 U15124 ( .A1(n15074), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12905) );
  OAI211_X1 U15125 ( .C1(n12907), .C2(n12952), .A(n12906), .B(n12905), .ZN(
        P3_U3457) );
  INV_X1 U15126 ( .A(n12909), .ZN(n12910) );
  OAI21_X1 U15127 ( .B1(n12911), .B2(n12952), .A(n12910), .ZN(P3_U3454) );
  INV_X1 U15128 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12913) );
  MUX2_X1 U15129 ( .A(n12913), .B(n12912), .S(n15076), .Z(n12914) );
  OAI21_X1 U15130 ( .B1(n12915), .B2(n12952), .A(n12914), .ZN(P3_U3453) );
  MUX2_X1 U15131 ( .A(n12917), .B(n12916), .S(n15076), .Z(n12918) );
  OAI21_X1 U15132 ( .B1(n12919), .B2(n12952), .A(n12918), .ZN(P3_U3452) );
  MUX2_X1 U15133 ( .A(n12921), .B(n12920), .S(n15076), .Z(n12922) );
  OAI21_X1 U15134 ( .B1(n12923), .B2(n12952), .A(n12922), .ZN(P3_U3451) );
  INV_X1 U15135 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12925) );
  MUX2_X1 U15136 ( .A(n12925), .B(n12924), .S(n15076), .Z(n12926) );
  OAI21_X1 U15137 ( .B1(n12927), .B2(n12952), .A(n12926), .ZN(P3_U3450) );
  INV_X1 U15138 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12929) );
  MUX2_X1 U15139 ( .A(n12929), .B(n12928), .S(n15076), .Z(n12930) );
  OAI21_X1 U15140 ( .B1(n12931), .B2(n12952), .A(n12930), .ZN(P3_U3449) );
  MUX2_X1 U15141 ( .A(n12933), .B(n12932), .S(n15076), .Z(n12934) );
  OAI21_X1 U15142 ( .B1(n12935), .B2(n12952), .A(n12934), .ZN(P3_U3448) );
  MUX2_X1 U15143 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12936), .S(n15076), .Z(
        n12937) );
  INV_X1 U15144 ( .A(n12937), .ZN(n12938) );
  OAI21_X1 U15145 ( .B1(n12939), .B2(n12952), .A(n12938), .ZN(P3_U3447) );
  INV_X1 U15146 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12941) );
  MUX2_X1 U15147 ( .A(n12941), .B(n12940), .S(n15076), .Z(n12942) );
  OAI21_X1 U15148 ( .B1(n12943), .B2(n12952), .A(n12942), .ZN(P3_U3446) );
  MUX2_X1 U15149 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12944), .S(n15076), .Z(
        P3_U3444) );
  INV_X1 U15150 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12946) );
  MUX2_X1 U15151 ( .A(n12946), .B(n12945), .S(n15076), .Z(n12947) );
  OAI21_X1 U15152 ( .B1(n12952), .B2(n12948), .A(n12947), .ZN(P3_U3441) );
  INV_X1 U15153 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12950) );
  MUX2_X1 U15154 ( .A(n12950), .B(n12949), .S(n15076), .Z(n12951) );
  OAI21_X1 U15155 ( .B1(n12953), .B2(n12952), .A(n12951), .ZN(P3_U3438) );
  MUX2_X1 U15156 ( .A(P3_D_REG_1__SCAN_IN), .B(n12954), .S(n12955), .Z(
        P3_U3377) );
  MUX2_X1 U15157 ( .A(P3_D_REG_0__SCAN_IN), .B(n12956), .S(n12955), .Z(
        P3_U3376) );
  INV_X1 U15158 ( .A(n12957), .ZN(n12963) );
  NOR4_X1 U15159 ( .A1(n12959), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12958), .A4(
        P3_U3151), .ZN(n12960) );
  AOI21_X1 U15160 ( .B1(n12961), .B2(SI_31_), .A(n12960), .ZN(n12962) );
  OAI21_X1 U15161 ( .B1(n12963), .B2(n12967), .A(n12962), .ZN(P3_U3264) );
  INV_X1 U15162 ( .A(n12964), .ZN(n12966) );
  OAI222_X1 U15163 ( .A1(n12968), .A2(n15211), .B1(n12967), .B2(n12966), .C1(
        n12965), .C2(P3_U3151), .ZN(P3_U3266) );
  XNOR2_X1 U15164 ( .A(n12970), .B(n12969), .ZN(n12977) );
  OR2_X1 U15165 ( .A1(n12971), .A2(n13076), .ZN(n12973) );
  OR2_X1 U15166 ( .A1(n13005), .A2(n13078), .ZN(n12972) );
  NAND2_X1 U15167 ( .A1(n12973), .A2(n12972), .ZN(n13245) );
  AOI22_X1 U15168 ( .A1(n13085), .A2(n13245), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12974) );
  OAI21_X1 U15169 ( .B1(n13249), .B2(n13087), .A(n12974), .ZN(n12975) );
  AOI21_X1 U15170 ( .B1(n13424), .B2(n13095), .A(n12975), .ZN(n12976) );
  OAI21_X1 U15171 ( .B1(n12977), .B2(n13091), .A(n12976), .ZN(P2_U3186) );
  XNOR2_X1 U15172 ( .A(n12978), .B(n12979), .ZN(n12985) );
  OAI22_X1 U15173 ( .A1(n12981), .A2(n13078), .B1(n12980), .B2(n13076), .ZN(
        n13308) );
  AOI22_X1 U15174 ( .A1(n13085), .A2(n13308), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12982) );
  OAI21_X1 U15175 ( .B1(n13306), .B2(n13087), .A(n12982), .ZN(n12983) );
  AOI21_X1 U15176 ( .B1(n13313), .B2(n13095), .A(n12983), .ZN(n12984) );
  OAI21_X1 U15177 ( .B1(n12985), .B2(n13091), .A(n12984), .ZN(P2_U3188) );
  INV_X1 U15178 ( .A(n12986), .ZN(n12987) );
  NOR2_X1 U15179 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  XNOR2_X1 U15180 ( .A(n12990), .B(n12989), .ZN(n12994) );
  AOI22_X1 U15181 ( .A1(n13109), .A2(n13065), .B1(n13064), .B2(n13111), .ZN(
        n13379) );
  NAND2_X1 U15182 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13199)
         );
  NAND2_X1 U15183 ( .A1(n13068), .A2(n13384), .ZN(n12991) );
  OAI211_X1 U15184 ( .C1(n13379), .C2(n13066), .A(n13199), .B(n12991), .ZN(
        n12992) );
  AOI21_X1 U15185 ( .B1(n13383), .B2(n13095), .A(n12992), .ZN(n12993) );
  OAI21_X1 U15186 ( .B1(n12994), .B2(n13091), .A(n12993), .ZN(P2_U3191) );
  XNOR2_X1 U15187 ( .A(n12996), .B(n12995), .ZN(n13002) );
  AND2_X1 U15188 ( .A1(n13107), .A2(n13065), .ZN(n12997) );
  AOI21_X1 U15189 ( .B1(n13109), .B2(n13064), .A(n12997), .ZN(n13345) );
  INV_X1 U15190 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12998) );
  OAI22_X1 U15191 ( .A1(n13345), .A2(n13066), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12998), .ZN(n12999) );
  AOI21_X1 U15192 ( .B1(n13349), .B2(n13068), .A(n12999), .ZN(n13001) );
  NAND2_X1 U15193 ( .A1(n13348), .A2(n13095), .ZN(n13000) );
  OAI211_X1 U15194 ( .C1(n13002), .C2(n13091), .A(n13001), .B(n13000), .ZN(
        P2_U3195) );
  XNOR2_X1 U15195 ( .A(n13004), .B(n13003), .ZN(n13012) );
  OR2_X1 U15196 ( .A1(n13005), .A2(n13076), .ZN(n13007) );
  NAND2_X1 U15197 ( .A1(n13105), .A2(n13064), .ZN(n13006) );
  NAND2_X1 U15198 ( .A1(n13007), .A2(n13006), .ZN(n13275) );
  AOI22_X1 U15199 ( .A1(n13085), .A2(n13275), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13008) );
  OAI21_X1 U15200 ( .B1(n13282), .B2(n13087), .A(n13008), .ZN(n13009) );
  AOI21_X1 U15201 ( .B1(n13010), .B2(n13095), .A(n13009), .ZN(n13011) );
  OAI21_X1 U15202 ( .B1(n13012), .B2(n13091), .A(n13011), .ZN(P2_U3197) );
  OAI21_X1 U15203 ( .B1(n13014), .B2(n13013), .A(n13025), .ZN(n13015) );
  NAND2_X1 U15204 ( .A1(n13015), .A2(n13060), .ZN(n13021) );
  OAI22_X1 U15205 ( .A1(n13017), .A2(n13066), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13016), .ZN(n13018) );
  AOI21_X1 U15206 ( .B1(n13019), .B2(n13068), .A(n13018), .ZN(n13020) );
  OAI211_X1 U15207 ( .C1(n13022), .C2(n13071), .A(n13021), .B(n13020), .ZN(
        P2_U3198) );
  AND3_X1 U15208 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(n13026) );
  OAI21_X1 U15209 ( .B1(n13027), .B2(n13026), .A(n13060), .ZN(n13032) );
  NAND2_X1 U15210 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13164)
         );
  OAI21_X1 U15211 ( .B1(n13028), .B2(n13066), .A(n13164), .ZN(n13029) );
  AOI21_X1 U15212 ( .B1(n13030), .B2(n13068), .A(n13029), .ZN(n13031) );
  OAI211_X1 U15213 ( .C1(n13033), .C2(n13071), .A(n13032), .B(n13031), .ZN(
        P2_U3200) );
  XNOR2_X1 U15214 ( .A(n13035), .B(n13034), .ZN(n13041) );
  OR2_X1 U15215 ( .A1(n13079), .A2(n13076), .ZN(n13037) );
  NAND2_X1 U15216 ( .A1(n13106), .A2(n13064), .ZN(n13036) );
  NAND2_X1 U15217 ( .A1(n13037), .A2(n13036), .ZN(n13290) );
  AOI22_X1 U15218 ( .A1(n13085), .A2(n13290), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13038) );
  OAI21_X1 U15219 ( .B1(n13299), .B2(n13087), .A(n13038), .ZN(n13039) );
  AOI21_X1 U15220 ( .B1(n13441), .B2(n13095), .A(n13039), .ZN(n13040) );
  OAI21_X1 U15221 ( .B1(n13041), .B2(n13091), .A(n13040), .ZN(P2_U3201) );
  OAI21_X1 U15222 ( .B1(n13044), .B2(n13043), .A(n13042), .ZN(n13045) );
  NAND2_X1 U15223 ( .A1(n13045), .A2(n13060), .ZN(n13051) );
  INV_X1 U15224 ( .A(n13046), .ZN(n13360) );
  AND2_X1 U15225 ( .A1(n13110), .A2(n13064), .ZN(n13047) );
  AOI21_X1 U15226 ( .B1(n13108), .B2(n13065), .A(n13047), .ZN(n13366) );
  INV_X1 U15227 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13048) );
  OAI22_X1 U15228 ( .A1(n13366), .A2(n13066), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13048), .ZN(n13049) );
  AOI21_X1 U15229 ( .B1(n13360), .B2(n13068), .A(n13049), .ZN(n13050) );
  OAI211_X1 U15230 ( .C1(n13362), .C2(n13071), .A(n13051), .B(n13050), .ZN(
        P2_U3205) );
  XNOR2_X1 U15231 ( .A(n13052), .B(n13053), .ZN(n13059) );
  NAND2_X1 U15232 ( .A1(n13108), .A2(n13064), .ZN(n13055) );
  NAND2_X1 U15233 ( .A1(n13106), .A2(n13065), .ZN(n13054) );
  NAND2_X1 U15234 ( .A1(n13055), .A2(n13054), .ZN(n13325) );
  AOI22_X1 U15235 ( .A1(n13325), .A2(n13085), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13056) );
  OAI21_X1 U15236 ( .B1(n13330), .B2(n13087), .A(n13056), .ZN(n13057) );
  AOI21_X1 U15237 ( .B1(n13332), .B2(n13095), .A(n13057), .ZN(n13058) );
  OAI21_X1 U15238 ( .B1(n13059), .B2(n13091), .A(n13058), .ZN(P2_U3207) );
  OAI211_X1 U15239 ( .C1(n13063), .C2(n13062), .A(n13061), .B(n13060), .ZN(
        n13070) );
  AOI22_X1 U15240 ( .A1(n13110), .A2(n13065), .B1(n13064), .B2(n13112), .ZN(
        n13392) );
  NAND2_X1 U15241 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14750)
         );
  OAI21_X1 U15242 ( .B1(n13392), .B2(n13066), .A(n14750), .ZN(n13067) );
  AOI21_X1 U15243 ( .B1(n13403), .B2(n13068), .A(n13067), .ZN(n13069) );
  OAI211_X1 U15244 ( .C1(n6936), .C2(n13071), .A(n13070), .B(n13069), .ZN(
        P2_U3210) );
  INV_X1 U15245 ( .A(n13072), .ZN(n13073) );
  AOI21_X1 U15246 ( .B1(n13075), .B2(n13074), .A(n13073), .ZN(n13084) );
  OAI22_X1 U15247 ( .A1(n13079), .A2(n13078), .B1(n13077), .B2(n13076), .ZN(
        n13260) );
  AOI22_X1 U15248 ( .A1(n13085), .A2(n13260), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13080) );
  OAI21_X1 U15249 ( .B1(n13267), .B2(n13087), .A(n13080), .ZN(n13081) );
  AOI21_X1 U15250 ( .B1(n13082), .B2(n13095), .A(n13081), .ZN(n13083) );
  OAI21_X1 U15251 ( .B1(n13084), .B2(n13091), .A(n13083), .ZN(P2_U3212) );
  AOI22_X1 U15252 ( .A1(n13085), .A2(n14421), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13086) );
  OAI21_X1 U15253 ( .B1(n13088), .B2(n13087), .A(n13086), .ZN(n13094) );
  AOI211_X1 U15254 ( .C1(n13089), .C2(n13092), .A(n13091), .B(n13090), .ZN(
        n13093) );
  AOI211_X1 U15255 ( .C1(n13096), .C2(n13095), .A(n13094), .B(n13093), .ZN(
        n13097) );
  INV_X1 U15256 ( .A(n13097), .ZN(P2_U3213) );
  MUX2_X1 U15257 ( .A(n13098), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13121), .Z(
        P2_U3562) );
  MUX2_X1 U15258 ( .A(n13099), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13121), .Z(
        P2_U3561) );
  MUX2_X1 U15259 ( .A(n13100), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13121), .Z(
        P2_U3560) );
  MUX2_X1 U15260 ( .A(n13101), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13121), .Z(
        P2_U3559) );
  MUX2_X1 U15261 ( .A(n13102), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13121), .Z(
        P2_U3558) );
  MUX2_X1 U15262 ( .A(n13103), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13121), .Z(
        P2_U3557) );
  MUX2_X1 U15263 ( .A(n13104), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13121), .Z(
        P2_U3556) );
  MUX2_X1 U15264 ( .A(n13105), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13121), .Z(
        P2_U3555) );
  MUX2_X1 U15265 ( .A(n13106), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13121), .Z(
        P2_U3554) );
  MUX2_X1 U15266 ( .A(n13107), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13121), .Z(
        P2_U3553) );
  MUX2_X1 U15267 ( .A(n13108), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13121), .Z(
        P2_U3552) );
  MUX2_X1 U15268 ( .A(n13109), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13121), .Z(
        P2_U3551) );
  INV_X1 U15269 ( .A(P2_U3947), .ZN(n13130) );
  MUX2_X1 U15270 ( .A(n13110), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13130), .Z(
        P2_U3550) );
  MUX2_X1 U15271 ( .A(n13111), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13121), .Z(
        P2_U3549) );
  MUX2_X1 U15272 ( .A(n13112), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13121), .Z(
        P2_U3548) );
  MUX2_X1 U15273 ( .A(n13113), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13130), .Z(
        P2_U3547) );
  MUX2_X1 U15274 ( .A(n13114), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13121), .Z(
        P2_U3546) );
  MUX2_X1 U15275 ( .A(n13115), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13130), .Z(
        P2_U3545) );
  MUX2_X1 U15276 ( .A(n13116), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13121), .Z(
        P2_U3544) );
  MUX2_X1 U15277 ( .A(n13117), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13130), .Z(
        P2_U3543) );
  MUX2_X1 U15278 ( .A(n13118), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13121), .Z(
        P2_U3542) );
  MUX2_X1 U15279 ( .A(n13119), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13121), .Z(
        P2_U3541) );
  MUX2_X1 U15280 ( .A(n13120), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13121), .Z(
        P2_U3540) );
  MUX2_X1 U15281 ( .A(n13122), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13121), .Z(
        P2_U3539) );
  MUX2_X1 U15282 ( .A(n13123), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13130), .Z(
        P2_U3538) );
  MUX2_X1 U15283 ( .A(n13124), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13130), .Z(
        P2_U3537) );
  MUX2_X1 U15284 ( .A(n13125), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13130), .Z(
        P2_U3536) );
  MUX2_X1 U15285 ( .A(n13126), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13130), .Z(
        P2_U3535) );
  MUX2_X1 U15286 ( .A(n13127), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13130), .Z(
        P2_U3534) );
  MUX2_X1 U15287 ( .A(n13128), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13130), .Z(
        P2_U3533) );
  MUX2_X1 U15288 ( .A(n13129), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13130), .Z(
        P2_U3532) );
  MUX2_X1 U15289 ( .A(n13131), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13130), .Z(
        P2_U3531) );
  NAND2_X1 U15290 ( .A1(n13133), .A2(n13132), .ZN(n13135) );
  MUX2_X1 U15291 ( .A(n13134), .B(P2_REG2_REG_12__SCAN_IN), .S(n13144), .Z(
        n13136) );
  AOI21_X1 U15292 ( .B1(n13137), .B2(n13135), .A(n13136), .ZN(n13151) );
  AND3_X1 U15293 ( .A1(n13137), .A2(n13136), .A3(n13135), .ZN(n13138) );
  OAI21_X1 U15294 ( .B1(n13151), .B2(n13138), .A(n14727), .ZN(n13150) );
  INV_X1 U15295 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n13140) );
  OAI21_X1 U15296 ( .B1(n14752), .B2(n13140), .A(n13139), .ZN(n13141) );
  AOI21_X1 U15297 ( .B1(n13144), .B2(n14741), .A(n13141), .ZN(n13149) );
  AOI21_X1 U15298 ( .B1(n13143), .B2(P2_REG1_REG_11__SCAN_IN), .A(n13142), 
        .ZN(n13146) );
  MUX2_X1 U15299 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8334), .S(n13144), .Z(
        n13145) );
  NOR2_X1 U15300 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  AND2_X1 U15301 ( .A1(n13146), .A2(n13145), .ZN(n13166) );
  OAI21_X1 U15302 ( .B1(n13147), .B2(n13166), .A(n14743), .ZN(n13148) );
  NAND3_X1 U15303 ( .A1(n13150), .A2(n13149), .A3(n13148), .ZN(P2_U3226) );
  AOI21_X1 U15304 ( .B1(n13134), .B2(n13167), .A(n13151), .ZN(n14698) );
  MUX2_X1 U15305 ( .A(n13152), .B(P2_REG2_REG_13__SCAN_IN), .S(n14693), .Z(
        n14697) );
  OAI21_X1 U15306 ( .B1(n13152), .B2(n14693), .A(n14696), .ZN(n13153) );
  NAND2_X1 U15307 ( .A1(n14710), .A2(n13153), .ZN(n13154) );
  XNOR2_X1 U15308 ( .A(n13153), .B(n13170), .ZN(n14709) );
  NAND2_X1 U15309 ( .A1(n14715), .A2(n13155), .ZN(n13156) );
  NAND2_X1 U15310 ( .A1(n14725), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13158) );
  OAI21_X1 U15311 ( .B1(n14725), .B2(P2_REG2_REG_16__SCAN_IN), .A(n13158), 
        .ZN(n13157) );
  INV_X1 U15312 ( .A(n13157), .ZN(n14730) );
  INV_X1 U15313 ( .A(n13158), .ZN(n13162) );
  AOI21_X1 U15314 ( .B1(n13189), .B2(P2_REG2_REG_17__SCAN_IN), .A(n13162), 
        .ZN(n13159) );
  OAI21_X1 U15315 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n13189), .A(n13159), 
        .ZN(n13163) );
  NAND2_X1 U15316 ( .A1(n13177), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13161) );
  INV_X1 U15317 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U15318 ( .A1(n13189), .A2(n13184), .ZN(n13160) );
  OAI211_X1 U15319 ( .C1(n14726), .C2(n13163), .A(n13183), .B(n14727), .ZN(
        n13182) );
  OAI21_X1 U15320 ( .B1(n14752), .B2(n6911), .A(n13164), .ZN(n13165) );
  AOI21_X1 U15321 ( .B1(n13177), .B2(n14741), .A(n13165), .ZN(n13181) );
  AOI21_X1 U15322 ( .B1(n8334), .B2(n13167), .A(n13166), .ZN(n14701) );
  MUX2_X1 U15323 ( .A(n13168), .B(P2_REG1_REG_13__SCAN_IN), .S(n14693), .Z(
        n14700) );
  NAND2_X1 U15324 ( .A1(n14701), .A2(n14700), .ZN(n14699) );
  OAI21_X1 U15325 ( .B1(n13168), .B2(n14693), .A(n14699), .ZN(n14707) );
  MUX2_X1 U15326 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13169), .S(n14710), .Z(
        n14706) );
  NAND2_X1 U15327 ( .A1(n14707), .A2(n14706), .ZN(n14705) );
  OAI21_X1 U15328 ( .B1(n13169), .B2(n13170), .A(n14705), .ZN(n13172) );
  NAND2_X1 U15329 ( .A1(n14715), .A2(n13172), .ZN(n13173) );
  XNOR2_X1 U15330 ( .A(n13172), .B(n13171), .ZN(n14719) );
  NAND2_X1 U15331 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14719), .ZN(n14718) );
  NAND2_X1 U15332 ( .A1(n13173), .A2(n14718), .ZN(n14732) );
  INV_X1 U15333 ( .A(n14732), .ZN(n13176) );
  XNOR2_X1 U15334 ( .A(n14725), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14731) );
  INV_X1 U15335 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13175) );
  OAI22_X1 U15336 ( .A1(n13176), .A2(n14731), .B1(n13175), .B2(n13174), .ZN(
        n13179) );
  AOI22_X1 U15337 ( .A1(n13177), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n13188), 
        .B2(n13189), .ZN(n13178) );
  NAND2_X1 U15338 ( .A1(n13178), .A2(n13179), .ZN(n13187) );
  OAI211_X1 U15339 ( .C1(n13179), .C2(n13178), .A(n13187), .B(n14743), .ZN(
        n13180) );
  NAND3_X1 U15340 ( .A1(n13182), .A2(n13181), .A3(n13180), .ZN(P2_U3231) );
  OAI21_X1 U15341 ( .B1(n13184), .B2(n13189), .A(n13183), .ZN(n13185) );
  NOR2_X1 U15342 ( .A1(n13185), .A2(n14740), .ZN(n13186) );
  NOR2_X1 U15343 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14739), .ZN(n14738) );
  OAI21_X1 U15344 ( .B1(n13189), .B2(n13188), .A(n13187), .ZN(n13190) );
  XOR2_X1 U15345 ( .A(n14740), .B(n13190), .Z(n14744) );
  NAND2_X1 U15346 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14744), .ZN(n14742) );
  NAND2_X1 U15347 ( .A1(n13190), .A2(n14740), .ZN(n13191) );
  NAND2_X1 U15348 ( .A1(n14742), .A2(n13191), .ZN(n13192) );
  XNOR2_X1 U15349 ( .A(n13192), .B(n13472), .ZN(n13195) );
  NOR2_X1 U15350 ( .A1(n13195), .A2(n14668), .ZN(n13193) );
  AOI211_X1 U15351 ( .C1(n13194), .C2(n14727), .A(n14741), .B(n13193), .ZN(
        n13198) );
  AOI22_X1 U15352 ( .A1(n13196), .A2(n14727), .B1(n14743), .B2(n13195), .ZN(
        n13197) );
  OAI211_X1 U15353 ( .C1(n13201), .C2(n14752), .A(n13200), .B(n13199), .ZN(
        P2_U3233) );
  XNOR2_X1 U15354 ( .A(n13209), .B(n8883), .ZN(n13202) );
  NAND2_X1 U15355 ( .A1(n13412), .A2(n13402), .ZN(n13207) );
  NOR2_X1 U15356 ( .A1(n13204), .A2(n13203), .ZN(n13415) );
  INV_X1 U15357 ( .A(n13415), .ZN(n13205) );
  NOR2_X1 U15358 ( .A1(n13411), .A2(n13205), .ZN(n13213) );
  AOI21_X1 U15359 ( .B1(n13411), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13213), 
        .ZN(n13206) );
  OAI211_X1 U15360 ( .C1(n13496), .C2(n13406), .A(n13207), .B(n13206), .ZN(
        P2_U3234) );
  INV_X1 U15361 ( .A(n13208), .ZN(n13211) );
  INV_X1 U15362 ( .A(n13209), .ZN(n13210) );
  AOI211_X1 U15363 ( .C1(n13212), .C2(n13211), .A(n13295), .B(n13210), .ZN(
        n13416) );
  NAND2_X1 U15364 ( .A1(n13416), .A2(n13402), .ZN(n13215) );
  AOI21_X1 U15365 ( .B1(n13411), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13213), 
        .ZN(n13214) );
  OAI211_X1 U15366 ( .C1(n13500), .C2(n13406), .A(n13215), .B(n13214), .ZN(
        P2_U3235) );
  INV_X1 U15367 ( .A(n13216), .ZN(n13226) );
  NAND2_X1 U15368 ( .A1(n13217), .A2(n13336), .ZN(n13225) );
  NOR2_X1 U15369 ( .A1(n13218), .A2(n13406), .ZN(n13222) );
  OAI22_X1 U15370 ( .A1(n13336), .A2(n13220), .B1(n13219), .B2(n13300), .ZN(
        n13221) );
  AOI211_X1 U15371 ( .C1(n13223), .C2(n13402), .A(n13222), .B(n13221), .ZN(
        n13224) );
  OAI211_X1 U15372 ( .C1(n13226), .C2(n13372), .A(n13225), .B(n13224), .ZN(
        P2_U3236) );
  OAI211_X1 U15373 ( .C1(n13502), .C2(n13248), .A(n12001), .B(n13230), .ZN(
        n13419) );
  OAI22_X1 U15374 ( .A1(n13502), .A2(n13406), .B1(n13336), .B2(n13231), .ZN(
        n13232) );
  AOI21_X1 U15375 ( .B1(n6633), .B2(n13402), .A(n13232), .ZN(n13243) );
  NAND2_X1 U15376 ( .A1(n13234), .A2(n13233), .ZN(n13235) );
  NAND3_X1 U15377 ( .A1(n13236), .A2(n14399), .A3(n13235), .ZN(n13239) );
  INV_X1 U15378 ( .A(n13237), .ZN(n13238) );
  OAI21_X1 U15379 ( .B1(n13240), .B2(n13300), .A(n13420), .ZN(n13241) );
  NAND2_X1 U15380 ( .A1(n13241), .A2(n13336), .ZN(n13242) );
  OAI211_X1 U15381 ( .C1(n13421), .C2(n13372), .A(n13243), .B(n13242), .ZN(
        P2_U3237) );
  XNOR2_X1 U15382 ( .A(n13244), .B(n13253), .ZN(n13246) );
  AOI21_X1 U15383 ( .B1(n13246), .B2(n14399), .A(n13245), .ZN(n13427) );
  NOR2_X1 U15384 ( .A1(n13252), .A2(n13266), .ZN(n13247) );
  INV_X1 U15385 ( .A(n13426), .ZN(n13257) );
  NOR2_X1 U15386 ( .A1(n13300), .A2(n13249), .ZN(n13250) );
  AOI21_X1 U15387 ( .B1(n13411), .B2(P2_REG2_REG_27__SCAN_IN), .A(n13250), 
        .ZN(n13251) );
  OAI21_X1 U15388 ( .B1(n13252), .B2(n13406), .A(n13251), .ZN(n13256) );
  OR2_X1 U15389 ( .A1(n13254), .A2(n13253), .ZN(n13423) );
  AND3_X1 U15390 ( .A1(n13423), .A2(n13422), .A3(n14417), .ZN(n13255) );
  AOI211_X1 U15391 ( .C1(n13257), .C2(n13402), .A(n13256), .B(n13255), .ZN(
        n13258) );
  OAI21_X1 U15392 ( .B1(n13411), .B2(n13427), .A(n13258), .ZN(P2_U3238) );
  XNOR2_X1 U15393 ( .A(n13259), .B(n13263), .ZN(n13262) );
  INV_X1 U15394 ( .A(n13260), .ZN(n13261) );
  OAI21_X1 U15395 ( .B1(n13262), .B2(n13393), .A(n13261), .ZN(n13430) );
  INV_X1 U15396 ( .A(n13430), .ZN(n13273) );
  XNOR2_X1 U15397 ( .A(n13264), .B(n13263), .ZN(n13432) );
  NOR2_X1 U15398 ( .A1(n13507), .A2(n13280), .ZN(n13265) );
  NOR2_X1 U15399 ( .A1(n13429), .A2(n14415), .ZN(n13271) );
  NOR2_X1 U15400 ( .A1(n13300), .A2(n13267), .ZN(n13268) );
  AOI21_X1 U15401 ( .B1(n13411), .B2(P2_REG2_REG_26__SCAN_IN), .A(n13268), 
        .ZN(n13269) );
  OAI21_X1 U15402 ( .B1(n13507), .B2(n13406), .A(n13269), .ZN(n13270) );
  AOI211_X1 U15403 ( .C1(n13432), .C2(n14417), .A(n13271), .B(n13270), .ZN(
        n13272) );
  OAI21_X1 U15404 ( .B1(n13411), .B2(n13273), .A(n13272), .ZN(P2_U3239) );
  XNOR2_X1 U15405 ( .A(n13274), .B(n13279), .ZN(n13277) );
  INV_X1 U15406 ( .A(n13275), .ZN(n13276) );
  OAI21_X1 U15407 ( .B1(n13277), .B2(n13393), .A(n13276), .ZN(n13436) );
  INV_X1 U15408 ( .A(n13436), .ZN(n13288) );
  OAI21_X1 U15409 ( .B1(n6586), .B2(n13279), .A(n13278), .ZN(n13438) );
  NOR2_X1 U15410 ( .A1(n13511), .A2(n13297), .ZN(n13281) );
  NOR2_X1 U15411 ( .A1(n13435), .A2(n14415), .ZN(n13286) );
  NOR2_X1 U15412 ( .A1(n13300), .A2(n13282), .ZN(n13283) );
  AOI21_X1 U15413 ( .B1(n13411), .B2(P2_REG2_REG_25__SCAN_IN), .A(n13283), 
        .ZN(n13284) );
  OAI21_X1 U15414 ( .B1(n13511), .B2(n13406), .A(n13284), .ZN(n13285) );
  AOI211_X1 U15415 ( .C1(n13438), .C2(n14417), .A(n13286), .B(n13285), .ZN(
        n13287) );
  OAI21_X1 U15416 ( .B1(n13411), .B2(n13288), .A(n13287), .ZN(P2_U3240) );
  XNOR2_X1 U15417 ( .A(n13289), .B(n13294), .ZN(n13292) );
  INV_X1 U15418 ( .A(n13290), .ZN(n13291) );
  OAI21_X1 U15419 ( .B1(n13292), .B2(n13393), .A(n13291), .ZN(n13443) );
  INV_X1 U15420 ( .A(n13443), .ZN(n13305) );
  XNOR2_X1 U15421 ( .A(n13293), .B(n13294), .ZN(n13445) );
  AND2_X1 U15422 ( .A1(n13441), .A2(n6555), .ZN(n13296) );
  OR3_X1 U15423 ( .A1(n13297), .A2(n13296), .A3(n13295), .ZN(n13442) );
  NAND2_X1 U15424 ( .A1(n13411), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13298) );
  OAI21_X1 U15425 ( .B1(n13300), .B2(n13299), .A(n13298), .ZN(n13301) );
  AOI21_X1 U15426 ( .B1(n13441), .B2(n14403), .A(n13301), .ZN(n13302) );
  OAI21_X1 U15427 ( .B1(n13442), .B2(n14415), .A(n13302), .ZN(n13303) );
  AOI21_X1 U15428 ( .B1(n13445), .B2(n14417), .A(n13303), .ZN(n13304) );
  OAI21_X1 U15429 ( .B1(n13305), .B2(n14420), .A(n13304), .ZN(P2_U3241) );
  INV_X1 U15430 ( .A(n13306), .ZN(n13311) );
  XNOR2_X1 U15431 ( .A(n13307), .B(n13316), .ZN(n13310) );
  INV_X1 U15432 ( .A(n13308), .ZN(n13309) );
  OAI21_X1 U15433 ( .B1(n13310), .B2(n13393), .A(n13309), .ZN(n13448) );
  AOI21_X1 U15434 ( .B1(n13311), .B2(n14402), .A(n13448), .ZN(n13320) );
  INV_X1 U15435 ( .A(n6555), .ZN(n13312) );
  AOI211_X1 U15436 ( .C1(n13313), .C2(n6492), .A(n13295), .B(n13312), .ZN(
        n13449) );
  INV_X1 U15437 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13314) );
  OAI22_X1 U15438 ( .A1(n13519), .A2(n13406), .B1(n13336), .B2(n13314), .ZN(
        n13315) );
  AOI21_X1 U15439 ( .B1(n13449), .B2(n13402), .A(n13315), .ZN(n13319) );
  XNOR2_X1 U15440 ( .A(n13317), .B(n13316), .ZN(n13450) );
  NAND2_X1 U15441 ( .A1(n13450), .A2(n14417), .ZN(n13318) );
  OAI211_X1 U15442 ( .C1(n13320), .C2(n14420), .A(n13319), .B(n13318), .ZN(
        P2_U3242) );
  OAI21_X1 U15443 ( .B1(n13322), .B2(n13323), .A(n13321), .ZN(n13455) );
  AOI21_X1 U15444 ( .B1(n13324), .B2(n13323), .A(n13393), .ZN(n13327) );
  AOI21_X1 U15445 ( .B1(n13327), .B2(n13326), .A(n13325), .ZN(n13454) );
  INV_X1 U15446 ( .A(n13454), .ZN(n13337) );
  INV_X1 U15447 ( .A(n13328), .ZN(n13347) );
  OAI211_X1 U15448 ( .C1(n6930), .C2(n13347), .A(n6492), .B(n12001), .ZN(
        n13453) );
  INV_X1 U15449 ( .A(n13330), .ZN(n13331) );
  AOI22_X1 U15450 ( .A1(n13411), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13331), 
        .B2(n14402), .ZN(n13334) );
  NAND2_X1 U15451 ( .A1(n13332), .A2(n14403), .ZN(n13333) );
  OAI211_X1 U15452 ( .C1(n13453), .C2(n14415), .A(n13334), .B(n13333), .ZN(
        n13335) );
  AOI21_X1 U15453 ( .B1(n13337), .B2(n13336), .A(n13335), .ZN(n13338) );
  OAI21_X1 U15454 ( .B1(n13372), .B2(n13455), .A(n13338), .ZN(P2_U3243) );
  XNOR2_X1 U15455 ( .A(n13340), .B(n13339), .ZN(n13461) );
  INV_X1 U15456 ( .A(n13461), .ZN(n13354) );
  OAI21_X1 U15457 ( .B1(n13343), .B2(n13342), .A(n13341), .ZN(n13344) );
  NAND2_X1 U15458 ( .A1(n13344), .A2(n14399), .ZN(n13346) );
  NAND2_X1 U15459 ( .A1(n13346), .A2(n13345), .ZN(n13459) );
  INV_X1 U15460 ( .A(n13348), .ZN(n13526) );
  AOI211_X1 U15461 ( .C1(n13348), .C2(n13357), .A(n13295), .B(n13347), .ZN(
        n13460) );
  NAND2_X1 U15462 ( .A1(n13460), .A2(n13402), .ZN(n13351) );
  AOI22_X1 U15463 ( .A1(n13349), .A2(n14402), .B1(n13411), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13350) );
  OAI211_X1 U15464 ( .C1(n13526), .C2(n13406), .A(n13351), .B(n13350), .ZN(
        n13352) );
  AOI21_X1 U15465 ( .B1(n13459), .B2(n13336), .A(n13352), .ZN(n13353) );
  OAI21_X1 U15466 ( .B1(n13354), .B2(n13372), .A(n13353), .ZN(P2_U3244) );
  XNOR2_X1 U15467 ( .A(n13356), .B(n13355), .ZN(n13468) );
  INV_X1 U15468 ( .A(n13381), .ZN(n13359) );
  INV_X1 U15469 ( .A(n13357), .ZN(n13358) );
  AOI211_X1 U15470 ( .C1(n13465), .C2(n13359), .A(n13295), .B(n13358), .ZN(
        n13464) );
  AOI22_X1 U15471 ( .A1(n13360), .A2(n14402), .B1(n13411), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n13361) );
  OAI21_X1 U15472 ( .B1(n13362), .B2(n13406), .A(n13361), .ZN(n13370) );
  OAI21_X1 U15473 ( .B1(n13365), .B2(n13364), .A(n13363), .ZN(n13368) );
  INV_X1 U15474 ( .A(n13366), .ZN(n13367) );
  AOI21_X1 U15475 ( .B1(n13368), .B2(n14399), .A(n13367), .ZN(n13467) );
  NOR2_X1 U15476 ( .A1(n13467), .A2(n13411), .ZN(n13369) );
  AOI211_X1 U15477 ( .C1(n13464), .C2(n13402), .A(n13370), .B(n13369), .ZN(
        n13371) );
  OAI21_X1 U15478 ( .B1(n13372), .B2(n13468), .A(n13371), .ZN(P2_U3245) );
  XNOR2_X1 U15479 ( .A(n13373), .B(n13377), .ZN(n13471) );
  INV_X1 U15480 ( .A(n13471), .ZN(n13390) );
  INV_X1 U15481 ( .A(n13374), .ZN(n13375) );
  AOI21_X1 U15482 ( .B1(n13377), .B2(n13376), .A(n13375), .ZN(n13380) );
  NAND2_X1 U15483 ( .A1(n13471), .A2(n14810), .ZN(n13378) );
  OAI211_X1 U15484 ( .C1(n13380), .C2(n13393), .A(n13379), .B(n13378), .ZN(
        n13469) );
  NAND2_X1 U15485 ( .A1(n13469), .A2(n13336), .ZN(n13388) );
  AOI211_X1 U15486 ( .C1(n13383), .C2(n13400), .A(n13295), .B(n13381), .ZN(
        n13470) );
  AOI22_X1 U15487 ( .A1(n13411), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13384), 
        .B2(n14402), .ZN(n13385) );
  OAI21_X1 U15488 ( .B1(n13532), .B2(n13406), .A(n13385), .ZN(n13386) );
  AOI21_X1 U15489 ( .B1(n13470), .B2(n13402), .A(n13386), .ZN(n13387) );
  OAI211_X1 U15490 ( .C1(n13390), .C2(n13389), .A(n13388), .B(n13387), .ZN(
        P2_U3246) );
  XNOR2_X1 U15491 ( .A(n13391), .B(n13398), .ZN(n13394) );
  OAI21_X1 U15492 ( .B1(n13394), .B2(n13393), .A(n13392), .ZN(n13475) );
  INV_X1 U15493 ( .A(n13475), .ZN(n13410) );
  INV_X1 U15494 ( .A(n13395), .ZN(n13396) );
  AOI21_X1 U15495 ( .B1(n13398), .B2(n13397), .A(n13396), .ZN(n13479) );
  INV_X1 U15496 ( .A(n13479), .ZN(n13408) );
  AOI21_X1 U15497 ( .B1(n13399), .B2(n13477), .A(n13295), .ZN(n13401) );
  AND2_X1 U15498 ( .A1(n13401), .A2(n13400), .ZN(n13476) );
  NAND2_X1 U15499 ( .A1(n13476), .A2(n13402), .ZN(n13405) );
  AOI22_X1 U15500 ( .A1(n13411), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13403), 
        .B2(n14402), .ZN(n13404) );
  OAI211_X1 U15501 ( .C1(n6936), .C2(n13406), .A(n13405), .B(n13404), .ZN(
        n13407) );
  AOI21_X1 U15502 ( .B1(n13408), .B2(n14417), .A(n13407), .ZN(n13409) );
  OAI21_X1 U15503 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(P2_U3247) );
  NOR2_X1 U15504 ( .A1(n13412), .A2(n13415), .ZN(n13493) );
  MUX2_X1 U15505 ( .A(n13413), .B(n13493), .S(n14842), .Z(n13414) );
  OAI21_X1 U15506 ( .B1(n13496), .B2(n13474), .A(n13414), .ZN(P2_U3530) );
  INV_X1 U15507 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13417) );
  NOR2_X1 U15508 ( .A1(n13416), .A2(n13415), .ZN(n13497) );
  MUX2_X1 U15509 ( .A(n13417), .B(n13497), .S(n14842), .Z(n13418) );
  OAI21_X1 U15510 ( .B1(n13500), .B2(n13474), .A(n13418), .ZN(P2_U3529) );
  NAND3_X1 U15511 ( .A1(n13423), .A2(n14816), .A3(n13422), .ZN(n13428) );
  NAND2_X1 U15512 ( .A1(n13424), .A2(n14819), .ZN(n13425) );
  NAND4_X1 U15513 ( .A1(n13428), .A2(n13427), .A3(n13426), .A4(n13425), .ZN(
        n13503) );
  MUX2_X1 U15514 ( .A(n13503), .B(P2_REG1_REG_27__SCAN_IN), .S(n8665), .Z(
        P2_U3526) );
  INV_X1 U15515 ( .A(n13429), .ZN(n13431) );
  AOI211_X1 U15516 ( .C1(n13432), .C2(n14816), .A(n13431), .B(n13430), .ZN(
        n13504) );
  MUX2_X1 U15517 ( .A(n13433), .B(n13504), .S(n14842), .Z(n13434) );
  OAI21_X1 U15518 ( .B1(n13507), .B2(n13474), .A(n13434), .ZN(P2_U3525) );
  INV_X1 U15519 ( .A(n13435), .ZN(n13437) );
  AOI211_X1 U15520 ( .C1(n14816), .C2(n13438), .A(n13437), .B(n13436), .ZN(
        n13508) );
  MUX2_X1 U15521 ( .A(n13439), .B(n13508), .S(n14842), .Z(n13440) );
  OAI21_X1 U15522 ( .B1(n13511), .B2(n13474), .A(n13440), .ZN(P2_U3524) );
  INV_X1 U15523 ( .A(n13441), .ZN(n13515) );
  INV_X1 U15524 ( .A(n13442), .ZN(n13444) );
  AOI211_X1 U15525 ( .C1(n13445), .C2(n14816), .A(n13444), .B(n13443), .ZN(
        n13512) );
  MUX2_X1 U15526 ( .A(n13446), .B(n13512), .S(n14842), .Z(n13447) );
  OAI21_X1 U15527 ( .B1(n13515), .B2(n13474), .A(n13447), .ZN(P2_U3523) );
  AOI211_X1 U15528 ( .C1(n14816), .C2(n13450), .A(n13449), .B(n13448), .ZN(
        n13516) );
  MUX2_X1 U15529 ( .A(n13451), .B(n13516), .S(n14842), .Z(n13452) );
  OAI21_X1 U15530 ( .B1(n13519), .B2(n13474), .A(n13452), .ZN(P2_U3522) );
  OAI211_X1 U15531 ( .C1(n13455), .C2(n13485), .A(n13454), .B(n13453), .ZN(
        n13456) );
  INV_X1 U15532 ( .A(n13456), .ZN(n13520) );
  MUX2_X1 U15533 ( .A(n13457), .B(n13520), .S(n14842), .Z(n13458) );
  OAI21_X1 U15534 ( .B1(n6930), .B2(n13474), .A(n13458), .ZN(P2_U3521) );
  INV_X1 U15535 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13462) );
  AOI211_X1 U15536 ( .C1(n13461), .C2(n14816), .A(n13460), .B(n13459), .ZN(
        n13523) );
  MUX2_X1 U15537 ( .A(n13462), .B(n13523), .S(n14842), .Z(n13463) );
  OAI21_X1 U15538 ( .B1(n13526), .B2(n13474), .A(n13463), .ZN(P2_U3520) );
  AOI21_X1 U15539 ( .B1(n14819), .B2(n13465), .A(n13464), .ZN(n13466) );
  OAI211_X1 U15540 ( .C1(n13468), .C2(n13485), .A(n13467), .B(n13466), .ZN(
        n13527) );
  MUX2_X1 U15541 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13527), .S(n14842), .Z(
        P2_U3519) );
  AOI211_X1 U15542 ( .C1(n14835), .C2(n13471), .A(n13470), .B(n13469), .ZN(
        n13528) );
  MUX2_X1 U15543 ( .A(n13472), .B(n13528), .S(n14842), .Z(n13473) );
  OAI21_X1 U15544 ( .B1(n13532), .B2(n13474), .A(n13473), .ZN(P2_U3518) );
  AOI211_X1 U15545 ( .C1(n14819), .C2(n13477), .A(n13476), .B(n13475), .ZN(
        n13478) );
  OAI21_X1 U15546 ( .B1(n13485), .B2(n13479), .A(n13478), .ZN(n13533) );
  MUX2_X1 U15547 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13533), .S(n14842), .Z(
        P2_U3517) );
  AOI211_X1 U15548 ( .C1(n14819), .C2(n13482), .A(n13481), .B(n13480), .ZN(
        n13483) );
  OAI21_X1 U15549 ( .B1(n13485), .B2(n13484), .A(n13483), .ZN(n13534) );
  MUX2_X1 U15550 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13534), .S(n14842), .Z(
        P2_U3516) );
  AOI211_X1 U15551 ( .C1(n14819), .C2(n13488), .A(n13487), .B(n13486), .ZN(
        n13492) );
  NAND3_X1 U15552 ( .A1(n13490), .A2(n14816), .A3(n13489), .ZN(n13491) );
  NAND2_X1 U15553 ( .A1(n13492), .A2(n13491), .ZN(n13535) );
  MUX2_X1 U15554 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13535), .S(n14842), .Z(
        P2_U3515) );
  MUX2_X1 U15555 ( .A(n13494), .B(n13493), .S(n14836), .Z(n13495) );
  OAI21_X1 U15556 ( .B1(n13496), .B2(n13531), .A(n13495), .ZN(P2_U3498) );
  INV_X1 U15557 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13498) );
  MUX2_X1 U15558 ( .A(n13498), .B(n13497), .S(n14836), .Z(n13499) );
  OAI21_X1 U15559 ( .B1(n13500), .B2(n13531), .A(n13499), .ZN(P2_U3497) );
  MUX2_X1 U15560 ( .A(n13503), .B(P2_REG0_REG_27__SCAN_IN), .S(n7143), .Z(
        P2_U3494) );
  MUX2_X1 U15561 ( .A(n13505), .B(n13504), .S(n14836), .Z(n13506) );
  OAI21_X1 U15562 ( .B1(n13507), .B2(n13531), .A(n13506), .ZN(P2_U3493) );
  MUX2_X1 U15563 ( .A(n13509), .B(n13508), .S(n14836), .Z(n13510) );
  OAI21_X1 U15564 ( .B1(n13511), .B2(n13531), .A(n13510), .ZN(P2_U3492) );
  MUX2_X1 U15565 ( .A(n13513), .B(n13512), .S(n14836), .Z(n13514) );
  OAI21_X1 U15566 ( .B1(n13515), .B2(n13531), .A(n13514), .ZN(P2_U3491) );
  MUX2_X1 U15567 ( .A(n13517), .B(n13516), .S(n14836), .Z(n13518) );
  OAI21_X1 U15568 ( .B1(n13519), .B2(n13531), .A(n13518), .ZN(P2_U3490) );
  MUX2_X1 U15569 ( .A(n13521), .B(n13520), .S(n14836), .Z(n13522) );
  OAI21_X1 U15570 ( .B1(n6930), .B2(n13531), .A(n13522), .ZN(P2_U3489) );
  INV_X1 U15571 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13524) );
  MUX2_X1 U15572 ( .A(n13524), .B(n13523), .S(n14836), .Z(n13525) );
  OAI21_X1 U15573 ( .B1(n13526), .B2(n13531), .A(n13525), .ZN(P2_U3488) );
  MUX2_X1 U15574 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13527), .S(n14836), .Z(
        P2_U3487) );
  INV_X1 U15575 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13529) );
  MUX2_X1 U15576 ( .A(n13529), .B(n13528), .S(n14836), .Z(n13530) );
  OAI21_X1 U15577 ( .B1(n13532), .B2(n13531), .A(n13530), .ZN(P2_U3486) );
  MUX2_X1 U15578 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13533), .S(n14836), .Z(
        P2_U3484) );
  MUX2_X1 U15579 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13534), .S(n14836), .Z(
        P2_U3481) );
  MUX2_X1 U15580 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13535), .S(n14836), .Z(
        P2_U3478) );
  INV_X1 U15581 ( .A(n13536), .ZN(n14151) );
  NOR4_X1 U15582 ( .A1(n6838), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8154), .A4(
        P2_U3088), .ZN(n13537) );
  AOI21_X1 U15583 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13543), .A(n13537), 
        .ZN(n13538) );
  OAI21_X1 U15584 ( .B1(n14151), .B2(n13552), .A(n13538), .ZN(P2_U3296) );
  INV_X1 U15585 ( .A(n13539), .ZN(n14153) );
  OAI222_X1 U15586 ( .A1(n13552), .A2(n14153), .B1(P2_U3088), .B2(n13541), 
        .C1(n13540), .C2(n13550), .ZN(P2_U3298) );
  AOI21_X1 U15587 ( .B1(n13543), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13542), 
        .ZN(n13544) );
  OAI21_X1 U15588 ( .B1(n13545), .B2(n13552), .A(n13544), .ZN(P2_U3299) );
  INV_X1 U15589 ( .A(n13546), .ZN(n14156) );
  OAI222_X1 U15590 ( .A1(n13550), .A2(n13548), .B1(n13559), .B2(n14156), .C1(
        n13547), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15591 ( .A(n13549), .ZN(n14159) );
  OAI222_X1 U15592 ( .A1(n13553), .A2(P2_U3088), .B1(n13552), .B2(n14159), 
        .C1(n13551), .C2(n13550), .ZN(P2_U3301) );
  INV_X1 U15593 ( .A(n13554), .ZN(n14162) );
  OAI222_X1 U15594 ( .A1(n13550), .A2(n13556), .B1(n13559), .B2(n14162), .C1(
        n13555), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15595 ( .A(n13557), .ZN(n14165) );
  OAI222_X1 U15596 ( .A1(n13550), .A2(n13560), .B1(n13559), .B2(n14165), .C1(
        n13558), .C2(P2_U3088), .ZN(P2_U3303) );
  MUX2_X1 U15597 ( .A(n13561), .B(n14663), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  AOI22_X1 U15598 ( .A1(n13681), .A2(n13702), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13565) );
  OAI21_X1 U15599 ( .B1(n13603), .B2(n14477), .A(n13565), .ZN(n13566) );
  AOI21_X1 U15600 ( .B1(n13567), .B2(n13695), .A(n13566), .ZN(n13568) );
  INV_X1 U15601 ( .A(n13570), .ZN(n13571) );
  NOR2_X1 U15602 ( .A1(n13572), .A2(n13571), .ZN(n13575) );
  INV_X1 U15603 ( .A(n13574), .ZN(n13628) );
  AOI21_X1 U15604 ( .B1(n13575), .B2(n13573), .A(n13628), .ZN(n13582) );
  NOR2_X1 U15605 ( .A1(n13943), .A2(n14634), .ZN(n14099) );
  NAND2_X1 U15606 ( .A1(n13706), .A2(n14006), .ZN(n13577) );
  NAND2_X1 U15607 ( .A1(n13704), .A2(n14008), .ZN(n13576) );
  NAND2_X1 U15608 ( .A1(n13577), .A2(n13576), .ZN(n14098) );
  AOI22_X1 U15609 ( .A1(n14098), .A2(n13658), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13578) );
  OAI21_X1 U15610 ( .B1(n14494), .B2(n13944), .A(n13578), .ZN(n13579) );
  AOI21_X1 U15611 ( .B1(n14099), .B2(n13580), .A(n13579), .ZN(n13581) );
  OAI21_X1 U15612 ( .B1(n13582), .B2(n14467), .A(n13581), .ZN(P1_U3216) );
  INV_X1 U15613 ( .A(n13583), .ZN(n13586) );
  OAI21_X1 U15614 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13588) );
  NAND3_X1 U15615 ( .A1(n13588), .A2(n14483), .A3(n13587), .ZN(n13592) );
  NOR2_X1 U15616 ( .A1(n14494), .A2(n14012), .ZN(n13590) );
  NAND2_X1 U15617 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13846)
         );
  OAI21_X1 U15618 ( .B1(n13598), .B2(n14478), .A(n13846), .ZN(n13589) );
  AOI211_X1 U15619 ( .C1(n13673), .C2(n14007), .A(n13590), .B(n13589), .ZN(
        n13591) );
  OAI211_X1 U15620 ( .C1(n6888), .C2(n13699), .A(n13592), .B(n13591), .ZN(
        P1_U3219) );
  INV_X1 U15621 ( .A(n13593), .ZN(n13594) );
  AOI21_X1 U15622 ( .B1(n13596), .B2(n13595), .A(n13594), .ZN(n13602) );
  OAI22_X1 U15623 ( .A1(n13598), .A2(n14021), .B1(n13597), .B2(n14045), .ZN(
        n13978) );
  AOI22_X1 U15624 ( .A1(n13978), .A2(n13658), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13599) );
  OAI21_X1 U15625 ( .B1(n14494), .B2(n13972), .A(n13599), .ZN(n13600) );
  AOI21_X1 U15626 ( .B1(n14109), .B2(n14490), .A(n13600), .ZN(n13601) );
  OAI21_X1 U15627 ( .B1(n13602), .B2(n14467), .A(n13601), .ZN(P1_U3223) );
  OAI22_X1 U15628 ( .A1(n13604), .A2(n14021), .B1(n13603), .B2(n14045), .ZN(
        n13905) );
  AOI22_X1 U15629 ( .A1(n13905), .A2(n13658), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13605) );
  OAI21_X1 U15630 ( .B1(n14494), .B2(n13908), .A(n13605), .ZN(n13613) );
  INV_X1 U15631 ( .A(n13607), .ZN(n13608) );
  NAND3_X1 U15632 ( .A1(n13606), .A2(n13609), .A3(n13608), .ZN(n13610) );
  AOI21_X1 U15633 ( .B1(n13611), .B2(n13610), .A(n14467), .ZN(n13612) );
  INV_X1 U15634 ( .A(n13614), .ZN(P1_U3225) );
  NAND2_X1 U15635 ( .A1(n13617), .A2(n13616), .ZN(n13618) );
  XNOR2_X1 U15636 ( .A(n13615), .B(n13618), .ZN(n13625) );
  AOI22_X1 U15637 ( .A1(n14007), .A2(n13681), .B1(P1_REG3_REG_17__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13620) );
  NAND2_X1 U15638 ( .A1(n13673), .A2(n13708), .ZN(n13619) );
  OAI211_X1 U15639 ( .C1(n14494), .C2(n13621), .A(n13620), .B(n13619), .ZN(
        n13622) );
  AOI21_X1 U15640 ( .B1(n13623), .B2(n14490), .A(n13622), .ZN(n13624) );
  OAI21_X1 U15641 ( .B1(n13625), .B2(n14467), .A(n13624), .ZN(P1_U3228) );
  NAND2_X1 U15642 ( .A1(n13928), .A2(n14124), .ZN(n14089) );
  NOR3_X1 U15643 ( .A1(n13628), .A2(n7158), .A3(n13627), .ZN(n13630) );
  INV_X1 U15644 ( .A(n13606), .ZN(n13629) );
  OAI21_X1 U15645 ( .B1(n13630), .B2(n13629), .A(n14483), .ZN(n13635) );
  INV_X1 U15646 ( .A(n13631), .ZN(n13927) );
  AOI22_X1 U15647 ( .A1(n13705), .A2(n14006), .B1(n14008), .B2(n13886), .ZN(
        n13921) );
  INV_X1 U15648 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13632) );
  OAI22_X1 U15649 ( .A1(n13921), .A2(n13692), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13632), .ZN(n13633) );
  AOI21_X1 U15650 ( .B1(n13927), .B2(n13695), .A(n13633), .ZN(n13634) );
  OAI211_X1 U15651 ( .C1(n13636), .C2(n14089), .A(n13635), .B(n13634), .ZN(
        P1_U3229) );
  XNOR2_X1 U15652 ( .A(n13637), .B(n13638), .ZN(n13644) );
  INV_X1 U15653 ( .A(n13989), .ZN(n13641) );
  NAND2_X1 U15654 ( .A1(n13984), .A2(n13673), .ZN(n13640) );
  AOI22_X1 U15655 ( .A1(n13681), .A2(n13983), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13639) );
  OAI211_X1 U15656 ( .C1(n14494), .C2(n13641), .A(n13640), .B(n13639), .ZN(
        n13642) );
  AOI21_X1 U15657 ( .B1(n14115), .B2(n14490), .A(n13642), .ZN(n13643) );
  OAI21_X1 U15658 ( .B1(n13644), .B2(n14467), .A(n13643), .ZN(P1_U3233) );
  OAI211_X1 U15659 ( .C1(n13647), .C2(n13646), .A(n13645), .B(n14483), .ZN(
        n13654) );
  INV_X1 U15660 ( .A(n13648), .ZN(n13652) );
  OAI22_X1 U15661 ( .A1(n13650), .A2(n13692), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13649), .ZN(n13651) );
  AOI21_X1 U15662 ( .B1(n13652), .B2(n13695), .A(n13651), .ZN(n13653) );
  OAI211_X1 U15663 ( .C1(n13655), .C2(n13699), .A(n13654), .B(n13653), .ZN(
        P1_U3234) );
  OAI22_X1 U15664 ( .A1(n13657), .A2(n14045), .B1(n13656), .B2(n14021), .ZN(
        n13961) );
  AOI22_X1 U15665 ( .A1(n13961), .A2(n13658), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13659) );
  OAI21_X1 U15666 ( .B1(n14494), .B2(n13963), .A(n13659), .ZN(n13665) );
  INV_X1 U15667 ( .A(n13660), .ZN(n13661) );
  NAND3_X1 U15668 ( .A1(n13593), .A2(n13662), .A3(n13661), .ZN(n13663) );
  AOI21_X1 U15669 ( .B1(n13573), .B2(n13663), .A(n14467), .ZN(n13664) );
  AOI211_X1 U15670 ( .C1(n14490), .C2(n14104), .A(n13665), .B(n13664), .ZN(
        n13666) );
  INV_X1 U15671 ( .A(n13666), .ZN(P1_U3235) );
  INV_X1 U15672 ( .A(n14125), .ZN(n14036) );
  OAI21_X1 U15673 ( .B1(n13668), .B2(n13667), .A(n13583), .ZN(n13669) );
  NAND2_X1 U15674 ( .A1(n13669), .A2(n14483), .ZN(n13675) );
  NOR2_X1 U15675 ( .A1(n14494), .A2(n14032), .ZN(n13672) );
  OAI21_X1 U15676 ( .B1(n14022), .B2(n14478), .A(n13670), .ZN(n13671) );
  AOI211_X1 U15677 ( .C1(n13673), .C2(n13707), .A(n13672), .B(n13671), .ZN(
        n13674) );
  OAI211_X1 U15678 ( .C1(n14036), .C2(n13699), .A(n13675), .B(n13674), .ZN(
        P1_U3238) );
  OAI21_X1 U15679 ( .B1(n13678), .B2(n13677), .A(n13676), .ZN(n13679) );
  NAND2_X1 U15680 ( .A1(n13679), .A2(n14483), .ZN(n13686) );
  INV_X1 U15681 ( .A(n13680), .ZN(n13890) );
  INV_X1 U15682 ( .A(n13886), .ZN(n13683) );
  AOI22_X1 U15683 ( .A1(n13681), .A2(n13887), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13682) );
  OAI21_X1 U15684 ( .B1(n13683), .B2(n14477), .A(n13682), .ZN(n13684) );
  AOI21_X1 U15685 ( .B1(n13890), .B2(n13695), .A(n13684), .ZN(n13685) );
  OAI211_X1 U15686 ( .C1(n13892), .C2(n13699), .A(n13686), .B(n13685), .ZN(
        P1_U3240) );
  OAI211_X1 U15687 ( .C1(n13690), .C2(n13689), .A(n13688), .B(n14483), .ZN(
        n13698) );
  OAI22_X1 U15688 ( .A1(n13693), .A2(n13692), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13691), .ZN(n13694) );
  AOI21_X1 U15689 ( .B1(n13696), .B2(n13695), .A(n13694), .ZN(n13697) );
  OAI211_X1 U15690 ( .C1(n13700), .C2(n13699), .A(n13698), .B(n13697), .ZN(
        P1_U3241) );
  MUX2_X1 U15691 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13851), .S(n13728), .Z(
        P1_U3591) );
  MUX2_X1 U15692 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13701), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15693 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13862), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15694 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13702), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15695 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13887), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15696 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13703), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15697 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13886), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15698 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13704), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15699 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13705), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15700 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13706), .S(n13728), .Z(
        P1_U3582) );
  MUX2_X1 U15701 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13983), .S(n13728), .Z(
        P1_U3581) );
  MUX2_X1 U15702 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14009), .S(n13728), .Z(
        P1_U3580) );
  MUX2_X1 U15703 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13984), .S(n13728), .Z(
        P1_U3579) );
  MUX2_X1 U15704 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14007), .S(n13728), .Z(
        P1_U3578) );
  MUX2_X1 U15705 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13707), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15706 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13708), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15707 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13709), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15708 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13710), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15709 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13711), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15710 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13712), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15711 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13713), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15712 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13714), .S(n13728), .Z(
        P1_U3570) );
  MUX2_X1 U15713 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13715), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15714 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13716), .S(n13728), .Z(
        P1_U3568) );
  MUX2_X1 U15715 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13717), .S(n13728), .Z(
        P1_U3567) );
  MUX2_X1 U15716 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13718), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15717 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13719), .S(n13728), .Z(
        P1_U3565) );
  MUX2_X1 U15718 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13720), .S(n13728), .Z(
        P1_U3564) );
  MUX2_X1 U15719 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n6478), .S(n13728), .Z(
        P1_U3563) );
  MUX2_X1 U15720 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13721), .S(n13728), .Z(
        P1_U3562) );
  MUX2_X1 U15721 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13722), .S(n13728), .Z(
        P1_U3561) );
  MUX2_X1 U15722 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13723), .S(n13728), .Z(
        P1_U3560) );
  AOI21_X1 U15723 ( .B1(n14546), .B2(n9793), .A(n8098), .ZN(n14545) );
  MUX2_X1 U15724 ( .A(n13725), .B(n13724), .S(n14157), .Z(n13727) );
  NAND2_X1 U15725 ( .A1(n13727), .A2(n13726), .ZN(n13729) );
  OAI211_X1 U15726 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14545), .A(n13729), .B(
        n13728), .ZN(n13771) );
  OAI22_X1 U15727 ( .A1(n14566), .A2(n6654), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13730), .ZN(n13731) );
  AOI21_X1 U15728 ( .B1(n13732), .B2(n14573), .A(n13731), .ZN(n13741) );
  NAND2_X1 U15729 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  NAND3_X1 U15730 ( .A1(n14560), .A2(n13744), .A3(n13735), .ZN(n13740) );
  OAI211_X1 U15731 ( .C1(n13738), .C2(n13737), .A(n14575), .B(n13736), .ZN(
        n13739) );
  NAND4_X1 U15732 ( .A1(n13771), .A2(n13741), .A3(n13740), .A4(n13739), .ZN(
        P1_U3245) );
  INV_X1 U15733 ( .A(n13767), .ZN(n13746) );
  NAND3_X1 U15734 ( .A1(n13744), .A2(n13743), .A3(n13742), .ZN(n13745) );
  NAND3_X1 U15735 ( .A1(n14560), .A2(n13746), .A3(n13745), .ZN(n13754) );
  OAI211_X1 U15736 ( .C1(n13749), .C2(n13748), .A(n14575), .B(n13747), .ZN(
        n13753) );
  AOI22_X1 U15737 ( .A1(n14570), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13752) );
  NAND2_X1 U15738 ( .A1(n14573), .A2(n13750), .ZN(n13751) );
  NAND4_X1 U15739 ( .A1(n13754), .A2(n13753), .A3(n13752), .A4(n13751), .ZN(
        P1_U3246) );
  INV_X1 U15740 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n13756) );
  OAI21_X1 U15741 ( .B1(n14566), .B2(n13756), .A(n13755), .ZN(n13757) );
  AOI21_X1 U15742 ( .B1(n13762), .B2(n14573), .A(n13757), .ZN(n13770) );
  OAI211_X1 U15743 ( .C1(n13760), .C2(n13759), .A(n14575), .B(n13758), .ZN(
        n13769) );
  INV_X1 U15744 ( .A(n13761), .ZN(n13764) );
  MUX2_X1 U15745 ( .A(n10402), .B(P1_REG2_REG_4__SCAN_IN), .S(n13762), .Z(
        n13763) );
  NAND2_X1 U15746 ( .A1(n13764), .A2(n13763), .ZN(n13766) );
  OAI211_X1 U15747 ( .C1(n13767), .C2(n13766), .A(n14560), .B(n13765), .ZN(
        n13768) );
  NAND4_X1 U15748 ( .A1(n13771), .A2(n13770), .A3(n13769), .A4(n13768), .ZN(
        P1_U3247) );
  NOR2_X1 U15749 ( .A1(n13838), .A2(n13772), .ZN(n13773) );
  AOI211_X1 U15750 ( .C1(n14570), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n13774), .B(
        n13773), .ZN(n13787) );
  OAI211_X1 U15751 ( .C1(n13777), .C2(n13776), .A(n14575), .B(n13775), .ZN(
        n13786) );
  MUX2_X1 U15752 ( .A(n10652), .B(P1_REG2_REG_6__SCAN_IN), .S(n13778), .Z(
        n13781) );
  INV_X1 U15753 ( .A(n13779), .ZN(n13780) );
  NAND2_X1 U15754 ( .A1(n13781), .A2(n13780), .ZN(n13783) );
  OAI211_X1 U15755 ( .C1(n13784), .C2(n13783), .A(n13782), .B(n14560), .ZN(
        n13785) );
  NAND3_X1 U15756 ( .A1(n13787), .A2(n13786), .A3(n13785), .ZN(P1_U3249) );
  MUX2_X1 U15757 ( .A(n10191), .B(P1_REG2_REG_10__SCAN_IN), .S(n13788), .Z(
        n13791) );
  INV_X1 U15758 ( .A(n13789), .ZN(n13790) );
  NAND2_X1 U15759 ( .A1(n13791), .A2(n13790), .ZN(n13793) );
  OAI211_X1 U15760 ( .C1(n13794), .C2(n13793), .A(n13792), .B(n14560), .ZN(
        n13804) );
  INV_X1 U15761 ( .A(n13795), .ZN(n13798) );
  NOR2_X1 U15762 ( .A1(n13838), .A2(n13796), .ZN(n13797) );
  AOI211_X1 U15763 ( .C1(n14570), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n13798), 
        .B(n13797), .ZN(n13803) );
  OAI211_X1 U15764 ( .C1(n13801), .C2(n13800), .A(n13799), .B(n14575), .ZN(
        n13802) );
  NAND3_X1 U15765 ( .A1(n13804), .A2(n13803), .A3(n13802), .ZN(P1_U3253) );
  NAND2_X1 U15766 ( .A1(n13809), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13805) );
  OAI21_X1 U15767 ( .B1(n13809), .B2(P1_REG2_REG_16__SCAN_IN), .A(n13805), 
        .ZN(n13807) );
  OAI211_X1 U15768 ( .C1(n13808), .C2(n13807), .A(n13806), .B(n14560), .ZN(
        n13817) );
  NAND2_X1 U15769 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14473)
         );
  INV_X1 U15770 ( .A(n14473), .ZN(n13811) );
  NOR2_X1 U15771 ( .A1(n13838), .A2(n13809), .ZN(n13810) );
  AOI211_X1 U15772 ( .C1(n14570), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n13811), 
        .B(n13810), .ZN(n13816) );
  OAI211_X1 U15773 ( .C1(n13814), .C2(n13813), .A(n13812), .B(n14575), .ZN(
        n13815) );
  NAND3_X1 U15774 ( .A1(n13817), .A2(n13816), .A3(n13815), .ZN(P1_U3259) );
  OAI211_X1 U15775 ( .C1(n13820), .C2(n13819), .A(n14560), .B(n13818), .ZN(
        n13829) );
  AND2_X1 U15776 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13823) );
  NOR2_X1 U15777 ( .A1(n13838), .A2(n13821), .ZN(n13822) );
  AOI211_X1 U15778 ( .C1(n14570), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13823), 
        .B(n13822), .ZN(n13828) );
  OAI211_X1 U15779 ( .C1(n13826), .C2(n13825), .A(n13824), .B(n14575), .ZN(
        n13827) );
  NAND3_X1 U15780 ( .A1(n13829), .A2(n13828), .A3(n13827), .ZN(P1_U3260) );
  NOR2_X1 U15781 ( .A1(n13831), .A2(n13830), .ZN(n13832) );
  XNOR2_X1 U15782 ( .A(n13832), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13842) );
  INV_X1 U15783 ( .A(n13842), .ZN(n13840) );
  NAND2_X1 U15784 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  NAND2_X1 U15785 ( .A1(n13836), .A2(n13835), .ZN(n13837) );
  XOR2_X1 U15786 ( .A(n13837), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13841) );
  OAI21_X1 U15787 ( .B1(n13841), .B2(n14579), .A(n13838), .ZN(n13839) );
  AOI21_X1 U15788 ( .B1(n13840), .B2(n14575), .A(n13839), .ZN(n13845) );
  AOI22_X1 U15789 ( .A1(n13842), .A2(n14575), .B1(n14560), .B2(n13841), .ZN(
        n13844) );
  MUX2_X1 U15790 ( .A(n13845), .B(n13844), .S(n13843), .Z(n13847) );
  OAI211_X1 U15791 ( .C1(n7210), .C2(n14566), .A(n13847), .B(n13846), .ZN(
        P1_U3262) );
  NAND2_X1 U15792 ( .A1(n14060), .A2(n13855), .ZN(n13854) );
  XOR2_X1 U15793 ( .A(n13854), .B(n14055), .Z(n13848) );
  NAND2_X1 U15794 ( .A1(n13848), .A2(n14126), .ZN(n14056) );
  NOR2_X1 U15795 ( .A1(n14047), .A2(n13849), .ZN(n13852) );
  INV_X1 U15796 ( .A(n14061), .ZN(n13850) );
  NAND2_X1 U15797 ( .A1(n13851), .A2(n13850), .ZN(n14058) );
  NOR2_X1 U15798 ( .A1(n14041), .A2(n14058), .ZN(n13857) );
  AOI211_X1 U15799 ( .C1(n14055), .C2(n14049), .A(n13852), .B(n13857), .ZN(
        n13853) );
  OAI21_X1 U15800 ( .B1(n14056), .B2(n13948), .A(n13853), .ZN(P1_U3263) );
  OAI211_X1 U15801 ( .C1(n14060), .C2(n13855), .A(n14126), .B(n13854), .ZN(
        n14059) );
  NOR2_X1 U15802 ( .A1(n14060), .A2(n14035), .ZN(n13856) );
  AOI211_X1 U15803 ( .C1(n14041), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13857), 
        .B(n13856), .ZN(n13858) );
  OAI21_X1 U15804 ( .B1(n13948), .B2(n14059), .A(n13858), .ZN(P1_U3264) );
  NAND2_X1 U15805 ( .A1(n13862), .A2(n14008), .ZN(n13864) );
  NAND2_X1 U15806 ( .A1(n13887), .A2(n14006), .ZN(n13863) );
  AOI21_X1 U15807 ( .B1(n14070), .B2(n13867), .A(n14509), .ZN(n13868) );
  NAND2_X1 U15808 ( .A1(n14070), .A2(n14049), .ZN(n13870) );
  NAND2_X1 U15809 ( .A1(n14041), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13869) );
  OAI211_X1 U15810 ( .C1(n14011), .C2(n13871), .A(n13870), .B(n13869), .ZN(
        n13876) );
  OAI21_X1 U15811 ( .B1(n13874), .B2(n13873), .A(n13872), .ZN(n14073) );
  NOR2_X1 U15812 ( .A1(n14073), .A2(n14019), .ZN(n13875) );
  OAI21_X1 U15813 ( .B1(n14041), .B2(n14072), .A(n13877), .ZN(P1_U3265) );
  XNOR2_X1 U15814 ( .A(n13878), .B(n13883), .ZN(n14083) );
  INV_X1 U15815 ( .A(n13880), .ZN(n13881) );
  AOI21_X1 U15816 ( .B1(n14079), .B2(n13907), .A(n13881), .ZN(n14080) );
  INV_X1 U15817 ( .A(n14080), .ZN(n13889) );
  OR3_X1 U15818 ( .A1(n13900), .A2(n13883), .A3(n13882), .ZN(n13884) );
  NAND2_X1 U15819 ( .A1(n13885), .A2(n13884), .ZN(n13888) );
  AOI222_X1 U15820 ( .A1(n13888), .A2(n14028), .B1(n13887), .B2(n14008), .C1(
        n13886), .C2(n14006), .ZN(n14082) );
  OAI21_X1 U15821 ( .B1(n14013), .B2(n13889), .A(n14082), .ZN(n13894) );
  AOI22_X1 U15822 ( .A1(n14041), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13890), 
        .B2(n14051), .ZN(n13891) );
  OAI21_X1 U15823 ( .B1(n13892), .B2(n14035), .A(n13891), .ZN(n13893) );
  AOI21_X1 U15824 ( .B1(n13894), .B2(n14047), .A(n13893), .ZN(n13895) );
  OAI21_X1 U15825 ( .B1(n14019), .B2(n14083), .A(n13895), .ZN(P1_U3267) );
  AOI21_X1 U15826 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n13899) );
  INV_X1 U15827 ( .A(n13899), .ZN(n14088) );
  INV_X1 U15828 ( .A(n13900), .ZN(n13904) );
  OAI21_X1 U15829 ( .B1(n6505), .B2(n13902), .A(n13901), .ZN(n13903) );
  NAND2_X1 U15830 ( .A1(n13904), .A2(n13903), .ZN(n13906) );
  AOI21_X1 U15831 ( .B1(n13906), .B2(n14028), .A(n13905), .ZN(n14087) );
  INV_X1 U15832 ( .A(n14087), .ZN(n13911) );
  AOI21_X1 U15833 ( .B1(n14084), .B2(n13925), .A(n13879), .ZN(n14085) );
  INV_X1 U15834 ( .A(n14085), .ZN(n13909) );
  OAI22_X1 U15835 ( .A1(n13909), .A2(n14013), .B1(n13908), .B2(n14011), .ZN(
        n13910) );
  OAI21_X1 U15836 ( .B1(n13911), .B2(n13910), .A(n14047), .ZN(n13913) );
  AOI22_X1 U15837 ( .A1(n14084), .A2(n14049), .B1(n14041), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U15838 ( .C1(n14088), .C2(n14019), .A(n13913), .B(n13912), .ZN(
        P1_U3268) );
  NAND2_X1 U15839 ( .A1(n13915), .A2(n13914), .ZN(n13916) );
  NAND2_X1 U15840 ( .A1(n13917), .A2(n13916), .ZN(n14092) );
  NAND2_X1 U15841 ( .A1(n13919), .A2(n13918), .ZN(n13920) );
  NAND2_X1 U15842 ( .A1(n13920), .A2(n14028), .ZN(n13922) );
  OAI21_X1 U15843 ( .B1(n6505), .B2(n13922), .A(n13921), .ZN(n13923) );
  AOI21_X1 U15844 ( .B1(n14092), .B2(n13924), .A(n13923), .ZN(n14094) );
  AOI21_X1 U15845 ( .B1(n13928), .B2(n13942), .A(n14509), .ZN(n13926) );
  NAND2_X1 U15846 ( .A1(n13926), .A2(n13925), .ZN(n14090) );
  AOI22_X1 U15847 ( .A1(n14041), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13927), 
        .B2(n14051), .ZN(n13930) );
  NAND2_X1 U15848 ( .A1(n13928), .A2(n14049), .ZN(n13929) );
  OAI211_X1 U15849 ( .C1(n14090), .C2(n13948), .A(n13930), .B(n13929), .ZN(
        n13931) );
  AOI21_X1 U15850 ( .B1(n14092), .B2(n13932), .A(n13931), .ZN(n13933) );
  OAI21_X1 U15851 ( .B1(n14094), .B2(n14041), .A(n13933), .ZN(P1_U3269) );
  INV_X1 U15852 ( .A(n13934), .ZN(n13935) );
  AOI21_X1 U15853 ( .B1(n13938), .B2(n13936), .A(n13935), .ZN(n14097) );
  OAI21_X1 U15854 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(n13940) );
  NAND2_X1 U15855 ( .A1(n13940), .A2(n14028), .ZN(n14101) );
  INV_X1 U15856 ( .A(n14098), .ZN(n13941) );
  AOI21_X1 U15857 ( .B1(n14101), .B2(n13941), .A(n14041), .ZN(n13950) );
  OAI211_X1 U15858 ( .C1(n13943), .C2(n6608), .A(n14126), .B(n13942), .ZN(
        n14100) );
  OAI22_X1 U15859 ( .A1(n14047), .A2(n13945), .B1(n13944), .B2(n14011), .ZN(
        n13946) );
  AOI21_X1 U15860 ( .B1(n6904), .B2(n14049), .A(n13946), .ZN(n13947) );
  OAI21_X1 U15861 ( .B1(n14100), .B2(n13948), .A(n13947), .ZN(n13949) );
  AOI211_X1 U15862 ( .C1(n14097), .C2(n13951), .A(n13950), .B(n13949), .ZN(
        n13952) );
  INV_X1 U15863 ( .A(n13952), .ZN(P1_U3270) );
  OAI21_X1 U15864 ( .B1(n13954), .B2(n13959), .A(n13953), .ZN(n13955) );
  INV_X1 U15865 ( .A(n13955), .ZN(n14108) );
  AOI21_X1 U15866 ( .B1(n14104), .B2(n13968), .A(n6608), .ZN(n14105) );
  AND2_X1 U15867 ( .A1(n13999), .A2(n14126), .ZN(n14050) );
  INV_X1 U15868 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n13956) );
  OAI22_X1 U15869 ( .A1(n13957), .A2(n14035), .B1(n13956), .B2(n14047), .ZN(
        n13958) );
  AOI21_X1 U15870 ( .B1(n14105), .B2(n14050), .A(n13958), .ZN(n13966) );
  XNOR2_X1 U15871 ( .A(n13960), .B(n13959), .ZN(n13962) );
  AOI21_X1 U15872 ( .B1(n13962), .B2(n14028), .A(n13961), .ZN(n14107) );
  OAI21_X1 U15873 ( .B1(n13963), .B2(n14011), .A(n14107), .ZN(n13964) );
  NAND2_X1 U15874 ( .A1(n13964), .A2(n14047), .ZN(n13965) );
  OAI211_X1 U15875 ( .C1(n14108), .C2(n14019), .A(n13966), .B(n13965), .ZN(
        P1_U3271) );
  XNOR2_X1 U15876 ( .A(n13967), .B(n13976), .ZN(n14113) );
  INV_X1 U15877 ( .A(n13987), .ZN(n13970) );
  INV_X1 U15878 ( .A(n13968), .ZN(n13969) );
  AOI21_X1 U15879 ( .B1(n14109), .B2(n13970), .A(n13969), .ZN(n14110) );
  NOR2_X1 U15880 ( .A1(n13971), .A2(n14035), .ZN(n13975) );
  OAI22_X1 U15881 ( .A1(n14047), .A2(n13973), .B1(n13972), .B2(n14011), .ZN(
        n13974) );
  AOI211_X1 U15882 ( .C1(n14110), .C2(n14050), .A(n13975), .B(n13974), .ZN(
        n13981) );
  XNOR2_X1 U15883 ( .A(n13977), .B(n13976), .ZN(n13979) );
  AOI21_X1 U15884 ( .B1(n13979), .B2(n14028), .A(n13978), .ZN(n14112) );
  OR2_X1 U15885 ( .A1(n14112), .A2(n14041), .ZN(n13980) );
  OAI211_X1 U15886 ( .C1(n14113), .C2(n14019), .A(n13981), .B(n13980), .ZN(
        P1_U3272) );
  OAI211_X1 U15887 ( .C1(n6595), .C2(n13993), .A(n13982), .B(n14028), .ZN(
        n13986) );
  AOI22_X1 U15888 ( .A1(n13984), .A2(n14006), .B1(n14008), .B2(n13983), .ZN(
        n13985) );
  AND2_X1 U15889 ( .A1(n13986), .A2(n13985), .ZN(n14117) );
  OAI21_X1 U15890 ( .B1(n6497), .B2(n13991), .A(n14126), .ZN(n13988) );
  NOR2_X1 U15891 ( .A1(n13988), .A2(n13987), .ZN(n14114) );
  AOI22_X1 U15892 ( .A1(n13989), .A2(n14051), .B1(n14041), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n13990) );
  OAI21_X1 U15893 ( .B1(n13991), .B2(n14035), .A(n13990), .ZN(n13998) );
  INV_X1 U15894 ( .A(n13992), .ZN(n14002) );
  OAI21_X1 U15895 ( .B1(n14002), .B2(n13994), .A(n13993), .ZN(n13996) );
  NAND2_X1 U15896 ( .A1(n13996), .A2(n13995), .ZN(n14118) );
  NOR2_X1 U15897 ( .A1(n14118), .A2(n14019), .ZN(n13997) );
  AOI211_X1 U15898 ( .C1(n14114), .C2(n13999), .A(n13998), .B(n13997), .ZN(
        n14000) );
  OAI21_X1 U15899 ( .B1(n14041), .B2(n14117), .A(n14000), .ZN(P1_U3273) );
  INV_X1 U15900 ( .A(n14001), .ZN(n14003) );
  AOI21_X1 U15901 ( .B1(n14003), .B2(n14005), .A(n14002), .ZN(n14123) );
  OAI21_X1 U15902 ( .B1(n6590), .B2(n14005), .A(n14004), .ZN(n14010) );
  AOI222_X1 U15903 ( .A1(n14010), .A2(n14028), .B1(n14009), .B2(n14008), .C1(
        n14007), .C2(n14006), .ZN(n14122) );
  INV_X1 U15904 ( .A(n14122), .ZN(n14016) );
  AOI21_X1 U15905 ( .B1(n14119), .B2(n14030), .A(n6497), .ZN(n14120) );
  INV_X1 U15906 ( .A(n14120), .ZN(n14014) );
  OAI22_X1 U15907 ( .A1(n14014), .A2(n14013), .B1(n14012), .B2(n14011), .ZN(
        n14015) );
  OAI21_X1 U15908 ( .B1(n14016), .B2(n14015), .A(n14047), .ZN(n14018) );
  AOI22_X1 U15909 ( .A1(n14119), .A2(n14049), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n14041), .ZN(n14017) );
  OAI211_X1 U15910 ( .C1(n14123), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        P1_U3274) );
  XOR2_X1 U15911 ( .A(n14020), .B(n14024), .Z(n14029) );
  OAI22_X1 U15912 ( .A1(n14022), .A2(n14045), .B1(n14463), .B2(n14021), .ZN(
        n14027) );
  XOR2_X1 U15913 ( .A(n14024), .B(n14023), .Z(n14131) );
  NOR2_X1 U15914 ( .A1(n14131), .A2(n14025), .ZN(n14026) );
  AOI211_X1 U15915 ( .C1(n14029), .C2(n14028), .A(n14027), .B(n14026), .ZN(
        n14129) );
  AOI21_X1 U15916 ( .B1(n14125), .B2(n14031), .A(n6889), .ZN(n14127) );
  INV_X1 U15917 ( .A(n14032), .ZN(n14033) );
  AOI22_X1 U15918 ( .A1(n14041), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14033), 
        .B2(n14051), .ZN(n14034) );
  OAI21_X1 U15919 ( .B1(n14036), .B2(n14035), .A(n14034), .ZN(n14039) );
  NOR2_X1 U15920 ( .A1(n14131), .A2(n14037), .ZN(n14038) );
  AOI211_X1 U15921 ( .C1(n14127), .C2(n14050), .A(n14039), .B(n14038), .ZN(
        n14040) );
  OAI21_X1 U15922 ( .B1(n14129), .B2(n14041), .A(n14040), .ZN(P1_U3275) );
  INV_X1 U15923 ( .A(n14042), .ZN(n14044) );
  NOR2_X1 U15924 ( .A1(n14043), .A2(n14168), .ZN(n14587) );
  NOR3_X1 U15925 ( .A1(n14582), .A2(n14044), .A3(n14587), .ZN(n14048) );
  NOR2_X1 U15926 ( .A1(n14046), .A2(n14045), .ZN(n14586) );
  OAI21_X1 U15927 ( .B1(n14048), .B2(n14586), .A(n14047), .ZN(n14054) );
  OAI21_X1 U15928 ( .B1(n14050), .B2(n14049), .A(n7408), .ZN(n14053) );
  AOI22_X1 U15929 ( .A1(n14041), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14051), .ZN(n14052) );
  NAND3_X1 U15930 ( .A1(n14054), .A2(n14053), .A3(n14052), .ZN(P1_U3293) );
  INV_X1 U15931 ( .A(n14055), .ZN(n14057) );
  OAI211_X1 U15932 ( .C1(n14057), .C2(n14634), .A(n14056), .B(n14058), .ZN(
        n14133) );
  MUX2_X1 U15933 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14133), .S(n14654), .Z(
        P1_U3559) );
  OAI211_X1 U15934 ( .C1(n14060), .C2(n14634), .A(n14059), .B(n14058), .ZN(
        n14134) );
  MUX2_X1 U15935 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14134), .S(n14654), .Z(
        P1_U3558) );
  NOR2_X1 U15936 ( .A1(n14062), .A2(n14061), .ZN(n14064) );
  MUX2_X1 U15937 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14135), .S(n14654), .Z(
        P1_U3557) );
  AOI21_X1 U15938 ( .B1(n14070), .B2(n14124), .A(n14069), .ZN(n14071) );
  OAI211_X1 U15939 ( .C1(n14073), .C2(n14583), .A(n14072), .B(n14071), .ZN(
        n14136) );
  MUX2_X1 U15940 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14136), .S(n14654), .Z(
        P1_U3556) );
  AOI21_X1 U15941 ( .B1(n14075), .B2(n14124), .A(n14074), .ZN(n14076) );
  OAI211_X1 U15942 ( .C1(n14078), .C2(n14130), .A(n14077), .B(n14076), .ZN(
        n14137) );
  MUX2_X1 U15943 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14137), .S(n14654), .Z(
        P1_U3555) );
  AOI22_X1 U15944 ( .A1(n14080), .A2(n14126), .B1(n14079), .B2(n14124), .ZN(
        n14081) );
  OAI211_X1 U15945 ( .C1(n14583), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        n14138) );
  MUX2_X1 U15946 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14138), .S(n14654), .Z(
        P1_U3554) );
  AOI22_X1 U15947 ( .A1(n14085), .A2(n14126), .B1(n14084), .B2(n14124), .ZN(
        n14086) );
  OAI211_X1 U15948 ( .C1(n14088), .C2(n14583), .A(n14087), .B(n14086), .ZN(
        n14139) );
  MUX2_X1 U15949 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14139), .S(n14654), .Z(
        P1_U3553) );
  INV_X1 U15950 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14095) );
  NAND2_X1 U15951 ( .A1(n14090), .A2(n14089), .ZN(n14091) );
  AOI21_X1 U15952 ( .B1(n14092), .B2(n14618), .A(n14091), .ZN(n14093) );
  AND2_X1 U15953 ( .A1(n14094), .A2(n14093), .ZN(n14140) );
  MUX2_X1 U15954 ( .A(n14095), .B(n14140), .S(n14654), .Z(n14096) );
  INV_X1 U15955 ( .A(n14096), .ZN(P1_U3552) );
  NAND2_X1 U15956 ( .A1(n14097), .A2(n14638), .ZN(n14103) );
  NOR2_X1 U15957 ( .A1(n14099), .A2(n14098), .ZN(n14102) );
  NAND4_X1 U15958 ( .A1(n14103), .A2(n14102), .A3(n14101), .A4(n14100), .ZN(
        n14142) );
  MUX2_X1 U15959 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14142), .S(n14654), .Z(
        P1_U3551) );
  AOI22_X1 U15960 ( .A1(n14105), .A2(n14126), .B1(n14104), .B2(n14124), .ZN(
        n14106) );
  OAI211_X1 U15961 ( .C1(n14108), .C2(n14583), .A(n14107), .B(n14106), .ZN(
        n14143) );
  MUX2_X1 U15962 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14143), .S(n14654), .Z(
        P1_U3550) );
  AOI22_X1 U15963 ( .A1(n14110), .A2(n14126), .B1(n14109), .B2(n14124), .ZN(
        n14111) );
  OAI211_X1 U15964 ( .C1(n14113), .C2(n14583), .A(n14112), .B(n14111), .ZN(
        n14144) );
  MUX2_X1 U15965 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14144), .S(n14654), .Z(
        P1_U3549) );
  AOI21_X1 U15966 ( .B1(n14115), .B2(n14124), .A(n14114), .ZN(n14116) );
  OAI211_X1 U15967 ( .C1(n14583), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n14145) );
  MUX2_X1 U15968 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14145), .S(n14654), .Z(
        P1_U3548) );
  AOI22_X1 U15969 ( .A1(n14120), .A2(n14126), .B1(n14119), .B2(n14124), .ZN(
        n14121) );
  OAI211_X1 U15970 ( .C1(n14123), .C2(n14583), .A(n14122), .B(n14121), .ZN(
        n14146) );
  MUX2_X1 U15971 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14146), .S(n14654), .Z(
        P1_U3547) );
  AOI22_X1 U15972 ( .A1(n14127), .A2(n14126), .B1(n14125), .B2(n14124), .ZN(
        n14128) );
  OAI211_X1 U15973 ( .C1(n14131), .C2(n14130), .A(n14129), .B(n14128), .ZN(
        n14147) );
  MUX2_X1 U15974 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14147), .S(n14654), .Z(
        P1_U3546) );
  MUX2_X1 U15975 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14132), .S(n14654), .Z(
        P1_U3537) );
  MUX2_X1 U15976 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14133), .S(n14641), .Z(
        P1_U3527) );
  MUX2_X1 U15977 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14134), .S(n14641), .Z(
        P1_U3526) );
  MUX2_X1 U15978 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14135), .S(n14641), .Z(
        P1_U3525) );
  MUX2_X1 U15979 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14136), .S(n14641), .Z(
        P1_U3524) );
  MUX2_X1 U15980 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14137), .S(n14641), .Z(
        P1_U3523) );
  MUX2_X1 U15981 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14138), .S(n14641), .Z(
        P1_U3522) );
  MUX2_X1 U15982 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14139), .S(n14641), .Z(
        P1_U3521) );
  INV_X1 U15983 ( .A(n14140), .ZN(n14141) );
  MUX2_X1 U15984 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14141), .S(n14641), .Z(
        P1_U3520) );
  MUX2_X1 U15985 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14142), .S(n14641), .Z(
        P1_U3519) );
  MUX2_X1 U15986 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14143), .S(n14641), .Z(
        P1_U3518) );
  MUX2_X1 U15987 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14144), .S(n14641), .Z(
        P1_U3517) );
  MUX2_X1 U15988 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14145), .S(n14641), .Z(
        P1_U3516) );
  MUX2_X1 U15989 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14146), .S(n14641), .Z(
        P1_U3515) );
  MUX2_X1 U15990 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14147), .S(n14641), .Z(
        P1_U3513) );
  NOR4_X1 U15991 ( .A1(n6738), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n7588), .ZN(n14148) );
  AOI21_X1 U15992 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14149), .A(n14148), 
        .ZN(n14150) );
  OAI21_X1 U15993 ( .B1(n14151), .B2(n14166), .A(n14150), .ZN(P1_U3324) );
  OAI222_X1 U15994 ( .A1(P1_U3086), .A2(n14154), .B1(n14166), .B2(n14153), 
        .C1(n14152), .C2(n14163), .ZN(P1_U3326) );
  OAI222_X1 U15995 ( .A1(P1_U3086), .A2(n14157), .B1(n14166), .B2(n14156), 
        .C1(n14155), .C2(n14163), .ZN(P1_U3328) );
  OAI222_X1 U15996 ( .A1(n14160), .A2(P1_U3086), .B1(n14166), .B2(n14159), 
        .C1(n14158), .C2(n14163), .ZN(P1_U3329) );
  OAI222_X1 U15997 ( .A1(P1_U3086), .A2(n8031), .B1(n14166), .B2(n14162), .C1(
        n14161), .C2(n14163), .ZN(P1_U3330) );
  OAI222_X1 U15998 ( .A1(P1_U3086), .A2(n14167), .B1(n14166), .B2(n14165), 
        .C1(n14164), .C2(n14163), .ZN(P1_U3331) );
  MUX2_X1 U15999 ( .A(n14169), .B(n14168), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16000 ( .A(n14170), .ZN(n14171) );
  MUX2_X1 U16001 ( .A(n14171), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16002 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14255) );
  INV_X1 U16003 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14259) );
  XNOR2_X1 U16004 ( .A(n14259), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n14257) );
  INV_X1 U16005 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14205) );
  INV_X1 U16006 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14203) );
  INV_X1 U16007 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14201) );
  INV_X1 U16008 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14198) );
  XNOR2_X1 U16009 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n14248) );
  INV_X1 U16010 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14196) );
  XNOR2_X1 U16011 ( .A(n14196), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14209) );
  INV_X1 U16012 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14191) );
  XNOR2_X1 U16013 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n14211) );
  INV_X1 U16014 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14189) );
  XNOR2_X1 U16015 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n14241) );
  INV_X1 U16016 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14184) );
  XNOR2_X1 U16017 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14235) );
  NAND2_X1 U16018 ( .A1(n14218), .A2(n14217), .ZN(n14172) );
  OAI21_X1 U16019 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n14173), .A(n14172), .ZN(
        n14216) );
  NAND2_X1 U16020 ( .A1(n14215), .A2(n14216), .ZN(n14174) );
  NAND2_X1 U16021 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14175), .ZN(n14176) );
  NAND2_X1 U16022 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14177), .ZN(n14179) );
  NAND2_X1 U16023 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14180), .ZN(n14182) );
  XNOR2_X1 U16024 ( .A(n14180), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14229) );
  NAND2_X1 U16025 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14185), .ZN(n14187) );
  XOR2_X1 U16026 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14185), .Z(n14238) );
  INV_X1 U16027 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14239) );
  NAND2_X1 U16028 ( .A1(n14238), .A2(n14239), .ZN(n14186) );
  NAND2_X1 U16029 ( .A1(n14187), .A2(n14186), .ZN(n14242) );
  NAND2_X1 U16030 ( .A1(n14241), .A2(n14242), .ZN(n14188) );
  NAND2_X1 U16031 ( .A1(n14211), .A2(n14212), .ZN(n14190) );
  NAND2_X1 U16032 ( .A1(n14191), .A2(n14192), .ZN(n14194) );
  XNOR2_X1 U16033 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14192), .ZN(n14210) );
  NAND2_X1 U16034 ( .A1(n14210), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n14193) );
  NAND2_X1 U16035 ( .A1(n14248), .A2(n14247), .ZN(n14197) );
  INV_X1 U16036 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U16037 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14199), .ZN(n14200) );
  XOR2_X1 U16038 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P3_ADDR_REG_14__SCAN_IN), 
        .Z(n14253) );
  NOR2_X1 U16039 ( .A1(n14254), .A2(n14253), .ZN(n14202) );
  AND2_X1 U16040 ( .A1(n14205), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n14204) );
  OAI22_X1 U16041 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14205), .B1(n14206), 
        .B2(n14204), .ZN(n14256) );
  XOR2_X1 U16042 ( .A(n14257), .B(n14256), .Z(n14542) );
  XNOR2_X1 U16043 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n14207) );
  XOR2_X1 U16044 ( .A(n14207), .B(n14206), .Z(n14539) );
  INV_X1 U16045 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14535) );
  INV_X1 U16046 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14530) );
  XOR2_X1 U16047 ( .A(n14209), .B(n14208), .Z(n14522) );
  XNOR2_X1 U16048 ( .A(n14210), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14287) );
  XNOR2_X1 U16049 ( .A(n14212), .B(n14211), .ZN(n14283) );
  XNOR2_X1 U16050 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14213), .ZN(n14214) );
  NAND2_X1 U16051 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14214), .ZN(n14228) );
  XOR2_X1 U16052 ( .A(n14214), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15290) );
  INV_X1 U16053 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14273) );
  XNOR2_X1 U16054 ( .A(n14216), .B(n14215), .ZN(n14271) );
  XNOR2_X1 U16055 ( .A(n14218), .B(n14217), .ZN(n14219) );
  NAND2_X1 U16056 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14219), .ZN(n14221) );
  AOI21_X1 U16057 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14876), .A(n14218), .ZN(
        n15293) );
  INV_X1 U16058 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15292) );
  NOR2_X1 U16059 ( .A1(n15293), .A2(n15292), .ZN(n15301) );
  XOR2_X1 U16060 ( .A(n14219), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15300) );
  NAND2_X1 U16061 ( .A1(n15301), .A2(n15300), .ZN(n14220) );
  NAND2_X1 U16062 ( .A1(n14221), .A2(n14220), .ZN(n14272) );
  NAND2_X1 U16063 ( .A1(n14271), .A2(n14272), .ZN(n14222) );
  NOR2_X1 U16064 ( .A1(n14271), .A2(n14272), .ZN(n14270) );
  AOI21_X1 U16065 ( .B1(n14273), .B2(n14222), .A(n14270), .ZN(n15297) );
  XNOR2_X1 U16066 ( .A(n14224), .B(n14223), .ZN(n15298) );
  NOR2_X1 U16067 ( .A1(n15297), .A2(n15298), .ZN(n14226) );
  INV_X1 U16068 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U16069 ( .A1(n15297), .A2(n15298), .ZN(n15296) );
  OAI21_X1 U16070 ( .B1(n14226), .B2(n14225), .A(n15296), .ZN(n15289) );
  NAND2_X1 U16071 ( .A1(n15290), .A2(n15289), .ZN(n14227) );
  NAND2_X1 U16072 ( .A1(n14228), .A2(n14227), .ZN(n14231) );
  XNOR2_X1 U16073 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14229), .ZN(n14230) );
  NOR2_X1 U16074 ( .A1(n14231), .A2(n14230), .ZN(n14233) );
  XNOR2_X1 U16075 ( .A(n14231), .B(n14230), .ZN(n15291) );
  NOR2_X1 U16076 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15291), .ZN(n14232) );
  NAND2_X1 U16077 ( .A1(n14234), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14237) );
  XNOR2_X1 U16078 ( .A(n14236), .B(n14235), .ZN(n14275) );
  XNOR2_X1 U16079 ( .A(n14239), .B(n14238), .ZN(n15295) );
  XNOR2_X1 U16080 ( .A(n14242), .B(n14241), .ZN(n14279) );
  NAND2_X1 U16081 ( .A1(n14283), .A2(n14282), .ZN(n14281) );
  OAI21_X1 U16082 ( .B1(n14244), .B2(n14243), .A(n14281), .ZN(n14286) );
  NOR2_X1 U16083 ( .A1(n14287), .A2(n14286), .ZN(n14246) );
  INV_X1 U16084 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U16085 ( .A1(n14287), .A2(n14286), .ZN(n14285) );
  XOR2_X1 U16086 ( .A(n14248), .B(n14247), .Z(n14250) );
  XNOR2_X1 U16087 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n14252) );
  XNOR2_X1 U16088 ( .A(n14252), .B(n14251), .ZN(n14529) );
  XNOR2_X1 U16089 ( .A(n14254), .B(n14253), .ZN(n14533) );
  NAND2_X1 U16090 ( .A1(n14539), .A2(n14538), .ZN(n14537) );
  NOR2_X1 U16091 ( .A1(n14257), .A2(n14256), .ZN(n14258) );
  AOI21_X1 U16092 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14259), .A(n14258), 
        .ZN(n14261) );
  XNOR2_X1 U16093 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14261), .ZN(n14262) );
  XNOR2_X1 U16094 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14262), .ZN(n14296) );
  XNOR2_X1 U16095 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n14265) );
  INV_X1 U16096 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U16097 ( .A1(n14261), .A2(n14260), .ZN(n14264) );
  NAND2_X1 U16098 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14262), .ZN(n14263) );
  NAND2_X1 U16099 ( .A1(n14264), .A2(n14263), .ZN(n15089) );
  XOR2_X1 U16100 ( .A(n14265), .B(n15089), .Z(n14266) );
  NOR2_X1 U16101 ( .A1(n14267), .A2(n14266), .ZN(n15086) );
  AOI21_X1 U16102 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14268) );
  OAI21_X1 U16103 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14268), 
        .ZN(U28) );
  AOI21_X1 U16104 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14269) );
  OAI21_X1 U16105 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14269), 
        .ZN(U29) );
  AOI21_X1 U16106 ( .B1(n14272), .B2(n14271), .A(n14270), .ZN(n14274) );
  XNOR2_X1 U16107 ( .A(n14274), .B(n14273), .ZN(SUB_1596_U61) );
  XOR2_X1 U16108 ( .A(n14276), .B(n14275), .Z(SUB_1596_U57) );
  OAI21_X1 U16109 ( .B1(n14279), .B2(n14278), .A(n14277), .ZN(n14280) );
  XNOR2_X1 U16110 ( .A(n14280), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  OAI21_X1 U16111 ( .B1(n14283), .B2(n14282), .A(n14281), .ZN(n14284) );
  XNOR2_X1 U16112 ( .A(n14284), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  OAI21_X1 U16113 ( .B1(n14287), .B2(n14286), .A(n14285), .ZN(n14288) );
  XNOR2_X1 U16114 ( .A(n14288), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI21_X1 U16115 ( .B1(n6896), .B2(n14634), .A(n14289), .ZN(n14291) );
  AOI211_X1 U16116 ( .C1(n14618), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14294) );
  INV_X1 U16117 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U16118 ( .A1(n14641), .A2(n14294), .B1(n14293), .B2(n14639), .ZN(
        P1_U3495) );
  AOI22_X1 U16119 ( .A1(n14654), .A2(n14294), .B1(n10325), .B2(n14651), .ZN(
        P1_U3540) );
  AOI21_X1 U16120 ( .B1(n14297), .B2(n14296), .A(n14295), .ZN(n14298) );
  XOR2_X1 U16121 ( .A(n14298), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  INV_X1 U16122 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U16123 ( .A1(n14944), .A2(n14299), .B1(n15021), .B2(
        P3_ADDR_REG_15__SCAN_IN), .ZN(n14313) );
  AOI21_X1 U16124 ( .B1(n12816), .B2(n14301), .A(n14300), .ZN(n14302) );
  INV_X1 U16125 ( .A(n14302), .ZN(n14311) );
  OAI21_X1 U16126 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14304), .A(n14303), 
        .ZN(n14310) );
  INV_X1 U16127 ( .A(n14305), .ZN(n14306) );
  OAI21_X1 U16128 ( .B1(n14308), .B2(n14307), .A(n14306), .ZN(n14309) );
  AOI222_X1 U16129 ( .A1(n14311), .A2(n14355), .B1(n15014), .B2(n14310), .C1(
        n14309), .C2(n15022), .ZN(n14312) );
  OAI211_X1 U16130 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n14314), .A(n14313), .B(
        n14312), .ZN(P3_U3197) );
  AOI22_X1 U16131 ( .A1(n14944), .A2(n14315), .B1(n15021), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U16132 ( .A1(n14316), .A2(n6623), .ZN(n14317) );
  XNOR2_X1 U16133 ( .A(n14318), .B(n14317), .ZN(n14322) );
  XNOR2_X1 U16134 ( .A(n14320), .B(n14319), .ZN(n14321) );
  AOI22_X1 U16135 ( .A1(n14322), .A2(n15022), .B1(n15014), .B2(n14321), .ZN(
        n14329) );
  NAND2_X1 U16136 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14328)
         );
  INV_X1 U16137 ( .A(n14323), .ZN(n14326) );
  OAI221_X1 U16138 ( .B1(n14326), .B2(n14325), .C1(n14326), .C2(n14324), .A(
        n14355), .ZN(n14327) );
  NAND4_X1 U16139 ( .A1(n14330), .A2(n14329), .A3(n14328), .A4(n14327), .ZN(
        P3_U3198) );
  AOI22_X1 U16140 ( .A1(n14944), .A2(n14331), .B1(n15021), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14345) );
  OAI21_X1 U16141 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14333), .A(n14332), 
        .ZN(n14338) );
  AOI211_X1 U16142 ( .C1(n14336), .C2(n14335), .A(n14334), .B(n15003), .ZN(
        n14337) );
  AOI21_X1 U16143 ( .B1(n15014), .B2(n14338), .A(n14337), .ZN(n14344) );
  NAND2_X1 U16144 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14343)
         );
  OAI221_X1 U16145 ( .B1(n14341), .B2(n14340), .C1(n14341), .C2(n14339), .A(
        n14355), .ZN(n14342) );
  NAND4_X1 U16146 ( .A1(n14345), .A2(n14344), .A3(n14343), .A4(n14342), .ZN(
        P3_U3199) );
  AOI22_X1 U16147 ( .A1(n14944), .A2(n14346), .B1(n15021), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14362) );
  XNOR2_X1 U16148 ( .A(n14348), .B(n14347), .ZN(n14354) );
  AOI21_X1 U16149 ( .B1(n14351), .B2(n14350), .A(n14349), .ZN(n14352) );
  NOR2_X1 U16150 ( .A1(n14352), .A2(n15003), .ZN(n14353) );
  AOI21_X1 U16151 ( .B1(n14354), .B2(n15014), .A(n14353), .ZN(n14361) );
  NAND2_X1 U16152 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14360)
         );
  OAI221_X1 U16153 ( .B1(n14358), .B2(n14357), .C1(n14358), .C2(n14356), .A(
        n14355), .ZN(n14359) );
  NAND4_X1 U16154 ( .A1(n14362), .A2(n14361), .A3(n14360), .A4(n14359), .ZN(
        P3_U3200) );
  OAI21_X1 U16155 ( .B1(n14364), .B2(n15068), .A(n14363), .ZN(n14365) );
  AOI21_X1 U16156 ( .B1(n14366), .B2(n15054), .A(n14365), .ZN(n14389) );
  AOI22_X1 U16157 ( .A1(n15085), .A2(n14389), .B1(n14367), .B2(n9553), .ZN(
        P3_U3474) );
  OAI21_X1 U16158 ( .B1(n14369), .B2(n15068), .A(n14368), .ZN(n14370) );
  AOI21_X1 U16159 ( .B1(n15054), .B2(n14371), .A(n14370), .ZN(n14390) );
  AOI22_X1 U16160 ( .A1(n15085), .A2(n14390), .B1(n12577), .B2(n9553), .ZN(
        P3_U3473) );
  NOR2_X1 U16161 ( .A1(n14373), .A2(n14372), .ZN(n14375) );
  AOI211_X1 U16162 ( .C1(n14383), .C2(n14376), .A(n14375), .B(n14374), .ZN(
        n14392) );
  INV_X1 U16163 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U16164 ( .A1(n15085), .A2(n14392), .B1(n14377), .B2(n9553), .ZN(
        P3_U3472) );
  OAI21_X1 U16165 ( .B1(n14379), .B2(n15068), .A(n14378), .ZN(n14380) );
  AOI21_X1 U16166 ( .B1(n14381), .B2(n15054), .A(n14380), .ZN(n14394) );
  AOI22_X1 U16167 ( .A1(n15085), .A2(n14394), .B1(n14382), .B2(n9553), .ZN(
        P3_U3471) );
  AOI22_X1 U16168 ( .A1(n14385), .A2(n15054), .B1(n14384), .B2(n14383), .ZN(
        n14386) );
  AND2_X1 U16169 ( .A1(n14387), .A2(n14386), .ZN(n14395) );
  INV_X1 U16170 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16171 ( .A1(n15085), .A2(n14395), .B1(n14388), .B2(n9553), .ZN(
        P3_U3470) );
  AOI22_X1 U16172 ( .A1(n15076), .A2(n14389), .B1(n9319), .B2(n15074), .ZN(
        P3_U3435) );
  AOI22_X1 U16173 ( .A1(n15076), .A2(n14390), .B1(n9301), .B2(n15074), .ZN(
        P3_U3432) );
  INV_X1 U16174 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U16175 ( .A1(n15076), .A2(n14392), .B1(n14391), .B2(n15074), .ZN(
        P3_U3429) );
  INV_X1 U16176 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U16177 ( .A1(n15076), .A2(n14394), .B1(n14393), .B2(n15074), .ZN(
        P3_U3426) );
  AOI22_X1 U16178 ( .A1(n15076), .A2(n14395), .B1(n9254), .B2(n15074), .ZN(
        P3_U3423) );
  XOR2_X1 U16179 ( .A(n14396), .B(n14406), .Z(n14400) );
  INV_X1 U16180 ( .A(n14397), .ZN(n14398) );
  AOI21_X1 U16181 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n14430) );
  AOI222_X1 U16182 ( .A1(n14412), .A2(n14403), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n13411), .C1(n14402), .C2(n14401), .ZN(n14419) );
  OR2_X1 U16183 ( .A1(n14405), .A2(n7132), .ZN(n14409) );
  NAND2_X1 U16184 ( .A1(n14407), .A2(n14406), .ZN(n14408) );
  AOI21_X1 U16185 ( .B1(n14412), .B2(n14411), .A(n13295), .ZN(n14414) );
  NAND2_X1 U16186 ( .A1(n14414), .A2(n14413), .ZN(n14428) );
  NOR2_X1 U16187 ( .A1(n14428), .A2(n14415), .ZN(n14416) );
  AOI21_X1 U16188 ( .B1(n14433), .B2(n14417), .A(n14416), .ZN(n14418) );
  OAI211_X1 U16189 ( .C1(n14420), .C2(n14430), .A(n14419), .B(n14418), .ZN(
        P2_U3251) );
  INV_X1 U16190 ( .A(n14421), .ZN(n14422) );
  OAI211_X1 U16191 ( .C1(n14424), .C2(n14828), .A(n14423), .B(n14422), .ZN(
        n14426) );
  AOI211_X1 U16192 ( .C1(n14816), .C2(n14427), .A(n14426), .B(n14425), .ZN(
        n14445) );
  AOI22_X1 U16193 ( .A1(n14842), .A2(n14445), .B1(n8379), .B2(n8665), .ZN(
        P2_U3514) );
  OAI21_X1 U16194 ( .B1(n14429), .B2(n14828), .A(n14428), .ZN(n14432) );
  INV_X1 U16195 ( .A(n14430), .ZN(n14431) );
  AOI211_X1 U16196 ( .C1(n14433), .C2(n14816), .A(n14432), .B(n14431), .ZN(
        n14447) );
  AOI22_X1 U16197 ( .A1(n14842), .A2(n14447), .B1(n13169), .B2(n8665), .ZN(
        P2_U3513) );
  OAI21_X1 U16198 ( .B1(n14435), .B2(n14828), .A(n14434), .ZN(n14437) );
  AOI211_X1 U16199 ( .C1(n14438), .C2(n14816), .A(n14437), .B(n14436), .ZN(
        n14449) );
  AOI22_X1 U16200 ( .A1(n14842), .A2(n14449), .B1(n13168), .B2(n8665), .ZN(
        P2_U3512) );
  OAI21_X1 U16201 ( .B1(n7308), .B2(n14828), .A(n14440), .ZN(n14441) );
  AOI21_X1 U16202 ( .B1(n14442), .B2(n14835), .A(n14441), .ZN(n14443) );
  AOI22_X1 U16203 ( .A1(n14842), .A2(n14451), .B1(n8334), .B2(n8665), .ZN(
        P2_U3511) );
  AOI22_X1 U16204 ( .A1(n14836), .A2(n14445), .B1(n8378), .B2(n7143), .ZN(
        P2_U3475) );
  INV_X1 U16205 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U16206 ( .A1(n14836), .A2(n14447), .B1(n14446), .B2(n7143), .ZN(
        P2_U3472) );
  INV_X1 U16207 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U16208 ( .A1(n14836), .A2(n14449), .B1(n14448), .B2(n7143), .ZN(
        P2_U3469) );
  INV_X1 U16209 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U16210 ( .A1(n14836), .A2(n14451), .B1(n14450), .B2(n7143), .ZN(
        P2_U3466) );
  OAI22_X1 U16211 ( .A1(n14462), .A2(n14478), .B1(n14477), .B2(n14452), .ZN(
        n14458) );
  NAND2_X1 U16212 ( .A1(n14454), .A2(n14453), .ZN(n14455) );
  AOI21_X1 U16213 ( .B1(n14456), .B2(n14455), .A(n14467), .ZN(n14457) );
  AOI211_X1 U16214 ( .C1(n14490), .C2(n14507), .A(n14458), .B(n14457), .ZN(
        n14460) );
  OAI211_X1 U16215 ( .C1(n14494), .C2(n14461), .A(n14460), .B(n14459), .ZN(
        P1_U3215) );
  OAI22_X1 U16216 ( .A1(n14463), .A2(n14478), .B1(n14477), .B2(n14462), .ZN(
        n14471) );
  INV_X1 U16217 ( .A(n13688), .ZN(n14466) );
  OAI21_X1 U16218 ( .B1(n14466), .B2(n14465), .A(n14464), .ZN(n14469) );
  AOI21_X1 U16219 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14470) );
  AOI211_X1 U16220 ( .C1(n14490), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        n14474) );
  OAI211_X1 U16221 ( .C1(n14494), .C2(n14475), .A(n14474), .B(n14473), .ZN(
        P1_U3226) );
  OAI22_X1 U16222 ( .A1(n14479), .A2(n14478), .B1(n14477), .B2(n14476), .ZN(
        n14488) );
  AOI21_X1 U16223 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n14484) );
  OAI21_X1 U16224 ( .B1(n14485), .B2(n14484), .A(n14483), .ZN(n14486) );
  INV_X1 U16225 ( .A(n14486), .ZN(n14487) );
  AOI211_X1 U16226 ( .C1(n14490), .C2(n14489), .A(n14488), .B(n14487), .ZN(
        n14492) );
  OAI211_X1 U16227 ( .C1(n14494), .C2(n14493), .A(n14492), .B(n14491), .ZN(
        P1_U3236) );
  NAND3_X1 U16228 ( .A1(n11653), .A2(n14495), .A3(n14638), .ZN(n14497) );
  OAI211_X1 U16229 ( .C1(n6890), .C2(n14634), .A(n14497), .B(n14496), .ZN(
        n14499) );
  NOR2_X1 U16230 ( .A1(n14499), .A2(n14498), .ZN(n14515) );
  AOI22_X1 U16231 ( .A1(n14654), .A2(n14515), .B1(n14500), .B2(n14651), .ZN(
        P1_U3545) );
  OAI211_X1 U16232 ( .C1(n14503), .C2(n14634), .A(n14502), .B(n14501), .ZN(
        n14504) );
  AOI211_X1 U16233 ( .C1(n14506), .C2(n14638), .A(n14505), .B(n14504), .ZN(
        n14517) );
  AOI22_X1 U16234 ( .A1(n14654), .A2(n14517), .B1(n11533), .B2(n14651), .ZN(
        P1_U3544) );
  INV_X1 U16235 ( .A(n14507), .ZN(n14508) );
  OAI22_X1 U16236 ( .A1(n14510), .A2(n14509), .B1(n14508), .B2(n14634), .ZN(
        n14511) );
  AOI211_X1 U16237 ( .C1(n14513), .C2(n14638), .A(n14512), .B(n14511), .ZN(
        n14519) );
  AOI22_X1 U16238 ( .A1(n14654), .A2(n14519), .B1(n7733), .B2(n14651), .ZN(
        P1_U3542) );
  INV_X1 U16239 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14514) );
  AOI22_X1 U16240 ( .A1(n14641), .A2(n14515), .B1(n14514), .B2(n14639), .ZN(
        P1_U3510) );
  INV_X1 U16241 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14516) );
  AOI22_X1 U16242 ( .A1(n14641), .A2(n14517), .B1(n14516), .B2(n14639), .ZN(
        P1_U3507) );
  INV_X1 U16243 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U16244 ( .A1(n14641), .A2(n14519), .B1(n14518), .B2(n14639), .ZN(
        P1_U3501) );
  AOI21_X1 U16245 ( .B1(n14522), .B2(n14521), .A(n14520), .ZN(n14523) );
  XOR2_X1 U16246 ( .A(n14523), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  NOR2_X1 U16247 ( .A1(n14525), .A2(n14524), .ZN(n14526) );
  XOR2_X1 U16248 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14526), .Z(SUB_1596_U68)
         );
  AOI21_X1 U16249 ( .B1(n14529), .B2(n14528), .A(n14527), .ZN(n14531) );
  XNOR2_X1 U16250 ( .A(n14531), .B(n14530), .ZN(SUB_1596_U67) );
  AOI21_X1 U16251 ( .B1(n14534), .B2(n14533), .A(n14532), .ZN(n14536) );
  XNOR2_X1 U16252 ( .A(n14536), .B(n14535), .ZN(SUB_1596_U66) );
  OAI21_X1 U16253 ( .B1(n14539), .B2(n14538), .A(n14537), .ZN(n14540) );
  XNOR2_X1 U16254 ( .A(n14540), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  OAI21_X1 U16255 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14544) );
  XNOR2_X1 U16256 ( .A(n14544), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  OAI21_X1 U16257 ( .B1(n14546), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14545), .ZN(
        n14548) );
  XNOR2_X1 U16258 ( .A(n14548), .B(n14547), .ZN(n14551) );
  AOI22_X1 U16259 ( .A1(n14570), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14549) );
  OAI21_X1 U16260 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(P1_U3243) );
  INV_X1 U16261 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14567) );
  MUX2_X1 U16262 ( .A(n10325), .B(P1_REG1_REG_12__SCAN_IN), .S(n14562), .Z(
        n14552) );
  NAND3_X1 U16263 ( .A1(n14554), .A2(n14553), .A3(n14552), .ZN(n14555) );
  NAND2_X1 U16264 ( .A1(n14556), .A2(n14555), .ZN(n14563) );
  OAI21_X1 U16265 ( .B1(n14559), .B2(n14558), .A(n14557), .ZN(n14561) );
  AOI222_X1 U16266 ( .A1(n14563), .A2(n14575), .B1(n14562), .B2(n14573), .C1(
        n14561), .C2(n14560), .ZN(n14565) );
  OAI211_X1 U16267 ( .C1(n14567), .C2(n14566), .A(n14565), .B(n14564), .ZN(
        P1_U3255) );
  AOI21_X1 U16268 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14569), .A(n14568), 
        .ZN(n14580) );
  AOI22_X1 U16269 ( .A1(n14570), .A2(P1_ADDR_REG_15__SCAN_IN), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(P1_U3086), .ZN(n14578) );
  OAI21_X1 U16270 ( .B1(n14572), .B2(n7758), .A(n14571), .ZN(n14576) );
  AOI22_X1 U16271 ( .A1(n14576), .A2(n14575), .B1(n14574), .B2(n14573), .ZN(
        n14577) );
  OAI211_X1 U16272 ( .C1(n14580), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        P1_U3258) );
  AND2_X1 U16273 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14581), .ZN(P1_U3294) );
  AND2_X1 U16274 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14581), .ZN(P1_U3295) );
  AND2_X1 U16275 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14581), .ZN(P1_U3296) );
  AND2_X1 U16276 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14581), .ZN(P1_U3297) );
  AND2_X1 U16277 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14581), .ZN(P1_U3298) );
  AND2_X1 U16278 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14581), .ZN(P1_U3299) );
  AND2_X1 U16279 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14581), .ZN(P1_U3300) );
  AND2_X1 U16280 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14581), .ZN(P1_U3301) );
  AND2_X1 U16281 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14581), .ZN(P1_U3302) );
  AND2_X1 U16282 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14581), .ZN(P1_U3303) );
  AND2_X1 U16283 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14581), .ZN(P1_U3304) );
  AND2_X1 U16284 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14581), .ZN(P1_U3305) );
  AND2_X1 U16285 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14581), .ZN(P1_U3306) );
  AND2_X1 U16286 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14581), .ZN(P1_U3307) );
  AND2_X1 U16287 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14581), .ZN(P1_U3308) );
  AND2_X1 U16288 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14581), .ZN(P1_U3309) );
  AND2_X1 U16289 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14581), .ZN(P1_U3310) );
  AND2_X1 U16290 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14581), .ZN(P1_U3311) );
  AND2_X1 U16291 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14581), .ZN(P1_U3312) );
  AND2_X1 U16292 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14581), .ZN(P1_U3313) );
  AND2_X1 U16293 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14581), .ZN(P1_U3314) );
  AND2_X1 U16294 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14581), .ZN(P1_U3315) );
  AND2_X1 U16295 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14581), .ZN(P1_U3316) );
  AND2_X1 U16296 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14581), .ZN(P1_U3317) );
  AND2_X1 U16297 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14581), .ZN(P1_U3318) );
  AND2_X1 U16298 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14581), .ZN(P1_U3319) );
  AND2_X1 U16299 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14581), .ZN(P1_U3320) );
  AND2_X1 U16300 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14581), .ZN(P1_U3321) );
  AND2_X1 U16301 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14581), .ZN(P1_U3322) );
  AND2_X1 U16302 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14581), .ZN(P1_U3323) );
  AOI21_X1 U16303 ( .B1(n14584), .B2(n14583), .A(n14582), .ZN(n14585) );
  AOI211_X1 U16304 ( .C1(n7408), .C2(n14587), .A(n14586), .B(n14585), .ZN(
        n14643) );
  INV_X1 U16305 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U16306 ( .A1(n14641), .A2(n14643), .B1(n14588), .B2(n14639), .ZN(
        P1_U3459) );
  OAI21_X1 U16307 ( .B1(n14590), .B2(n14634), .A(n14589), .ZN(n14592) );
  AOI211_X1 U16308 ( .C1(n14618), .C2(n14593), .A(n14592), .B(n14591), .ZN(
        n14645) );
  INV_X1 U16309 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14594) );
  AOI22_X1 U16310 ( .A1(n14641), .A2(n14645), .B1(n14594), .B2(n14639), .ZN(
        P1_U3462) );
  INV_X1 U16311 ( .A(n14595), .ZN(n14603) );
  INV_X1 U16312 ( .A(n14596), .ZN(n14600) );
  INV_X1 U16313 ( .A(n14597), .ZN(n14598) );
  NAND4_X1 U16314 ( .A1(n14601), .A2(n14600), .A3(n14599), .A4(n14598), .ZN(
        n14602) );
  AOI21_X1 U16315 ( .B1(n14603), .B2(n14638), .A(n14602), .ZN(n14646) );
  AOI22_X1 U16316 ( .A1(n14641), .A2(n14646), .B1(n7539), .B2(n14639), .ZN(
        P1_U3471) );
  INV_X1 U16317 ( .A(n14604), .ZN(n14606) );
  AOI211_X1 U16318 ( .C1(n14607), .C2(n14618), .A(n14606), .B(n14605), .ZN(
        n14608) );
  AND2_X1 U16319 ( .A1(n14609), .A2(n14608), .ZN(n14647) );
  INV_X1 U16320 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14610) );
  AOI22_X1 U16321 ( .A1(n14641), .A2(n14647), .B1(n14610), .B2(n14639), .ZN(
        P1_U3474) );
  INV_X1 U16322 ( .A(n14611), .ZN(n14613) );
  NAND3_X1 U16323 ( .A1(n14614), .A2(n14613), .A3(n14612), .ZN(n14616) );
  AOI211_X1 U16324 ( .C1(n14617), .C2(n14638), .A(n14616), .B(n14615), .ZN(
        n14648) );
  AOI22_X1 U16325 ( .A1(n14641), .A2(n14648), .B1(n6739), .B2(n14639), .ZN(
        P1_U3477) );
  NAND2_X1 U16326 ( .A1(n14619), .A2(n14618), .ZN(n14621) );
  OAI211_X1 U16327 ( .C1(n14622), .C2(n14634), .A(n14621), .B(n14620), .ZN(
        n14623) );
  NOR2_X1 U16328 ( .A1(n14624), .A2(n14623), .ZN(n14649) );
  INV_X1 U16329 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14625) );
  AOI22_X1 U16330 ( .A1(n14641), .A2(n14649), .B1(n14625), .B2(n14639), .ZN(
        P1_U3480) );
  OR2_X1 U16331 ( .A1(n14627), .A2(n14626), .ZN(n14629) );
  AOI211_X1 U16332 ( .C1(n14638), .C2(n14630), .A(n14629), .B(n14628), .ZN(
        n14650) );
  INV_X1 U16333 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14631) );
  AOI22_X1 U16334 ( .A1(n14641), .A2(n14650), .B1(n14631), .B2(n14639), .ZN(
        P1_U3483) );
  OAI211_X1 U16335 ( .C1(n14635), .C2(n14634), .A(n14633), .B(n14632), .ZN(
        n14636) );
  AOI21_X1 U16336 ( .B1(n14638), .B2(n14637), .A(n14636), .ZN(n14653) );
  INV_X1 U16337 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16338 ( .A1(n14641), .A2(n14653), .B1(n14640), .B2(n14639), .ZN(
        P1_U3489) );
  INV_X1 U16339 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14642) );
  AOI22_X1 U16340 ( .A1(n14654), .A2(n14643), .B1(n14642), .B2(n14651), .ZN(
        P1_U3528) );
  AOI22_X1 U16341 ( .A1(n14654), .A2(n14645), .B1(n14644), .B2(n14651), .ZN(
        P1_U3529) );
  AOI22_X1 U16342 ( .A1(n14654), .A2(n14646), .B1(n7541), .B2(n14651), .ZN(
        P1_U3532) );
  AOI22_X1 U16343 ( .A1(n14654), .A2(n14647), .B1(n9805), .B2(n14651), .ZN(
        P1_U3533) );
  AOI22_X1 U16344 ( .A1(n14654), .A2(n14648), .B1(n9808), .B2(n14651), .ZN(
        P1_U3534) );
  AOI22_X1 U16345 ( .A1(n14654), .A2(n14649), .B1(n9810), .B2(n14651), .ZN(
        P1_U3535) );
  AOI22_X1 U16346 ( .A1(n14654), .A2(n14650), .B1(n7624), .B2(n14651), .ZN(
        P1_U3536) );
  AOI22_X1 U16347 ( .A1(n14654), .A2(n14653), .B1(n14652), .B2(n14651), .ZN(
        P1_U3538) );
  NOR2_X1 U16348 ( .A1(n14724), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16349 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14727), .B1(n14743), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16350 ( .A1(n14724), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14657) );
  OAI22_X1 U16351 ( .A1(n14747), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14668), .ZN(n14655) );
  OAI21_X1 U16352 ( .B1(n14741), .B2(n14655), .A(n14663), .ZN(n14656) );
  OAI211_X1 U16353 ( .C1(n14663), .C2(n14658), .A(n14657), .B(n14656), .ZN(
        P2_U3214) );
  INV_X1 U16354 ( .A(n14659), .ZN(n14661) );
  OAI21_X1 U16355 ( .B1(n14661), .B2(n14660), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14662) );
  OAI21_X1 U16356 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14662), .ZN(n14676) );
  INV_X1 U16357 ( .A(n14663), .ZN(n14664) );
  NOR2_X1 U16358 ( .A1(n14664), .A2(n8158), .ZN(n14667) );
  OAI211_X1 U16359 ( .C1(n14667), .C2(n14666), .A(n14727), .B(n14665), .ZN(
        n14675) );
  AOI211_X1 U16360 ( .C1(n14671), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14672) );
  INV_X1 U16361 ( .A(n14672), .ZN(n14674) );
  NAND2_X1 U16362 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14724), .ZN(n14673) );
  NAND4_X1 U16363 ( .A1(n14676), .A2(n14675), .A3(n14674), .A4(n14673), .ZN(
        P2_U3215) );
  INV_X1 U16364 ( .A(n14677), .ZN(n14678) );
  OAI21_X1 U16365 ( .B1(n14694), .B2(n14679), .A(n14678), .ZN(n14680) );
  AOI21_X1 U16366 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14724), .A(n14680), .ZN(
        n14690) );
  AOI211_X1 U16367 ( .C1(n14683), .C2(n14682), .A(n14681), .B(n14747), .ZN(
        n14684) );
  INV_X1 U16368 ( .A(n14684), .ZN(n14689) );
  OAI211_X1 U16369 ( .C1(n14687), .C2(n14686), .A(n14743), .B(n14685), .ZN(
        n14688) );
  NAND3_X1 U16370 ( .A1(n14690), .A2(n14689), .A3(n14688), .ZN(P2_U3217) );
  INV_X1 U16371 ( .A(n14691), .ZN(n14692) );
  OAI21_X1 U16372 ( .B1(n14694), .B2(n14693), .A(n14692), .ZN(n14695) );
  AOI21_X1 U16373 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14724), .A(n14695), 
        .ZN(n14704) );
  OAI211_X1 U16374 ( .C1(n14698), .C2(n14697), .A(n14696), .B(n14727), .ZN(
        n14703) );
  OAI211_X1 U16375 ( .C1(n14701), .C2(n14700), .A(n14699), .B(n14743), .ZN(
        n14702) );
  NAND3_X1 U16376 ( .A1(n14704), .A2(n14703), .A3(n14702), .ZN(P2_U3227) );
  AOI22_X1 U16377 ( .A1(n14724), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14714) );
  OAI211_X1 U16378 ( .C1(n14707), .C2(n14706), .A(n14705), .B(n14743), .ZN(
        n14713) );
  OAI211_X1 U16379 ( .C1(n14709), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14708), 
        .B(n14727), .ZN(n14712) );
  NAND2_X1 U16380 ( .A1(n14741), .A2(n14710), .ZN(n14711) );
  NAND4_X1 U16381 ( .A1(n14714), .A2(n14713), .A3(n14712), .A4(n14711), .ZN(
        P2_U3228) );
  AOI22_X1 U16382 ( .A1(n14724), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14723) );
  NAND2_X1 U16383 ( .A1(n14741), .A2(n14715), .ZN(n14722) );
  OAI211_X1 U16384 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14717), .A(n14727), 
        .B(n14716), .ZN(n14721) );
  OAI211_X1 U16385 ( .C1(n14719), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14743), 
        .B(n14718), .ZN(n14720) );
  NAND4_X1 U16386 ( .A1(n14723), .A2(n14722), .A3(n14721), .A4(n14720), .ZN(
        P2_U3229) );
  AOI22_X1 U16387 ( .A1(n14724), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n14737) );
  NAND2_X1 U16388 ( .A1(n14741), .A2(n14725), .ZN(n14736) );
  INV_X1 U16389 ( .A(n14726), .ZN(n14728) );
  OAI211_X1 U16390 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14735) );
  XNOR2_X1 U16391 ( .A(n14732), .B(n14731), .ZN(n14733) );
  NAND2_X1 U16392 ( .A1(n14733), .A2(n14743), .ZN(n14734) );
  NAND4_X1 U16393 ( .A1(n14737), .A2(n14736), .A3(n14735), .A4(n14734), .ZN(
        P2_U3230) );
  INV_X1 U16394 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14753) );
  AOI21_X1 U16395 ( .B1(n14739), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14738), 
        .ZN(n14748) );
  NAND2_X1 U16396 ( .A1(n14741), .A2(n14740), .ZN(n14746) );
  OAI211_X1 U16397 ( .C1(n14744), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14743), 
        .B(n14742), .ZN(n14745) );
  OAI211_X1 U16398 ( .C1(n14748), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        n14749) );
  INV_X1 U16399 ( .A(n14749), .ZN(n14751) );
  OAI211_X1 U16400 ( .C1(n14753), .C2(n14752), .A(n14751), .B(n14750), .ZN(
        P2_U3232) );
  INV_X1 U16401 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n14755) );
  NOR2_X1 U16402 ( .A1(n14786), .A2(n14755), .ZN(P2_U3266) );
  INV_X1 U16403 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n14756) );
  NOR2_X1 U16404 ( .A1(n14786), .A2(n14756), .ZN(P2_U3267) );
  INV_X1 U16405 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14757) );
  NOR2_X1 U16406 ( .A1(n14786), .A2(n14757), .ZN(P2_U3268) );
  INV_X1 U16407 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14758) );
  NOR2_X1 U16408 ( .A1(n14786), .A2(n14758), .ZN(P2_U3269) );
  INV_X1 U16409 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14759) );
  NOR2_X1 U16410 ( .A1(n14769), .A2(n14759), .ZN(P2_U3270) );
  INV_X1 U16411 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14760) );
  NOR2_X1 U16412 ( .A1(n14769), .A2(n14760), .ZN(P2_U3271) );
  INV_X1 U16413 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14761) );
  NOR2_X1 U16414 ( .A1(n14769), .A2(n14761), .ZN(P2_U3272) );
  INV_X1 U16415 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14762) );
  NOR2_X1 U16416 ( .A1(n14769), .A2(n14762), .ZN(P2_U3273) );
  INV_X1 U16417 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14763) );
  NOR2_X1 U16418 ( .A1(n14769), .A2(n14763), .ZN(P2_U3274) );
  INV_X1 U16419 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14764) );
  NOR2_X1 U16420 ( .A1(n14769), .A2(n14764), .ZN(P2_U3275) );
  INV_X1 U16421 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14765) );
  NOR2_X1 U16422 ( .A1(n14769), .A2(n14765), .ZN(P2_U3276) );
  INV_X1 U16423 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14766) );
  NOR2_X1 U16424 ( .A1(n14769), .A2(n14766), .ZN(P2_U3277) );
  INV_X1 U16425 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14767) );
  NOR2_X1 U16426 ( .A1(n14769), .A2(n14767), .ZN(P2_U3278) );
  INV_X1 U16427 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14768) );
  NOR2_X1 U16428 ( .A1(n14769), .A2(n14768), .ZN(P2_U3279) );
  INV_X1 U16429 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14770) );
  NOR2_X1 U16430 ( .A1(n14786), .A2(n14770), .ZN(P2_U3280) );
  INV_X1 U16431 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14771) );
  NOR2_X1 U16432 ( .A1(n14786), .A2(n14771), .ZN(P2_U3281) );
  INV_X1 U16433 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14772) );
  NOR2_X1 U16434 ( .A1(n14786), .A2(n14772), .ZN(P2_U3282) );
  INV_X1 U16435 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14773) );
  NOR2_X1 U16436 ( .A1(n14786), .A2(n14773), .ZN(P2_U3283) );
  INV_X1 U16437 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14774) );
  NOR2_X1 U16438 ( .A1(n14786), .A2(n14774), .ZN(P2_U3284) );
  INV_X1 U16439 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14775) );
  NOR2_X1 U16440 ( .A1(n14786), .A2(n14775), .ZN(P2_U3285) );
  INV_X1 U16441 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14776) );
  NOR2_X1 U16442 ( .A1(n14786), .A2(n14776), .ZN(P2_U3286) );
  INV_X1 U16443 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14777) );
  NOR2_X1 U16444 ( .A1(n14786), .A2(n14777), .ZN(P2_U3287) );
  INV_X1 U16445 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14778) );
  NOR2_X1 U16446 ( .A1(n14786), .A2(n14778), .ZN(P2_U3288) );
  INV_X1 U16447 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14779) );
  NOR2_X1 U16448 ( .A1(n14786), .A2(n14779), .ZN(P2_U3289) );
  INV_X1 U16449 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14780) );
  NOR2_X1 U16450 ( .A1(n14786), .A2(n14780), .ZN(P2_U3290) );
  INV_X1 U16451 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14781) );
  NOR2_X1 U16452 ( .A1(n14786), .A2(n14781), .ZN(P2_U3291) );
  INV_X1 U16453 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14782) );
  NOR2_X1 U16454 ( .A1(n14786), .A2(n14782), .ZN(P2_U3292) );
  INV_X1 U16455 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14783) );
  NOR2_X1 U16456 ( .A1(n14786), .A2(n14783), .ZN(P2_U3293) );
  INV_X1 U16457 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14784) );
  NOR2_X1 U16458 ( .A1(n14786), .A2(n14784), .ZN(P2_U3294) );
  INV_X1 U16459 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14785) );
  NOR2_X1 U16460 ( .A1(n14786), .A2(n14785), .ZN(P2_U3295) );
  MUX2_X1 U16461 ( .A(P2_D_REG_0__SCAN_IN), .B(n14787), .S(n14786), .Z(
        P2_U3416) );
  AOI22_X1 U16462 ( .A1(n14791), .A2(n14790), .B1(n14789), .B2(n14788), .ZN(
        P2_U3417) );
  INV_X1 U16463 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14792) );
  AOI22_X1 U16464 ( .A1(n14836), .A2(n14793), .B1(n14792), .B2(n7143), .ZN(
        P2_U3430) );
  INV_X1 U16465 ( .A(n14798), .ZN(n14800) );
  AOI211_X1 U16466 ( .C1(n14819), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14797) );
  OAI21_X1 U16467 ( .B1(n14805), .B2(n14798), .A(n14797), .ZN(n14799) );
  AOI21_X1 U16468 ( .B1(n14810), .B2(n14800), .A(n14799), .ZN(n14837) );
  INV_X1 U16469 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16470 ( .A1(n14836), .A2(n14837), .B1(n14801), .B2(n7143), .ZN(
        P2_U3445) );
  AOI21_X1 U16471 ( .B1(n14819), .B2(n14803), .A(n14802), .ZN(n14804) );
  OAI21_X1 U16472 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14807) );
  AOI211_X1 U16473 ( .C1(n14810), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        n14838) );
  INV_X1 U16474 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U16475 ( .A1(n14836), .A2(n14838), .B1(n14811), .B2(n7143), .ZN(
        P2_U3448) );
  OAI21_X1 U16476 ( .B1(n14813), .B2(n14828), .A(n14812), .ZN(n14815) );
  AOI211_X1 U16477 ( .C1(n14817), .C2(n14816), .A(n14815), .B(n14814), .ZN(
        n14839) );
  INV_X1 U16478 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14818) );
  AOI22_X1 U16479 ( .A1(n14836), .A2(n14839), .B1(n14818), .B2(n7143), .ZN(
        P2_U3451) );
  AND2_X1 U16480 ( .A1(n14820), .A2(n14819), .ZN(n14821) );
  OR2_X1 U16481 ( .A1(n14822), .A2(n14821), .ZN(n14823) );
  AOI21_X1 U16482 ( .B1(n14824), .B2(n14835), .A(n14823), .ZN(n14825) );
  AND2_X1 U16483 ( .A1(n14826), .A2(n14825), .ZN(n14840) );
  AOI22_X1 U16484 ( .A1(n14836), .A2(n14840), .B1(n8270), .B2(n7143), .ZN(
        P2_U3454) );
  OAI21_X1 U16485 ( .B1(n14829), .B2(n14828), .A(n14827), .ZN(n14833) );
  OAI21_X1 U16486 ( .B1(n14831), .B2(n10023), .A(n14830), .ZN(n14832) );
  AOI211_X1 U16487 ( .C1(n14835), .C2(n14834), .A(n14833), .B(n14832), .ZN(
        n14841) );
  AOI22_X1 U16488 ( .A1(n14836), .A2(n14841), .B1(n8311), .B2(n7143), .ZN(
        P2_U3463) );
  AOI22_X1 U16489 ( .A1(n14842), .A2(n14837), .B1(n8229), .B2(n8665), .ZN(
        P2_U3504) );
  AOI22_X1 U16490 ( .A1(n14842), .A2(n14838), .B1(n8242), .B2(n8665), .ZN(
        P2_U3505) );
  AOI22_X1 U16491 ( .A1(n14842), .A2(n14839), .B1(n9884), .B2(n8665), .ZN(
        P2_U3506) );
  AOI22_X1 U16492 ( .A1(n14842), .A2(n14840), .B1(n8274), .B2(n8665), .ZN(
        P2_U3507) );
  AOI22_X1 U16493 ( .A1(n14842), .A2(n14841), .B1(n8316), .B2(n8665), .ZN(
        P2_U3510) );
  NOR2_X1 U16494 ( .A1(P3_U3897), .A2(n15021), .ZN(P3_U3150) );
  OAI211_X1 U16495 ( .C1(n14845), .C2(n14844), .A(n14843), .B(n14857), .ZN(
        n14850) );
  AOI21_X1 U16496 ( .B1(n14848), .B2(n14847), .A(n14846), .ZN(n14849) );
  OAI211_X1 U16497 ( .C1(n14852), .C2(n14851), .A(n14850), .B(n14849), .ZN(
        n14853) );
  INV_X1 U16498 ( .A(n14853), .ZN(n14854) );
  OAI21_X1 U16499 ( .B1(n14867), .B2(n14855), .A(n14854), .ZN(P3_U3153) );
  INV_X1 U16500 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n14885) );
  OAI22_X1 U16501 ( .A1(n15052), .A2(n14856), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14885), .ZN(n14863) );
  OAI211_X1 U16502 ( .C1(n14860), .C2(n14859), .A(n14858), .B(n14857), .ZN(
        n14861) );
  INV_X1 U16503 ( .A(n14861), .ZN(n14862) );
  AOI211_X1 U16504 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14866) );
  OAI21_X1 U16505 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n14867), .A(n14866), .ZN(
        P3_U3158) );
  OAI21_X1 U16506 ( .B1(n14869), .B2(P3_IR_REG_0__SCAN_IN), .A(n14868), .ZN(
        n14871) );
  NAND3_X1 U16507 ( .A1(n15028), .A2(n14913), .A3(n15003), .ZN(n14870) );
  NAND2_X1 U16508 ( .A1(n14871), .A2(n14870), .ZN(n14875) );
  OAI22_X1 U16509 ( .A1(n15018), .A2(n6746), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14872), .ZN(n14873) );
  INV_X1 U16510 ( .A(n14873), .ZN(n14874) );
  OAI211_X1 U16511 ( .C1(n14876), .C2(n14953), .A(n14875), .B(n14874), .ZN(
        P3_U3182) );
  NOR2_X1 U16512 ( .A1(n14877), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U16513 ( .A1(n14879), .A2(n14878), .ZN(n14895) );
  AND3_X1 U16514 ( .A1(n14882), .A2(n14881), .A3(n14880), .ZN(n14883) );
  OAI21_X1 U16515 ( .B1(n14884), .B2(n14883), .A(n15022), .ZN(n14888) );
  NOR2_X1 U16516 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14885), .ZN(n14886) );
  AOI21_X1 U16517 ( .B1(n15021), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n14886), .ZN(
        n14887) );
  OAI211_X1 U16518 ( .C1(n15018), .C2(n14889), .A(n14888), .B(n14887), .ZN(
        n14890) );
  INV_X1 U16519 ( .A(n14890), .ZN(n14894) );
  XNOR2_X1 U16520 ( .A(n14891), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n14892) );
  NAND2_X1 U16521 ( .A1(n15014), .A2(n14892), .ZN(n14893) );
  OAI211_X1 U16522 ( .C1(n14895), .C2(n15028), .A(n14894), .B(n14893), .ZN(
        P3_U3185) );
  AOI21_X1 U16523 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(n14916) );
  AOI21_X1 U16524 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14906) );
  INV_X1 U16525 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15151) );
  NOR2_X1 U16526 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15151), .ZN(n14904) );
  NOR2_X1 U16527 ( .A1(n15018), .A2(n14902), .ZN(n14903) );
  AOI211_X1 U16528 ( .C1(n15021), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n14904), .B(
        n14903), .ZN(n14905) );
  OAI21_X1 U16529 ( .B1(n14906), .B2(n15003), .A(n14905), .ZN(n14907) );
  INV_X1 U16530 ( .A(n14907), .ZN(n14915) );
  INV_X1 U16531 ( .A(n14908), .ZN(n14909) );
  AOI21_X1 U16532 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14912) );
  OR2_X1 U16533 ( .A1(n14913), .A2(n14912), .ZN(n14914) );
  OAI211_X1 U16534 ( .C1(n14916), .C2(n15028), .A(n14915), .B(n14914), .ZN(
        P3_U3186) );
  AOI21_X1 U16535 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14933) );
  NOR2_X1 U16536 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15191), .ZN(n14927) );
  NOR2_X1 U16537 ( .A1(n14921), .A2(n14920), .ZN(n14922) );
  XNOR2_X1 U16538 ( .A(n14923), .B(n14922), .ZN(n14925) );
  OAI22_X1 U16539 ( .A1(n14925), .A2(n15003), .B1(n14924), .B2(n15018), .ZN(
        n14926) );
  AOI211_X1 U16540 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15021), .A(n14927), .B(
        n14926), .ZN(n14932) );
  OAI21_X1 U16541 ( .B1(n14929), .B2(P3_REG1_REG_5__SCAN_IN), .A(n14928), .ZN(
        n14930) );
  NAND2_X1 U16542 ( .A1(n15014), .A2(n14930), .ZN(n14931) );
  OAI211_X1 U16543 ( .C1(n14933), .C2(n15028), .A(n14932), .B(n14931), .ZN(
        P3_U3187) );
  NAND2_X1 U16544 ( .A1(n14935), .A2(n14934), .ZN(n14936) );
  XNOR2_X1 U16545 ( .A(n14937), .B(n14936), .ZN(n14938) );
  NOR2_X1 U16546 ( .A1(n14938), .A2(n15003), .ZN(n14950) );
  AOI21_X1 U16547 ( .B1(n14941), .B2(n14940), .A(n14939), .ZN(n14948) );
  OAI21_X1 U16548 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14943), .A(n14942), .ZN(
        n14946) );
  AOI22_X1 U16549 ( .A1(n14946), .A2(n15014), .B1(n14945), .B2(n14944), .ZN(
        n14947) );
  OAI21_X1 U16550 ( .B1(n14948), .B2(n15028), .A(n14947), .ZN(n14949) );
  NOR2_X1 U16551 ( .A1(n14950), .A2(n14949), .ZN(n14952) );
  OAI211_X1 U16552 ( .C1(n14954), .C2(n14953), .A(n14952), .B(n14951), .ZN(
        P3_U3191) );
  AOI21_X1 U16553 ( .B1(n9253), .B2(n14956), .A(n14955), .ZN(n14971) );
  OAI21_X1 U16554 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n14958), .A(n14957), 
        .ZN(n14964) );
  AND2_X1 U16555 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n14960) );
  AOI21_X1 U16556 ( .B1(n15021), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n14960), 
        .ZN(n14961) );
  OAI21_X1 U16557 ( .B1(n15018), .B2(n14962), .A(n14961), .ZN(n14963) );
  AOI21_X1 U16558 ( .B1(n14964), .B2(n15014), .A(n14963), .ZN(n14970) );
  AOI21_X1 U16559 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n14968) );
  OR2_X1 U16560 ( .A1(n14968), .A2(n15003), .ZN(n14969) );
  OAI211_X1 U16561 ( .C1(n14971), .C2(n15028), .A(n14970), .B(n14969), .ZN(
        P3_U3193) );
  AOI21_X1 U16562 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14989) );
  OAI21_X1 U16563 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n14983) );
  NOR2_X1 U16564 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14978), .ZN(n14979) );
  AOI21_X1 U16565 ( .B1(n15021), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n14979), 
        .ZN(n14980) );
  OAI21_X1 U16566 ( .B1(n15018), .B2(n14981), .A(n14980), .ZN(n14982) );
  AOI21_X1 U16567 ( .B1(n14983), .B2(n15014), .A(n14982), .ZN(n14988) );
  OAI211_X1 U16568 ( .C1(n14986), .C2(n14985), .A(n14984), .B(n15022), .ZN(
        n14987) );
  OAI211_X1 U16569 ( .C1(n14989), .C2(n15028), .A(n14988), .B(n14987), .ZN(
        P3_U3194) );
  AOI21_X1 U16570 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n15007) );
  OAI21_X1 U16571 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n14994), .A(n14993), 
        .ZN(n14999) );
  INV_X1 U16572 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15250) );
  NOR2_X1 U16573 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15250), .ZN(n14995) );
  AOI21_X1 U16574 ( .B1(n15021), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n14995), 
        .ZN(n14996) );
  OAI21_X1 U16575 ( .B1(n15018), .B2(n14997), .A(n14996), .ZN(n14998) );
  AOI21_X1 U16576 ( .B1(n14999), .B2(n15014), .A(n14998), .ZN(n15006) );
  AOI21_X1 U16577 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15004) );
  OR2_X1 U16578 ( .A1(n15004), .A2(n15003), .ZN(n15005) );
  OAI211_X1 U16579 ( .C1(n15007), .C2(n15028), .A(n15006), .B(n15005), .ZN(
        P3_U3195) );
  AOI21_X1 U16580 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15029) );
  OAI21_X1 U16581 ( .B1(n15013), .B2(n15012), .A(n15011), .ZN(n15015) );
  AND2_X1 U16582 ( .A1(n15015), .A2(n15014), .ZN(n15020) );
  OAI21_X1 U16583 ( .B1(n15018), .B2(n15017), .A(n15016), .ZN(n15019) );
  AOI211_X1 U16584 ( .C1(P3_ADDR_REG_14__SCAN_IN), .C2(n15021), .A(n15020), 
        .B(n15019), .ZN(n15027) );
  OAI211_X1 U16585 ( .C1(n15025), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        n15026) );
  OAI211_X1 U16586 ( .C1(n15029), .C2(n15028), .A(n15027), .B(n15026), .ZN(
        P3_U3196) );
  XNOR2_X1 U16587 ( .A(n15030), .B(n15036), .ZN(n15049) );
  NOR2_X1 U16588 ( .A1(n15031), .A2(n15068), .ZN(n15048) );
  INV_X1 U16589 ( .A(n15048), .ZN(n15035) );
  INV_X1 U16590 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15033) );
  OAI22_X1 U16591 ( .A1(n15035), .A2(n15034), .B1(n15033), .B2(n15032), .ZN(
        n15043) );
  XNOR2_X1 U16592 ( .A(n15036), .B(n9596), .ZN(n15037) );
  OAI222_X1 U16593 ( .A1(n15042), .A2(n15041), .B1(n15040), .B2(n15039), .C1(
        n15038), .C2(n15037), .ZN(n15047) );
  AOI211_X1 U16594 ( .C1(n15044), .C2(n15049), .A(n15043), .B(n15047), .ZN(
        n15046) );
  AOI22_X1 U16595 ( .A1(n12844), .A2(n10046), .B1(n15046), .B2(n15045), .ZN(
        P3_U3232) );
  AOI211_X1 U16596 ( .C1(n15054), .C2(n15049), .A(n15048), .B(n15047), .ZN(
        n15077) );
  INV_X1 U16597 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15050) );
  AOI22_X1 U16598 ( .A1(n15076), .A2(n15077), .B1(n15050), .B2(n15074), .ZN(
        P3_U3393) );
  OAI21_X1 U16599 ( .B1(n15052), .B2(n15068), .A(n15051), .ZN(n15053) );
  AOI21_X1 U16600 ( .B1(n15055), .B2(n15054), .A(n15053), .ZN(n15078) );
  INV_X1 U16601 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U16602 ( .A1(n15076), .A2(n15078), .B1(n15056), .B2(n15074), .ZN(
        P3_U3399) );
  NOR2_X1 U16603 ( .A1(n15057), .A2(n15068), .ZN(n15059) );
  AOI211_X1 U16604 ( .C1(n15060), .C2(n15072), .A(n15059), .B(n15058), .ZN(
        n15080) );
  INV_X1 U16605 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15061) );
  AOI22_X1 U16606 ( .A1(n15076), .A2(n15080), .B1(n15061), .B2(n15074), .ZN(
        P3_U3408) );
  NOR2_X1 U16607 ( .A1(n15062), .A2(n15068), .ZN(n15064) );
  AOI211_X1 U16608 ( .C1(n15065), .C2(n15072), .A(n15064), .B(n15063), .ZN(
        n15082) );
  INV_X1 U16609 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U16610 ( .A1(n15076), .A2(n15082), .B1(n15066), .B2(n15074), .ZN(
        P3_U3414) );
  INV_X1 U16611 ( .A(n15067), .ZN(n15073) );
  NOR2_X1 U16612 ( .A1(n15069), .A2(n15068), .ZN(n15071) );
  AOI211_X1 U16613 ( .C1(n15073), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        n15084) );
  INV_X1 U16614 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U16615 ( .A1(n15076), .A2(n15084), .B1(n15075), .B2(n15074), .ZN(
        P3_U3417) );
  AOI22_X1 U16616 ( .A1(n15085), .A2(n15077), .B1(n10168), .B2(n9553), .ZN(
        P3_U3460) );
  AOI22_X1 U16617 ( .A1(n15085), .A2(n15078), .B1(n10433), .B2(n9553), .ZN(
        P3_U3462) );
  AOI22_X1 U16618 ( .A1(n15085), .A2(n15080), .B1(n15079), .B2(n9553), .ZN(
        P3_U3465) );
  AOI22_X1 U16619 ( .A1(n15085), .A2(n15082), .B1(n15081), .B2(n9553), .ZN(
        P3_U3467) );
  AOI22_X1 U16620 ( .A1(n15085), .A2(n15084), .B1(n15083), .B2(n9553), .ZN(
        P3_U3468) );
  NOR2_X1 U16621 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n15086), .ZN(n15087) );
  NOR2_X1 U16622 ( .A1(n15088), .A2(n15087), .ZN(n15288) );
  AND2_X1 U16623 ( .A1(n11525), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n15090) );
  OAI22_X1 U16624 ( .A1(n15090), .A2(n15089), .B1(P3_ADDR_REG_18__SCAN_IN), 
        .B2(n11525), .ZN(n15286) );
  OAI22_X1 U16625 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        keyinput_g59), .B2(P3_REG3_REG_2__SCAN_IN), .ZN(n15091) );
  AOI221_X1 U16626 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput_g59), .A(n15091), .ZN(n15098) );
  OAI22_X1 U16627 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        keyinput_g14), .B2(SI_18_), .ZN(n15092) );
  AOI221_X1 U16628 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        SI_18_), .C2(keyinput_g14), .A(n15092), .ZN(n15097) );
  OAI22_X1 U16629 ( .A1(SI_27_), .A2(keyinput_g5), .B1(SI_20_), .B2(
        keyinput_g12), .ZN(n15093) );
  AOI221_X1 U16630 ( .B1(SI_27_), .B2(keyinput_g5), .C1(keyinput_g12), .C2(
        SI_20_), .A(n15093), .ZN(n15096) );
  OAI22_X1 U16631 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .ZN(n15094) );
  AOI221_X1 U16632 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g49), .C2(P3_REG3_REG_5__SCAN_IN), .A(n15094), .ZN(n15095) );
  NAND4_X1 U16633 ( .A1(n15098), .A2(n15097), .A3(n15096), .A4(n15095), .ZN(
        n15125) );
  OAI22_X1 U16634 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        keyinput_g23), .B2(SI_9_), .ZN(n15099) );
  AOI221_X1 U16635 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_9_), .C2(keyinput_g23), .A(n15099), .ZN(n15105) );
  OAI22_X1 U16636 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        keyinput_g11), .B2(SI_21_), .ZN(n15100) );
  AOI221_X1 U16637 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_21_), .C2(keyinput_g11), .A(n15100), .ZN(n15104) );
  OAI22_X1 U16638 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        keyinput_g43), .B2(P3_REG3_REG_8__SCAN_IN), .ZN(n15101) );
  AOI221_X1 U16639 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n15101), .ZN(n15103) );
  XNOR2_X1 U16640 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n15102)
         );
  NAND4_X1 U16641 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        n15124) );
  OAI22_X1 U16642 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(SI_10_), 
        .B2(keyinput_g22), .ZN(n15106) );
  AOI221_X1 U16643 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        keyinput_g22), .C2(SI_10_), .A(n15106), .ZN(n15113) );
  OAI22_X1 U16644 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        keyinput_g40), .B2(P3_REG3_REG_3__SCAN_IN), .ZN(n15107) );
  AOI221_X1 U16645 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n15107), .ZN(n15112) );
  OAI22_X1 U16646 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        keyinput_g44), .B2(P3_REG3_REG_1__SCAN_IN), .ZN(n15108) );
  AOI221_X1 U16647 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n15108), .ZN(n15111) );
  OAI22_X1 U16648 ( .A1(SI_17_), .A2(keyinput_g15), .B1(keyinput_g17), .B2(
        SI_15_), .ZN(n15109) );
  AOI221_X1 U16649 ( .B1(SI_17_), .B2(keyinput_g15), .C1(SI_15_), .C2(
        keyinput_g17), .A(n15109), .ZN(n15110) );
  NAND4_X1 U16650 ( .A1(n15113), .A2(n15112), .A3(n15111), .A4(n15110), .ZN(
        n15123) );
  OAI22_X1 U16651 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n15114) );
  AOI221_X1 U16652 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        keyinput_g33), .C2(P3_RD_REG_SCAN_IN), .A(n15114), .ZN(n15121) );
  OAI22_X1 U16653 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_30_), .B2(
        keyinput_g2), .ZN(n15115) );
  AOI221_X1 U16654 ( .B1(SI_0_), .B2(keyinput_g32), .C1(keyinput_g2), .C2(
        SI_30_), .A(n15115), .ZN(n15120) );
  OAI22_X1 U16655 ( .A1(SI_28_), .A2(keyinput_g4), .B1(keyinput_g60), .B2(
        P3_REG3_REG_18__SCAN_IN), .ZN(n15116) );
  AOI221_X1 U16656 ( .B1(SI_28_), .B2(keyinput_g4), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n15116), .ZN(n15119)
         );
  OAI22_X1 U16657 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        SI_31_), .B2(keyinput_g1), .ZN(n15117) );
  AOI221_X1 U16658 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        keyinput_g1), .C2(SI_31_), .A(n15117), .ZN(n15118) );
  NAND4_X1 U16659 ( .A1(n15121), .A2(n15120), .A3(n15119), .A4(n15118), .ZN(
        n15122) );
  OR4_X1 U16660 ( .A1(n15125), .A2(n15124), .A3(n15123), .A4(n15122), .ZN(
        n15281) );
  AOI22_X1 U16661 ( .A1(n15127), .A2(keyinput_g18), .B1(n12207), .B2(
        keyinput_g38), .ZN(n15126) );
  OAI221_X1 U16662 ( .B1(n15127), .B2(keyinput_g18), .C1(n12207), .C2(
        keyinput_g38), .A(n15126), .ZN(n15149) );
  INV_X1 U16663 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U16664 ( .A1(n15216), .A2(keyinput_g53), .B1(keyinput_g20), .B2(
        n15176), .ZN(n15128) );
  OAI221_X1 U16665 ( .B1(n15216), .B2(keyinput_g53), .C1(n15176), .C2(
        keyinput_g20), .A(n15128), .ZN(n15148) );
  INV_X1 U16666 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15187) );
  INV_X1 U16667 ( .A(SI_22_), .ZN(n15130) );
  AOI22_X1 U16668 ( .A1(n15187), .A2(keyinput_g39), .B1(keyinput_g10), .B2(
        n15130), .ZN(n15129) );
  OAI221_X1 U16669 ( .B1(n15187), .B2(keyinput_g39), .C1(n15130), .C2(
        keyinput_g10), .A(n15129), .ZN(n15147) );
  INV_X1 U16670 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15132) );
  AOI22_X1 U16671 ( .A1(n15132), .A2(keyinput_g0), .B1(n15219), .B2(
        keyinput_g57), .ZN(n15131) );
  OAI221_X1 U16672 ( .B1(n15132), .B2(keyinput_g0), .C1(n15219), .C2(
        keyinput_g57), .A(n15131), .ZN(n15145) );
  AOI22_X1 U16673 ( .A1(n15186), .A2(keyinput_g6), .B1(keyinput_g7), .B2(
        n15221), .ZN(n15133) );
  OAI221_X1 U16674 ( .B1(n15186), .B2(keyinput_g6), .C1(n15221), .C2(
        keyinput_g7), .A(n15133), .ZN(n15144) );
  XNOR2_X1 U16675 ( .A(SI_6_), .B(keyinput_g26), .ZN(n15137) );
  XNOR2_X1 U16676 ( .A(SI_8_), .B(keyinput_g24), .ZN(n15136) );
  XNOR2_X1 U16677 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n15135)
         );
  XNOR2_X1 U16678 ( .A(SI_1_), .B(keyinput_g31), .ZN(n15134) );
  NAND4_X1 U16679 ( .A1(n15137), .A2(n15136), .A3(n15135), .A4(n15134), .ZN(
        n15143) );
  XNOR2_X1 U16680 ( .A(SI_5_), .B(keyinput_g27), .ZN(n15141) );
  XNOR2_X1 U16681 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n15140)
         );
  XNOR2_X1 U16682 ( .A(SI_7_), .B(keyinput_g25), .ZN(n15139) );
  XNOR2_X1 U16683 ( .A(SI_3_), .B(keyinput_g29), .ZN(n15138) );
  NAND4_X1 U16684 ( .A1(n15141), .A2(n15140), .A3(n15139), .A4(n15138), .ZN(
        n15142) );
  OR4_X1 U16685 ( .A1(n15145), .A2(n15144), .A3(n15143), .A4(n15142), .ZN(
        n15146) );
  NOR4_X1 U16686 ( .A1(n15149), .A2(n15148), .A3(n15147), .A4(n15146), .ZN(
        n15171) );
  AOI22_X1 U16687 ( .A1(n15194), .A2(keyinput_g16), .B1(n11289), .B2(
        keyinput_g8), .ZN(n15150) );
  OAI221_X1 U16688 ( .B1(n15194), .B2(keyinput_g16), .C1(n11289), .C2(
        keyinput_g8), .A(n15150), .ZN(n15157) );
  XNOR2_X1 U16689 ( .A(keyinput_g63), .B(P3_REG3_REG_15__SCAN_IN), .ZN(n15155)
         );
  XNOR2_X1 U16690 ( .A(keyinput_g56), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n15154)
         );
  XNOR2_X1 U16691 ( .A(keyinput_g9), .B(SI_23_), .ZN(n15153) );
  XNOR2_X1 U16692 ( .A(keyinput_g52), .B(P3_REG3_REG_4__SCAN_IN), .ZN(n15152)
         );
  NAND4_X1 U16693 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15156) );
  NOR2_X1 U16694 ( .A1(n15157), .A2(n15156), .ZN(n15170) );
  AOI22_X1 U16695 ( .A1(n15175), .A2(keyinput_g19), .B1(n15195), .B2(
        keyinput_g37), .ZN(n15158) );
  OAI221_X1 U16696 ( .B1(n15175), .B2(keyinput_g19), .C1(n15195), .C2(
        keyinput_g37), .A(n15158), .ZN(n15162) );
  AOI22_X1 U16697 ( .A1(n15160), .A2(keyinput_g13), .B1(n15192), .B2(
        keyinput_g35), .ZN(n15159) );
  OAI221_X1 U16698 ( .B1(n15160), .B2(keyinput_g13), .C1(n15192), .C2(
        keyinput_g35), .A(n15159), .ZN(n15161) );
  NOR2_X1 U16699 ( .A1(n15162), .A2(n15161), .ZN(n15169) );
  AOI22_X1 U16700 ( .A1(n15211), .A2(keyinput_g3), .B1(n15213), .B2(
        keyinput_g21), .ZN(n15163) );
  OAI221_X1 U16701 ( .B1(n15211), .B2(keyinput_g3), .C1(n15213), .C2(
        keyinput_g21), .A(n15163), .ZN(n15167) );
  INV_X1 U16702 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16703 ( .A1(n15165), .A2(keyinput_g30), .B1(n15183), .B2(
        keyinput_g48), .ZN(n15164) );
  OAI221_X1 U16704 ( .B1(n15165), .B2(keyinput_g30), .C1(n15183), .C2(
        keyinput_g48), .A(n15164), .ZN(n15166) );
  NOR2_X1 U16705 ( .A1(n15167), .A2(n15166), .ZN(n15168) );
  NAND4_X1 U16706 ( .A1(n15171), .A2(n15170), .A3(n15169), .A4(n15168), .ZN(
        n15280) );
  INV_X1 U16707 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U16708 ( .A1(n15173), .A2(keyinput_f45), .B1(n12207), .B2(
        keyinput_f38), .ZN(n15172) );
  OAI221_X1 U16709 ( .B1(n15173), .B2(keyinput_f45), .C1(n12207), .C2(
        keyinput_f38), .A(n15172), .ZN(n15181) );
  AOI22_X1 U16710 ( .A1(n15176), .A2(keyinput_f20), .B1(n15175), .B2(
        keyinput_f19), .ZN(n15174) );
  OAI221_X1 U16711 ( .B1(n15176), .B2(keyinput_f20), .C1(n15175), .C2(
        keyinput_f19), .A(n15174), .ZN(n15180) );
  XNOR2_X1 U16712 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_f44), .ZN(n15178)
         );
  XNOR2_X1 U16713 ( .A(keyinput_f1), .B(SI_31_), .ZN(n15177) );
  NAND2_X1 U16714 ( .A1(n15178), .A2(n15177), .ZN(n15179) );
  NOR3_X1 U16715 ( .A1(n15181), .A2(n15180), .A3(n15179), .ZN(n15209) );
  AOI22_X1 U16716 ( .A1(n15184), .A2(keyinput_f4), .B1(keyinput_f48), .B2(
        n15183), .ZN(n15182) );
  OAI221_X1 U16717 ( .B1(n15184), .B2(keyinput_f4), .C1(n15183), .C2(
        keyinput_f48), .A(n15182), .ZN(n15189) );
  AOI22_X1 U16718 ( .A1(n15187), .A2(keyinput_f39), .B1(keyinput_f6), .B2(
        n15186), .ZN(n15185) );
  OAI221_X1 U16719 ( .B1(n15187), .B2(keyinput_f39), .C1(n15186), .C2(
        keyinput_f6), .A(n15185), .ZN(n15188) );
  NOR2_X1 U16720 ( .A1(n15189), .A2(n15188), .ZN(n15208) );
  AOI22_X1 U16721 ( .A1(n15192), .A2(keyinput_f35), .B1(keyinput_f49), .B2(
        n15191), .ZN(n15190) );
  OAI221_X1 U16722 ( .B1(n15192), .B2(keyinput_f35), .C1(n15191), .C2(
        keyinput_f49), .A(n15190), .ZN(n15197) );
  AOI22_X1 U16723 ( .A1(n15195), .A2(keyinput_f37), .B1(keyinput_f16), .B2(
        n15194), .ZN(n15193) );
  OAI221_X1 U16724 ( .B1(n15195), .B2(keyinput_f37), .C1(n15194), .C2(
        keyinput_f16), .A(n15193), .ZN(n15196) );
  NOR2_X1 U16725 ( .A1(n15197), .A2(n15196), .ZN(n15207) );
  AOI22_X1 U16726 ( .A1(n9452), .A2(keyinput_f47), .B1(keyinput_f59), .B2(
        n15199), .ZN(n15198) );
  OAI221_X1 U16727 ( .B1(n9452), .B2(keyinput_f47), .C1(n15199), .C2(
        keyinput_f59), .A(n15198), .ZN(n15205) );
  XNOR2_X1 U16728 ( .A(SI_19_), .B(keyinput_f13), .ZN(n15203) );
  XNOR2_X1 U16729 ( .A(SI_8_), .B(keyinput_f24), .ZN(n15202) );
  XNOR2_X1 U16730 ( .A(SI_14_), .B(keyinput_f18), .ZN(n15201) );
  XNOR2_X1 U16731 ( .A(SI_1_), .B(keyinput_f31), .ZN(n15200) );
  NAND4_X1 U16732 ( .A1(n15203), .A2(n15202), .A3(n15201), .A4(n15200), .ZN(
        n15204) );
  NOR2_X1 U16733 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  NAND4_X1 U16734 ( .A1(n15209), .A2(n15208), .A3(n15207), .A4(n15206), .ZN(
        n15232) );
  OAI22_X1 U16735 ( .A1(n9758), .A2(keyinput_f32), .B1(n15211), .B2(
        keyinput_f3), .ZN(n15210) );
  AOI221_X1 U16736 ( .B1(n9758), .B2(keyinput_f32), .C1(keyinput_f3), .C2(
        n15211), .A(n15210), .ZN(n15230) );
  AOI22_X1 U16737 ( .A1(n10934), .A2(keyinput_f9), .B1(keyinput_f21), .B2(
        n15213), .ZN(n15212) );
  OAI221_X1 U16738 ( .B1(n10934), .B2(keyinput_f9), .C1(n15213), .C2(
        keyinput_f21), .A(n15212), .ZN(n15226) );
  AOI22_X1 U16739 ( .A1(n15216), .A2(keyinput_f53), .B1(keyinput_f2), .B2(
        n15215), .ZN(n15214) );
  OAI221_X1 U16740 ( .B1(n15216), .B2(keyinput_f53), .C1(n15215), .C2(
        keyinput_f2), .A(n15214), .ZN(n15225) );
  AOI22_X1 U16741 ( .A1(n15219), .A2(keyinput_f57), .B1(keyinput_f5), .B2(
        n15218), .ZN(n15217) );
  OAI221_X1 U16742 ( .B1(n15219), .B2(keyinput_f57), .C1(n15218), .C2(
        keyinput_f5), .A(n15217), .ZN(n15224) );
  AOI22_X1 U16743 ( .A1(n15222), .A2(keyinput_f62), .B1(keyinput_f7), .B2(
        n15221), .ZN(n15220) );
  OAI221_X1 U16744 ( .B1(n15222), .B2(keyinput_f62), .C1(n15221), .C2(
        keyinput_f7), .A(n15220), .ZN(n15223) );
  NOR4_X1 U16745 ( .A1(n15226), .A2(n15225), .A3(n15224), .A4(n15223), .ZN(
        n15229) );
  XNOR2_X1 U16746 ( .A(SI_24_), .B(keyinput_f8), .ZN(n15228) );
  XNOR2_X1 U16747 ( .A(keyinput_f33), .B(P3_RD_REG_SCAN_IN), .ZN(n15227) );
  NAND4_X1 U16748 ( .A1(n15230), .A2(n15229), .A3(n15228), .A4(n15227), .ZN(
        n15231) );
  NOR2_X1 U16749 ( .A1(n15232), .A2(n15231), .ZN(n15246) );
  AOI22_X1 U16750 ( .A1(SI_18_), .A2(keyinput_f14), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n15233) );
  OAI221_X1 U16751 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n15233), .ZN(n15240)
         );
  AOI22_X1 U16752 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n15234) );
  OAI221_X1 U16753 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n15234), .ZN(n15239)
         );
  AOI22_X1 U16754 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n15235) );
  OAI221_X1 U16755 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n15235), .ZN(n15238)
         );
  AOI22_X1 U16756 ( .A1(SI_15_), .A2(keyinput_f17), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n15236) );
  OAI221_X1 U16757 ( .B1(SI_15_), .B2(keyinput_f17), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n15236), .ZN(n15237) );
  NOR4_X1 U16758 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15245) );
  OAI22_X1 U16759 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        keyinput_f26), .B2(SI_6_), .ZN(n15241) );
  AOI221_X1 U16760 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(SI_6_), .C2(keyinput_f26), .A(n15241), .ZN(n15244) );
  OAI22_X1 U16761 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n15242) );
  AOI221_X1 U16762 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        keyinput_f43), .C2(P3_REG3_REG_8__SCAN_IN), .A(n15242), .ZN(n15243) );
  AND4_X1 U16763 ( .A1(n15246), .A2(n15245), .A3(n15244), .A4(n15243), .ZN(
        n15273) );
  AOI22_X1 U16764 ( .A1(SI_2_), .A2(keyinput_f30), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n15247) );
  OAI221_X1 U16765 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_21_), .C2(
        keyinput_f11), .A(n15247), .ZN(n15257) );
  AOI22_X1 U16766 ( .A1(SI_5_), .A2(keyinput_f27), .B1(SI_7_), .B2(
        keyinput_f25), .ZN(n15248) );
  OAI221_X1 U16767 ( .B1(SI_5_), .B2(keyinput_f27), .C1(SI_7_), .C2(
        keyinput_f25), .A(n15248), .ZN(n15256) );
  AOI22_X1 U16768 ( .A1(n15251), .A2(keyinput_f41), .B1(keyinput_f56), .B2(
        n15250), .ZN(n15249) );
  OAI221_X1 U16769 ( .B1(n15251), .B2(keyinput_f41), .C1(n15250), .C2(
        keyinput_f56), .A(n15249), .ZN(n15255) );
  AOI22_X1 U16770 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(n15253), .B2(keyinput_f15), .ZN(n15252) );
  OAI221_X1 U16771 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        n15253), .C2(keyinput_f15), .A(n15252), .ZN(n15254) );
  NOR4_X1 U16772 ( .A1(n15257), .A2(n15256), .A3(n15255), .A4(n15254), .ZN(
        n15272) );
  AOI22_X1 U16773 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n15258) );
  OAI221_X1 U16774 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n15258), .ZN(n15265)
         );
  AOI22_X1 U16775 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(SI_22_), 
        .B2(keyinput_f10), .ZN(n15259) );
  OAI221_X1 U16776 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(SI_22_), 
        .C2(keyinput_f10), .A(n15259), .ZN(n15264) );
  AOI22_X1 U16777 ( .A1(SI_3_), .A2(keyinput_f29), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n15260) );
  OAI221_X1 U16778 ( .B1(SI_3_), .B2(keyinput_f29), .C1(SI_20_), .C2(
        keyinput_f12), .A(n15260), .ZN(n15263) );
  AOI22_X1 U16779 ( .A1(SI_10_), .A2(keyinput_f22), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n15261) );
  OAI221_X1 U16780 ( .B1(SI_10_), .B2(keyinput_f22), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n15261), .ZN(n15262)
         );
  NOR4_X1 U16781 ( .A1(n15265), .A2(n15264), .A3(n15263), .A4(n15262), .ZN(
        n15268) );
  OAI22_X1 U16782 ( .A1(SI_9_), .A2(keyinput_f23), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(keyinput_f54), .ZN(n15266) );
  AOI221_X1 U16783 ( .B1(SI_9_), .B2(keyinput_f23), .C1(keyinput_f54), .C2(
        P3_REG3_REG_0__SCAN_IN), .A(n15266), .ZN(n15267) );
  OAI211_X1 U16784 ( .C1(n15270), .C2(keyinput_f55), .A(n15268), .B(n15267), 
        .ZN(n15269) );
  AOI21_X1 U16785 ( .B1(n15270), .B2(keyinput_f55), .A(n15269), .ZN(n15271) );
  NAND3_X1 U16786 ( .A1(n15273), .A2(n15272), .A3(n15271), .ZN(n15276) );
  AOI21_X1 U16787 ( .B1(keyinput_f28), .B2(n15276), .A(keyinput_g28), .ZN(
        n15278) );
  INV_X1 U16788 ( .A(keyinput_f28), .ZN(n15275) );
  INV_X1 U16789 ( .A(keyinput_g28), .ZN(n15274) );
  AOI21_X1 U16790 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(n15277) );
  MUX2_X1 U16791 ( .A(n15278), .B(n15277), .S(SI_4_), .Z(n15279) );
  OAI21_X1 U16792 ( .B1(n15281), .B2(n15280), .A(n15279), .ZN(n15284) );
  XNOR2_X1 U16793 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15282) );
  XNOR2_X1 U16794 ( .A(n15282), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15283) );
  XNOR2_X1 U16795 ( .A(n15284), .B(n15283), .ZN(n15285) );
  XOR2_X1 U16796 ( .A(n15286), .B(n15285), .Z(n15287) );
  XNOR2_X1 U16797 ( .A(n15288), .B(n15287), .ZN(SUB_1596_U4) );
  XOR2_X1 U16798 ( .A(n15290), .B(n15289), .Z(SUB_1596_U59) );
  XNOR2_X1 U16799 ( .A(n15291), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16800 ( .B1(n15293), .B2(n15292), .A(n15301), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16801 ( .A(n15295), .B(n15294), .ZN(SUB_1596_U56) );
  OAI21_X1 U16802 ( .B1(n15298), .B2(n15297), .A(n15296), .ZN(n15299) );
  XNOR2_X1 U16803 ( .A(n15299), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16804 ( .A(n15301), .B(n15300), .Z(SUB_1596_U5) );
  NAND2_X1 U7283 ( .A1(n14858), .A2(n7368), .ZN(n10829) );
  CLKBUF_X1 U7280 ( .A(n8884), .Z(n6645) );
  CLKBUF_X1 U7281 ( .A(n9165), .Z(n9382) );
  CLKBUF_X1 U7282 ( .A(n12009), .Z(n6637) );
  CLKBUF_X1 U7306 ( .A(n10480), .Z(n6641) );
  CLKBUF_X1 U7338 ( .A(n8864), .Z(n6681) );
  OAI21_X1 U7422 ( .B1(n9604), .B2(n12551), .A(n10829), .ZN(n10969) );
  AOI22_X1 U7530 ( .A1(n10969), .A2(n10970), .B1(n9605), .B2(n12419), .ZN(
        n11027) );
  NOR2_X1 U7563 ( .A1(n9586), .A2(n12524), .ZN(n9590) );
  OR2_X1 U7656 ( .A1(n11772), .A2(n11771), .ZN(n15308) );
endmodule

