

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575;

  AOI21_X1 U3661 ( .B1(n6193), .B2(n5322), .A(n5961), .ZN(n5966) );
  INV_X1 U3662 ( .A(n7426), .ZN(n7412) );
  INV_X2 U3663 ( .A(n4049), .ZN(n6447) );
  NAND2_X1 U3664 ( .A1(n4773), .A2(n4772), .ZN(n4847) );
  INV_X1 U3665 ( .A(n5024), .ZN(n5322) );
  CLKBUF_X2 U3666 ( .A(n3829), .Z(n3629) );
  CLKBUF_X2 U3667 ( .A(n3837), .Z(n3800) );
  NAND4_X1 U3668 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n5454)
         );
  AND2_X2 U3669 ( .A1(n3649), .A2(n6960), .ZN(n3837) );
  AOI21_X1 U3670 ( .B1(n3826), .B2(INSTQUEUE_REG_1__1__SCAN_IN), .A(n3731), 
        .ZN(n3732) );
  NAND2_X2 U3671 ( .A1(n5024), .A2(n5924), .ZN(n5947) );
  NAND2_X1 U3672 ( .A1(n3760), .A2(n3763), .ZN(n4142) );
  OR2_X1 U3673 ( .A1(n6184), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3870) );
  OR2_X1 U3674 ( .A1(n5623), .A2(n5284), .ZN(n4282) );
  AND2_X1 U3675 ( .A1(n6083), .A2(n6082), .ZN(n6156) );
  CLKBUF_X3 U3676 ( .A(n3759), .Z(n3634) );
  AND2_X2 U3677 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6960) );
  INV_X1 U3678 ( .A(n7428), .ZN(n7396) );
  BUF_X2 U3679 ( .A(n4905), .Z(n3627) );
  NAND4_X1 U3680 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n4905)
         );
  NAND2_X1 U3681 ( .A1(n3914), .A2(n3913), .ZN(n3953) );
  OAI21_X1 U3682 ( .B1(n7246), .B2(STATE2_REG_0__SCAN_IN), .A(n3912), .ZN(
        n3914) );
  CLKBUF_X1 U3683 ( .A(n6157), .Z(n6546) );
  OAI21_X1 U3684 ( .B1(n6477), .B2(n6551), .A(n6157), .ZN(n6441) );
  AND2_X1 U3685 ( .A1(n6085), .A2(n6084), .ZN(n6432) );
  NAND2_X1 U3686 ( .A1(n4073), .A2(n3636), .ZN(n6060) );
  OR2_X1 U3687 ( .A1(n6128), .A2(n6079), .ZN(n6083) );
  CLKBUF_X1 U3688 ( .A(n6128), .Z(n6446) );
  NAND2_X1 U3689 ( .A1(n4313), .A2(n4312), .ZN(n5699) );
  AND2_X1 U3690 ( .A1(n5846), .A2(n6466), .ZN(n4057) );
  OR2_X1 U3691 ( .A1(n4030), .A2(n4029), .ZN(n4036) );
  OR2_X2 U3692 ( .A1(n4042), .A2(n4041), .ZN(n4049) );
  OR2_X1 U3693 ( .A1(n3993), .A2(n4029), .ZN(n4000) );
  NAND2_X1 U3694 ( .A1(n3992), .A2(n4018), .ZN(n3993) );
  NAND2_X2 U3695 ( .A1(n6392), .A2(n4783), .ZN(n6391) );
  BUF_X2 U3696 ( .A(n4249), .Z(n5187) );
  AND2_X2 U3697 ( .A1(n4694), .A2(n4813), .ZN(n4811) );
  NAND2_X2 U3699 ( .A1(n7118), .A2(n6119), .ZN(n6357) );
  NAND2_X1 U3700 ( .A1(n3896), .A2(n3895), .ZN(n5167) );
  NAND2_X1 U3701 ( .A1(n5269), .A2(n5268), .ZN(n5326) );
  CLKBUF_X1 U3702 ( .A(n4631), .Z(n7436) );
  XNOR2_X1 U3703 ( .A(n4847), .B(n4774), .ZN(n5522) );
  NAND2_X1 U3704 ( .A1(n5948), .A2(n5322), .ZN(n5963) );
  INV_X2 U3705 ( .A(n4775), .ZN(n5924) );
  NAND2_X1 U3706 ( .A1(n3631), .A2(n3633), .ZN(n4775) );
  BUF_X2 U3707 ( .A(n3757), .Z(n4915) );
  AND4_X1 U3708 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3756)
         );
  CLKBUF_X2 U3709 ( .A(n3856), .Z(n3635) );
  INV_X2 U3710 ( .A(n6489), .ZN(n3628) );
  BUF_X2 U3711 ( .A(n3683), .Z(n5980) );
  AND4_X1 U3712 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3753)
         );
  NAND2_X2 U3713 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7525), .ZN(n7071) );
  AND4_X1 U3714 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3755)
         );
  AND4_X1 U3715 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3754)
         );
  BUF_X2 U3716 ( .A(n3799), .Z(n5972) );
  BUF_X2 U3717 ( .A(n3828), .Z(n5975) );
  CLKBUF_X1 U3718 ( .A(n3830), .Z(n3677) );
  CLKBUF_X2 U3719 ( .A(n3740), .Z(n4419) );
  OR2_X2 U3720 ( .A1(n7522), .A2(STATE_REG_2__SCAN_IN), .ZN(n7056) );
  AND2_X2 U3721 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5435), .ZN(n7167) );
  BUF_X2 U3722 ( .A(n3826), .Z(n3630) );
  BUF_X2 U3723 ( .A(n3855), .Z(n5973) );
  BUF_X2 U3724 ( .A(n3808), .Z(n5983) );
  AND2_X2 U3725 ( .A1(n5602), .A2(n7161), .ZN(n7205) );
  NOR2_X2 U3726 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U3727 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3631)
         );
  NAND4_X1 U3728 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3632)
         );
  NAND2_X2 U3729 ( .A1(n3818), .A2(n3817), .ZN(n3887) );
  NAND4_X1 U3730 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3633)
         );
  NOR2_X2 U3731 ( .A1(n5326), .A2(n5325), .ZN(n5584) );
  NOR2_X2 U3732 ( .A1(n6288), .A2(n6090), .ZN(n6261) );
  OR2_X2 U3733 ( .A1(n6329), .A2(n6290), .ZN(n6288) );
  INV_X1 U3734 ( .A(n4568), .ZN(n4546) );
  AND2_X1 U3735 ( .A1(n3776), .A2(n4755), .ZN(n4654) );
  AND2_X1 U3736 ( .A1(n4693), .A2(n5454), .ZN(n3759) );
  INV_X1 U3737 ( .A(n3627), .ZN(n4693) );
  AND2_X1 U3738 ( .A1(n4276), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4242)
         );
  NAND2_X1 U3740 ( .A1(n3991), .A2(n3990), .ZN(n4018) );
  AND2_X1 U3741 ( .A1(n6464), .A2(n4060), .ZN(n4064) );
  NAND2_X1 U3742 ( .A1(n4028), .A2(n4084), .ZN(n4042) );
  AND2_X1 U3743 ( .A1(n4922), .A2(n3627), .ZN(n4084) );
  NAND2_X1 U3744 ( .A1(n3768), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3924) );
  INV_X1 U3745 ( .A(n4279), .ZN(n5999) );
  NAND2_X1 U3746 ( .A1(n4388), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4392)
         );
  NOR2_X2 U3747 ( .A1(n4282), .A2(n5283), .ZN(n5625) );
  NOR2_X1 U3748 ( .A1(n4274), .A2(n4144), .ZN(n4276) );
  INV_X1 U3749 ( .A(n4246), .ZN(n4262) );
  NAND2_X1 U3750 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4262), .ZN(n4274)
         );
  AND2_X1 U3752 ( .A1(n4654), .A2(n3788), .ZN(n4777) );
  NAND2_X1 U3753 ( .A1(n4652), .A2(n3784), .ZN(n3817) );
  AND2_X1 U3754 ( .A1(n5120), .A2(n5233), .ZN(n5128) );
  AND2_X1 U3755 ( .A1(n7390), .A2(n5446), .ZN(n7426) );
  NAND2_X1 U3756 ( .A1(n5031), .A2(n3954), .ZN(n3977) );
  NAND2_X1 U3757 ( .A1(n4085), .A2(n4084), .ZN(n4127) );
  AND2_X1 U3758 ( .A1(n5909), .A2(n4058), .ZN(n6464) );
  OR2_X2 U3759 ( .A1(n3700), .A2(n3699), .ZN(n3763) );
  INV_X1 U3760 ( .A(n5628), .ZN(n5592) );
  OR2_X1 U3761 ( .A1(n7165), .A2(n5436), .ZN(n7390) );
  OR2_X1 U3762 ( .A1(n6196), .A2(n4737), .ZN(n4757) );
  AOI21_X1 U3763 ( .B1(n4240), .B2(n4546), .A(n4239), .ZN(n5623) );
  OR2_X1 U3764 ( .A1(n4392), .A2(n6417), .ZN(n4374) );
  AND2_X1 U3765 ( .A1(n4148), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4388)
         );
  NAND2_X1 U3766 ( .A1(n4404), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4408)
         );
  AND2_X1 U3767 ( .A1(n6152), .A2(n6105), .ZN(n6286) );
  OR2_X1 U3768 ( .A1(n6323), .A2(n6322), .ZN(n6325) );
  NOR2_X1 U3769 ( .A1(n4519), .A2(n4530), .ZN(n4516) );
  NAND2_X1 U3770 ( .A1(n4516), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4515)
         );
  NOR2_X1 U3771 ( .A1(n4369), .A2(n5863), .ZN(n4564) );
  NAND2_X1 U3772 ( .A1(n4354), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4369)
         );
  NAND2_X1 U3773 ( .A1(n5725), .A2(n5724), .ZN(n5723) );
  AND2_X1 U3774 ( .A1(n4298), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4314)
         );
  INV_X1 U3775 ( .A(n5578), .ZN(n4313) );
  AOI21_X1 U3776 ( .B1(n4245), .B2(n4546), .A(n4244), .ZN(n5284) );
  AOI21_X1 U3777 ( .B1(n4281), .B2(n4546), .A(n4280), .ZN(n5021) );
  INV_X1 U3778 ( .A(n3993), .ZN(n4281) );
  AOI21_X1 U3779 ( .B1(n5233), .B2(n4546), .A(n4265), .ZN(n4887) );
  AND2_X1 U3780 ( .A1(n6024), .A2(n6023), .ZN(n6191) );
  NAND2_X1 U3781 ( .A1(n6326), .A2(n6327), .ZN(n6329) );
  AND2_X1 U3782 ( .A1(n6125), .A2(n6544), .ZN(n6326) );
  AND2_X1 U3783 ( .A1(n6132), .A2(n6124), .ZN(n6125) );
  NOR2_X2 U3784 ( .A1(n6334), .A2(n6133), .ZN(n6132) );
  OR2_X1 U3785 ( .A1(n5913), .A2(n5912), .ZN(n6301) );
  NOR2_X2 U3786 ( .A1(n6301), .A2(n6300), .ZN(n6350) );
  CLKBUF_X1 U3787 ( .A(n5845), .Z(n5847) );
  AND3_X1 U3788 ( .A1(n4878), .A2(n5939), .A3(n4877), .ZN(n4879) );
  INV_X1 U3789 ( .A(n4870), .ZN(n4868) );
  INV_X1 U3790 ( .A(n4871), .ZN(n4869) );
  NAND2_X1 U3791 ( .A1(n3770), .A2(n3769), .ZN(n3818) );
  OR2_X1 U3792 ( .A1(n3924), .A2(n4787), .ZN(n3770) );
  NAND2_X1 U3793 ( .A1(n3892), .A2(n3891), .ZN(n3895) );
  OR2_X1 U3794 ( .A1(n3924), .A2(n6074), .ZN(n3892) );
  INV_X1 U3795 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4787) );
  CLKBUF_X1 U3796 ( .A(n3640), .Z(n6963) );
  AND2_X1 U3797 ( .A1(n5292), .A2(n5756), .ZN(n5295) );
  AND2_X1 U3798 ( .A1(n5757), .A2(n5756), .ZN(n5765) );
  AND4_X1 U3799 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3734)
         );
  AND4_X1 U3800 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3733)
         );
  BUF_X1 U3801 ( .A(n3763), .Z(n4922) );
  AND2_X1 U3802 ( .A1(n7390), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U3803 ( .A1(n5458), .A2(n5457), .ZN(n7415) );
  INV_X1 U3804 ( .A(n7105), .ZN(n7114) );
  NAND2_X1 U3805 ( .A1(n4842), .A2(n4780), .ZN(n6392) );
  OR2_X1 U3806 ( .A1(n6000), .A2(n6401), .ZN(n5439) );
  NOR2_X1 U3807 ( .A1(n6146), .A2(n6145), .ZN(n7529) );
  AND2_X1 U3808 ( .A1(n6343), .A2(n6342), .ZN(n7526) );
  AND2_X1 U3809 ( .A1(n6347), .A2(n6299), .ZN(n7116) );
  INV_X1 U3810 ( .A(n7132), .ZN(n7147) );
  AND2_X1 U3811 ( .A1(n6237), .A2(n6236), .ZN(n6507) );
  AOI21_X1 U3812 ( .B1(n6087), .B2(n4049), .A(n6086), .ZN(n6089) );
  AOI21_X1 U3813 ( .B1(n6432), .B2(n6531), .A(n6477), .ZN(n6086) );
  OR2_X1 U3814 ( .A1(n6156), .A2(n6155), .ZN(n6547) );
  AND2_X1 U3815 ( .A1(n4663), .A2(n4643), .ZN(n7238) );
  INV_X1 U3816 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6175) );
  INV_X1 U3817 ( .A(n5187), .ZN(n5178) );
  INV_X1 U3818 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6074) );
  AND2_X1 U3819 ( .A1(n5182), .A2(n5038), .ZN(n5365) );
  INV_X1 U3820 ( .A(n5194), .ZN(n5229) );
  AND2_X1 U3821 ( .A1(n6261), .A2(n6260), .ZN(n6249) );
  NAND2_X1 U3822 ( .A1(n6350), .A2(n6349), .ZN(n5893) );
  INV_X1 U3823 ( .A(n6447), .ZN(n6477) );
  INV_X1 U3824 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3923) );
  AND2_X1 U3825 ( .A1(n6356), .A2(n4576), .ZN(n6049) );
  OR2_X1 U3826 ( .A1(n6395), .A2(n4074), .ZN(n3636) );
  INV_X1 U3827 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3881) );
  NAND2_X1 U3828 ( .A1(n4926), .A2(n3633), .ZN(n4768) );
  NAND2_X1 U3829 ( .A1(n5376), .A2(n5475), .ZN(n3637) );
  AND4_X1 U3830 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3638)
         );
  AND4_X1 U3831 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3639)
         );
  INV_X1 U3832 ( .A(n3975), .ZN(n3976) );
  OR2_X1 U3833 ( .A1(n3814), .A2(n3813), .ZN(n3916) );
  INV_X1 U3834 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U3835 ( .A1(n4142), .A2(n4899), .ZN(n3701) );
  INV_X1 U3836 ( .A(n3953), .ZN(n3954) );
  INV_X1 U3837 ( .A(n4127), .ZN(n4134) );
  OR2_X1 U3838 ( .A1(n3964), .A2(n3963), .ZN(n3994) );
  AND2_X1 U3839 ( .A1(n3758), .A2(n6119), .ZN(n3761) );
  AND2_X1 U3840 ( .A1(n5454), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4089) );
  OR2_X1 U3841 ( .A1(n4018), .A2(n4017), .ZN(n4028) );
  NOR2_X1 U3842 ( .A1(n4577), .A2(n6048), .ZN(n4149) );
  AND2_X1 U3843 ( .A1(n4147), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4404)
         );
  NOR2_X1 U3844 ( .A1(n4293), .A2(n4145), .ZN(n4298) );
  INV_X1 U3845 ( .A(n3764), .ZN(n3760) );
  INV_X1 U3846 ( .A(n6130), .ZN(n6078) );
  OR2_X1 U3847 ( .A1(n4142), .A2(n4768), .ZN(n4715) );
  AND2_X1 U3848 ( .A1(n4089), .A2(n3764), .ZN(n4085) );
  NAND2_X1 U3849 ( .A1(n3899), .A2(n3898), .ZN(n4137) );
  OR2_X1 U3850 ( .A1(n3664), .A2(n3663), .ZN(n3764) );
  INV_X1 U3851 ( .A(n6194), .ZN(n5960) );
  INV_X1 U3852 ( .A(n3763), .ZN(n6120) );
  AND4_X1 U3853 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3735)
         );
  OR2_X1 U3854 ( .A1(n4374), .A2(n6239), .ZN(n4577) );
  AND2_X1 U3855 ( .A1(n4564), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4537)
         );
  AND2_X1 U3856 ( .A1(n4330), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4354)
         );
  NOR2_X1 U3857 ( .A1(n6416), .A2(n4076), .ZN(n4077) );
  NAND2_X1 U3858 ( .A1(n5924), .A2(n5322), .ZN(n5956) );
  INV_X1 U3859 ( .A(n5830), .ZN(n5732) );
  OR2_X1 U3860 ( .A1(n5327), .A2(n7099), .ZN(n5325) );
  NAND2_X1 U3861 ( .A1(n4000), .A2(n3999), .ZN(n4002) );
  INV_X1 U3862 ( .A(n3703), .ZN(n6962) );
  NAND2_X1 U3863 ( .A1(n3787), .A2(n4594), .ZN(n4631) );
  NAND2_X1 U3864 ( .A1(n5032), .A2(n7161), .ZN(n3942) );
  AND3_X1 U3865 ( .A1(n5233), .A2(n5288), .A3(n5062), .ZN(n5761) );
  AND3_X1 U3866 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7161), .A3(n4898), .ZN(
        n4927) );
  NOR2_X2 U3867 ( .A1(n4647), .A2(n3785), .ZN(n4618) );
  NOR2_X1 U3868 ( .A1(n4482), .A2(n6450), .ZN(n4446) );
  AND2_X1 U3869 ( .A1(n6119), .A2(n4915), .ZN(n6118) );
  NOR2_X1 U3870 ( .A1(n6050), .A2(n4585), .ZN(n6189) );
  AND2_X1 U3871 ( .A1(n6356), .A2(n6104), .ZN(n6152) );
  NAND2_X1 U3872 ( .A1(n4537), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4519)
         );
  OR2_X1 U3873 ( .A1(n5723), .A2(n4371), .ZN(n4372) );
  AND2_X1 U3874 ( .A1(n4314), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4330)
         );
  NAND2_X1 U3875 ( .A1(n5625), .A2(n5318), .ZN(n5578) );
  NAND2_X1 U3876 ( .A1(n4139), .A2(n4138), .ZN(n6202) );
  INV_X1 U3877 ( .A(n6024), .ZN(n6252) );
  NAND2_X1 U3878 ( .A1(n5853), .A2(n5852), .ZN(n5913) );
  NAND2_X1 U3879 ( .A1(n4869), .A2(n4868), .ZN(n4880) );
  AND3_X1 U3880 ( .A1(n3783), .A2(n3782), .A3(n3781), .ZN(n3784) );
  NAND2_X1 U3881 ( .A1(n3930), .A2(n3929), .ZN(n5165) );
  OR2_X1 U3882 ( .A1(n6202), .A2(n4732), .ZN(n6069) );
  OR2_X1 U3883 ( .A1(n5234), .A2(n5233), .ZN(n5369) );
  NAND2_X1 U3884 ( .A1(n3942), .A2(n3941), .ZN(n5031) );
  INV_X1 U3885 ( .A(n5761), .ZN(n5816) );
  AND2_X1 U3886 ( .A1(n4940), .A2(n5187), .ZN(n5062) );
  OR2_X1 U3887 ( .A1(n5592), .A2(n5379), .ZN(n5535) );
  NAND2_X1 U3888 ( .A1(n4618), .A2(n5454), .ZN(n6197) );
  NAND2_X1 U3889 ( .A1(n4483), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4482)
         );
  AND2_X1 U3890 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4146), .ZN(n4483)
         );
  AND2_X1 U3891 ( .A1(n7390), .A2(n5440), .ZN(n7428) );
  AND2_X1 U3892 ( .A1(n6014), .A2(n5452), .ZN(n7409) );
  OR2_X1 U3893 ( .A1(n5893), .A2(n5894), .ZN(n6336) );
  BUF_X1 U3894 ( .A(n4775), .Z(n5962) );
  NAND2_X1 U3895 ( .A1(n6049), .A2(n6051), .ZN(n6050) );
  AND2_X1 U3896 ( .A1(n6392), .A2(n6121), .ZN(n7539) );
  INV_X1 U3897 ( .A(n5454), .ZN(n4668) );
  INV_X1 U3898 ( .A(n6152), .ZN(n6323) );
  AOI21_X1 U3899 ( .B1(n6348), .B2(n6347), .A(n6346), .ZN(n7348) );
  XNOR2_X1 U3900 ( .A(n5723), .B(n4371), .ZN(n5860) );
  NAND2_X1 U3901 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4293)
         );
  OR2_X1 U3902 ( .A1(n6202), .A2(n7499), .ZN(n4690) );
  INV_X1 U3903 ( .A(n7152), .ZN(n7143) );
  OR2_X1 U3904 ( .A1(n6063), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U3905 ( .A1(n4072), .A2(n4071), .ZN(n6424) );
  OR2_X1 U3906 ( .A1(n4067), .A2(n4066), .ZN(n6131) );
  INV_X1 U3907 ( .A(n6584), .ZN(n7239) );
  INV_X1 U3908 ( .A(n5369), .ZN(n5373) );
  OR3_X1 U3909 ( .A1(n5335), .A2(n3637), .A3(n5334), .ZN(n5361) );
  AND2_X1 U3910 ( .A1(n5128), .A2(n6180), .ZN(n5818) );
  OR3_X1 U3911 ( .A1(n4985), .A2(n3637), .A3(n4984), .ZN(n5011) );
  AND2_X1 U3912 ( .A1(n5094), .A2(n5038), .ZN(n5117) );
  AND2_X1 U3913 ( .A1(n4900), .A2(n6180), .ZN(n7571) );
  OR2_X1 U3914 ( .A1(n4690), .A2(n6197), .ZN(n4691) );
  INV_X1 U3915 ( .A(n7403), .ZN(n7418) );
  INV_X1 U3916 ( .A(n7409), .ZN(n7431) );
  AND2_X1 U3917 ( .A1(n4758), .A2(n7473), .ZN(n7118) );
  OAI21_X1 U3918 ( .B1(n6286), .B2(n6107), .A(n6265), .ZN(n6378) );
  OAI21_X1 U3919 ( .B1(n6117), .B2(n6146), .A(n6116), .ZN(n7397) );
  NOR2_X1 U3920 ( .A1(n7167), .A2(n4669), .ZN(n6992) );
  OR2_X1 U3921 ( .A1(n4690), .A2(n4667), .ZN(n7024) );
  OR2_X1 U3922 ( .A1(n4690), .A2(n7447), .ZN(n7433) );
  NAND2_X1 U3923 ( .A1(n5373), .A2(n6180), .ZN(n5687) );
  NAND2_X1 U3924 ( .A1(n5063), .A2(n6180), .ZN(n5368) );
  OR2_X1 U3925 ( .A1(n5298), .A2(n5288), .ZN(n5511) );
  OR2_X1 U3926 ( .A1(n5121), .A2(n6180), .ZN(n5507) );
  INV_X1 U3927 ( .A(n4982), .ZN(n5017) );
  NOR2_X2 U3928 ( .A1(n3642), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4726)
         );
  NOR2_X4 U3929 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6961) );
  AND2_X2 U3930 ( .A1(n4726), .A2(n6961), .ZN(n3740) );
  INV_X1 U3931 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3640) );
  NOR2_X2 U3932 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n3640), .ZN(n3648)
         );
  AND2_X2 U3933 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5162) );
  AND2_X2 U3934 ( .A1(n3648), .A2(n5162), .ZN(n3835) );
  AOI22_X1 U3935 ( .A1(n3740), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3646) );
  AND2_X2 U3936 ( .A1(n3648), .A2(n3649), .ZN(n3827) );
  AND2_X2 U3937 ( .A1(n4726), .A2(n6960), .ZN(n3829) );
  AOI22_X1 U3938 ( .A1(n3827), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3645) );
  INV_X1 U3939 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3641) );
  NOR2_X2 U3940 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n3641), .ZN(n3647)
         );
  AND2_X2 U3941 ( .A1(n3647), .A2(n5162), .ZN(n3901) );
  AND2_X2 U3942 ( .A1(n3642), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3650)
         );
  AND2_X2 U3943 ( .A1(n3650), .A2(n6960), .ZN(n3830) );
  AOI22_X1 U3944 ( .A1(n3901), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3644) );
  AND2_X2 U3945 ( .A1(n3647), .A2(n3650), .ZN(n3828) );
  AND2_X2 U3946 ( .A1(n6961), .A2(n5162), .ZN(n3838) );
  AOI22_X1 U3947 ( .A1(n3828), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3643) );
  AND2_X2 U3948 ( .A1(n3647), .A2(n4726), .ZN(n3856) );
  AND2_X2 U3949 ( .A1(n3647), .A2(n3649), .ZN(n3826) );
  AOI22_X1 U3950 ( .A1(n3856), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3654) );
  AND2_X2 U3951 ( .A1(n4726), .A2(n3648), .ZN(n3836) );
  AOI22_X1 U3952 ( .A1(n3836), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3653) );
  AND2_X2 U3953 ( .A1(n3648), .A2(n3650), .ZN(n3805) );
  AND2_X2 U3954 ( .A1(n3649), .A2(n6961), .ZN(n3855) );
  AOI22_X1 U3955 ( .A1(n3805), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3652) );
  AND2_X2 U3956 ( .A1(n3650), .A2(n6961), .ZN(n3799) );
  AND2_X2 U3957 ( .A1(n6960), .A2(n5162), .ZN(n3808) );
  AOI22_X1 U3958 ( .A1(n3799), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3651) );
  NAND2_X2 U3959 ( .A1(n3639), .A2(n3638), .ZN(n3757) );
  INV_X2 U3960 ( .A(n3757), .ZN(n4656) );
  AOI22_X1 U3961 ( .A1(n3740), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U3962 ( .A1(n3827), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U3963 ( .A1(n3901), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U3964 ( .A1(n3828), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U3965 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3664)
         );
  AOI22_X1 U3966 ( .A1(n3856), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U3967 ( .A1(n3836), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U3968 ( .A1(n3805), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U3969 ( .A1(n3799), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U3970 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3663)
         );
  AOI22_X1 U3971 ( .A1(n3856), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U3972 ( .A1(n3836), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U3973 ( .A1(n3740), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U3974 ( .A1(n3830), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U3975 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3674)
         );
  AOI22_X1 U3976 ( .A1(n3829), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        INSTQUEUE_REG_13__7__SCAN_IN), .B2(n3901), .ZN(n3672) );
  AOI22_X1 U3977 ( .A1(n3827), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3828), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U3978 ( .A1(n3855), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U3979 ( .A1(n3835), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U3980 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3673)
         );
  OR2_X2 U3981 ( .A1(n3674), .A2(n3673), .ZN(n6119) );
  NAND3_X1 U3982 ( .A1(n4656), .A2(n3764), .A3(n6119), .ZN(n3703) );
  BUF_X1 U3983 ( .A(n3835), .Z(n3675) );
  AOI22_X1 U3984 ( .A1(n4419), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3682) );
  BUF_X1 U3985 ( .A(n3827), .Z(n3676) );
  AOI22_X1 U3986 ( .A1(n3676), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3681) );
  BUF_X1 U3987 ( .A(n3901), .Z(n3807) );
  AOI22_X1 U3988 ( .A1(n3807), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3680) );
  BUF_X1 U3989 ( .A(n3838), .Z(n3678) );
  AOI22_X1 U3990 ( .A1(n3828), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U3991 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3690)
         );
  AOI22_X1 U3992 ( .A1(n3856), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U3994 ( .A1(n3683), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3687) );
  BUF_X1 U3995 ( .A(n3805), .Z(n3684) );
  AOI22_X1 U3996 ( .A1(n3684), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U3997 ( .A1(n3799), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U3998 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3689)
         );
  OR2_X2 U3999 ( .A1(n3690), .A2(n3689), .ZN(n4899) );
  AOI22_X1 U4000 ( .A1(n3836), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4001 ( .A1(n3740), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4002 ( .A1(n3805), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4003 ( .A1(n3799), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4004 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3700)
         );
  AOI22_X1 U4005 ( .A1(n3835), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4006 ( .A1(n3827), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4007 ( .A1(n3856), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4008 ( .A1(n3828), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3695) );
  NAND4_X1 U4009 ( .A1(n3698), .A2(n3697), .A3(n3696), .A4(n3695), .ZN(n3699)
         );
  NOR2_X1 U4010 ( .A1(n4899), .A2(n6120), .ZN(n3846) );
  NAND2_X1 U4011 ( .A1(n3703), .A2(n3846), .ZN(n3702) );
  NAND2_X1 U4012 ( .A1(n3702), .A2(n3701), .ZN(n3715) );
  NAND2_X1 U4013 ( .A1(n4656), .A2(n3763), .ZN(n4781) );
  AOI22_X1 U4014 ( .A1(n3740), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4015 ( .A1(n3827), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4016 ( .A1(n3901), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4017 ( .A1(n3828), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4018 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3713)
         );
  AOI22_X1 U4019 ( .A1(n3856), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4020 ( .A1(n3836), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4021 ( .A1(n3805), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4022 ( .A1(n3799), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4023 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3712)
         );
  OR2_X2 U4024 ( .A1(n3713), .A2(n3712), .ZN(n4926) );
  NAND2_X1 U4025 ( .A1(n4781), .A2(n4926), .ZN(n3780) );
  OAI21_X1 U4026 ( .B1(n6962), .B2(n6118), .A(n3780), .ZN(n3714) );
  NOR2_X1 U4027 ( .A1(n3715), .A2(n3714), .ZN(n4595) );
  NAND2_X1 U4028 ( .A1(n3740), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U4029 ( .A1(n3835), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3718)
         );
  NAND2_X1 U4030 ( .A1(n3828), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3717) );
  NAND2_X1 U4031 ( .A1(n3901), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3716)
         );
  NAND2_X1 U4032 ( .A1(n3836), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3723)
         );
  NAND2_X1 U4033 ( .A1(n3856), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3722) );
  NAND2_X1 U4034 ( .A1(n3805), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U4035 ( .A1(n3837), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4036 ( .A1(n3829), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3727)
         );
  NAND2_X1 U4037 ( .A1(n3827), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4038 ( .A1(n3830), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4039 ( .A1(n3838), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3724)
         );
  NAND2_X1 U4040 ( .A1(n3855), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4041 ( .A1(n3808), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3729)
         );
  NAND2_X1 U4042 ( .A1(n3799), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3728) );
  NAND3_X1 U4043 ( .A1(n3730), .A2(n3729), .A3(n3728), .ZN(n3731) );
  NAND2_X1 U4044 ( .A1(n4595), .A2(n4693), .ZN(n3786) );
  NAND2_X1 U4045 ( .A1(n3856), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3739) );
  NAND2_X1 U4046 ( .A1(n3836), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3738)
         );
  NAND2_X1 U4047 ( .A1(n3826), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4048 ( .A1(n3837), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4049 ( .A1(n3740), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4050 ( .A1(n3835), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3743)
         );
  NAND2_X1 U4051 ( .A1(n3901), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3742)
         );
  NAND2_X1 U4052 ( .A1(n3830), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4053 ( .A1(n3827), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4054 ( .A1(n3829), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3747)
         );
  NAND2_X1 U4055 ( .A1(n3828), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4056 ( .A1(n3838), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3745)
         );
  NAND2_X1 U4057 ( .A1(n3805), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3752) );
  NAND2_X1 U4058 ( .A1(n3799), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3751) );
  NAND2_X1 U4059 ( .A1(n3855), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3750) );
  NAND2_X1 U4060 ( .A1(n3808), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3749)
         );
  NAND2_X1 U4061 ( .A1(n3786), .A2(n4668), .ZN(n3772) );
  NAND2_X1 U4062 ( .A1(n6120), .A2(n3757), .ZN(n3758) );
  OAI211_X1 U4063 ( .C1(n4142), .C2(n4915), .A(n3761), .B(n4926), .ZN(n3775)
         );
  OR2_X2 U4064 ( .A1(n3775), .A2(n4899), .ZN(n4647) );
  INV_X1 U4065 ( .A(n4647), .ZN(n3767) );
  NAND2_X1 U4066 ( .A1(n3761), .A2(n4753), .ZN(n4619) );
  INV_X1 U4067 ( .A(STATE_REG_2__SCAN_IN), .ZN(n3762) );
  XNOR2_X1 U4068 ( .A(n3762), .B(STATE_REG_1__SCAN_IN), .ZN(n7509) );
  NOR2_X1 U4069 ( .A1(n3627), .A2(n7509), .ZN(n3789) );
  NAND2_X1 U4070 ( .A1(n4781), .A2(n3764), .ZN(n3773) );
  OAI211_X1 U4071 ( .C1(n3789), .C2(n4922), .A(n4715), .B(n3773), .ZN(n3765)
         );
  AOI21_X1 U4072 ( .B1(n3634), .B2(n4619), .A(n3765), .ZN(n3766) );
  NAND3_X1 U4073 ( .A1(n3772), .A2(n3767), .A3(n3766), .ZN(n3768) );
  INV_X1 U4074 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7487) );
  AND2_X1 U4075 ( .A1(n7487), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4140) );
  NOR2_X1 U4076 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7481) );
  INV_X1 U4077 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U4078 ( .A1(n7481), .A2(n7161), .ZN(n4587) );
  MUX2_X1 U4079 ( .A(n4140), .B(n4587), .S(n6175), .Z(n3769) );
  AND2_X1 U4080 ( .A1(n4084), .A2(n4753), .ZN(n3771) );
  OR2_X1 U4081 ( .A1(n3772), .A2(n3771), .ZN(n4652) );
  INV_X1 U4082 ( .A(n3773), .ZN(n3774) );
  OAI21_X1 U4083 ( .B1(n3775), .B2(n3774), .A(n3627), .ZN(n3783) );
  NOR2_X1 U4084 ( .A1(n4926), .A2(n5454), .ZN(n3776) );
  INV_X1 U4085 ( .A(n4899), .ZN(n4755) );
  NAND2_X1 U4086 ( .A1(n4654), .A2(n6962), .ZN(n3779) );
  NAND2_X1 U4087 ( .A1(n7481), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3777) );
  AOI21_X1 U4088 ( .B1(n4899), .B2(n5454), .A(n3777), .ZN(n3778) );
  AND3_X1 U4089 ( .A1(n3779), .A2(n3778), .A3(n4715), .ZN(n3782) );
  OAI21_X1 U4090 ( .B1(n4619), .B2(n3780), .A(n3634), .ZN(n3781) );
  INV_X1 U4091 ( .A(n3887), .ZN(n3798) );
  OR2_X1 U4092 ( .A1(n3924), .A2(n6963), .ZN(n3792) );
  NAND2_X1 U4093 ( .A1(n4753), .A2(n4656), .ZN(n3785) );
  INV_X1 U4094 ( .A(n3786), .ZN(n3787) );
  NOR2_X1 U4095 ( .A1(n4142), .A2(n5454), .ZN(n4594) );
  NOR2_X1 U4096 ( .A1(n4922), .A2(n3627), .ZN(n3788) );
  NAND2_X1 U4097 ( .A1(n4777), .A2(n6118), .ZN(n4633) );
  OAI211_X1 U4098 ( .C1(n3789), .C2(n6197), .A(n4631), .B(n4633), .ZN(n3790)
         );
  NAND2_X1 U4099 ( .A1(n3790), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3794) );
  INV_X1 U4100 ( .A(n4587), .ZN(n3928) );
  INV_X1 U4101 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U4102 ( .A1(n5381), .A2(n6175), .ZN(n3791) );
  NAND2_X1 U4103 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5064) );
  AND2_X1 U4104 ( .A1(n3791), .A2(n5064), .ZN(n5529) );
  INV_X1 U4105 ( .A(n4140), .ZN(n3927) );
  AOI22_X1 U4106 ( .A1(n3928), .A2(n5529), .B1(n3927), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3793) );
  NAND3_X1 U4107 ( .A1(n3792), .A2(n3794), .A3(n3793), .ZN(n3885) );
  INV_X1 U4108 ( .A(n3793), .ZN(n3796) );
  INV_X1 U4109 ( .A(n3794), .ZN(n3795) );
  OAI21_X1 U4110 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3796), .A(n3795), 
        .ZN(n3797) );
  NAND2_X2 U4111 ( .A1(n3885), .A2(n3797), .ZN(n3884) );
  XNOR2_X2 U4112 ( .A(n3798), .B(n3884), .ZN(n4892) );
  NAND2_X1 U4113 ( .A1(n4892), .A2(n7161), .ZN(n3816) );
  NAND2_X1 U4114 ( .A1(n4753), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4115 ( .A1(n3635), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4116 ( .A1(n4419), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3803) );
  BUF_X1 U4117 ( .A(n3830), .Z(n5982) );
  AOI22_X1 U4118 ( .A1(n3629), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4119 ( .A1(n5973), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4120 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3814)
         );
  INV_X1 U4121 ( .A(n3805), .ZN(n3806) );
  INV_X1 U4122 ( .A(n3806), .ZN(n3900) );
  AOI22_X1 U4123 ( .A1(n3683), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4124 ( .A1(n3807), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5981), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4125 ( .A1(n4557), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4126 ( .A1(n5975), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4127 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  INV_X1 U4128 ( .A(n3916), .ZN(n3819) );
  OR2_X1 U4129 ( .A1(n3899), .A2(n3819), .ZN(n3815) );
  NAND2_X1 U4130 ( .A1(n3816), .A2(n3815), .ZN(n3823) );
  OAI21_X2 U4131 ( .B1(n3818), .B2(n3817), .A(n3887), .ZN(n6184) );
  OR2_X1 U4132 ( .A1(n5454), .A2(n7161), .ZN(n3898) );
  OAI21_X1 U4133 ( .B1(n3819), .B2(n3898), .A(n3899), .ZN(n3820) );
  AOI21_X1 U4134 ( .B1(INSTQUEUE_REG_0__1__SCAN_IN), .B2(n4085), .A(n3820), 
        .ZN(n3821) );
  NAND2_X1 U4135 ( .A1(n3870), .A2(n3821), .ZN(n3822) );
  AND2_X2 U4136 ( .A1(n3823), .A2(n3822), .ZN(n3913) );
  INV_X1 U4137 ( .A(n3913), .ZN(n3825) );
  OR2_X1 U4138 ( .A1(n3823), .A2(n3822), .ZN(n3824) );
  AND2_X2 U4139 ( .A1(n3825), .A2(n3824), .ZN(n4249) );
  NAND2_X1 U4140 ( .A1(n4249), .A2(n4084), .ZN(n3850) );
  AOI22_X1 U4141 ( .A1(n3635), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3834) );
  BUF_X1 U4142 ( .A(n3827), .Z(n5981) );
  AOI22_X1 U4143 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5981), .B1(n5975), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4144 ( .A1(n3629), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4145 ( .A1(n5972), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4146 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3844)
         );
  BUF_X1 U4147 ( .A(n4419), .Z(n5971) );
  BUF_X1 U4148 ( .A(n3835), .Z(n4557) );
  AOI22_X1 U4149 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5971), .B1(n4557), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4150 ( .A1(n3683), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3841) );
  CLKBUF_X1 U4151 ( .A(n3901), .Z(n4226) );
  AOI22_X1 U4153 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4226), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4154 ( .A1(n3900), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4155 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3843)
         );
  OR2_X1 U4156 ( .A1(n3844), .A2(n3843), .ZN(n3915) );
  INV_X1 U4157 ( .A(n3915), .ZN(n3845) );
  XNOR2_X1 U4158 ( .A(n3845), .B(n3916), .ZN(n3848) );
  INV_X1 U4159 ( .A(n3846), .ZN(n3847) );
  AOI21_X1 U4160 ( .B1(n3848), .B2(n3634), .A(n3847), .ZN(n3849) );
  NAND2_X1 U4161 ( .A1(n3850), .A2(n3849), .ZN(n3880) );
  NAND2_X1 U4162 ( .A1(n3880), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4791)
         );
  NAND2_X1 U4163 ( .A1(n4085), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3865) );
  AOI21_X1 U4164 ( .B1(n4668), .B2(n3915), .A(n7161), .ZN(n3863) );
  AOI22_X1 U4165 ( .A1(n3683), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4166 ( .A1(n4419), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4167 ( .A1(n4557), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4168 ( .A1(n5982), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3851) );
  NAND4_X1 U4169 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3862)
         );
  AOI22_X1 U4170 ( .A1(n5981), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4171 ( .A1(n3629), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4172 ( .A1(n3900), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4173 ( .A1(n3635), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4174 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  OR2_X1 U4175 ( .A1(n3862), .A2(n3861), .ZN(n4043) );
  NAND2_X1 U4176 ( .A1(n4753), .A2(n4043), .ZN(n4039) );
  AND2_X1 U4177 ( .A1(n3863), .A2(n4039), .ZN(n3864) );
  NAND2_X1 U4178 ( .A1(n3865), .A2(n3864), .ZN(n3871) );
  INV_X1 U4179 ( .A(n3899), .ZN(n3868) );
  INV_X1 U4180 ( .A(n4043), .ZN(n3866) );
  XNOR2_X1 U4181 ( .A(n3866), .B(n3915), .ZN(n3867) );
  NAND2_X1 U4182 ( .A1(n3868), .A2(n3867), .ZN(n3872) );
  AND2_X1 U4183 ( .A1(n3871), .A2(n3872), .ZN(n3869) );
  NAND2_X1 U4184 ( .A1(n3870), .A2(n3869), .ZN(n3876) );
  INV_X1 U4185 ( .A(n3871), .ZN(n3874) );
  INV_X1 U4186 ( .A(n3872), .ZN(n3873) );
  NAND2_X1 U4187 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  NAND2_X2 U4188 ( .A1(n3876), .A2(n3875), .ZN(n6180) );
  NAND2_X1 U4189 ( .A1(n6180), .A2(n4084), .ZN(n3879) );
  INV_X1 U4190 ( .A(n3634), .ZN(n7169) );
  NAND2_X1 U4191 ( .A1(n4668), .A2(n4926), .ZN(n3917) );
  OAI21_X1 U4192 ( .B1(n7169), .B2(n3915), .A(n3917), .ZN(n3877) );
  INV_X1 U4193 ( .A(n3877), .ZN(n3878) );
  NAND2_X1 U4194 ( .A1(n3879), .A2(n3878), .ZN(n4616) );
  NAND2_X1 U4195 ( .A1(n4616), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4794)
         );
  NAND2_X1 U4196 ( .A1(n4791), .A2(n4794), .ZN(n3883) );
  INV_X1 U4197 ( .A(n3880), .ZN(n3882) );
  NAND2_X1 U4198 ( .A1(n3882), .A2(n3881), .ZN(n4792) );
  NAND2_X1 U4199 ( .A1(n3883), .A2(n4792), .ZN(n3921) );
  INV_X1 U4200 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4849) );
  OR2_X2 U4201 ( .A1(n3921), .A2(n4849), .ZN(n7120) );
  INV_X1 U4202 ( .A(n3884), .ZN(n3888) );
  INV_X1 U4203 ( .A(n3885), .ZN(n3886) );
  AOI21_X2 U4204 ( .B1(n3888), .B2(n3887), .A(n3886), .ZN(n3896) );
  INV_X1 U4205 ( .A(n3896), .ZN(n3894) );
  INV_X1 U4206 ( .A(n5064), .ZN(n3889) );
  AND2_X1 U4207 ( .A1(n3889), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4893)
         );
  INV_X1 U4208 ( .A(n4893), .ZN(n3925) );
  INV_X1 U4209 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U4210 ( .A1(n5064), .A2(n7462), .ZN(n3890) );
  AND2_X1 U4211 ( .A1(n3925), .A2(n3890), .ZN(n4987) );
  AOI22_X1 U4212 ( .A1(n4987), .A2(n3928), .B1(n3927), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3891) );
  INV_X1 U4213 ( .A(n3895), .ZN(n3893) );
  NAND2_X1 U4214 ( .A1(n3894), .A2(n3893), .ZN(n3897) );
  NAND2_X2 U4215 ( .A1(n3897), .A2(n5167), .ZN(n7246) );
  AOI22_X1 U4216 ( .A1(n3900), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4217 ( .A1(n4226), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4218 ( .A1(n5981), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4219 ( .A1(n5980), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4220 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3911)
         );
  AOI22_X1 U4221 ( .A1(n3635), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4222 ( .A1(n5972), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4223 ( .A1(n5982), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4224 ( .A1(n5971), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4225 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3910)
         );
  OR2_X1 U4226 ( .A1(n3911), .A2(n3910), .ZN(n3943) );
  AOI22_X1 U4227 ( .A1(n4137), .A2(n3943), .B1(n4085), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3912) );
  OR2_X1 U4228 ( .A1(n3914), .A2(n3913), .ZN(n4939) );
  NAND2_X2 U4229 ( .A1(n4939), .A2(n3953), .ZN(n4890) );
  INV_X1 U4230 ( .A(n4890), .ZN(n3920) );
  NAND2_X1 U4231 ( .A1(n3916), .A2(n3915), .ZN(n3945) );
  XNOR2_X1 U4232 ( .A(n3945), .B(n3943), .ZN(n3918) );
  OAI21_X1 U4233 ( .B1(n3918), .B2(n7169), .A(n3917), .ZN(n3919) );
  AOI21_X1 U4234 ( .B1(n3920), .B2(n4084), .A(n3919), .ZN(n7122) );
  NAND2_X1 U4235 ( .A1(n3921), .A2(n4849), .ZN(n7119) );
  INV_X1 U4236 ( .A(n7119), .ZN(n3922) );
  AOI21_X2 U4237 ( .B1(n7120), .B2(n7122), .A(n3922), .ZN(n3949) );
  NAND2_X1 U4238 ( .A1(n3949), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4860)
         );
  OR2_X1 U4239 ( .A1(n3924), .A2(n3923), .ZN(n3930) );
  INV_X1 U4240 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4112) );
  NAND2_X1 U4241 ( .A1(n4893), .A2(n4112), .ZN(n5289) );
  NAND2_X1 U4242 ( .A1(n3925), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3926) );
  NAND2_X1 U4243 ( .A1(n5289), .A2(n3926), .ZN(n5336) );
  AOI22_X1 U4244 ( .A1(n5336), .A2(n3928), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3927), .ZN(n3929) );
  XNOR2_X2 U4245 ( .A(n5167), .B(n5165), .ZN(n5032) );
  AOI22_X1 U4246 ( .A1(n4419), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4247 ( .A1(n5981), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4248 ( .A1(n4226), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4249 ( .A1(n5975), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4250 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3940)
         );
  AOI22_X1 U4251 ( .A1(n3635), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4252 ( .A1(n5980), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4253 ( .A1(n3900), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4254 ( .A1(n5972), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3935) );
  NAND4_X1 U4255 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3939)
         );
  OR2_X1 U4256 ( .A1(n3940), .A2(n3939), .ZN(n3967) );
  AOI22_X1 U4257 ( .A1(n4137), .A2(n3967), .B1(n4085), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3941) );
  XNOR2_X2 U4258 ( .A(n5031), .B(n3953), .ZN(n5233) );
  INV_X1 U4259 ( .A(n3943), .ZN(n3944) );
  NAND2_X1 U4260 ( .A1(n3945), .A2(n3944), .ZN(n3968) );
  INV_X1 U4261 ( .A(n3967), .ZN(n3946) );
  XNOR2_X1 U4262 ( .A(n3968), .B(n3946), .ZN(n3947) );
  AND2_X1 U4263 ( .A1(n3947), .A2(n3634), .ZN(n3948) );
  AOI21_X1 U4264 ( .B1(n5233), .B2(n4084), .A(n3948), .ZN(n4861) );
  NAND2_X1 U4265 ( .A1(n4860), .A2(n4861), .ZN(n3952) );
  INV_X1 U4266 ( .A(n3949), .ZN(n3951) );
  INV_X1 U4267 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4268 ( .A1(n3951), .A2(n3950), .ZN(n4859) );
  NAND2_X1 U4269 ( .A1(n3952), .A2(n4859), .ZN(n4876) );
  AOI22_X1 U4270 ( .A1(n4419), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4271 ( .A1(n5981), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4272 ( .A1(n4226), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4273 ( .A1(n5975), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4274 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3964)
         );
  AOI22_X1 U4275 ( .A1(n3635), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4276 ( .A1(n5980), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4277 ( .A1(n3900), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4278 ( .A1(n5972), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4279 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3963)
         );
  NAND2_X1 U4280 ( .A1(n4137), .A2(n3994), .ZN(n3966) );
  NAND2_X1 U4281 ( .A1(n4085), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U4282 ( .A1(n3966), .A2(n3965), .ZN(n3975) );
  XNOR2_X1 U4283 ( .A(n3977), .B(n3975), .ZN(n4266) );
  NAND2_X1 U4284 ( .A1(n4266), .A2(n4084), .ZN(n3971) );
  NAND2_X1 U4285 ( .A1(n3968), .A2(n3967), .ZN(n3996) );
  XNOR2_X1 U4286 ( .A(n3996), .B(n3994), .ZN(n3969) );
  NAND2_X1 U4287 ( .A1(n3969), .A2(n3634), .ZN(n3970) );
  NAND2_X1 U4288 ( .A1(n3971), .A2(n3970), .ZN(n3972) );
  XNOR2_X1 U4289 ( .A(n3972), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4875)
         );
  INV_X1 U4290 ( .A(n3972), .ZN(n3974) );
  INV_X1 U4291 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3973) );
  OAI22_X1 U4292 ( .A1(n4876), .A2(n4875), .B1(n3974), .B2(n3973), .ZN(n7125)
         );
  NOR2_X2 U4293 ( .A1(n3977), .A2(n3976), .ZN(n3991) );
  AOI22_X1 U4294 ( .A1(n3635), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4295 ( .A1(n5980), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4296 ( .A1(n4226), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4297 ( .A1(n4419), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4298 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3987)
         );
  AOI22_X1 U4299 ( .A1(n5981), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4300 ( .A1(n4557), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4301 ( .A1(n5972), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4302 ( .A1(n3677), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4303 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  OR2_X1 U4304 ( .A1(n3987), .A2(n3986), .ZN(n3997) );
  NAND2_X1 U4305 ( .A1(n4137), .A2(n3997), .ZN(n3989) );
  NAND2_X1 U4306 ( .A1(n4085), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3988) );
  NAND2_X1 U4307 ( .A1(n3989), .A2(n3988), .ZN(n3990) );
  OR2_X1 U4308 ( .A1(n3991), .A2(n3990), .ZN(n3992) );
  INV_X1 U4309 ( .A(n4084), .ZN(n4029) );
  INV_X1 U4310 ( .A(n3994), .ZN(n3995) );
  NOR2_X1 U4311 ( .A1(n3996), .A2(n3995), .ZN(n3998) );
  NAND2_X1 U4312 ( .A1(n3998), .A2(n3997), .ZN(n4031) );
  OAI211_X1 U4313 ( .C1(n3998), .C2(n3997), .A(n4031), .B(n3634), .ZN(n3999)
         );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4001) );
  XNOR2_X1 U4315 ( .A(n4002), .B(n4001), .ZN(n7127) );
  NAND2_X1 U4316 ( .A1(n7125), .A2(n7127), .ZN(n4004) );
  NAND2_X1 U4317 ( .A1(n4002), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4003)
         );
  NAND2_X1 U4318 ( .A1(n4004), .A2(n4003), .ZN(n5262) );
  AOI22_X1 U4319 ( .A1(n4419), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4320 ( .A1(n5981), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4321 ( .A1(n4226), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4322 ( .A1(n5975), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4323 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4014)
         );
  AOI22_X1 U4324 ( .A1(n3635), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4325 ( .A1(n5980), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4326 ( .A1(n3900), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4327 ( .A1(n5972), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4328 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  OR2_X1 U4329 ( .A1(n4014), .A2(n4013), .ZN(n4032) );
  NAND2_X1 U4330 ( .A1(n4137), .A2(n4032), .ZN(n4016) );
  NAND2_X1 U4331 ( .A1(n4085), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4015) );
  AND2_X1 U4332 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  NAND2_X1 U4333 ( .A1(n4018), .A2(n4017), .ZN(n4245) );
  INV_X1 U4334 ( .A(n4245), .ZN(n4019) );
  OR2_X1 U4335 ( .A1(n4042), .A2(n4019), .ZN(n4022) );
  XNOR2_X1 U4336 ( .A(n4031), .B(n4032), .ZN(n4020) );
  NAND2_X1 U4337 ( .A1(n4020), .A2(n3634), .ZN(n4021) );
  NAND2_X1 U4338 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  OR2_X1 U4339 ( .A1(n4023), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5260)
         );
  NAND2_X1 U4340 ( .A1(n5262), .A2(n5260), .ZN(n4024) );
  NAND2_X1 U4341 ( .A1(n4023), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5259)
         );
  NAND2_X1 U4342 ( .A1(n4024), .A2(n5259), .ZN(n7138) );
  NAND2_X1 U4343 ( .A1(n4137), .A2(n4043), .ZN(n4026) );
  NAND2_X1 U4344 ( .A1(n4085), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U4345 ( .A1(n4026), .A2(n4025), .ZN(n4027) );
  XNOR2_X2 U4346 ( .A(n4028), .B(n4027), .ZN(n4240) );
  INV_X1 U4347 ( .A(n4240), .ZN(n4030) );
  INV_X1 U4348 ( .A(n4031), .ZN(n4033) );
  NAND2_X1 U4349 ( .A1(n4033), .A2(n4032), .ZN(n4045) );
  XNOR2_X1 U4350 ( .A(n4045), .B(n4043), .ZN(n4034) );
  NAND2_X1 U4351 ( .A1(n4034), .A2(n3634), .ZN(n4035) );
  NAND2_X1 U4352 ( .A1(n4036), .A2(n4035), .ZN(n4037) );
  INV_X1 U4353 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7209) );
  XNOR2_X1 U4354 ( .A(n4037), .B(n7209), .ZN(n7137) );
  NAND2_X1 U4355 ( .A1(n7138), .A2(n7137), .ZN(n7136) );
  NAND2_X1 U4356 ( .A1(n4037), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4038)
         );
  NAND2_X1 U4357 ( .A1(n7136), .A2(n4038), .ZN(n5416) );
  INV_X1 U4358 ( .A(n4039), .ZN(n4040) );
  NAND2_X1 U4359 ( .A1(n4040), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4360 ( .A1(n3634), .A2(n4043), .ZN(n4044) );
  OR2_X1 U4361 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  NAND2_X1 U4362 ( .A1(n4049), .A2(n4046), .ZN(n4047) );
  INV_X1 U4363 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5428) );
  XNOR2_X1 U4364 ( .A(n4047), .B(n5428), .ZN(n5415) );
  NAND2_X1 U4365 ( .A1(n5416), .A2(n5415), .ZN(n5414) );
  NAND2_X1 U4366 ( .A1(n4047), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U4367 ( .A1(n5414), .A2(n4048), .ZN(n5692) );
  XNOR2_X1 U4368 ( .A(n6395), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5691)
         );
  NAND2_X1 U4369 ( .A1(n5692), .A2(n5691), .ZN(n5748) );
  NAND2_X1 U4370 ( .A1(n6447), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5747)
         );
  INV_X1 U4371 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n7212) );
  OR2_X1 U4372 ( .A1(n4049), .A2(n7212), .ZN(n5827) );
  INV_X1 U4373 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6948) );
  OR2_X1 U4374 ( .A1(n4049), .A2(n6948), .ZN(n5824) );
  AND2_X1 U4375 ( .A1(n5827), .A2(n5824), .ZN(n5868) );
  INV_X4 U4376 ( .A(n6447), .ZN(n6395) );
  INV_X1 U4377 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6955) );
  OR2_X1 U4378 ( .A1(n6395), .A2(n6955), .ZN(n5873) );
  AND2_X1 U4379 ( .A1(n5868), .A2(n5873), .ZN(n4050) );
  AND2_X1 U4380 ( .A1(n5747), .A2(n4050), .ZN(n4051) );
  NAND2_X1 U4381 ( .A1(n5748), .A2(n4051), .ZN(n4055) );
  NAND2_X1 U4382 ( .A1(n6395), .A2(n7212), .ZN(n5825) );
  NAND2_X1 U4383 ( .A1(n6395), .A2(n6948), .ZN(n5870) );
  NAND2_X1 U4384 ( .A1(n5825), .A2(n5870), .ZN(n4053) );
  NAND2_X1 U4385 ( .A1(n6395), .A2(n6955), .ZN(n5872) );
  INV_X1 U4386 ( .A(n5872), .ZN(n4052) );
  NOR2_X1 U4387 ( .A1(n4053), .A2(n4052), .ZN(n4054) );
  NAND2_X1 U4388 ( .A1(n4055), .A2(n4054), .ZN(n5845) );
  XNOR2_X1 U4389 ( .A(n6477), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5846)
         );
  NAND2_X1 U4390 ( .A1(n6447), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U4391 ( .A1(n6447), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4056) );
  AND2_X1 U4392 ( .A1(n6475), .A2(n4056), .ZN(n6466) );
  NAND2_X1 U4393 ( .A1(n5845), .A2(n4057), .ZN(n4061) );
  INV_X1 U4394 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U4395 ( .A1(n6395), .A2(n5848), .ZN(n5909) );
  INV_X1 U4396 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U4397 ( .A1(n6395), .A2(n5922), .ZN(n4058) );
  INV_X1 U4398 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6580) );
  AND2_X1 U4399 ( .A1(n6395), .A2(n6580), .ZN(n6467) );
  INV_X1 U4400 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5887) );
  AND2_X1 U4401 ( .A1(n6395), .A2(n5887), .ZN(n4059) );
  NOR2_X1 U4402 ( .A1(n6467), .A2(n4059), .ZN(n4060) );
  NAND2_X1 U4403 ( .A1(n4061), .A2(n4064), .ZN(n6454) );
  INV_X1 U4404 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5881) );
  INV_X1 U4405 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5923) );
  AND3_X1 U4406 ( .A1(n5887), .A2(n5881), .A3(n5923), .ZN(n4062) );
  AOI21_X1 U4407 ( .B1(n6454), .B2(n4062), .A(n6395), .ZN(n4067) );
  NAND2_X1 U4408 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6026) );
  INV_X1 U4409 ( .A(n6026), .ZN(n4063) );
  NAND2_X1 U4410 ( .A1(n4064), .A2(n4063), .ZN(n4065) );
  NOR2_X1 U4411 ( .A1(n5845), .A2(n4065), .ZN(n4066) );
  NAND2_X1 U4412 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6035) );
  AND2_X1 U4413 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6080) );
  AND2_X1 U4414 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U4415 ( .A1(n6080), .A2(n6040), .ZN(n6430) );
  OAI21_X1 U4416 ( .B1(n6035), .B2(n6430), .A(n6395), .ZN(n4068) );
  NAND2_X1 U4417 ( .A1(n6131), .A2(n4068), .ZN(n4072) );
  NOR2_X1 U4418 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6084) );
  NOR2_X1 U4419 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4069) );
  INV_X1 U4420 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6088) );
  INV_X1 U4421 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6531) );
  NAND4_X1 U4422 ( .A1(n6084), .A2(n4069), .A3(n6088), .A4(n6531), .ZN(n4070)
         );
  NAND2_X1 U4423 ( .A1(n6447), .A2(n4070), .ZN(n4071) );
  INV_X1 U4424 ( .A(n6424), .ZN(n4073) );
  INV_X1 U4425 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4074) );
  NAND2_X1 U4426 ( .A1(n6395), .A2(n4074), .ZN(n4075) );
  NAND2_X1 U4427 ( .A1(n6060), .A2(n4075), .ZN(n6416) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6414) );
  AND2_X1 U4429 ( .A1(n4049), .A2(n6414), .ZN(n4076) );
  INV_X1 U4430 ( .A(n4077), .ZN(n6406) );
  INV_X1 U4431 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6505) );
  AND2_X1 U4432 ( .A1(n4049), .A2(n6505), .ZN(n4078) );
  NOR2_X2 U4433 ( .A1(n6406), .A2(n4078), .ZN(n6063) );
  INV_X1 U4434 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4079) );
  NAND2_X1 U4435 ( .A1(n6505), .A2(n4079), .ZN(n6042) );
  NOR2_X1 U4436 ( .A1(n6042), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4080)
         );
  NOR2_X1 U4437 ( .A1(n6395), .A2(n4080), .ZN(n6058) );
  OAI22_X1 U4438 ( .A1(n6063), .A2(n6058), .B1(n6447), .B2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4082) );
  INV_X1 U4439 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6096) );
  XNOR2_X1 U4440 ( .A(n6477), .B(n6096), .ZN(n4081) );
  XNOR2_X1 U4441 ( .A(n4082), .B(n4081), .ZN(n6103) );
  XNOR2_X1 U4442 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4101) );
  NAND2_X1 U4443 ( .A1(n6175), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4099) );
  XNOR2_X1 U4444 ( .A(n4101), .B(n4099), .ZN(n4600) );
  INV_X1 U4445 ( .A(n4085), .ZN(n4124) );
  NAND2_X1 U4446 ( .A1(n4137), .A2(n3627), .ZN(n4083) );
  OAI211_X1 U4447 ( .C1(n4600), .C2(n4124), .A(n4083), .B(n4922), .ZN(n4096)
         );
  NAND2_X1 U4448 ( .A1(n4600), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4086) );
  NAND2_X1 U4449 ( .A1(n4127), .A2(n4086), .ZN(n4095) );
  OAI21_X1 U4450 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6175), .A(n4099), 
        .ZN(n4087) );
  INV_X1 U4451 ( .A(n4087), .ZN(n4088) );
  NAND2_X1 U4452 ( .A1(n4137), .A2(n4088), .ZN(n4093) );
  NAND2_X1 U4453 ( .A1(n4142), .A2(n4088), .ZN(n4090) );
  NAND2_X1 U4454 ( .A1(n4090), .A2(n4089), .ZN(n4092) );
  NAND2_X1 U4455 ( .A1(n6120), .A2(n5454), .ZN(n4091) );
  NAND2_X1 U4456 ( .A1(n4091), .A2(n4693), .ZN(n4114) );
  AOI22_X1 U4457 ( .A1(n4127), .A2(n4093), .B1(n4092), .B2(n4114), .ZN(n4094)
         );
  OAI21_X1 U4458 ( .B1(n4096), .B2(n4095), .A(n4094), .ZN(n4098) );
  NAND2_X1 U4459 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  NAND2_X1 U4460 ( .A1(n4098), .A2(n4097), .ZN(n4107) );
  MUX2_X1 U4461 ( .A(n7462), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4108) );
  INV_X1 U4462 ( .A(n4108), .ZN(n4104) );
  INV_X1 U4463 ( .A(n4099), .ZN(n4100) );
  NAND2_X1 U4464 ( .A1(n4101), .A2(n4100), .ZN(n4103) );
  NAND2_X1 U4465 ( .A1(n5381), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4102) );
  NAND2_X1 U4466 ( .A1(n4103), .A2(n4102), .ZN(n4109) );
  XNOR2_X1 U4467 ( .A(n4104), .B(n4109), .ZN(n4597) );
  NAND2_X1 U4468 ( .A1(n4137), .A2(n4597), .ZN(n4105) );
  OAI211_X1 U4469 ( .C1(n4597), .C2(n4124), .A(n4105), .B(n4114), .ZN(n4106)
         );
  NAND2_X1 U4470 ( .A1(n4107), .A2(n4106), .ZN(n4119) );
  NAND2_X1 U4471 ( .A1(n4109), .A2(n4108), .ZN(n4111) );
  NAND2_X1 U4472 ( .A1(n7462), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4110) );
  NAND2_X1 U4473 ( .A1(n4111), .A2(n4110), .ZN(n4122) );
  MUX2_X1 U4474 ( .A(n4112), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4121) );
  INV_X1 U4475 ( .A(n4121), .ZN(n4113) );
  XNOR2_X1 U4476 ( .A(n4122), .B(n4113), .ZN(n4598) );
  INV_X1 U4477 ( .A(n4114), .ZN(n4115) );
  NAND3_X1 U4478 ( .A1(n4137), .A2(n4115), .A3(n4597), .ZN(n4116) );
  OAI21_X1 U4479 ( .B1(n4127), .B2(n4598), .A(n4116), .ZN(n4117) );
  INV_X1 U4480 ( .A(n4117), .ZN(n4118) );
  NAND2_X1 U4481 ( .A1(n4119), .A2(n4118), .ZN(n4126) );
  NOR2_X1 U4482 ( .A1(n3923), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4120)
         );
  AOI21_X1 U4483 ( .B1(n4122), .B2(n4121), .A(n4120), .ZN(n4133) );
  INV_X1 U4484 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5171) );
  AND2_X1 U4485 ( .A1(n5171), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4131)
         );
  NAND2_X1 U4486 ( .A1(n4133), .A2(n4131), .ZN(n4596) );
  NAND2_X1 U4487 ( .A1(n4596), .A2(n4598), .ZN(n4123) );
  NAND2_X1 U4488 ( .A1(n4124), .A2(n4123), .ZN(n4125) );
  NAND2_X1 U4489 ( .A1(n4126), .A2(n4125), .ZN(n4130) );
  INV_X1 U4490 ( .A(n4596), .ZN(n4128) );
  AOI22_X1 U4491 ( .A1(n4134), .A2(n4128), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7161), .ZN(n4129) );
  NAND2_X1 U4492 ( .A1(n4130), .A2(n4129), .ZN(n4136) );
  INV_X1 U4493 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U4494 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6991), .ZN(n4132) );
  AOI21_X1 U4495 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4602) );
  NAND2_X1 U4496 ( .A1(n4134), .A2(n4602), .ZN(n4135) );
  NAND2_X1 U4497 ( .A1(n4136), .A2(n4135), .ZN(n4139) );
  NAND2_X1 U4498 ( .A1(n4137), .A2(n4602), .ZN(n4138) );
  NAND2_X1 U4499 ( .A1(n4140), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7499) );
  NAND2_X1 U4500 ( .A1(n6962), .A2(n4922), .ZN(n4653) );
  AND2_X1 U4501 ( .A1(n4653), .A2(n4668), .ZN(n4141) );
  NOR2_X1 U4502 ( .A1(n4647), .A2(n4141), .ZN(n4632) );
  INV_X1 U4503 ( .A(n4142), .ZN(n4143) );
  NAND2_X1 U4504 ( .A1(n4632), .A2(n4143), .ZN(n7447) );
  OR2_X1 U4505 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5997) );
  NAND2_X1 U4506 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U4507 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4144) );
  INV_X1 U4508 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4145) );
  INV_X1 U4509 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5863) );
  INV_X1 U4510 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4530) );
  INV_X1 U4511 ( .A(n4515), .ZN(n4146) );
  INV_X1 U4512 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U4513 ( .A1(n4446), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4450)
         );
  INV_X1 U4514 ( .A(n4450), .ZN(n4147) );
  INV_X1 U4515 ( .A(n4408), .ZN(n4148) );
  INV_X1 U4516 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6417) );
  INV_X1 U4517 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6239) );
  INV_X1 U4518 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U4519 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6000)
         );
  INV_X1 U4520 ( .A(n4149), .ZN(n4150) );
  INV_X1 U4521 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U4522 ( .A1(n4150), .A2(n6218), .ZN(n4151) );
  NAND2_X1 U4523 ( .A1(n6000), .A2(n4151), .ZN(n6217) );
  AOI22_X1 U4524 ( .A1(n3676), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U4525 ( .A1(n4226), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U4526 ( .A1(n5980), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U4527 ( .A1(n3675), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U4528 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4161)
         );
  AOI22_X1 U4529 ( .A1(n3635), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U4530 ( .A1(n5971), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U4531 ( .A1(n3684), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U4532 ( .A1(n3629), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4156) );
  NAND4_X1 U4533 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4160)
         );
  NOR2_X1 U4534 ( .A1(n4161), .A2(n4160), .ZN(n4376) );
  AOI22_X1 U4535 ( .A1(n5980), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4536 ( .A1(n3675), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4537 ( .A1(n3900), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4538 ( .A1(n5975), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U4539 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4171)
         );
  AOI22_X1 U4540 ( .A1(n5971), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4541 ( .A1(n5981), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4542 ( .A1(n3635), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U4543 ( .A1(n5972), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U4544 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4170)
         );
  NOR2_X1 U4545 ( .A1(n4171), .A2(n4170), .ZN(n4394) );
  AOI22_X1 U4546 ( .A1(n5980), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4547 ( .A1(n5971), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4548 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4226), .B1(n3629), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U4549 ( .A1(n5973), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4172) );
  NAND4_X1 U4550 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4181)
         );
  AOI22_X1 U4551 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3900), .B1(n5972), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U4552 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n5981), .B1(n5982), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U4553 ( .A1(n3635), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U4554 ( .A1(n5975), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4176) );
  NAND4_X1 U4555 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4180)
         );
  NOR2_X1 U4556 ( .A1(n4181), .A2(n4180), .ZN(n4409) );
  AOI22_X1 U4557 ( .A1(n3635), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U4558 ( .A1(n5972), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U4559 ( .A1(n3900), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U4560 ( .A1(n3629), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4182) );
  NAND4_X1 U4561 ( .A1(n4185), .A2(n4184), .A3(n4183), .A4(n4182), .ZN(n4191)
         );
  AOI22_X1 U4562 ( .A1(n5971), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4563 ( .A1(n5981), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U4564 ( .A1(n5980), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4565 ( .A1(n4557), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U4566 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4190)
         );
  NOR2_X1 U4567 ( .A1(n4191), .A2(n4190), .ZN(n4410) );
  OR2_X1 U4568 ( .A1(n4409), .A2(n4410), .ZN(n4400) );
  AOI22_X1 U4569 ( .A1(n4557), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U4570 ( .A1(n3630), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U4571 ( .A1(n3900), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U4572 ( .A1(n5980), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4192) );
  NAND4_X1 U4573 ( .A1(n4195), .A2(n4194), .A3(n4193), .A4(n4192), .ZN(n4201)
         );
  AOI22_X1 U4574 ( .A1(n3635), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4575 ( .A1(n5975), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U4576 ( .A1(n5981), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4197) );
  INV_X1 U4577 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U4578 ( .A1(n5971), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4196) );
  NAND4_X1 U4579 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(n4200)
         );
  NOR2_X1 U4580 ( .A1(n4201), .A2(n4200), .ZN(n4399) );
  OR2_X1 U4581 ( .A1(n4400), .A2(n4399), .ZN(n4393) );
  NOR2_X1 U4582 ( .A1(n4394), .A2(n4393), .ZN(n4383) );
  AOI22_X1 U4583 ( .A1(n5971), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U4584 ( .A1(n5981), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U4585 ( .A1(n4226), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4586 ( .A1(n5975), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U4587 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4211)
         );
  AOI22_X1 U4588 ( .A1(n3635), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4589 ( .A1(n5980), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4590 ( .A1(n3900), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U4591 ( .A1(n5972), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4206) );
  NAND4_X1 U4592 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4210)
         );
  OR2_X1 U4593 ( .A1(n4211), .A2(n4210), .ZN(n4382) );
  NAND2_X1 U4594 ( .A1(n4383), .A2(n4382), .ZN(n4377) );
  NOR2_X1 U4595 ( .A1(n4376), .A2(n4377), .ZN(n4580) );
  AOI22_X1 U4596 ( .A1(n3635), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U4597 ( .A1(n5980), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U4598 ( .A1(n3684), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U4599 ( .A1(n5972), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4212) );
  NAND4_X1 U4600 ( .A1(n4215), .A2(n4214), .A3(n4213), .A4(n4212), .ZN(n4221)
         );
  AOI22_X1 U4601 ( .A1(n5971), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U4602 ( .A1(n5981), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U4603 ( .A1(n4226), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U4604 ( .A1(n5975), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4216) );
  NAND4_X1 U4605 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4220)
         );
  OR2_X1 U4606 ( .A1(n4221), .A2(n4220), .ZN(n4579) );
  NAND2_X1 U4607 ( .A1(n4580), .A2(n4579), .ZN(n5969) );
  AOI22_X1 U4608 ( .A1(n3635), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U4609 ( .A1(n5980), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4610 ( .A1(n5981), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U4611 ( .A1(n5982), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4222) );
  NAND4_X1 U4612 ( .A1(n4225), .A2(n4224), .A3(n4223), .A4(n4222), .ZN(n4232)
         );
  AOI22_X1 U4613 ( .A1(n5971), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U4614 ( .A1(n3629), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U4615 ( .A1(n4557), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U4616 ( .A1(n3684), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4227) );
  NAND4_X1 U4617 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4231)
         );
  NOR2_X1 U4618 ( .A1(n4232), .A2(n4231), .ZN(n5970) );
  XNOR2_X1 U4619 ( .A(n5969), .B(n5970), .ZN(n4235) );
  NAND2_X1 U4620 ( .A1(n6962), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5992) );
  INV_X1 U4621 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5995) );
  AOI21_X1 U4622 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5995), .A(n6001), 
        .ZN(n4234) );
  NOR2_X1 U4623 ( .A1(n6119), .A2(n5995), .ZN(n4533) );
  INV_X1 U4624 ( .A(n4533), .ZN(n4279) );
  NAND2_X1 U4625 ( .A1(n5999), .A2(EAX_REG_29__SCAN_IN), .ZN(n4233) );
  OAI211_X1 U4626 ( .C1(n4235), .C2(n5992), .A(n4234), .B(n4233), .ZN(n4236)
         );
  OAI21_X1 U4627 ( .B1(n5997), .B2(n6217), .A(n4236), .ZN(n4585) );
  NAND2_X1 U4628 ( .A1(n4656), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4568) );
  OR2_X1 U4629 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4237) );
  NAND2_X1 U4630 ( .A1(n4237), .A2(n4293), .ZN(n7305) );
  NAND2_X1 U4631 ( .A1(n5995), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4531) );
  INV_X1 U4632 ( .A(n4531), .ZN(n5968) );
  AOI22_X1 U4633 ( .A1(n7305), .A2(n6001), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4238) );
  OAI21_X1 U4634 ( .B1(n4279), .B2(n7007), .A(n4238), .ZN(n4239) );
  NOR2_X1 U4635 ( .A1(n4276), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4241)
         );
  OR2_X1 U4636 ( .A1(n4242), .A2(n4241), .ZN(n7292) );
  INV_X1 U4637 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4699) );
  INV_X1 U4638 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7286) );
  OAI22_X1 U4639 ( .A1(n4279), .A2(n4699), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7286), .ZN(n4243) );
  MUX2_X1 U4640 ( .A(n7292), .B(n4243), .S(n5997), .Z(n4244) );
  OAI21_X1 U4641 ( .B1(n4890), .B2(n4568), .A(n4531), .ZN(n4260) );
  NAND2_X1 U4642 ( .A1(n6118), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4269) );
  INV_X1 U4643 ( .A(n5997), .ZN(n6001) );
  OAI21_X1 U4644 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4246), .ZN(n7247) );
  AOI22_X1 U4645 ( .A1(n5968), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6001), 
        .B2(n7247), .ZN(n4248) );
  NAND2_X1 U4646 ( .A1(n5999), .A2(EAX_REG_2__SCAN_IN), .ZN(n4247) );
  OAI211_X1 U4647 ( .C1(n4269), .C2(n6074), .A(n4248), .B(n4247), .ZN(n4259)
         );
  NAND2_X1 U4648 ( .A1(n4260), .A2(n4259), .ZN(n4258) );
  NAND2_X1 U4649 ( .A1(n5187), .A2(n4546), .ZN(n4254) );
  AOI22_X1 U4650 ( .A1(n5999), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5995), .ZN(n4252) );
  INV_X1 U4651 ( .A(n4269), .ZN(n4250) );
  NAND2_X1 U4652 ( .A1(n4250), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4251) );
  AND2_X1 U4653 ( .A1(n4252), .A2(n4251), .ZN(n4253) );
  NAND2_X1 U4654 ( .A1(n4254), .A2(n4253), .ZN(n4767) );
  OAI21_X1 U4655 ( .B1(n6180), .B2(n4915), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4255) );
  NAND2_X1 U4656 ( .A1(n4255), .A2(n4279), .ZN(n4752) );
  OR2_X1 U4657 ( .A1(n6184), .A2(n4568), .ZN(n4257) );
  AOI22_X1 U4658 ( .A1(n5999), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n5995), .ZN(n4256) );
  OAI211_X1 U4659 ( .C1(n4269), .C2(n4787), .A(n4257), .B(n4256), .ZN(n4751)
         );
  MUX2_X1 U4660 ( .A(n6001), .B(n4752), .S(n4751), .Z(n4766) );
  NAND2_X1 U4661 ( .A1(n4767), .A2(n4766), .ZN(n4845) );
  NAND2_X1 U4662 ( .A1(n4258), .A2(n4845), .ZN(n4261) );
  OR2_X1 U4663 ( .A1(n4260), .A2(n4259), .ZN(n4843) );
  NAND2_X1 U4664 ( .A1(n4261), .A2(n4843), .ZN(n4886) );
  OAI21_X1 U4665 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4262), .A(n4274), 
        .ZN(n5590) );
  AOI22_X1 U4666 ( .A1(n6001), .A2(n5590), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U4667 ( .A1(n5999), .A2(EAX_REG_3__SCAN_IN), .ZN(n4263) );
  OAI211_X1 U4668 ( .C1(n4269), .C2(n3923), .A(n4264), .B(n4263), .ZN(n4265)
         );
  NOR2_X2 U4669 ( .A1(n4886), .A2(n4887), .ZN(n5019) );
  NAND2_X1 U4670 ( .A1(n4266), .A2(n4546), .ZN(n4273) );
  NAND2_X1 U4671 ( .A1(n5995), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4268)
         );
  NAND2_X1 U4672 ( .A1(n4533), .A2(EAX_REG_4__SCAN_IN), .ZN(n4267) );
  OAI211_X1 U4673 ( .C1(n4269), .C2(n5171), .A(n4268), .B(n4267), .ZN(n4271)
         );
  XNOR2_X1 U4674 ( .A(n4274), .B(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n7263) );
  NOR2_X1 U4675 ( .A1(n7263), .A2(n5997), .ZN(n4270) );
  AOI21_X1 U4676 ( .B1(n4271), .B2(n5997), .A(n4270), .ZN(n4272) );
  NAND2_X1 U4677 ( .A1(n4273), .A2(n4272), .ZN(n5018) );
  NAND2_X1 U4678 ( .A1(n5019), .A2(n5018), .ZN(n5022) );
  INV_X1 U4679 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4697) );
  INV_X1 U4680 ( .A(n4274), .ZN(n4275) );
  AOI21_X1 U4681 ( .B1(n4275), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4277) );
  OR2_X1 U4682 ( .A1(n4277), .A2(n4276), .ZN(n7284) );
  AOI22_X1 U4683 ( .A1(n7284), .A2(n6001), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4278) );
  OAI21_X1 U4684 ( .B1(n4279), .B2(n4697), .A(n4278), .ZN(n4280) );
  OR2_X2 U4685 ( .A1(n5022), .A2(n5021), .ZN(n5283) );
  AOI22_X1 U4686 ( .A1(n3635), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U4687 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n5971), .B1(n4226), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U4688 ( .A1(n5980), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U4689 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n5981), .B1(n5974), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4283) );
  NAND4_X1 U4690 ( .A1(n4286), .A2(n4285), .A3(n4284), .A4(n4283), .ZN(n4292)
         );
  AOI22_X1 U4691 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5975), .B1(n3629), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4290) );
  AOI22_X1 U4692 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4557), .B1(n5982), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4289) );
  AOI22_X1 U4693 ( .A1(n3900), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4288) );
  AOI22_X1 U4694 ( .A1(n5972), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4287) );
  NAND4_X1 U4695 ( .A1(n4290), .A2(n4289), .A3(n4288), .A4(n4287), .ZN(n4291)
         );
  NOR2_X1 U4696 ( .A1(n4292), .A2(n4291), .ZN(n4297) );
  INV_X1 U4697 ( .A(n4293), .ZN(n4294) );
  XNOR2_X1 U4698 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4294), .ZN(n5612) );
  AOI22_X1 U4699 ( .A1(n6001), .A2(n5612), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U4700 ( .A1(n4533), .A2(EAX_REG_8__SCAN_IN), .ZN(n4295) );
  OAI211_X1 U4701 ( .C1(n4568), .C2(n4297), .A(n4296), .B(n4295), .ZN(n5318)
         );
  XOR2_X1 U4702 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4298), .Z(n5693) );
  AOI22_X1 U4703 ( .A1(n3900), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4302) );
  AOI22_X1 U4704 ( .A1(n3629), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U4705 ( .A1(n4226), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U4706 ( .A1(n4419), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4299) );
  NAND4_X1 U4707 ( .A1(n4302), .A2(n4301), .A3(n4300), .A4(n4299), .ZN(n4308)
         );
  AOI22_X1 U4708 ( .A1(n3635), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U4709 ( .A1(n5980), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U4710 ( .A1(n4557), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U4711 ( .A1(n5981), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4303) );
  NAND4_X1 U4712 ( .A1(n4306), .A2(n4305), .A3(n4304), .A4(n4303), .ZN(n4307)
         );
  OR2_X1 U4713 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  AOI22_X1 U4714 ( .A1(n4546), .A2(n4309), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4311) );
  NAND2_X1 U4715 ( .A1(n4533), .A2(EAX_REG_9__SCAN_IN), .ZN(n4310) );
  OAI211_X1 U4716 ( .C1(n5693), .C2(n5997), .A(n4311), .B(n4310), .ZN(n4312)
         );
  INV_X1 U4717 ( .A(n4312), .ZN(n5579) );
  XNOR2_X1 U4718 ( .A(n4314), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5751)
         );
  NAND2_X1 U4719 ( .A1(n5751), .A2(n6001), .ZN(n4329) );
  AOI22_X1 U4720 ( .A1(n4419), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U4721 ( .A1(n5981), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U4722 ( .A1(n3635), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U4723 ( .A1(n3900), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4315) );
  NAND4_X1 U4724 ( .A1(n4318), .A2(n4317), .A3(n4316), .A4(n4315), .ZN(n4324)
         );
  AOI22_X1 U4725 ( .A1(n5980), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4726 ( .A1(n4226), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4727 ( .A1(n5972), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U4728 ( .A1(n5975), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4319) );
  NAND4_X1 U4729 ( .A1(n4322), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(n4323)
         );
  OAI21_X1 U4730 ( .B1(n4324), .B2(n4323), .A(n4546), .ZN(n4327) );
  NAND2_X1 U4731 ( .A1(n4533), .A2(EAX_REG_10__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U4732 ( .A1(n5968), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4325)
         );
  AND3_X1 U4733 ( .A1(n4327), .A2(n4326), .A3(n4325), .ZN(n4328) );
  AND2_X1 U4734 ( .A1(n4329), .A2(n4328), .ZN(n5700) );
  NOR2_X2 U4735 ( .A1(n5699), .A2(n5700), .ZN(n5720) );
  XOR2_X1 U4736 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4330), .Z(n7312) );
  AOI22_X1 U4737 ( .A1(n3635), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4738 ( .A1(n3676), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U4739 ( .A1(n4419), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U4740 ( .A1(n3900), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4331) );
  NAND4_X1 U4741 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(n4340)
         );
  AOI22_X1 U4742 ( .A1(n4557), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4743 ( .A1(n5980), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U4744 ( .A1(n5975), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4745 ( .A1(n5972), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4335) );
  NAND4_X1 U4746 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(n4339)
         );
  OR2_X1 U4747 ( .A1(n4340), .A2(n4339), .ZN(n4341) );
  AOI22_X1 U4748 ( .A1(n4546), .A2(n4341), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U4749 ( .A1(n5999), .A2(EAX_REG_11__SCAN_IN), .ZN(n4342) );
  OAI211_X1 U4750 ( .C1(n7312), .C2(n5997), .A(n4343), .B(n4342), .ZN(n5719)
         );
  AND2_X2 U4751 ( .A1(n5720), .A2(n5719), .ZN(n5725) );
  AOI22_X1 U4752 ( .A1(n5971), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U4753 ( .A1(n3901), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4754 ( .A1(n3635), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U4755 ( .A1(n3684), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4344) );
  NAND4_X1 U4756 ( .A1(n4347), .A2(n4346), .A3(n4345), .A4(n4344), .ZN(n4353)
         );
  AOI22_X1 U4757 ( .A1(n5980), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4351) );
  AOI22_X1 U4758 ( .A1(n3629), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4759 ( .A1(n5972), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4760 ( .A1(n3676), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4348) );
  NAND4_X1 U4761 ( .A1(n4351), .A2(n4350), .A3(n4349), .A4(n4348), .ZN(n4352)
         );
  NOR2_X1 U4762 ( .A1(n4353), .A2(n4352), .ZN(n4357) );
  XNOR2_X1 U4763 ( .A(n4354), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5876)
         );
  NAND2_X1 U4764 ( .A1(n5876), .A2(n6001), .ZN(n4356) );
  AOI22_X1 U4765 ( .A1(n5999), .A2(EAX_REG_12__SCAN_IN), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4355) );
  OAI211_X1 U4766 ( .C1(n4357), .C2(n4568), .A(n4356), .B(n4355), .ZN(n5724)
         );
  AOI22_X1 U4767 ( .A1(n3676), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U4768 ( .A1(n3807), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U4769 ( .A1(n5980), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U4770 ( .A1(n3675), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4358) );
  NAND4_X1 U4771 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(n4367)
         );
  AOI22_X1 U4772 ( .A1(n3635), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4773 ( .A1(n5971), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4774 ( .A1(n3684), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U4775 ( .A1(n3629), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4362) );
  NAND4_X1 U4776 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4366)
         );
  OR2_X1 U4777 ( .A1(n4367), .A2(n4366), .ZN(n4368) );
  NAND2_X1 U4778 ( .A1(n4546), .A2(n4368), .ZN(n4371) );
  XNOR2_X1 U4779 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4369), .ZN(n7322)
         );
  OAI22_X1 U4780 ( .A1(n5997), .A2(n7322), .B1(n4531), .B2(n5863), .ZN(n4370)
         );
  AOI21_X1 U4781 ( .B1(n5999), .B2(EAX_REG_13__SCAN_IN), .A(n4370), .ZN(n5859)
         );
  OR2_X2 U4782 ( .A1(n5860), .A2(n5859), .ZN(n4373) );
  NAND2_X4 U4783 ( .A1(n4373), .A2(n4372), .ZN(n6356) );
  NAND2_X1 U4784 ( .A1(n4374), .A2(n6239), .ZN(n4375) );
  NAND2_X1 U4785 ( .A1(n4577), .A2(n4375), .ZN(n6410) );
  XNOR2_X1 U4786 ( .A(n4377), .B(n4376), .ZN(n4380) );
  AOI21_X1 U4787 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5995), .A(n6001), 
        .ZN(n4379) );
  NAND2_X1 U4788 ( .A1(n5999), .A2(EAX_REG_27__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U4789 ( .C1(n4380), .C2(n5992), .A(n4379), .B(n4378), .ZN(n4381)
         );
  OAI21_X1 U4790 ( .B1(n5997), .B2(n6410), .A(n4381), .ZN(n6234) );
  INV_X1 U4791 ( .A(n6234), .ZN(n4575) );
  XNOR2_X1 U4792 ( .A(n4392), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6421)
         );
  AOI21_X1 U4793 ( .B1(n6417), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4386) );
  XNOR2_X1 U4794 ( .A(n4383), .B(n4382), .ZN(n4384) );
  NOR2_X1 U4795 ( .A1(n4384), .A2(n5992), .ZN(n4385) );
  AOI211_X1 U4796 ( .C1(n5999), .C2(EAX_REG_26__SCAN_IN), .A(n4386), .B(n4385), 
        .ZN(n4387) );
  AOI21_X1 U4797 ( .B1(n6001), .B2(n6421), .A(n4387), .ZN(n6248) );
  INV_X1 U4798 ( .A(n4388), .ZN(n4390) );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U4800 ( .A1(n4390), .A2(n4389), .ZN(n4391) );
  NAND2_X1 U4801 ( .A1(n4392), .A2(n4391), .ZN(n6426) );
  XNOR2_X1 U4802 ( .A(n4394), .B(n4393), .ZN(n4397) );
  AOI21_X1 U4803 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5995), .A(n6001), 
        .ZN(n4396) );
  NAND2_X1 U4804 ( .A1(n5999), .A2(EAX_REG_25__SCAN_IN), .ZN(n4395) );
  OAI211_X1 U4805 ( .C1(n4397), .C2(n5992), .A(n4396), .B(n4395), .ZN(n4398)
         );
  OAI21_X1 U4806 ( .B1(n5997), .B2(n6426), .A(n4398), .ZN(n6264) );
  INV_X1 U4807 ( .A(n6264), .ZN(n4574) );
  XNOR2_X1 U4808 ( .A(n4400), .B(n4399), .ZN(n4403) );
  AOI22_X1 U4809 ( .A1(n5999), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5968), .ZN(n4402) );
  XOR2_X1 U4810 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .B(n4408), .Z(n6279) );
  NAND2_X1 U4811 ( .A1(n6279), .A2(n6001), .ZN(n4401) );
  OAI211_X1 U4812 ( .C1(n4403), .C2(n5992), .A(n4402), .B(n4401), .ZN(n6107)
         );
  INV_X1 U4813 ( .A(n4404), .ZN(n4406) );
  INV_X1 U4814 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U4815 ( .A1(n4406), .A2(n4405), .ZN(n4407) );
  NAND2_X1 U4816 ( .A1(n4408), .A2(n4407), .ZN(n6436) );
  XNOR2_X1 U4817 ( .A(n4410), .B(n4409), .ZN(n4413) );
  AOI21_X1 U4818 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5995), .A(n6001), 
        .ZN(n4412) );
  NAND2_X1 U4819 ( .A1(n5999), .A2(EAX_REG_23__SCAN_IN), .ZN(n4411) );
  OAI211_X1 U4820 ( .C1(n4413), .C2(n5992), .A(n4412), .B(n4411), .ZN(n4414)
         );
  OAI21_X1 U4821 ( .B1(n5997), .B2(n6436), .A(n4414), .ZN(n6287) );
  AOI22_X1 U4822 ( .A1(n3635), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U4823 ( .A1(n3676), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U4824 ( .A1(n4557), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U4825 ( .A1(n5972), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4415) );
  NAND4_X1 U4826 ( .A1(n4418), .A2(n4417), .A3(n4416), .A4(n4415), .ZN(n4425)
         );
  AOI22_X1 U4827 ( .A1(n4419), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4423) );
  AOI22_X1 U4828 ( .A1(n5980), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4422) );
  AOI22_X1 U4829 ( .A1(n3900), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U4830 ( .A1(n3629), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4420) );
  NAND4_X1 U4831 ( .A1(n4423), .A2(n4422), .A3(n4421), .A4(n4420), .ZN(n4424)
         );
  NOR2_X1 U4832 ( .A1(n4425), .A2(n4424), .ZN(n4429) );
  NAND2_X1 U4833 ( .A1(n5995), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4426)
         );
  NAND2_X1 U4834 ( .A1(n5997), .A2(n4426), .ZN(n4427) );
  AOI21_X1 U4835 ( .B1(n5999), .B2(EAX_REG_22__SCAN_IN), .A(n4427), .ZN(n4428)
         );
  OAI21_X1 U4836 ( .B1(n5992), .B2(n4429), .A(n4428), .ZN(n4431) );
  XNOR2_X1 U4837 ( .A(n4450), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n7427)
         );
  NAND2_X1 U4838 ( .A1(n7427), .A2(n6001), .ZN(n4430) );
  NAND2_X1 U4839 ( .A1(n4431), .A2(n4430), .ZN(n6322) );
  NOR2_X1 U4840 ( .A1(n6287), .A2(n6322), .ZN(n6105) );
  AND2_X1 U4841 ( .A1(n6107), .A2(n6105), .ZN(n4573) );
  AOI22_X1 U4842 ( .A1(n3635), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U4843 ( .A1(n3676), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U4844 ( .A1(n3629), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U4845 ( .A1(n3684), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4432) );
  NAND4_X1 U4846 ( .A1(n4435), .A2(n4434), .A3(n4433), .A4(n4432), .ZN(n4441)
         );
  AOI22_X1 U4847 ( .A1(n5971), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U4848 ( .A1(n5980), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U4849 ( .A1(n5982), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U4850 ( .A1(n3675), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4436) );
  NAND4_X1 U4851 ( .A1(n4439), .A2(n4438), .A3(n4437), .A4(n4436), .ZN(n4440)
         );
  NOR2_X1 U4852 ( .A1(n4441), .A2(n4440), .ZN(n4445) );
  INV_X1 U4853 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7502) );
  OAI21_X1 U4854 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n7502), .A(n5995), 
        .ZN(n4442) );
  INV_X1 U4855 ( .A(n4442), .ZN(n4443) );
  AOI21_X1 U4856 ( .B1(n5999), .B2(EAX_REG_21__SCAN_IN), .A(n4443), .ZN(n4444)
         );
  OAI21_X1 U4857 ( .B1(n5992), .B2(n4445), .A(n4444), .ZN(n4452) );
  INV_X1 U4858 ( .A(n4446), .ZN(n4448) );
  INV_X1 U4859 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U4860 ( .A1(n4448), .A2(n4447), .ZN(n4449) );
  NAND2_X1 U4861 ( .A1(n4450), .A2(n4449), .ZN(n7413) );
  OR2_X1 U4862 ( .A1(n7413), .A2(n5997), .ZN(n4451) );
  AND2_X1 U4863 ( .A1(n4452), .A2(n4451), .ZN(n6153) );
  AOI22_X1 U4864 ( .A1(n5980), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3684), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4456) );
  AOI22_X1 U4865 ( .A1(n5971), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U4866 ( .A1(n3676), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U4867 ( .A1(n3629), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4453) );
  NAND4_X1 U4868 ( .A1(n4456), .A2(n4455), .A3(n4454), .A4(n4453), .ZN(n4462)
         );
  AOI22_X1 U4869 ( .A1(n3635), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4460) );
  AOI22_X1 U4870 ( .A1(n5973), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4459) );
  AOI22_X1 U4871 ( .A1(n4226), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U4872 ( .A1(n5972), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4457) );
  NAND4_X1 U4873 ( .A1(n4460), .A2(n4459), .A3(n4458), .A4(n4457), .ZN(n4461)
         );
  NOR2_X1 U4874 ( .A1(n4462), .A2(n4461), .ZN(n4465) );
  OAI21_X1 U4875 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6450), .A(n5997), .ZN(
        n4463) );
  AOI21_X1 U4876 ( .B1(n5999), .B2(EAX_REG_20__SCAN_IN), .A(n4463), .ZN(n4464)
         );
  OAI21_X1 U4877 ( .B1(n5992), .B2(n4465), .A(n4464), .ZN(n4467) );
  XNOR2_X1 U4878 ( .A(n4482), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7399)
         );
  NAND2_X1 U4879 ( .A1(n7399), .A2(n6001), .ZN(n4466) );
  AND2_X1 U4880 ( .A1(n4467), .A2(n4466), .ZN(n6117) );
  AOI22_X1 U4881 ( .A1(n3635), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U4882 ( .A1(n5971), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5975), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U4883 ( .A1(n4557), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4469) );
  AOI22_X1 U4884 ( .A1(n5973), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4468) );
  NAND4_X1 U4885 ( .A1(n4471), .A2(n4470), .A3(n4469), .A4(n4468), .ZN(n4477)
         );
  AOI22_X1 U4886 ( .A1(n5980), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4475) );
  AOI22_X1 U4887 ( .A1(n3629), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U4888 ( .A1(n4226), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U4889 ( .A1(n5981), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4472) );
  NAND4_X1 U4890 ( .A1(n4475), .A2(n4474), .A3(n4473), .A4(n4472), .ZN(n4476)
         );
  NOR2_X1 U4891 ( .A1(n4477), .A2(n4476), .ZN(n4481) );
  NAND2_X1 U4892 ( .A1(n5995), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4478)
         );
  NAND2_X1 U4893 ( .A1(n5997), .A2(n4478), .ZN(n4479) );
  AOI21_X1 U4894 ( .B1(n4533), .B2(EAX_REG_19__SCAN_IN), .A(n4479), .ZN(n4480)
         );
  OAI21_X1 U4895 ( .B1(n5992), .B2(n4481), .A(n4480), .ZN(n4485) );
  OAI21_X1 U4896 ( .B1(n4483), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n4482), 
        .ZN(n7389) );
  OR2_X1 U4897 ( .A1(n7389), .A2(n5997), .ZN(n4484) );
  NAND2_X1 U4898 ( .A1(n4485), .A2(n4484), .ZN(n6144) );
  INV_X1 U4899 ( .A(n6144), .ZN(n4572) );
  AOI22_X1 U4900 ( .A1(n5980), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U4901 ( .A1(n4226), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5981), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4488) );
  AOI22_X1 U4902 ( .A1(n4557), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U4903 ( .A1(n5975), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4486) );
  NAND4_X1 U4904 ( .A1(n4489), .A2(n4488), .A3(n4487), .A4(n4486), .ZN(n4495)
         );
  AOI22_X1 U4905 ( .A1(n3900), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U4906 ( .A1(n3629), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U4907 ( .A1(n3635), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U4908 ( .A1(n5971), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4490) );
  NAND4_X1 U4909 ( .A1(n4493), .A2(n4492), .A3(n4491), .A4(n4490), .ZN(n4494)
         );
  NOR2_X1 U4910 ( .A1(n4495), .A2(n4494), .ZN(n4498) );
  INV_X1 U4911 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6459) );
  AOI21_X1 U4912 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6459), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4496) );
  AOI21_X1 U4913 ( .B1(n4533), .B2(EAX_REG_18__SCAN_IN), .A(n4496), .ZN(n4497)
         );
  OAI21_X1 U4914 ( .B1(n5992), .B2(n4498), .A(n4497), .ZN(n4500) );
  XNOR2_X1 U4915 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4515), .ZN(n7375)
         );
  NAND2_X1 U4916 ( .A1(n7375), .A2(n6001), .ZN(n4499) );
  NAND2_X1 U4917 ( .A1(n4500), .A2(n4499), .ZN(n6333) );
  INV_X1 U4918 ( .A(n6333), .ZN(n4571) );
  AOI22_X1 U4919 ( .A1(n3635), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U4920 ( .A1(n5980), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U4921 ( .A1(n5971), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U4922 ( .A1(n3676), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4501) );
  NAND4_X1 U4923 ( .A1(n4504), .A2(n4503), .A3(n4502), .A4(n4501), .ZN(n4510)
         );
  AOI22_X1 U4924 ( .A1(n4226), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4508) );
  AOI22_X1 U4925 ( .A1(n5973), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U4926 ( .A1(n5975), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U4927 ( .A1(n5972), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4505) );
  NAND4_X1 U4928 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(n4509)
         );
  NOR2_X1 U4929 ( .A1(n4510), .A2(n4509), .ZN(n4514) );
  NAND2_X1 U4930 ( .A1(n5995), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4511)
         );
  NAND2_X1 U4931 ( .A1(n5997), .A2(n4511), .ZN(n4512) );
  AOI21_X1 U4932 ( .B1(n4533), .B2(EAX_REG_17__SCAN_IN), .A(n4512), .ZN(n4513)
         );
  OAI21_X1 U4933 ( .B1(n5992), .B2(n4514), .A(n4513), .ZN(n4518) );
  OAI21_X1 U4934 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4516), .A(n4515), 
        .ZN(n7362) );
  OR2_X1 U4935 ( .A1(n5997), .A2(n7362), .ZN(n4517) );
  AND2_X1 U4936 ( .A1(n4518), .A2(n4517), .ZN(n6341) );
  XNOR2_X1 U4937 ( .A(n4519), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n7352)
         );
  INV_X1 U4938 ( .A(n7352), .ZN(n6472) );
  AOI22_X1 U4939 ( .A1(n3630), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U4940 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4226), .B1(n5971), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U4941 ( .A1(n5981), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U4942 ( .A1(n4557), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4520) );
  NAND4_X1 U4943 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4529)
         );
  AOI22_X1 U4944 ( .A1(n3635), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5980), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U4945 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3629), .B1(n5972), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U4946 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5973), .B1(n3800), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U4947 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4524) );
  NAND4_X1 U4948 ( .A1(n4527), .A2(n4526), .A3(n4525), .A4(n4524), .ZN(n4528)
         );
  NOR2_X1 U4949 ( .A1(n4529), .A2(n4528), .ZN(n4535) );
  NOR2_X1 U4950 ( .A1(n4531), .A2(n4530), .ZN(n4532) );
  AOI21_X1 U4951 ( .B1(n4533), .B2(EAX_REG_16__SCAN_IN), .A(n4532), .ZN(n4534)
         );
  OAI21_X1 U4952 ( .B1(n5992), .B2(n4535), .A(n4534), .ZN(n4536) );
  AOI21_X1 U4953 ( .B1(n6472), .B2(n6001), .A(n4536), .ZN(n6348) );
  INV_X1 U4954 ( .A(n6348), .ZN(n4570) );
  XNOR2_X1 U4955 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4537), .ZN(n6481)
         );
  AOI22_X1 U4956 ( .A1(n3635), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U4957 ( .A1(n5971), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5981), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4540) );
  AOI22_X1 U4958 ( .A1(n3900), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U4959 ( .A1(n5980), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4538) );
  NAND4_X1 U4960 ( .A1(n4541), .A2(n4540), .A3(n4539), .A4(n4538), .ZN(n4548)
         );
  AOI22_X1 U4961 ( .A1(n4557), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U4962 ( .A1(n3629), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U4963 ( .A1(n5973), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U4964 ( .A1(n5975), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4542) );
  NAND4_X1 U4965 ( .A1(n4545), .A2(n4544), .A3(n4543), .A4(n4542), .ZN(n4547)
         );
  OAI21_X1 U4966 ( .B1(n4548), .B2(n4547), .A(n4546), .ZN(n4551) );
  NAND2_X1 U4967 ( .A1(n5999), .A2(EAX_REG_15__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U4968 ( .A1(n5968), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4549)
         );
  NAND3_X1 U4969 ( .A1(n4551), .A2(n4550), .A3(n4549), .ZN(n4552) );
  AOI21_X1 U4970 ( .B1(n6481), .B2(n6001), .A(n4552), .ZN(n6298) );
  INV_X1 U4971 ( .A(n6298), .ZN(n4569) );
  AOI22_X1 U4972 ( .A1(n5980), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U4973 ( .A1(n4226), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5981), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U4974 ( .A1(n5972), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3800), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U4975 ( .A1(n5971), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4553) );
  NAND4_X1 U4976 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(n4563)
         );
  AOI22_X1 U4977 ( .A1(n3900), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4557), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U4978 ( .A1(n3629), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5982), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U4979 ( .A1(n3635), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U4980 ( .A1(n5975), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4558) );
  NAND4_X1 U4981 ( .A1(n4561), .A2(n4560), .A3(n4559), .A4(n4558), .ZN(n4562)
         );
  NOR2_X1 U4982 ( .A1(n4563), .A2(n4562), .ZN(n4567) );
  XNOR2_X1 U4983 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4564), .ZN(n7336)
         );
  AOI22_X1 U4984 ( .A1(n6001), .A2(n7336), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U4985 ( .A1(n5999), .A2(EAX_REG_14__SCAN_IN), .ZN(n4565) );
  OAI211_X1 U4986 ( .C1(n4568), .C2(n4567), .A(n4566), .B(n4565), .ZN(n6355)
         );
  AND2_X1 U4987 ( .A1(n4569), .A2(n6355), .ZN(n6297) );
  AND2_X1 U4988 ( .A1(n4570), .A2(n6297), .ZN(n6340) );
  AND2_X1 U4989 ( .A1(n6341), .A2(n6340), .ZN(n6330) );
  AND2_X1 U4990 ( .A1(n4571), .A2(n6330), .ZN(n6143) );
  AND2_X1 U4991 ( .A1(n4572), .A2(n6143), .ZN(n6114) );
  AND2_X1 U4992 ( .A1(n6117), .A2(n6114), .ZN(n6115) );
  AND2_X1 U4993 ( .A1(n6153), .A2(n6115), .ZN(n6104) );
  AND2_X1 U4994 ( .A1(n4573), .A2(n6104), .ZN(n6106) );
  AND2_X1 U4995 ( .A1(n4574), .A2(n6106), .ZN(n6246) );
  AND2_X1 U4996 ( .A1(n6248), .A2(n6246), .ZN(n6233) );
  AND2_X1 U4997 ( .A1(n4575), .A2(n6233), .ZN(n4576) );
  INV_X1 U4998 ( .A(n4577), .ZN(n4578) );
  XOR2_X1 U4999 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n4578), .Z(n6227) );
  OAI21_X1 U5000 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6048), .A(n5997), .ZN(
        n4583) );
  XNOR2_X1 U5001 ( .A(n4580), .B(n4579), .ZN(n4581) );
  NOR2_X1 U5002 ( .A1(n4581), .A2(n5992), .ZN(n4582) );
  AOI211_X1 U5003 ( .C1(n5999), .C2(EAX_REG_28__SCAN_IN), .A(n4583), .B(n4582), 
        .ZN(n4584) );
  AOI21_X1 U5004 ( .B1(n6001), .B2(n6227), .A(n4584), .ZN(n6051) );
  AOI21_X1 U5005 ( .B1(n4585), .B2(n6050), .A(n6189), .ZN(n6309) );
  NOR2_X2 U5006 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5756) );
  NOR2_X1 U5007 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7487), .ZN(n5435) );
  NAND2_X1 U5008 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5435), .ZN(n7163) );
  INV_X1 U5009 ( .A(n7163), .ZN(n4586) );
  NAND2_X1 U5010 ( .A1(n5756), .A2(n4586), .ZN(n6489) );
  INV_X1 U5011 ( .A(n5756), .ZN(n5379) );
  NAND2_X1 U5012 ( .A1(n5379), .A2(n4587), .ZN(n7166) );
  NAND2_X1 U5013 ( .A1(n7166), .A2(n7161), .ZN(n4588) );
  NAND2_X1 U5014 ( .A1(n7433), .A2(n4588), .ZN(n7132) );
  NAND2_X1 U5015 ( .A1(n7161), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U5016 ( .A1(n7502), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5017 ( .A1(n4590), .A2(n4589), .ZN(n4760) );
  NAND2_X1 U5018 ( .A1(n7132), .A2(n4760), .ZN(n7152) );
  AND2_X1 U5019 ( .A1(n5756), .A2(n7487), .ZN(n5602) );
  INV_X1 U5020 ( .A(n7205), .ZN(n7213) );
  INV_X1 U5021 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7065) );
  NOR2_X1 U5022 ( .A1(n7213), .A2(n7065), .ZN(n6099) );
  AOI21_X1 U5023 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6099), 
        .ZN(n4591) );
  OAI21_X1 U5024 ( .B1(n7152), .B2(n6217), .A(n4591), .ZN(n4592) );
  AOI21_X1 U5025 ( .B1(n6309), .B2(n3628), .A(n4592), .ZN(n4593) );
  OAI21_X1 U5026 ( .B1(n6103), .B2(n7433), .A(n4593), .ZN(U2957) );
  NOR2_X1 U5027 ( .A1(n5454), .A2(n3627), .ZN(n5437) );
  INV_X1 U5028 ( .A(n5437), .ZN(n4606) );
  AND2_X1 U5029 ( .A1(n4595), .A2(n4594), .ZN(n6200) );
  AND3_X1 U5030 ( .A1(n4598), .A2(n4597), .A3(n4596), .ZN(n4599) );
  AND2_X1 U5031 ( .A1(n4600), .A2(n4599), .ZN(n4601) );
  OR2_X1 U5032 ( .A1(n4602), .A2(n4601), .ZN(n6199) );
  INV_X1 U5033 ( .A(n6199), .ZN(n4603) );
  NAND2_X1 U5034 ( .A1(n6200), .A2(n4603), .ZN(n4604) );
  AND2_X1 U5035 ( .A1(n6197), .A2(n4604), .ZN(n4605) );
  AOI21_X1 U5036 ( .B1(n6202), .B2(n4606), .A(n4605), .ZN(n6207) );
  INV_X1 U5037 ( .A(n6207), .ZN(n4607) );
  OAI21_X1 U5038 ( .B1(n4607), .B2(n7499), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4609) );
  NOR2_X1 U5039 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n7495) );
  NAND3_X1 U5040 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7495), .A3(n4732), .ZN(
        n4608) );
  NAND2_X1 U5041 ( .A1(n4609), .A2(n4608), .ZN(U2790) );
  NOR2_X1 U5042 ( .A1(n6199), .A2(n7499), .ZN(n4610) );
  NAND2_X1 U5043 ( .A1(n6200), .A2(n4610), .ZN(n4613) );
  INV_X1 U5044 ( .A(n4613), .ZN(n4612) );
  INV_X1 U5045 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7524) );
  INV_X1 U5046 ( .A(n5602), .ZN(n4611) );
  OAI211_X1 U5047 ( .C1(n4612), .C2(n7524), .A(n4691), .B(n4611), .ZN(U2788)
         );
  NAND2_X1 U5048 ( .A1(n4691), .A2(n4613), .ZN(n7165) );
  INV_X1 U5049 ( .A(n7165), .ZN(n4615) );
  AND2_X1 U5050 ( .A1(n4668), .A2(n3627), .ZN(n5442) );
  OR2_X1 U5051 ( .A1(n5442), .A2(n3634), .ZN(n6205) );
  OAI21_X1 U5052 ( .B1(n5602), .B2(READREQUEST_REG_SCAN_IN), .A(n4615), .ZN(
        n4614) );
  OAI21_X1 U5053 ( .B1(n4615), .B2(n6205), .A(n4614), .ZN(U3474) );
  OAI21_X1 U5054 ( .B1(n4616), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4794), 
        .ZN(n4763) );
  INV_X1 U5055 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U5056 ( .A1(n7509), .A2(n7158), .ZN(n7159) );
  INV_X1 U5057 ( .A(n7159), .ZN(n5453) );
  NOR2_X1 U5058 ( .A1(n3627), .A2(n5453), .ZN(n4617) );
  OR3_X1 U5059 ( .A1(n6202), .A2(READY_N), .A3(n4617), .ZN(n4748) );
  INV_X1 U5060 ( .A(n4736), .ZN(n4717) );
  INV_X1 U5061 ( .A(n6200), .ZN(n4622) );
  MUX2_X1 U5062 ( .A(n4693), .B(n4619), .S(n4781), .Z(n4620) );
  NAND2_X1 U5063 ( .A1(n4620), .A2(n5454), .ZN(n4650) );
  NAND2_X1 U5064 ( .A1(n4632), .A2(n4650), .ZN(n4621) );
  NAND2_X1 U5065 ( .A1(n4622), .A2(n4621), .ZN(n4744) );
  NAND2_X1 U5066 ( .A1(n3627), .A2(n7159), .ZN(n4623) );
  NOR2_X1 U5067 ( .A1(READY_N), .A2(n6199), .ZN(n4739) );
  NAND3_X1 U5068 ( .A1(n4623), .A2(n4739), .A3(n4899), .ZN(n4624) );
  AND2_X1 U5069 ( .A1(n4744), .A2(n4624), .ZN(n4626) );
  AND2_X1 U5070 ( .A1(n6962), .A2(n3627), .ZN(n4659) );
  NAND2_X1 U5071 ( .A1(n6202), .A2(n4659), .ZN(n4625) );
  OAI211_X1 U5072 ( .C1(n4748), .C2(n4717), .A(n4626), .B(n4625), .ZN(n4627)
         );
  INV_X1 U5073 ( .A(n7499), .ZN(n7473) );
  NAND2_X1 U5074 ( .A1(n4627), .A2(n7473), .ZN(n4630) );
  OAI21_X1 U5075 ( .B1(n6118), .B2(n4668), .A(n4755), .ZN(n4628) );
  OR2_X1 U5076 ( .A1(n4690), .A2(n4628), .ZN(n4629) );
  NAND2_X1 U5077 ( .A1(n4630), .A2(n4629), .ZN(n4663) );
  NAND2_X1 U5078 ( .A1(n4632), .A2(n5437), .ZN(n4738) );
  AND2_X1 U5079 ( .A1(n7447), .A2(n4738), .ZN(n6198) );
  NOR2_X1 U5080 ( .A1(n4633), .A2(n4753), .ZN(n4634) );
  AOI21_X1 U5081 ( .B1(n4736), .B2(n5924), .A(n4634), .ZN(n4635) );
  NAND3_X1 U5082 ( .A1(n7436), .A2(n6198), .A3(n4635), .ZN(n4636) );
  NAND2_X1 U5083 ( .A1(n4663), .A2(n4636), .ZN(n6584) );
  INV_X1 U5084 ( .A(n4926), .ZN(n4637) );
  NAND2_X1 U5085 ( .A1(n4637), .A2(n3632), .ZN(n4769) );
  INV_X1 U5086 ( .A(n5963), .ZN(n5952) );
  INV_X1 U5087 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7195) );
  INV_X1 U5088 ( .A(n4769), .ZN(n4770) );
  NAND2_X1 U5089 ( .A1(n4769), .A2(EBX_REG_0__SCAN_IN), .ZN(n4640) );
  INV_X1 U5090 ( .A(n4768), .ZN(n5024) );
  INV_X1 U5091 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5092 ( .A1(n4768), .A2(n4638), .ZN(n4639) );
  NAND2_X1 U5093 ( .A1(n4640), .A2(n4639), .ZN(n4774) );
  INV_X1 U5094 ( .A(n4774), .ZN(n4641) );
  AOI21_X1 U5095 ( .B1(n5952), .B2(n7195), .A(n4641), .ZN(n5459) );
  NAND2_X1 U5096 ( .A1(n4736), .A2(n3634), .ZN(n7477) );
  NAND3_X1 U5097 ( .A1(n4777), .A2(n4753), .A3(n6118), .ZN(n4642) );
  NAND2_X1 U5098 ( .A1(n7477), .A2(n4642), .ZN(n4643) );
  NAND2_X1 U5099 ( .A1(n7205), .A2(REIP_REG_0__SCAN_IN), .ZN(n4762) );
  INV_X1 U5100 ( .A(n4762), .ZN(n4645) );
  OR2_X1 U5101 ( .A1(n4663), .A2(n7205), .ZN(n7184) );
  AND2_X1 U5102 ( .A1(n6200), .A2(n3627), .ZN(n6964) );
  NAND2_X1 U5103 ( .A1(n4663), .A2(n6964), .ZN(n4865) );
  AOI21_X1 U5104 ( .B1(n7184), .B2(n4865), .A(n7195), .ZN(n4644) );
  AOI211_X1 U5105 ( .C1(n5459), .C2(n7238), .A(n4645), .B(n4644), .ZN(n4665)
         );
  NAND2_X1 U5106 ( .A1(n6118), .A2(n4668), .ZN(n4646) );
  AOI22_X1 U5107 ( .A1(n4654), .A2(n3627), .B1(n4646), .B2(n4899), .ZN(n4649)
         );
  NAND2_X1 U5108 ( .A1(n4647), .A2(n5963), .ZN(n4648) );
  AND3_X1 U5109 ( .A1(n4650), .A2(n4649), .A3(n4648), .ZN(n4651) );
  NAND2_X1 U5110 ( .A1(n4652), .A2(n4651), .ZN(n4719) );
  INV_X1 U5111 ( .A(n4653), .ZN(n4655) );
  NAND2_X1 U5112 ( .A1(n4655), .A2(n4654), .ZN(n5152) );
  NAND2_X1 U5113 ( .A1(n4777), .A2(n4656), .ZN(n4657) );
  OAI211_X1 U5114 ( .C1(n4715), .C2(n5454), .A(n5152), .B(n4657), .ZN(n4658)
         );
  NOR2_X1 U5115 ( .A1(n4719), .A2(n4658), .ZN(n4661) );
  NAND2_X1 U5116 ( .A1(n4661), .A2(n4659), .ZN(n6196) );
  INV_X1 U5117 ( .A(n6196), .ZN(n4660) );
  NAND2_X1 U5118 ( .A1(n4663), .A2(n4660), .ZN(n6036) );
  INV_X1 U5119 ( .A(n6036), .ZN(n7197) );
  INV_X1 U5120 ( .A(n4661), .ZN(n4662) );
  NAND2_X1 U5121 ( .A1(n4663), .A2(n4662), .ZN(n4863) );
  INV_X1 U5122 ( .A(n4863), .ZN(n4664) );
  OAI21_X1 U5123 ( .B1(n7197), .B2(n4664), .A(n7195), .ZN(n7183) );
  OAI211_X1 U5124 ( .C1(n4763), .C2(n6584), .A(n4665), .B(n7183), .ZN(U3018)
         );
  INV_X1 U5125 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4671) );
  INV_X1 U5126 ( .A(n7477), .ZN(n4666) );
  OAI21_X1 U5127 ( .B1(n6964), .B2(n4666), .A(n5453), .ZN(n4667) );
  OR2_X1 U5128 ( .A1(n7024), .A2(n4668), .ZN(n4808) );
  INV_X1 U5129 ( .A(n7024), .ZN(n4669) );
  AOI22_X1 U5130 ( .A1(n7167), .A2(UWORD_REG_7__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4670) );
  OAI21_X1 U5131 ( .B1(n4671), .B2(n4808), .A(n4670), .ZN(U2900) );
  INV_X1 U5132 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5133 ( .A1(n7167), .A2(UWORD_REG_5__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4672) );
  OAI21_X1 U5134 ( .B1(n4673), .B2(n4808), .A(n4672), .ZN(U2902) );
  INV_X1 U5135 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U5136 ( .A1(n7167), .A2(UWORD_REG_4__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4674) );
  OAI21_X1 U5137 ( .B1(n4675), .B2(n4808), .A(n4674), .ZN(U2903) );
  INV_X1 U5138 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4677) );
  AOI22_X1 U5139 ( .A1(n7167), .A2(UWORD_REG_9__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4676) );
  OAI21_X1 U5140 ( .B1(n4677), .B2(n4808), .A(n4676), .ZN(U2898) );
  INV_X1 U5141 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U5142 ( .A1(n7167), .A2(UWORD_REG_6__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4678) );
  OAI21_X1 U5143 ( .B1(n4679), .B2(n4808), .A(n4678), .ZN(U2901) );
  INV_X1 U5144 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5145 ( .A1(n7167), .A2(UWORD_REG_13__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4680) );
  OAI21_X1 U5146 ( .B1(n4681), .B2(n4808), .A(n4680), .ZN(U2894) );
  INV_X1 U5147 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5148 ( .A1(n7167), .A2(UWORD_REG_10__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4682) );
  OAI21_X1 U5149 ( .B1(n4683), .B2(n4808), .A(n4682), .ZN(U2897) );
  INV_X1 U5150 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U5151 ( .A1(n7167), .A2(UWORD_REG_11__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4684) );
  OAI21_X1 U5152 ( .B1(n4685), .B2(n4808), .A(n4684), .ZN(U2896) );
  INV_X1 U5153 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5154 ( .A1(n7167), .A2(UWORD_REG_12__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4686) );
  OAI21_X1 U5155 ( .B1(n4687), .B2(n4808), .A(n4686), .ZN(U2895) );
  INV_X1 U5156 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5157 ( .A1(n7167), .A2(UWORD_REG_8__SCAN_IN), .B1(n6992), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4688) );
  OAI21_X1 U5158 ( .B1(n4689), .B2(n4808), .A(n4688), .ZN(U2899) );
  OR2_X1 U5159 ( .A1(n4690), .A2(n7477), .ZN(n4813) );
  INV_X1 U5160 ( .A(n4691), .ZN(n4692) );
  INV_X1 U5161 ( .A(READY_N), .ZN(n7513) );
  NAND2_X1 U5162 ( .A1(n4692), .A2(n7513), .ZN(n4694) );
  OR2_X1 U5163 ( .A1(n4694), .A2(n4693), .ZN(n4842) );
  INV_X1 U5164 ( .A(n4842), .ZN(n4810) );
  NAND2_X1 U5165 ( .A1(n4810), .A2(DATAI_7_), .ZN(n4839) );
  NAND2_X1 U5166 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4811), .ZN(n4695) );
  OAI211_X1 U5167 ( .C1(n4813), .C2(n7007), .A(n4839), .B(n4695), .ZN(U2946)
         );
  NAND2_X1 U5168 ( .A1(n4810), .A2(DATAI_5_), .ZN(n4711) );
  NAND2_X1 U5169 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4811), .ZN(n4696) );
  OAI211_X1 U5170 ( .C1(n4813), .C2(n4697), .A(n4711), .B(n4696), .ZN(U2944)
         );
  NAND2_X1 U5171 ( .A1(n4810), .A2(DATAI_6_), .ZN(n4817) );
  NAND2_X1 U5172 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4811), .ZN(n4698) );
  OAI211_X1 U5173 ( .C1(n4813), .C2(n4699), .A(n4817), .B(n4698), .ZN(U2945)
         );
  NAND2_X1 U5174 ( .A1(n4810), .A2(DATAI_1_), .ZN(n4823) );
  INV_X2 U5175 ( .A(n4813), .ZN(n4840) );
  AOI22_X1 U5176 ( .A1(n4840), .A2(EAX_REG_17__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5177 ( .A1(n4823), .A2(n4700), .ZN(U2925) );
  NAND2_X1 U5178 ( .A1(n4810), .A2(DATAI_3_), .ZN(n4713) );
  AOI22_X1 U5179 ( .A1(n4840), .A2(EAX_REG_19__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5180 ( .A1(n4713), .A2(n4701), .ZN(U2927) );
  NAND2_X1 U5181 ( .A1(n4810), .A2(DATAI_12_), .ZN(n4827) );
  AOI22_X1 U5182 ( .A1(n4840), .A2(EAX_REG_12__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5183 ( .A1(n4827), .A2(n4702), .ZN(U2951) );
  NAND2_X1 U5184 ( .A1(n4810), .A2(DATAI_14_), .ZN(n4831) );
  AOI22_X1 U5185 ( .A1(n4840), .A2(EAX_REG_14__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U5186 ( .A1(n4831), .A2(n4703), .ZN(U2953) );
  NAND2_X1 U5187 ( .A1(n4810), .A2(DATAI_4_), .ZN(n4815) );
  AOI22_X1 U5188 ( .A1(n4840), .A2(EAX_REG_4__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U5189 ( .A1(n4815), .A2(n4704), .ZN(U2943) );
  NAND2_X1 U5190 ( .A1(n4810), .A2(DATAI_2_), .ZN(n4837) );
  AOI22_X1 U5191 ( .A1(n4840), .A2(EAX_REG_18__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5192 ( .A1(n4837), .A2(n4705), .ZN(U2926) );
  NAND2_X1 U5193 ( .A1(n4810), .A2(DATAI_0_), .ZN(n4833) );
  AOI22_X1 U5194 ( .A1(n4840), .A2(EAX_REG_16__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4706) );
  NAND2_X1 U5195 ( .A1(n4833), .A2(n4706), .ZN(U2924) );
  NAND2_X1 U5196 ( .A1(n4810), .A2(DATAI_10_), .ZN(n4835) );
  AOI22_X1 U5197 ( .A1(n4840), .A2(EAX_REG_10__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5198 ( .A1(n4835), .A2(n4707), .ZN(U2949) );
  NAND2_X1 U5199 ( .A1(n4810), .A2(DATAI_9_), .ZN(n4821) );
  AOI22_X1 U5200 ( .A1(n4840), .A2(EAX_REG_9__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U5201 ( .A1(n4821), .A2(n4708), .ZN(U2948) );
  NAND2_X1 U5202 ( .A1(n4810), .A2(DATAI_8_), .ZN(n4819) );
  AOI22_X1 U5203 ( .A1(n4840), .A2(EAX_REG_8__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5204 ( .A1(n4819), .A2(n4709), .ZN(U2947) );
  AOI22_X1 U5205 ( .A1(n4840), .A2(EAX_REG_21__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5206 ( .A1(n4711), .A2(n4710), .ZN(U2929) );
  AOI22_X1 U5207 ( .A1(n4840), .A2(EAX_REG_3__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5208 ( .A1(n4713), .A2(n4712), .ZN(U2942) );
  NAND2_X1 U5209 ( .A1(n4810), .A2(DATAI_11_), .ZN(n4825) );
  AOI22_X1 U5210 ( .A1(n4840), .A2(EAX_REG_11__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U5211 ( .A1(n4825), .A2(n4714), .ZN(U2950) );
  INV_X1 U5212 ( .A(n4777), .ZN(n4716) );
  NAND4_X1 U5213 ( .A1(n7436), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4718)
         );
  NOR2_X1 U5214 ( .A1(n4719), .A2(n4718), .ZN(n5149) );
  INV_X1 U5215 ( .A(n5149), .ZN(n6959) );
  NAND2_X1 U5216 ( .A1(n5032), .A2(n6959), .ZN(n4731) );
  AOI21_X1 U5217 ( .B1(n6960), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3923), 
        .ZN(n4720) );
  NOR2_X1 U5218 ( .A1(n3677), .A2(n4720), .ZN(n4733) );
  NAND2_X1 U5219 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5220 ( .A1(n6964), .A2(n4721), .ZN(n4725) );
  NAND2_X1 U5221 ( .A1(n6196), .A2(n4738), .ZN(n5155) );
  INV_X1 U5222 ( .A(n6960), .ZN(n6073) );
  NAND2_X1 U5223 ( .A1(n6073), .A2(n6074), .ZN(n4723) );
  INV_X1 U5224 ( .A(n4721), .ZN(n4722) );
  AOI22_X1 U5225 ( .A1(n5155), .A2(n4723), .B1(n6964), .B2(n4722), .ZN(n4724)
         );
  MUX2_X1 U5226 ( .A(n4725), .B(n4724), .S(n3923), .Z(n4728) );
  NAND2_X1 U5227 ( .A1(n6073), .A2(n4726), .ZN(n4727) );
  OAI211_X1 U5228 ( .C1(n4733), .C2(n5152), .A(n4728), .B(n4727), .ZN(n4729)
         );
  INV_X1 U5229 ( .A(n4729), .ZN(n4730) );
  NAND2_X1 U5230 ( .A1(n4731), .A2(n4730), .ZN(n5148) );
  INV_X1 U5231 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4732) );
  INV_X1 U5232 ( .A(n6069), .ZN(n7494) );
  INV_X1 U5233 ( .A(n4733), .ZN(n4734) );
  AOI22_X1 U5234 ( .A1(n5148), .A2(n7481), .B1(n7494), .B2(n4734), .ZN(n4750)
         );
  INV_X1 U5235 ( .A(n6197), .ZN(n4735) );
  OAI22_X1 U5236 ( .A1(n6964), .A2(n4736), .B1(n5453), .B2(n4735), .ZN(n4747)
         );
  INV_X1 U5237 ( .A(n6202), .ZN(n4737) );
  OR2_X1 U5238 ( .A1(n6202), .A2(n4738), .ZN(n4742) );
  INV_X1 U5239 ( .A(n7436), .ZN(n4740) );
  NAND2_X1 U5240 ( .A1(n4740), .A2(n4739), .ZN(n4741) );
  NAND2_X1 U5241 ( .A1(n4742), .A2(n4741), .ZN(n4779) );
  NAND2_X1 U5242 ( .A1(n5442), .A2(n4755), .ZN(n4743) );
  NAND2_X1 U5243 ( .A1(n4744), .A2(n4743), .ZN(n4745) );
  NOR2_X1 U5244 ( .A1(n4779), .A2(n4745), .ZN(n4746) );
  OAI211_X1 U5245 ( .C1(n4748), .C2(n4747), .A(n4757), .B(n4746), .ZN(n7456)
         );
  INV_X1 U5246 ( .A(n7456), .ZN(n5158) );
  NOR2_X1 U5247 ( .A1(n5995), .A2(n7487), .ZN(n7484) );
  NAND2_X1 U5248 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7484), .ZN(n7491) );
  INV_X1 U5249 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7443) );
  OAI22_X1 U5250 ( .A1(n5158), .A2(n7499), .B1(n7491), .B2(n7443), .ZN(n7437)
         );
  AOI21_X1 U5251 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7161), .A(n7437), .ZN(
        n6076) );
  NAND2_X1 U5252 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6076), .ZN(n4749) );
  OAI21_X1 U5253 ( .B1(n4750), .B2(n6076), .A(n4749), .ZN(U3456) );
  XNOR2_X1 U5254 ( .A(n4752), .B(n4751), .ZN(n5462) );
  INV_X1 U5255 ( .A(n6119), .ZN(n6185) );
  AND3_X1 U5256 ( .A1(n6185), .A2(n4753), .A3(n4915), .ZN(n4776) );
  NOR2_X1 U5257 ( .A1(n4926), .A2(n4922), .ZN(n4754) );
  NAND4_X1 U5258 ( .A1(n4776), .A2(n4755), .A3(n5924), .A4(n4754), .ZN(n4756)
         );
  NAND2_X1 U5259 ( .A1(n4757), .A2(n4756), .ZN(n4758) );
  NAND2_X1 U5260 ( .A1(n7118), .A2(n6185), .ZN(n7105) );
  INV_X1 U5261 ( .A(n7118), .ZN(n6338) );
  AOI22_X1 U5262 ( .A1(n7114), .A2(n5459), .B1(EBX_REG_0__SCAN_IN), .B2(n6338), 
        .ZN(n4759) );
  OAI21_X1 U5263 ( .B1(n5462), .B2(n6357), .A(n4759), .ZN(U2859) );
  OAI21_X1 U5264 ( .B1(n7147), .B2(n4760), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4761) );
  OAI211_X1 U5265 ( .C1(n4763), .C2(n7433), .A(n4762), .B(n4761), .ZN(n4764)
         );
  INV_X1 U5266 ( .A(n4764), .ZN(n4765) );
  OAI21_X1 U5267 ( .B1(n6489), .B2(n5462), .A(n4765), .ZN(U2986) );
  OAI21_X1 U5268 ( .B1(n4767), .B2(n4766), .A(n4845), .ZN(n5524) );
  MUX2_X1 U5269 ( .A(n5947), .B(n4769), .S(EBX_REG_1__SCAN_IN), .Z(n4773) );
  NAND2_X1 U5270 ( .A1(n4770), .A2(n4775), .ZN(n5939) );
  NAND2_X1 U5271 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4775), .ZN(n4771)
         );
  AND2_X1 U5272 ( .A1(n5939), .A2(n4771), .ZN(n4772) );
  XNOR2_X1 U5273 ( .A(n5522), .B(n5962), .ZN(n7179) );
  OAI222_X1 U5274 ( .A1(n5524), .A2(n6357), .B1(n7118), .B2(n5519), .C1(n7179), 
        .C2(n7105), .ZN(U2858) );
  AND2_X1 U5275 ( .A1(n4777), .A2(n4776), .ZN(n4778) );
  OAI21_X1 U5276 ( .B1(n4779), .B2(n4778), .A(n7473), .ZN(n4780) );
  NAND2_X1 U5277 ( .A1(n4781), .A2(n6119), .ZN(n4783) );
  INV_X1 U5278 ( .A(n4783), .ZN(n4782) );
  NAND2_X1 U5279 ( .A1(n6392), .A2(n4782), .ZN(n6394) );
  INV_X1 U5280 ( .A(DATAI_0_), .ZN(n6387) );
  INV_X1 U5281 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6995) );
  OAI222_X1 U5282 ( .A1(n6394), .A2(n6387), .B1(n6392), .B2(n6995), .C1(n6391), 
        .C2(n5462), .ZN(U2891) );
  INV_X1 U5283 ( .A(DATAI_1_), .ZN(n4904) );
  INV_X1 U5284 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6997) );
  OAI222_X1 U5285 ( .A1(n4904), .A2(n6394), .B1(n6392), .B2(n6997), .C1(n6391), 
        .C2(n5524), .ZN(U2890) );
  OR2_X1 U5286 ( .A1(n6184), .A2(n5149), .ZN(n4785) );
  NAND2_X1 U5287 ( .A1(n6962), .A2(n4787), .ZN(n4784) );
  NAND2_X1 U5288 ( .A1(n4785), .A2(n4784), .ZN(n7455) );
  OAI22_X1 U5289 ( .A1(n6069), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n7487), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4786) );
  AOI21_X1 U5290 ( .B1(n7455), .B2(n7481), .A(n4786), .ZN(n4790) );
  NAND2_X1 U5291 ( .A1(n6964), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7453) );
  INV_X1 U5292 ( .A(n7481), .ZN(n6971) );
  INV_X1 U5293 ( .A(n6076), .ZN(n7441) );
  OAI22_X1 U5294 ( .A1(n7453), .A2(n6971), .B1(n4787), .B2(n7441), .ZN(n4788)
         );
  INV_X1 U5295 ( .A(n4788), .ZN(n4789) );
  OAI21_X1 U5296 ( .B1(n4790), .B2(n6076), .A(n4789), .ZN(U3461) );
  NAND2_X1 U5297 ( .A1(n4792), .A2(n4791), .ZN(n4793) );
  XOR2_X1 U5298 ( .A(n4794), .B(n4793), .Z(n7181) );
  INV_X1 U5299 ( .A(n7433), .ZN(n7148) );
  NAND2_X1 U5300 ( .A1(n7181), .A2(n7148), .ZN(n4798) );
  INV_X1 U5301 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U5302 ( .A1(n7205), .A2(REIP_REG_1__SCAN_IN), .ZN(n7177) );
  OAI21_X1 U5303 ( .B1(n7132), .B2(n4796), .A(n7177), .ZN(n4795) );
  AOI21_X1 U5304 ( .B1(n7143), .B2(n4796), .A(n4795), .ZN(n4797) );
  OAI211_X1 U5305 ( .C1(n6489), .C2(n5524), .A(n4798), .B(n4797), .ZN(U2985)
         );
  INV_X1 U5306 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U5307 ( .A1(n7167), .A2(UWORD_REG_14__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4799) );
  OAI21_X1 U5308 ( .B1(n4800), .B2(n4808), .A(n4799), .ZN(U2893) );
  INV_X1 U5309 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5310 ( .A1(n7167), .A2(UWORD_REG_0__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4801) );
  OAI21_X1 U5311 ( .B1(n4802), .B2(n4808), .A(n4801), .ZN(U2907) );
  INV_X1 U5312 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5313 ( .A1(n7167), .A2(UWORD_REG_1__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4803) );
  OAI21_X1 U5314 ( .B1(n4804), .B2(n4808), .A(n4803), .ZN(U2906) );
  INV_X1 U5315 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4806) );
  AOI22_X1 U5316 ( .A1(n7167), .A2(UWORD_REG_2__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4805) );
  OAI21_X1 U5317 ( .B1(n4806), .B2(n4808), .A(n4805), .ZN(U2905) );
  INV_X1 U5318 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4809) );
  AOI22_X1 U5319 ( .A1(n7167), .A2(UWORD_REG_3__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4807) );
  OAI21_X1 U5320 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(U2904) );
  INV_X1 U5321 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U5322 ( .A1(n4810), .A2(DATAI_13_), .ZN(n4829) );
  NAND2_X1 U5323 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n4811), .ZN(n4812) );
  OAI211_X1 U5324 ( .C1(n4813), .C2(n7019), .A(n4829), .B(n4812), .ZN(U2952)
         );
  AOI22_X1 U5325 ( .A1(n4840), .A2(EAX_REG_20__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4814) );
  NAND2_X1 U5326 ( .A1(n4815), .A2(n4814), .ZN(U2928) );
  AOI22_X1 U5327 ( .A1(n4840), .A2(EAX_REG_22__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4816) );
  NAND2_X1 U5328 ( .A1(n4817), .A2(n4816), .ZN(U2930) );
  AOI22_X1 U5329 ( .A1(n4840), .A2(EAX_REG_24__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4818) );
  NAND2_X1 U5330 ( .A1(n4819), .A2(n4818), .ZN(U2932) );
  AOI22_X1 U5331 ( .A1(n4840), .A2(EAX_REG_25__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U5332 ( .A1(n4821), .A2(n4820), .ZN(U2933) );
  AOI22_X1 U5333 ( .A1(n4840), .A2(EAX_REG_1__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U5334 ( .A1(n4823), .A2(n4822), .ZN(U2940) );
  AOI22_X1 U5335 ( .A1(n4840), .A2(EAX_REG_27__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5336 ( .A1(n4825), .A2(n4824), .ZN(U2935) );
  AOI22_X1 U5337 ( .A1(n4840), .A2(EAX_REG_28__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U5338 ( .A1(n4827), .A2(n4826), .ZN(U2936) );
  AOI22_X1 U5339 ( .A1(n4840), .A2(EAX_REG_29__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U5340 ( .A1(n4829), .A2(n4828), .ZN(U2937) );
  AOI22_X1 U5341 ( .A1(n4840), .A2(EAX_REG_30__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5342 ( .A1(n4831), .A2(n4830), .ZN(U2938) );
  AOI22_X1 U5343 ( .A1(n4840), .A2(EAX_REG_0__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U5344 ( .A1(n4833), .A2(n4832), .ZN(U2939) );
  AOI22_X1 U5345 ( .A1(n4840), .A2(EAX_REG_26__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5346 ( .A1(n4835), .A2(n4834), .ZN(U2934) );
  AOI22_X1 U5347 ( .A1(n4840), .A2(EAX_REG_2__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U5348 ( .A1(n4837), .A2(n4836), .ZN(U2941) );
  AOI22_X1 U5349 ( .A1(n4840), .A2(EAX_REG_23__SCAN_IN), .B1(n4811), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4838) );
  NAND2_X1 U5350 ( .A1(n4839), .A2(n4838), .ZN(U2931) );
  INV_X1 U5351 ( .A(DATAI_15_), .ZN(n6390) );
  AOI22_X1 U5352 ( .A1(n4840), .A2(EAX_REG_15__SCAN_IN), .B1(n4811), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4841) );
  OAI21_X1 U5353 ( .B1(n4842), .B2(n6390), .A(n4841), .ZN(U2954) );
  INV_X1 U5354 ( .A(n4843), .ZN(n4846) );
  INV_X1 U5355 ( .A(n4886), .ZN(n4844) );
  AOI21_X1 U5356 ( .B1(n4846), .B2(n4845), .A(n4844), .ZN(n7255) );
  INV_X1 U5357 ( .A(n7255), .ZN(n4889) );
  INV_X1 U5358 ( .A(n4847), .ZN(n4848) );
  AOI21_X2 U5359 ( .B1(n5522), .B2(n5924), .A(n4848), .ZN(n4855) );
  OR2_X1 U5360 ( .A1(n5947), .A2(EBX_REG_2__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5361 ( .A1(n5948), .A2(n4849), .ZN(n4851) );
  INV_X1 U5362 ( .A(EBX_REG_2__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U5363 ( .A1(n5924), .A2(n7252), .ZN(n4850) );
  NAND3_X1 U5364 ( .A1(n4851), .A2(n5322), .A3(n4850), .ZN(n4852) );
  NAND2_X1 U5365 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  NAND2_X1 U5366 ( .A1(n4855), .A2(n4854), .ZN(n4871) );
  OR2_X1 U5367 ( .A1(n4855), .A2(n4854), .ZN(n4856) );
  NAND2_X1 U5368 ( .A1(n4871), .A2(n4856), .ZN(n7258) );
  INV_X1 U5369 ( .A(n7258), .ZN(n4857) );
  AOI22_X1 U5370 ( .A1(n7114), .A2(n4857), .B1(EBX_REG_2__SCAN_IN), .B2(n6338), 
        .ZN(n4858) );
  OAI21_X1 U5371 ( .B1(n4889), .B2(n6357), .A(n4858), .ZN(U2857) );
  NAND2_X1 U5372 ( .A1(n4860), .A2(n4859), .ZN(n4862) );
  XNOR2_X1 U5373 ( .A(n4862), .B(n4861), .ZN(n4938) );
  AOI21_X1 U5374 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4866) );
  INV_X1 U5375 ( .A(n4866), .ZN(n7193) );
  NAND2_X1 U5376 ( .A1(n4865), .A2(n4863), .ZN(n6029) );
  NAND2_X1 U5377 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7194) );
  OR2_X1 U5378 ( .A1(n4863), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4864)
         );
  NAND2_X1 U5379 ( .A1(n4864), .A2(n7184), .ZN(n5839) );
  AOI21_X1 U5380 ( .B1(n6029), .B2(n7194), .A(n5839), .ZN(n7203) );
  OAI21_X1 U5381 ( .B1(n6036), .B2(n7193), .A(n7203), .ZN(n5263) );
  NAND2_X1 U5382 ( .A1(n4865), .A2(n7195), .ZN(n7176) );
  NAND2_X1 U5383 ( .A1(n6029), .A2(n7176), .ZN(n6566) );
  INV_X1 U5384 ( .A(n7194), .ZN(n5425) );
  AOI21_X1 U5385 ( .B1(n6946), .B2(n5425), .A(n7197), .ZN(n5423) );
  NOR2_X1 U5386 ( .A1(n4866), .A2(n5423), .ZN(n4882) );
  AOI22_X1 U5387 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n5263), .B1(n4882), 
        .B2(n3950), .ZN(n4874) );
  MUX2_X1 U5388 ( .A(n5956), .B(n5322), .S(EBX_REG_3__SCAN_IN), .Z(n4867) );
  OAI21_X1 U5389 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5963), .A(n4867), 
        .ZN(n4870) );
  NAND2_X1 U5390 ( .A1(n4871), .A2(n4870), .ZN(n4872) );
  AND2_X1 U5391 ( .A1(n4880), .A2(n4872), .ZN(n5589) );
  AND2_X1 U5392 ( .A1(n7205), .A2(REIP_REG_3__SCAN_IN), .ZN(n4934) );
  AOI21_X1 U5393 ( .B1(n7238), .B2(n5589), .A(n4934), .ZN(n4873) );
  OAI211_X1 U5394 ( .C1(n4938), .C2(n6584), .A(n4874), .B(n4873), .ZN(U3015)
         );
  XNOR2_X1 U5395 ( .A(n4876), .B(n4875), .ZN(n5282) );
  INV_X1 U5396 ( .A(n7238), .ZN(n7215) );
  MUX2_X1 U5397 ( .A(n5947), .B(n5948), .S(EBX_REG_4__SCAN_IN), .Z(n4878) );
  NAND2_X1 U5398 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n5962), .ZN(n4877)
         );
  OR2_X2 U5399 ( .A1(n4880), .A2(n4879), .ZN(n5027) );
  NAND2_X1 U5400 ( .A1(n4880), .A2(n4879), .ZN(n4881) );
  NAND2_X1 U5401 ( .A1(n5027), .A2(n4881), .ZN(n7262) );
  NAND2_X1 U5402 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5264) );
  OAI211_X1 U5403 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4882), .B(n5264), .ZN(n4883) );
  INV_X1 U5404 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7272) );
  OR2_X1 U5405 ( .A1(n7213), .A2(n7272), .ZN(n5277) );
  OAI211_X1 U5406 ( .C1(n7215), .C2(n7262), .A(n4883), .B(n5277), .ZN(n4884)
         );
  AOI21_X1 U5407 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n5263), .A(n4884), 
        .ZN(n4885) );
  OAI21_X1 U5408 ( .B1(n5282), .B2(n6584), .A(n4885), .ZN(U3014) );
  AOI21_X1 U5409 ( .B1(n4887), .B2(n4886), .A(n5019), .ZN(n5600) );
  INV_X1 U5410 ( .A(n5600), .ZN(n5060) );
  AOI22_X1 U5411 ( .A1(n7114), .A2(n5589), .B1(EBX_REG_3__SCAN_IN), .B2(n6338), 
        .ZN(n4888) );
  OAI21_X1 U5412 ( .B1(n5060), .B2(n6357), .A(n4888), .ZN(U2856) );
  INV_X1 U5413 ( .A(DATAI_2_), .ZN(n6384) );
  INV_X1 U5414 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6999) );
  OAI222_X1 U5415 ( .A1(n6394), .A2(n6384), .B1(n6392), .B2(n6999), .C1(n6391), 
        .C2(n4889), .ZN(U2889) );
  INV_X1 U5416 ( .A(n5031), .ZN(n4891) );
  NOR2_X1 U5417 ( .A1(n4891), .A2(n4890), .ZN(n5094) );
  AND2_X1 U5418 ( .A1(n5094), .A2(n5187), .ZN(n4900) );
  NAND2_X1 U5419 ( .A1(n5756), .A2(n7502), .ZN(n5629) );
  OAI21_X1 U5420 ( .B1(n4900), .B2(n6489), .A(n5629), .ZN(n4895) );
  INV_X1 U5421 ( .A(n5032), .ZN(n5628) );
  INV_X1 U5422 ( .A(n6184), .ZN(n4941) );
  AND2_X1 U5423 ( .A1(n5592), .A2(n4941), .ZN(n5122) );
  INV_X1 U5424 ( .A(n4892), .ZN(n5518) );
  OR2_X1 U5425 ( .A1(n7246), .A2(n5518), .ZN(n5534) );
  INV_X1 U5426 ( .A(n5534), .ZN(n5290) );
  AND2_X1 U5427 ( .A1(n4893), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4928)
         );
  AOI21_X1 U5428 ( .B1(n5122), .B2(n5290), .A(n4928), .ZN(n4897) );
  NOR3_X1 U5429 ( .A1(n4112), .A2(n7462), .A3(n5381), .ZN(n4896) );
  OAI21_X1 U5430 ( .B1(n7495), .B2(n7484), .A(n6069), .ZN(n4898) );
  NAND2_X1 U5431 ( .A1(n7161), .A2(n4898), .ZN(n5175) );
  AOI21_X1 U5432 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6175), .A(n5175), .ZN(
        n5294) );
  OAI21_X1 U5433 ( .B1(n5756), .B2(n4896), .A(n5294), .ZN(n4894) );
  AOI21_X1 U5434 ( .B1(n4895), .B2(n4897), .A(n4894), .ZN(n4933) );
  INV_X1 U5435 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4903) );
  INV_X1 U5436 ( .A(n4896), .ZN(n5192) );
  OAI22_X1 U5437 ( .A1(n4897), .A2(n5379), .B1(n5192), .B2(n5995), .ZN(n4929)
         );
  NOR2_X1 U5438 ( .A1(n6384), .A2(n5175), .ZN(n5568) );
  NAND2_X1 U5439 ( .A1(n4927), .A2(n4899), .ZN(n5657) );
  INV_X1 U5440 ( .A(n5657), .ZN(n5797) );
  AOI22_X1 U5441 ( .A1(n4929), .A2(n5568), .B1(n5797), .B2(n4928), .ZN(n4902)
         );
  INV_X1 U5442 ( .A(n6180), .ZN(n5288) );
  NAND2_X1 U5443 ( .A1(n4900), .A2(n5288), .ZN(n5194) );
  AND2_X1 U5444 ( .A1(n3628), .A2(DATAI_26_), .ZN(n5801) );
  NAND2_X1 U5445 ( .A1(n3628), .A2(DATAI_18_), .ZN(n5799) );
  INV_X1 U5446 ( .A(n5799), .ZN(n5659) );
  AOI22_X1 U5447 ( .A1(n5229), .A2(n5801), .B1(n7571), .B2(n5659), .ZN(n4901)
         );
  OAI211_X1 U5448 ( .C1(n4933), .C2(n4903), .A(n4902), .B(n4901), .ZN(U3142)
         );
  INV_X1 U5449 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4908) );
  NOR2_X1 U5450 ( .A1(n4904), .A2(n5175), .ZN(n7550) );
  NAND2_X1 U5451 ( .A1(n4927), .A2(n3627), .ZN(n5663) );
  INV_X1 U5452 ( .A(n5663), .ZN(n7551) );
  AOI22_X1 U5453 ( .A1(n4929), .A2(n7550), .B1(n7551), .B2(n4928), .ZN(n4907)
         );
  AND2_X1 U5454 ( .A1(n3628), .A2(DATAI_25_), .ZN(n7553) );
  NAND2_X1 U5455 ( .A1(n3628), .A2(DATAI_17_), .ZN(n5771) );
  INV_X1 U5456 ( .A(n5771), .ZN(n7552) );
  AOI22_X1 U5457 ( .A1(n5229), .A2(n7553), .B1(n7571), .B2(n7552), .ZN(n4906)
         );
  OAI211_X1 U5458 ( .C1(n4933), .C2(n4908), .A(n4907), .B(n4906), .ZN(U3141)
         );
  INV_X1 U5459 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4911) );
  NOR2_X1 U5460 ( .A1(n6387), .A2(n5175), .ZN(n7543) );
  NAND2_X1 U5461 ( .A1(n4927), .A2(n3632), .ZN(n5646) );
  INV_X1 U5462 ( .A(n5646), .ZN(n7544) );
  AOI22_X1 U5463 ( .A1(n4929), .A2(n7543), .B1(n7544), .B2(n4928), .ZN(n4910)
         );
  AND2_X1 U5464 ( .A1(n3628), .A2(DATAI_24_), .ZN(n7546) );
  NAND2_X1 U5465 ( .A1(n3628), .A2(DATAI_16_), .ZN(n5776) );
  INV_X1 U5466 ( .A(n5776), .ZN(n7545) );
  AOI22_X1 U5467 ( .A1(n5229), .A2(n7546), .B1(n7571), .B2(n7545), .ZN(n4909)
         );
  OAI211_X1 U5468 ( .C1(n4933), .C2(n4911), .A(n4910), .B(n4909), .ZN(U3140)
         );
  INV_X1 U5469 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4914) );
  INV_X1 U5470 ( .A(DATAI_7_), .ZN(n6381) );
  NOR2_X1 U5471 ( .A1(n6381), .A2(n5175), .ZN(n5541) );
  NAND2_X1 U5472 ( .A1(n4927), .A2(n6119), .ZN(n5668) );
  INV_X1 U5473 ( .A(n5668), .ZN(n5804) );
  AOI22_X1 U5474 ( .A1(n4929), .A2(n5541), .B1(n5804), .B2(n4928), .ZN(n4913)
         );
  AND2_X1 U5475 ( .A1(n3628), .A2(DATAI_31_), .ZN(n5808) );
  NAND2_X1 U5476 ( .A1(n3628), .A2(DATAI_23_), .ZN(n5806) );
  INV_X1 U5477 ( .A(n5806), .ZN(n5670) );
  AOI22_X1 U5478 ( .A1(n5229), .A2(n5808), .B1(n7571), .B2(n5670), .ZN(n4912)
         );
  OAI211_X1 U5479 ( .C1(n4933), .C2(n4914), .A(n4913), .B(n4912), .ZN(U3147)
         );
  INV_X1 U5480 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4918) );
  INV_X1 U5481 ( .A(DATAI_6_), .ZN(n5287) );
  NOR2_X1 U5482 ( .A1(n5287), .A2(n5175), .ZN(n5536) );
  NAND2_X1 U5483 ( .A1(n4927), .A2(n4915), .ZN(n5640) );
  INV_X1 U5484 ( .A(n5640), .ZN(n5813) );
  AOI22_X1 U5485 ( .A1(n4929), .A2(n5536), .B1(n5813), .B2(n4928), .ZN(n4917)
         );
  AND2_X1 U5486 ( .A1(n3628), .A2(DATAI_30_), .ZN(n5819) );
  NAND2_X1 U5487 ( .A1(n3628), .A2(DATAI_22_), .ZN(n5815) );
  INV_X1 U5488 ( .A(n5815), .ZN(n5642) );
  AOI22_X1 U5489 ( .A1(n5229), .A2(n5819), .B1(n7571), .B2(n5642), .ZN(n4916)
         );
  OAI211_X1 U5490 ( .C1(n4933), .C2(n4918), .A(n4917), .B(n4916), .ZN(U3146)
         );
  INV_X1 U5491 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4921) );
  INV_X1 U5492 ( .A(DATAI_4_), .ZN(n5030) );
  NOR2_X1 U5493 ( .A1(n5030), .A2(n5175), .ZN(n7557) );
  NAND2_X1 U5494 ( .A1(n4927), .A2(n3764), .ZN(n5674) );
  INV_X1 U5495 ( .A(n5674), .ZN(n7558) );
  AOI22_X1 U5496 ( .A1(n4929), .A2(n7557), .B1(n7558), .B2(n4928), .ZN(n4920)
         );
  AND2_X1 U5497 ( .A1(n3628), .A2(DATAI_28_), .ZN(n7560) );
  NAND2_X1 U5498 ( .A1(n3628), .A2(DATAI_20_), .ZN(n5781) );
  INV_X1 U5499 ( .A(n5781), .ZN(n7559) );
  AOI22_X1 U5500 ( .A1(n5229), .A2(n7560), .B1(n7571), .B2(n7559), .ZN(n4919)
         );
  OAI211_X1 U5501 ( .C1(n4933), .C2(n4921), .A(n4920), .B(n4919), .ZN(U3144)
         );
  INV_X1 U5502 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4925) );
  INV_X1 U5503 ( .A(DATAI_5_), .ZN(n5058) );
  NOR2_X1 U5504 ( .A1(n5058), .A2(n5175), .ZN(n7564) );
  NAND2_X1 U5505 ( .A1(n4927), .A2(n4922), .ZN(n5681) );
  INV_X1 U5506 ( .A(n5681), .ZN(n7567) );
  AOI22_X1 U5507 ( .A1(n4929), .A2(n7564), .B1(n7567), .B2(n4928), .ZN(n4924)
         );
  AND2_X1 U5508 ( .A1(n3628), .A2(DATAI_29_), .ZN(n7570) );
  NAND2_X1 U5509 ( .A1(n3628), .A2(DATAI_21_), .ZN(n5793) );
  INV_X1 U5510 ( .A(n5793), .ZN(n7568) );
  AOI22_X1 U5511 ( .A1(n5229), .A2(n7570), .B1(n7571), .B2(n7568), .ZN(n4923)
         );
  OAI211_X1 U5512 ( .C1(n4933), .C2(n4925), .A(n4924), .B(n4923), .ZN(U3145)
         );
  INV_X1 U5513 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4932) );
  INV_X1 U5514 ( .A(DATAI_3_), .ZN(n5061) );
  NOR2_X1 U5515 ( .A1(n5061), .A2(n5175), .ZN(n5554) );
  NAND2_X1 U5516 ( .A1(n4927), .A2(n4926), .ZN(n5651) );
  INV_X1 U5517 ( .A(n5651), .ZN(n5785) );
  AOI22_X1 U5518 ( .A1(n4929), .A2(n5554), .B1(n5785), .B2(n4928), .ZN(n4931)
         );
  AND2_X1 U5519 ( .A1(n3628), .A2(DATAI_27_), .ZN(n5789) );
  NAND2_X1 U5520 ( .A1(n3628), .A2(DATAI_19_), .ZN(n5787) );
  INV_X1 U5521 ( .A(n5787), .ZN(n5653) );
  AOI22_X1 U5522 ( .A1(n5229), .A2(n5789), .B1(n7571), .B2(n5653), .ZN(n4930)
         );
  OAI211_X1 U5523 ( .C1(n4933), .C2(n4932), .A(n4931), .B(n4930), .ZN(U3143)
         );
  AOI21_X1 U5524 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4934), 
        .ZN(n4935) );
  OAI21_X1 U5525 ( .B1(n5590), .B2(n7152), .A(n4935), .ZN(n4936) );
  AOI21_X1 U5526 ( .B1(n5600), .B2(n3628), .A(n4936), .ZN(n4937) );
  OAI21_X1 U5527 ( .B1(n4938), .B2(n7433), .A(n4937), .ZN(U2983) );
  INV_X1 U5528 ( .A(n5233), .ZN(n5066) );
  INV_X1 U5529 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U5530 ( .A1(n5062), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5065) );
  OAI21_X1 U5531 ( .B1(n5066), .B2(n5065), .A(n5756), .ZN(n4946) );
  INV_X1 U5532 ( .A(n4946), .ZN(n4944) );
  AND2_X1 U5533 ( .A1(n4892), .A2(n7246), .ZN(n5637) );
  AND2_X1 U5534 ( .A1(n5637), .A2(n5032), .ZN(n5763) );
  NAND3_X1 U5535 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7462), .ZN(n5762) );
  NOR2_X1 U5536 ( .A1(n6175), .A2(n5762), .ZN(n4975) );
  AOI21_X1 U5537 ( .B1(n5763), .B2(n4941), .A(n4975), .ZN(n4945) );
  INV_X1 U5538 ( .A(n5762), .ZN(n4942) );
  OAI21_X1 U5539 ( .B1(n5756), .B2(n4942), .A(n5294), .ZN(n4943) );
  AOI21_X1 U5540 ( .B1(n4944), .B2(n4945), .A(n4943), .ZN(n4981) );
  INV_X1 U5541 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U5542 ( .A1(n4946), .A2(n4945), .B1(n5762), .B2(n5995), .ZN(n4978)
         );
  AND3_X1 U5543 ( .A1(n5233), .A2(n5062), .A3(n6180), .ZN(n4982) );
  AOI22_X1 U5544 ( .A1(n5761), .A2(n7546), .B1(n7544), .B2(n4975), .ZN(n4947)
         );
  OAI21_X1 U5545 ( .B1(n5776), .B2(n5017), .A(n4947), .ZN(n4948) );
  AOI21_X1 U5546 ( .B1(n4978), .B2(n7543), .A(n4948), .ZN(n4949) );
  OAI21_X1 U5547 ( .B1(n4981), .B2(n4950), .A(n4949), .ZN(U3108) );
  INV_X1 U5548 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U5549 ( .A1(n5761), .A2(n7553), .B1(n7551), .B2(n4975), .ZN(n4951)
         );
  OAI21_X1 U5550 ( .B1(n5771), .B2(n5017), .A(n4951), .ZN(n4952) );
  AOI21_X1 U5551 ( .B1(n4978), .B2(n7550), .A(n4952), .ZN(n4953) );
  OAI21_X1 U5552 ( .B1(n4981), .B2(n4954), .A(n4953), .ZN(U3109) );
  INV_X1 U5553 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4958) );
  AOI22_X1 U5554 ( .A1(n5761), .A2(n5808), .B1(n5804), .B2(n4975), .ZN(n4955)
         );
  OAI21_X1 U5555 ( .B1(n5806), .B2(n5017), .A(n4955), .ZN(n4956) );
  AOI21_X1 U5556 ( .B1(n4978), .B2(n5541), .A(n4956), .ZN(n4957) );
  OAI21_X1 U5557 ( .B1(n4981), .B2(n4958), .A(n4957), .ZN(U3115) );
  INV_X1 U5558 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4962) );
  AOI22_X1 U5559 ( .A1(n5761), .A2(n7560), .B1(n7558), .B2(n4975), .ZN(n4959)
         );
  OAI21_X1 U5560 ( .B1(n5781), .B2(n5017), .A(n4959), .ZN(n4960) );
  AOI21_X1 U5561 ( .B1(n4978), .B2(n7557), .A(n4960), .ZN(n4961) );
  OAI21_X1 U5562 ( .B1(n4981), .B2(n4962), .A(n4961), .ZN(U3112) );
  INV_X1 U5563 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4966) );
  AOI22_X1 U5564 ( .A1(n5761), .A2(n5789), .B1(n5785), .B2(n4975), .ZN(n4963)
         );
  OAI21_X1 U5565 ( .B1(n5787), .B2(n5017), .A(n4963), .ZN(n4964) );
  AOI21_X1 U5566 ( .B1(n4978), .B2(n5554), .A(n4964), .ZN(n4965) );
  OAI21_X1 U5567 ( .B1(n4981), .B2(n4966), .A(n4965), .ZN(U3111) );
  INV_X1 U5568 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4970) );
  AOI22_X1 U5569 ( .A1(n5761), .A2(n5801), .B1(n5797), .B2(n4975), .ZN(n4967)
         );
  OAI21_X1 U5570 ( .B1(n5799), .B2(n5017), .A(n4967), .ZN(n4968) );
  AOI21_X1 U5571 ( .B1(n4978), .B2(n5568), .A(n4968), .ZN(n4969) );
  OAI21_X1 U5572 ( .B1(n4981), .B2(n4970), .A(n4969), .ZN(U3110) );
  INV_X1 U5573 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U5574 ( .A1(n5761), .A2(n7570), .B1(n7567), .B2(n4975), .ZN(n4971)
         );
  OAI21_X1 U5575 ( .B1(n5793), .B2(n5017), .A(n4971), .ZN(n4972) );
  AOI21_X1 U5576 ( .B1(n4978), .B2(n7564), .A(n4972), .ZN(n4973) );
  OAI21_X1 U5577 ( .B1(n4981), .B2(n4974), .A(n4973), .ZN(U3113) );
  INV_X1 U5578 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4980) );
  AOI22_X1 U5579 ( .A1(n5761), .A2(n5819), .B1(n5813), .B2(n4975), .ZN(n4976)
         );
  OAI21_X1 U5580 ( .B1(n5815), .B2(n5017), .A(n4976), .ZN(n4977) );
  AOI21_X1 U5581 ( .B1(n4978), .B2(n5536), .A(n4977), .ZN(n4979) );
  OAI21_X1 U5582 ( .B1(n4981), .B2(n4980), .A(n4979), .ZN(U3114) );
  INV_X1 U5583 ( .A(n7553), .ZN(n5667) );
  OR2_X1 U5584 ( .A1(n7246), .A2(n4892), .ZN(n5033) );
  NAND2_X1 U5585 ( .A1(n5033), .A2(n5756), .ZN(n5330) );
  NOR2_X1 U5586 ( .A1(n5187), .A2(n6180), .ZN(n5038) );
  AOI211_X1 U5587 ( .C1(n5535), .C2(n5330), .A(n4982), .B(n5117), .ZN(n4985)
         );
  INV_X1 U5588 ( .A(n5175), .ZN(n5376) );
  INV_X1 U5589 ( .A(n4987), .ZN(n4983) );
  NAND2_X1 U5590 ( .A1(n4983), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5475) );
  NAND3_X1 U5591 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5381), .ZN(n5097) );
  NOR2_X1 U5592 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5097), .ZN(n4986)
         );
  INV_X1 U5593 ( .A(n5629), .ZN(n5469) );
  NAND2_X1 U5594 ( .A1(n5033), .A2(n5469), .ZN(n5333) );
  INV_X1 U5595 ( .A(n5529), .ZN(n5238) );
  NAND2_X1 U5596 ( .A1(n5336), .A2(n5238), .ZN(n5476) );
  NAND2_X1 U5597 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5476), .ZN(n5466) );
  OAI211_X1 U5598 ( .C1(n4732), .C2(n4986), .A(n5333), .B(n5466), .ZN(n4984)
         );
  NAND2_X1 U5599 ( .A1(n5011), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4992)
         );
  INV_X1 U5600 ( .A(n4986), .ZN(n5013) );
  NAND2_X1 U5601 ( .A1(n5592), .A2(n5756), .ZN(n5527) );
  OR2_X1 U5602 ( .A1(n5527), .A2(n5033), .ZN(n4989) );
  NAND2_X1 U5603 ( .A1(n4987), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5533) );
  OR2_X1 U5604 ( .A1(n5476), .A2(n5533), .ZN(n4988) );
  AND2_X1 U5605 ( .A1(n4989), .A2(n4988), .ZN(n5012) );
  INV_X1 U5606 ( .A(n7550), .ZN(n5774) );
  OAI22_X1 U5607 ( .A1(n5663), .A2(n5013), .B1(n5012), .B2(n5774), .ZN(n4990)
         );
  AOI21_X1 U5608 ( .B1(n5117), .B2(n7552), .A(n4990), .ZN(n4991) );
  OAI211_X1 U5609 ( .C1(n5017), .C2(n5667), .A(n4992), .B(n4991), .ZN(U3117)
         );
  INV_X1 U5610 ( .A(n7570), .ZN(n5688) );
  NAND2_X1 U5611 ( .A1(n5011), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4995)
         );
  INV_X1 U5612 ( .A(n7564), .ZN(n5796) );
  OAI22_X1 U5613 ( .A1(n5681), .A2(n5013), .B1(n5012), .B2(n5796), .ZN(n4993)
         );
  AOI21_X1 U5614 ( .B1(n5117), .B2(n7568), .A(n4993), .ZN(n4994) );
  OAI211_X1 U5615 ( .C1(n5017), .C2(n5688), .A(n4995), .B(n4994), .ZN(U3121)
         );
  INV_X1 U5616 ( .A(n7546), .ZN(n5650) );
  NAND2_X1 U5617 ( .A1(n5011), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4998)
         );
  INV_X1 U5618 ( .A(n7543), .ZN(n5779) );
  OAI22_X1 U5619 ( .A1(n5646), .A2(n5013), .B1(n5012), .B2(n5779), .ZN(n4996)
         );
  AOI21_X1 U5620 ( .B1(n5117), .B2(n7545), .A(n4996), .ZN(n4997) );
  OAI211_X1 U5621 ( .C1(n5017), .C2(n5650), .A(n4998), .B(n4997), .ZN(U3116)
         );
  INV_X1 U5622 ( .A(n5801), .ZN(n5662) );
  NAND2_X1 U5623 ( .A1(n5011), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5001)
         );
  INV_X1 U5624 ( .A(n5568), .ZN(n5803) );
  OAI22_X1 U5625 ( .A1(n5657), .A2(n5013), .B1(n5012), .B2(n5803), .ZN(n4999)
         );
  AOI21_X1 U5626 ( .B1(n5117), .B2(n5659), .A(n4999), .ZN(n5000) );
  OAI211_X1 U5627 ( .C1(n5017), .C2(n5662), .A(n5001), .B(n5000), .ZN(U3118)
         );
  INV_X1 U5628 ( .A(n5808), .ZN(n5673) );
  NAND2_X1 U5629 ( .A1(n5011), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5004)
         );
  INV_X1 U5630 ( .A(n5541), .ZN(n5810) );
  OAI22_X1 U5631 ( .A1(n5668), .A2(n5013), .B1(n5012), .B2(n5810), .ZN(n5002)
         );
  AOI21_X1 U5632 ( .B1(n5117), .B2(n5670), .A(n5002), .ZN(n5003) );
  OAI211_X1 U5633 ( .C1(n5017), .C2(n5673), .A(n5004), .B(n5003), .ZN(U3123)
         );
  INV_X1 U5634 ( .A(n5819), .ZN(n5645) );
  NAND2_X1 U5635 ( .A1(n5011), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5007)
         );
  INV_X1 U5636 ( .A(n5536), .ZN(n5821) );
  OAI22_X1 U5637 ( .A1(n5640), .A2(n5013), .B1(n5012), .B2(n5821), .ZN(n5005)
         );
  AOI21_X1 U5638 ( .B1(n5117), .B2(n5642), .A(n5005), .ZN(n5006) );
  OAI211_X1 U5639 ( .C1(n5017), .C2(n5645), .A(n5007), .B(n5006), .ZN(U3122)
         );
  INV_X1 U5640 ( .A(n5789), .ZN(n5656) );
  NAND2_X1 U5641 ( .A1(n5011), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5010)
         );
  INV_X1 U5642 ( .A(n5554), .ZN(n5791) );
  OAI22_X1 U5643 ( .A1(n5651), .A2(n5013), .B1(n5012), .B2(n5791), .ZN(n5008)
         );
  AOI21_X1 U5644 ( .B1(n5117), .B2(n5653), .A(n5008), .ZN(n5009) );
  OAI211_X1 U5645 ( .C1(n5017), .C2(n5656), .A(n5010), .B(n5009), .ZN(U3119)
         );
  INV_X1 U5646 ( .A(n7560), .ZN(n5678) );
  NAND2_X1 U5647 ( .A1(n5011), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5016)
         );
  INV_X1 U5648 ( .A(n7557), .ZN(n5784) );
  OAI22_X1 U5649 ( .A1(n5674), .A2(n5013), .B1(n5012), .B2(n5784), .ZN(n5014)
         );
  AOI21_X1 U5650 ( .B1(n5117), .B2(n7559), .A(n5014), .ZN(n5015) );
  OAI211_X1 U5651 ( .C1(n5017), .C2(n5678), .A(n5016), .B(n5015), .ZN(U3120)
         );
  INV_X1 U5652 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5020) );
  OAI21_X1 U5653 ( .B1(n5019), .B2(n5018), .A(n5022), .ZN(n7266) );
  OAI222_X1 U5654 ( .A1(n7262), .A2(n7105), .B1(n7118), .B2(n5020), .C1(n7266), 
        .C2(n6357), .ZN(U2855) );
  NAND2_X1 U5655 ( .A1(n5022), .A2(n5021), .ZN(n5023) );
  AND2_X1 U5656 ( .A1(n5283), .A2(n5023), .ZN(n7279) );
  INV_X1 U5657 ( .A(n7279), .ZN(n5059) );
  MUX2_X1 U5658 ( .A(n5956), .B(n5322), .S(EBX_REG_5__SCAN_IN), .Z(n5025) );
  OAI21_X1 U5659 ( .B1(n5963), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n5025), 
        .ZN(n5026) );
  NOR2_X4 U5660 ( .A1(n5027), .A2(n5026), .ZN(n5269) );
  AND2_X1 U5661 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  NOR2_X1 U5662 ( .A1(n5269), .A2(n5028), .ZN(n7273) );
  AOI22_X1 U5663 ( .A1(n7114), .A2(n7273), .B1(EBX_REG_5__SCAN_IN), .B2(n6338), 
        .ZN(n5029) );
  OAI21_X1 U5664 ( .B1(n5059), .B2(n6357), .A(n5029), .ZN(U2854) );
  INV_X1 U5665 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U5666 ( .A1(n6394), .A2(n5030), .B1(n6392), .B2(n7003), .C1(n6391), 
        .C2(n7266), .ZN(U2887) );
  NOR2_X1 U5667 ( .A1(n4890), .A2(n5031), .ZN(n5182) );
  NOR2_X1 U5668 ( .A1(n5187), .A2(n5288), .ZN(n5092) );
  NAND2_X1 U5669 ( .A1(n5182), .A2(n5092), .ZN(n5571) );
  OR2_X1 U5670 ( .A1(n5032), .A2(n6184), .ZN(n5371) );
  INV_X1 U5671 ( .A(n5371), .ZN(n5291) );
  INV_X1 U5672 ( .A(n5033), .ZN(n5338) );
  NAND3_X1 U5673 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4112), .A3(n5381), .ZN(n5331) );
  NOR2_X1 U5674 ( .A1(n6175), .A2(n5331), .ZN(n5055) );
  AOI21_X1 U5675 ( .B1(n5291), .B2(n5338), .A(n5055), .ZN(n5037) );
  NAND2_X1 U5676 ( .A1(n5178), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5177) );
  INV_X1 U5677 ( .A(n5177), .ZN(n5093) );
  AOI21_X1 U5678 ( .B1(n5182), .B2(n5093), .A(n5379), .ZN(n5035) );
  AOI22_X1 U5679 ( .A1(n5037), .A2(n5035), .B1(n5379), .B2(n5331), .ZN(n5034)
         );
  NAND2_X1 U5680 ( .A1(n5294), .A2(n5034), .ZN(n5054) );
  INV_X1 U5681 ( .A(n5035), .ZN(n5036) );
  OAI22_X1 U5682 ( .A1(n5037), .A2(n5036), .B1(n5995), .B2(n5331), .ZN(n5053)
         );
  AOI22_X1 U5683 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5054), .B1(n5541), 
        .B2(n5053), .ZN(n5040) );
  AOI22_X1 U5684 ( .A1(n5365), .A2(n5808), .B1(n5804), .B2(n5055), .ZN(n5039)
         );
  OAI211_X1 U5685 ( .C1(n5806), .C2(n5571), .A(n5040), .B(n5039), .ZN(U3067)
         );
  AOI22_X1 U5686 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5054), .B1(n7564), 
        .B2(n5053), .ZN(n5042) );
  AOI22_X1 U5687 ( .A1(n5365), .A2(n7570), .B1(n7567), .B2(n5055), .ZN(n5041)
         );
  OAI211_X1 U5688 ( .C1(n5793), .C2(n5571), .A(n5042), .B(n5041), .ZN(U3065)
         );
  AOI22_X1 U5689 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5054), .B1(n5554), 
        .B2(n5053), .ZN(n5044) );
  AOI22_X1 U5690 ( .A1(n5365), .A2(n5789), .B1(n5785), .B2(n5055), .ZN(n5043)
         );
  OAI211_X1 U5691 ( .C1(n5787), .C2(n5571), .A(n5044), .B(n5043), .ZN(U3063)
         );
  AOI22_X1 U5692 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5054), .B1(n5568), 
        .B2(n5053), .ZN(n5046) );
  AOI22_X1 U5693 ( .A1(n5365), .A2(n5801), .B1(n5797), .B2(n5055), .ZN(n5045)
         );
  OAI211_X1 U5694 ( .C1(n5799), .C2(n5571), .A(n5046), .B(n5045), .ZN(U3062)
         );
  AOI22_X1 U5695 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5054), .B1(n7550), 
        .B2(n5053), .ZN(n5048) );
  AOI22_X1 U5696 ( .A1(n5365), .A2(n7553), .B1(n7551), .B2(n5055), .ZN(n5047)
         );
  OAI211_X1 U5697 ( .C1(n5771), .C2(n5571), .A(n5048), .B(n5047), .ZN(U3061)
         );
  AOI22_X1 U5698 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5054), .B1(n7543), 
        .B2(n5053), .ZN(n5050) );
  AOI22_X1 U5699 ( .A1(n5365), .A2(n7546), .B1(n7544), .B2(n5055), .ZN(n5049)
         );
  OAI211_X1 U5700 ( .C1(n5776), .C2(n5571), .A(n5050), .B(n5049), .ZN(U3060)
         );
  AOI22_X1 U5701 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5054), .B1(n5536), 
        .B2(n5053), .ZN(n5052) );
  AOI22_X1 U5702 ( .A1(n5365), .A2(n5819), .B1(n5813), .B2(n5055), .ZN(n5051)
         );
  OAI211_X1 U5703 ( .C1(n5815), .C2(n5571), .A(n5052), .B(n5051), .ZN(U3066)
         );
  AOI22_X1 U5704 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5054), .B1(n7557), 
        .B2(n5053), .ZN(n5057) );
  AOI22_X1 U5705 ( .A1(n5365), .A2(n7560), .B1(n7558), .B2(n5055), .ZN(n5056)
         );
  OAI211_X1 U5706 ( .C1(n5781), .C2(n5571), .A(n5057), .B(n5056), .ZN(U3064)
         );
  OAI222_X1 U5707 ( .A1(n5059), .A2(n6391), .B1(n6394), .B2(n5058), .C1(n6392), 
        .C2(n4697), .ZN(U2886) );
  INV_X1 U5708 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7001) );
  OAI222_X1 U5709 ( .A1(n5061), .A2(n6394), .B1(n6392), .B2(n7001), .C1(n6391), 
        .C2(n5060), .ZN(U2888) );
  NAND2_X1 U5710 ( .A1(n5066), .A2(n5062), .ZN(n5072) );
  INV_X1 U5711 ( .A(n5072), .ZN(n5063) );
  NAND2_X1 U5712 ( .A1(n4112), .A2(n7462), .ZN(n5370) );
  NOR2_X1 U5713 ( .A1(n5064), .A2(n5370), .ZN(n5089) );
  AOI21_X1 U5714 ( .B1(n5291), .B2(n5637), .A(n5089), .ZN(n5070) );
  INV_X1 U5715 ( .A(n5065), .ZN(n5067) );
  AOI21_X1 U5716 ( .B1(n5067), .B2(n5066), .A(n5379), .ZN(n5069) );
  INV_X1 U5717 ( .A(n5370), .ZN(n5382) );
  NAND2_X1 U5718 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5382), .ZN(n5632) );
  AOI22_X1 U5719 ( .A1(n5070), .A2(n5069), .B1(n5379), .B2(n5632), .ZN(n5068)
         );
  NAND2_X1 U5720 ( .A1(n5294), .A2(n5068), .ZN(n5088) );
  INV_X1 U5721 ( .A(n5069), .ZN(n5071) );
  OAI22_X1 U5722 ( .A1(n5071), .A2(n5070), .B1(n5995), .B2(n5632), .ZN(n5087)
         );
  AOI22_X1 U5723 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5088), .B1(n7543), 
        .B2(n5087), .ZN(n5074) );
  NOR2_X2 U5724 ( .A1(n5072), .A2(n6180), .ZN(n5684) );
  AOI22_X1 U5725 ( .A1(n5684), .A2(n7546), .B1(n7544), .B2(n5089), .ZN(n5073)
         );
  OAI211_X1 U5726 ( .C1(n5776), .C2(n5368), .A(n5074), .B(n5073), .ZN(U3044)
         );
  AOI22_X1 U5727 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5088), .B1(n5568), 
        .B2(n5087), .ZN(n5076) );
  AOI22_X1 U5728 ( .A1(n5684), .A2(n5801), .B1(n5797), .B2(n5089), .ZN(n5075)
         );
  OAI211_X1 U5729 ( .C1(n5799), .C2(n5368), .A(n5076), .B(n5075), .ZN(U3046)
         );
  AOI22_X1 U5730 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5088), .B1(n5536), 
        .B2(n5087), .ZN(n5078) );
  AOI22_X1 U5731 ( .A1(n5684), .A2(n5819), .B1(n5813), .B2(n5089), .ZN(n5077)
         );
  OAI211_X1 U5732 ( .C1(n5815), .C2(n5368), .A(n5078), .B(n5077), .ZN(U3050)
         );
  AOI22_X1 U5733 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5088), .B1(n5554), 
        .B2(n5087), .ZN(n5080) );
  AOI22_X1 U5734 ( .A1(n5684), .A2(n5789), .B1(n5785), .B2(n5089), .ZN(n5079)
         );
  OAI211_X1 U5735 ( .C1(n5787), .C2(n5368), .A(n5080), .B(n5079), .ZN(U3047)
         );
  AOI22_X1 U5736 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5088), .B1(n5541), 
        .B2(n5087), .ZN(n5082) );
  AOI22_X1 U5737 ( .A1(n5684), .A2(n5808), .B1(n5804), .B2(n5089), .ZN(n5081)
         );
  OAI211_X1 U5738 ( .C1(n5806), .C2(n5368), .A(n5082), .B(n5081), .ZN(U3051)
         );
  AOI22_X1 U5739 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5088), .B1(n7564), 
        .B2(n5087), .ZN(n5084) );
  AOI22_X1 U5740 ( .A1(n5684), .A2(n7570), .B1(n7567), .B2(n5089), .ZN(n5083)
         );
  OAI211_X1 U5741 ( .C1(n5793), .C2(n5368), .A(n5084), .B(n5083), .ZN(U3049)
         );
  AOI22_X1 U5742 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5088), .B1(n7557), 
        .B2(n5087), .ZN(n5086) );
  AOI22_X1 U5743 ( .A1(n5684), .A2(n7560), .B1(n7558), .B2(n5089), .ZN(n5085)
         );
  OAI211_X1 U5744 ( .C1(n5781), .C2(n5368), .A(n5086), .B(n5085), .ZN(U3048)
         );
  AOI22_X1 U5745 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5088), .B1(n7550), 
        .B2(n5087), .ZN(n5091) );
  AOI22_X1 U5746 ( .A1(n5684), .A2(n7553), .B1(n7551), .B2(n5089), .ZN(n5090)
         );
  OAI211_X1 U5747 ( .C1(n5771), .C2(n5368), .A(n5091), .B(n5090), .ZN(U3045)
         );
  NAND2_X1 U5748 ( .A1(n5094), .A2(n5092), .ZN(n5227) );
  NOR2_X1 U5749 ( .A1(n6175), .A2(n5097), .ZN(n5116) );
  AOI21_X1 U5750 ( .B1(n5122), .B2(n5338), .A(n5116), .ZN(n5099) );
  AND2_X1 U5751 ( .A1(n5094), .A2(n5093), .ZN(n5181) );
  NOR2_X1 U5752 ( .A1(n5181), .A2(n5379), .ZN(n5096) );
  AOI22_X1 U5753 ( .A1(n5099), .A2(n5096), .B1(n5379), .B2(n5097), .ZN(n5095)
         );
  NAND2_X1 U5754 ( .A1(n5294), .A2(n5095), .ZN(n5115) );
  INV_X1 U5755 ( .A(n5096), .ZN(n5098) );
  OAI22_X1 U5756 ( .A1(n5099), .A2(n5098), .B1(n5995), .B2(n5097), .ZN(n5114)
         );
  AOI22_X1 U5757 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5115), .B1(n7564), 
        .B2(n5114), .ZN(n5101) );
  AOI22_X1 U5758 ( .A1(n5117), .A2(n7570), .B1(n7567), .B2(n5116), .ZN(n5100)
         );
  OAI211_X1 U5759 ( .C1(n5793), .C2(n5227), .A(n5101), .B(n5100), .ZN(U3129)
         );
  AOI22_X1 U5760 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5115), .B1(n7543), 
        .B2(n5114), .ZN(n5103) );
  AOI22_X1 U5761 ( .A1(n5117), .A2(n7546), .B1(n7544), .B2(n5116), .ZN(n5102)
         );
  OAI211_X1 U5762 ( .C1(n5776), .C2(n5227), .A(n5103), .B(n5102), .ZN(U3124)
         );
  AOI22_X1 U5763 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5115), .B1(n5554), 
        .B2(n5114), .ZN(n5105) );
  AOI22_X1 U5764 ( .A1(n5117), .A2(n5789), .B1(n5785), .B2(n5116), .ZN(n5104)
         );
  OAI211_X1 U5765 ( .C1(n5787), .C2(n5227), .A(n5105), .B(n5104), .ZN(U3127)
         );
  AOI22_X1 U5766 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5115), .B1(n5541), 
        .B2(n5114), .ZN(n5107) );
  AOI22_X1 U5767 ( .A1(n5117), .A2(n5808), .B1(n5804), .B2(n5116), .ZN(n5106)
         );
  OAI211_X1 U5768 ( .C1(n5806), .C2(n5227), .A(n5107), .B(n5106), .ZN(U3131)
         );
  AOI22_X1 U5769 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5115), .B1(n5536), 
        .B2(n5114), .ZN(n5109) );
  AOI22_X1 U5770 ( .A1(n5117), .A2(n5819), .B1(n5813), .B2(n5116), .ZN(n5108)
         );
  OAI211_X1 U5771 ( .C1(n5815), .C2(n5227), .A(n5109), .B(n5108), .ZN(U3130)
         );
  AOI22_X1 U5772 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5115), .B1(n5568), 
        .B2(n5114), .ZN(n5111) );
  AOI22_X1 U5773 ( .A1(n5117), .A2(n5801), .B1(n5797), .B2(n5116), .ZN(n5110)
         );
  OAI211_X1 U5774 ( .C1(n5799), .C2(n5227), .A(n5111), .B(n5110), .ZN(U3126)
         );
  AOI22_X1 U5775 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5115), .B1(n7550), 
        .B2(n5114), .ZN(n5113) );
  AOI22_X1 U5776 ( .A1(n5117), .A2(n7553), .B1(n7551), .B2(n5116), .ZN(n5112)
         );
  OAI211_X1 U5777 ( .C1(n5771), .C2(n5227), .A(n5113), .B(n5112), .ZN(U3125)
         );
  AOI22_X1 U5778 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5115), .B1(n7557), 
        .B2(n5114), .ZN(n5119) );
  AOI22_X1 U5779 ( .A1(n5117), .A2(n7560), .B1(n7558), .B2(n5116), .ZN(n5118)
         );
  OAI211_X1 U5780 ( .C1(n5781), .C2(n5227), .A(n5119), .B(n5118), .ZN(U3128)
         );
  NAND2_X1 U5781 ( .A1(n4890), .A2(n5178), .ZN(n5234) );
  INV_X1 U5782 ( .A(n5234), .ZN(n5120) );
  INV_X1 U5783 ( .A(n5128), .ZN(n5121) );
  NOR3_X1 U5784 ( .A1(n4112), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5465) );
  OAI21_X1 U5785 ( .B1(n5121), .B2(n7502), .A(n5756), .ZN(n5126) );
  INV_X1 U5786 ( .A(n5126), .ZN(n5123) );
  NAND2_X1 U5787 ( .A1(n7246), .A2(n5518), .ZN(n5474) );
  INV_X1 U5788 ( .A(n5474), .ZN(n5468) );
  INV_X1 U5789 ( .A(n5465), .ZN(n5125) );
  NOR2_X1 U5790 ( .A1(n6175), .A2(n5125), .ZN(n5145) );
  AOI21_X1 U5791 ( .B1(n5122), .B2(n5468), .A(n5145), .ZN(n5127) );
  NAND2_X1 U5792 ( .A1(n5123), .A2(n5127), .ZN(n5124) );
  OAI211_X1 U5793 ( .C1(n5756), .C2(n5465), .A(n5294), .B(n5124), .ZN(n5144)
         );
  OAI22_X1 U5794 ( .A1(n5127), .A2(n5126), .B1(n5995), .B2(n5125), .ZN(n5143)
         );
  AOI22_X1 U5795 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5144), .B1(n5568), 
        .B2(n5143), .ZN(n5130) );
  AOI22_X1 U5796 ( .A1(n5818), .A2(n5659), .B1(n5797), .B2(n5145), .ZN(n5129)
         );
  OAI211_X1 U5797 ( .C1(n5662), .C2(n5507), .A(n5130), .B(n5129), .ZN(U3094)
         );
  AOI22_X1 U5798 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5144), .B1(n5554), 
        .B2(n5143), .ZN(n5132) );
  AOI22_X1 U5799 ( .A1(n5818), .A2(n5653), .B1(n5785), .B2(n5145), .ZN(n5131)
         );
  OAI211_X1 U5800 ( .C1(n5656), .C2(n5507), .A(n5132), .B(n5131), .ZN(U3095)
         );
  AOI22_X1 U5801 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5144), .B1(n5541), 
        .B2(n5143), .ZN(n5134) );
  AOI22_X1 U5802 ( .A1(n5818), .A2(n5670), .B1(n5804), .B2(n5145), .ZN(n5133)
         );
  OAI211_X1 U5803 ( .C1(n5673), .C2(n5507), .A(n5134), .B(n5133), .ZN(U3099)
         );
  AOI22_X1 U5804 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5144), .B1(n7550), 
        .B2(n5143), .ZN(n5136) );
  AOI22_X1 U5805 ( .A1(n5818), .A2(n7552), .B1(n7551), .B2(n5145), .ZN(n5135)
         );
  OAI211_X1 U5806 ( .C1(n5667), .C2(n5507), .A(n5136), .B(n5135), .ZN(U3093)
         );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5144), .B1(n7543), 
        .B2(n5143), .ZN(n5138) );
  AOI22_X1 U5808 ( .A1(n5818), .A2(n7545), .B1(n7544), .B2(n5145), .ZN(n5137)
         );
  OAI211_X1 U5809 ( .C1(n5650), .C2(n5507), .A(n5138), .B(n5137), .ZN(U3092)
         );
  AOI22_X1 U5810 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5144), .B1(n7564), 
        .B2(n5143), .ZN(n5140) );
  AOI22_X1 U5811 ( .A1(n5818), .A2(n7568), .B1(n7567), .B2(n5145), .ZN(n5139)
         );
  OAI211_X1 U5812 ( .C1(n5688), .C2(n5507), .A(n5140), .B(n5139), .ZN(U3097)
         );
  AOI22_X1 U5813 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5144), .B1(n5536), 
        .B2(n5143), .ZN(n5142) );
  AOI22_X1 U5814 ( .A1(n5818), .A2(n5642), .B1(n5813), .B2(n5145), .ZN(n5141)
         );
  OAI211_X1 U5815 ( .C1(n5645), .C2(n5507), .A(n5142), .B(n5141), .ZN(U3098)
         );
  AOI22_X1 U5816 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5144), .B1(n7557), 
        .B2(n5143), .ZN(n5147) );
  AOI22_X1 U5817 ( .A1(n5818), .A2(n7559), .B1(n7558), .B2(n5145), .ZN(n5146)
         );
  OAI211_X1 U5818 ( .C1(n5678), .C2(n5507), .A(n5147), .B(n5146), .ZN(U3096)
         );
  MUX2_X1 U5819 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5148), .S(n7456), 
        .Z(n7467) );
  OR2_X1 U5820 ( .A1(n7246), .A2(n5149), .ZN(n5157) );
  XNOR2_X1 U5821 ( .A(n6960), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5154)
         );
  XNOR2_X1 U5822 ( .A(n6963), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5150)
         );
  NAND2_X1 U5823 ( .A1(n6964), .A2(n5150), .ZN(n5151) );
  OAI21_X1 U5824 ( .B1(n5154), .B2(n5152), .A(n5151), .ZN(n5153) );
  AOI21_X1 U5825 ( .B1(n5155), .B2(n5154), .A(n5153), .ZN(n5156) );
  NAND2_X1 U5826 ( .A1(n5157), .A2(n5156), .ZN(n6070) );
  NAND2_X1 U5827 ( .A1(n6070), .A2(n7456), .ZN(n5160) );
  NAND2_X1 U5828 ( .A1(n5158), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U5829 ( .A1(n5160), .A2(n5159), .ZN(n7463) );
  NAND3_X1 U5830 ( .A1(n7467), .A2(n7487), .A3(n7463), .ZN(n5164) );
  NOR2_X1 U5831 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7487), .ZN(n5161) );
  NAND2_X1 U5832 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  AND2_X1 U5833 ( .A1(n5164), .A2(n5163), .ZN(n7452) );
  OR2_X1 U5834 ( .A1(n7452), .A2(n6961), .ZN(n5174) );
  MUX2_X1 U5835 ( .A(n7456), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5172) );
  INV_X1 U5836 ( .A(n5165), .ZN(n5166) );
  OR2_X1 U5837 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  XNOR2_X1 U5838 ( .A(n5168), .B(n5171), .ZN(n7435) );
  OR2_X1 U5839 ( .A1(n7436), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5169) );
  OR2_X1 U5840 ( .A1(n7435), .A2(n5169), .ZN(n5170) );
  OAI21_X1 U5841 ( .B1(n5172), .B2(n5171), .A(n5170), .ZN(n7450) );
  INV_X1 U5842 ( .A(n7450), .ZN(n5173) );
  NAND2_X1 U5843 ( .A1(n5174), .A2(n5173), .ZN(n7490) );
  NOR2_X1 U5844 ( .A1(n7490), .A2(FLUSH_REG_SCAN_IN), .ZN(n5176) );
  OAI21_X1 U5845 ( .B1(n5176), .B2(n7491), .A(n5175), .ZN(n6990) );
  OAI21_X1 U5846 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7487), .A(n6990), .ZN(
        n6183) );
  INV_X1 U5847 ( .A(n6990), .ZN(n6177) );
  NOR2_X1 U5848 ( .A1(n6177), .A2(n5379), .ZN(n6181) );
  OAI21_X1 U5849 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5178), .A(n5177), .ZN(
        n5179) );
  AOI22_X1 U5850 ( .A1(n6181), .A2(n5179), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6177), .ZN(n5180) );
  OAI21_X1 U5851 ( .B1(n5518), .B2(n6183), .A(n5180), .ZN(U3464) );
  INV_X1 U5852 ( .A(n5181), .ZN(n5184) );
  OAI21_X1 U5853 ( .B1(n4890), .B2(n7502), .A(n5233), .ZN(n5183) );
  NAND2_X1 U5854 ( .A1(n5182), .A2(n5187), .ZN(n5298) );
  OR2_X1 U5855 ( .A1(n5298), .A2(n7502), .ZN(n5292) );
  NAND3_X1 U5856 ( .A1(n5184), .A2(n5183), .A3(n5292), .ZN(n5185) );
  AOI22_X1 U5857 ( .A1(n6181), .A2(n5185), .B1(n6177), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5186) );
  OAI21_X1 U5858 ( .B1(n5628), .B2(n6183), .A(n5186), .ZN(U3462) );
  INV_X1 U5859 ( .A(n6181), .ZN(n5190) );
  NAND2_X1 U5860 ( .A1(n5187), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5188) );
  XNOR2_X1 U5861 ( .A(n4890), .B(n5188), .ZN(n5189) );
  OAI222_X1 U5862 ( .A1(n6183), .A2(n7246), .B1(n6990), .B2(n7462), .C1(n5190), 
        .C2(n5189), .ZN(U3463) );
  NAND2_X1 U5863 ( .A1(n5534), .A2(n5756), .ZN(n5526) );
  INV_X1 U5864 ( .A(n5227), .ZN(n5191) );
  AOI21_X1 U5865 ( .B1(n5535), .B2(n5526), .A(n5191), .ZN(n5195) );
  NOR2_X1 U5866 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5192), .ZN(n5225)
         );
  NAND2_X1 U5867 ( .A1(n5534), .A2(n5469), .ZN(n5530) );
  NAND2_X1 U5868 ( .A1(n5529), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U5869 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5758), .ZN(n5767) );
  OAI211_X1 U5870 ( .C1(n4732), .C2(n5225), .A(n5530), .B(n5767), .ZN(n5193)
         );
  AOI211_X2 U5871 ( .C1(n5195), .C2(n5194), .A(n3637), .B(n5193), .ZN(n5232)
         );
  INV_X1 U5872 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5199) );
  OAI22_X1 U5873 ( .A1(n5527), .A2(n5534), .B1(n5758), .B2(n5533), .ZN(n5224)
         );
  AOI22_X1 U5874 ( .A1(n5804), .A2(n5225), .B1(n5541), .B2(n5224), .ZN(n5196)
         );
  OAI21_X1 U5875 ( .B1(n5227), .B2(n5673), .A(n5196), .ZN(n5197) );
  AOI21_X1 U5876 ( .B1(n5229), .B2(n5670), .A(n5197), .ZN(n5198) );
  OAI21_X1 U5877 ( .B1(n5232), .B2(n5199), .A(n5198), .ZN(U3139) );
  INV_X1 U5878 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5203) );
  AOI22_X1 U5879 ( .A1(n7558), .A2(n5225), .B1(n7557), .B2(n5224), .ZN(n5200)
         );
  OAI21_X1 U5880 ( .B1(n5227), .B2(n5678), .A(n5200), .ZN(n5201) );
  AOI21_X1 U5881 ( .B1(n5229), .B2(n7559), .A(n5201), .ZN(n5202) );
  OAI21_X1 U5882 ( .B1(n5232), .B2(n5203), .A(n5202), .ZN(U3136) );
  INV_X1 U5883 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5207) );
  AOI22_X1 U5884 ( .A1(n5797), .A2(n5225), .B1(n5568), .B2(n5224), .ZN(n5204)
         );
  OAI21_X1 U5885 ( .B1(n5227), .B2(n5662), .A(n5204), .ZN(n5205) );
  AOI21_X1 U5886 ( .B1(n5229), .B2(n5659), .A(n5205), .ZN(n5206) );
  OAI21_X1 U5887 ( .B1(n5232), .B2(n5207), .A(n5206), .ZN(U3134) );
  INV_X1 U5888 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5211) );
  AOI22_X1 U5889 ( .A1(n7567), .A2(n5225), .B1(n7564), .B2(n5224), .ZN(n5208)
         );
  OAI21_X1 U5890 ( .B1(n5227), .B2(n5688), .A(n5208), .ZN(n5209) );
  AOI21_X1 U5891 ( .B1(n5229), .B2(n7568), .A(n5209), .ZN(n5210) );
  OAI21_X1 U5892 ( .B1(n5232), .B2(n5211), .A(n5210), .ZN(U3137) );
  INV_X1 U5893 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5215) );
  AOI22_X1 U5894 ( .A1(n7551), .A2(n5225), .B1(n7550), .B2(n5224), .ZN(n5212)
         );
  OAI21_X1 U5895 ( .B1(n5227), .B2(n5667), .A(n5212), .ZN(n5213) );
  AOI21_X1 U5896 ( .B1(n5229), .B2(n7552), .A(n5213), .ZN(n5214) );
  OAI21_X1 U5897 ( .B1(n5232), .B2(n5215), .A(n5214), .ZN(U3133) );
  INV_X1 U5898 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5219) );
  AOI22_X1 U5899 ( .A1(n5785), .A2(n5225), .B1(n5554), .B2(n5224), .ZN(n5216)
         );
  OAI21_X1 U5900 ( .B1(n5227), .B2(n5656), .A(n5216), .ZN(n5217) );
  AOI21_X1 U5901 ( .B1(n5229), .B2(n5653), .A(n5217), .ZN(n5218) );
  OAI21_X1 U5902 ( .B1(n5232), .B2(n5219), .A(n5218), .ZN(U3135) );
  INV_X1 U5903 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5223) );
  AOI22_X1 U5904 ( .A1(n7544), .A2(n5225), .B1(n7543), .B2(n5224), .ZN(n5220)
         );
  OAI21_X1 U5905 ( .B1(n5227), .B2(n5650), .A(n5220), .ZN(n5221) );
  AOI21_X1 U5906 ( .B1(n5229), .B2(n7545), .A(n5221), .ZN(n5222) );
  OAI21_X1 U5907 ( .B1(n5232), .B2(n5223), .A(n5222), .ZN(U3132) );
  INV_X1 U5908 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5231) );
  AOI22_X1 U5909 ( .A1(n5813), .A2(n5225), .B1(n5536), .B2(n5224), .ZN(n5226)
         );
  OAI21_X1 U5910 ( .B1(n5227), .B2(n5645), .A(n5226), .ZN(n5228) );
  AOI21_X1 U5911 ( .B1(n5229), .B2(n5642), .A(n5228), .ZN(n5230) );
  OAI21_X1 U5912 ( .B1(n5232), .B2(n5231), .A(n5230), .ZN(U3138) );
  NOR2_X2 U5913 ( .A1(n5369), .A2(n6180), .ZN(n7569) );
  OAI21_X1 U5914 ( .B1(n7571), .B2(n7569), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5237) );
  NAND2_X1 U5915 ( .A1(n5474), .A2(n5756), .ZN(n5463) );
  NAND2_X1 U5916 ( .A1(n5527), .A2(n5463), .ZN(n5236) );
  NOR3_X1 U5917 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n5370), .ZN(n7566) );
  AND2_X1 U5918 ( .A1(n5533), .A2(n5376), .ZN(n5769) );
  OAI21_X1 U5919 ( .B1(n5529), .B2(n5336), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n5332) );
  OAI211_X1 U5920 ( .C1(n7566), .C2(n4732), .A(n5769), .B(n5332), .ZN(n5235)
         );
  AOI21_X1 U5921 ( .B1(n5237), .B2(n5236), .A(n5235), .ZN(n7575) );
  INV_X1 U5922 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5245) );
  INV_X1 U5923 ( .A(n7566), .ZN(n5254) );
  OR2_X1 U5924 ( .A1(n5535), .A2(n5474), .ZN(n5241) );
  INV_X1 U5925 ( .A(n5475), .ZN(n5760) );
  INV_X1 U5926 ( .A(n5336), .ZN(n5239) );
  NAND3_X1 U5927 ( .A1(n5760), .A2(n5239), .A3(n5238), .ZN(n5240) );
  AND2_X1 U5928 ( .A1(n5241), .A2(n5240), .ZN(n7542) );
  OAI22_X1 U5929 ( .A1(n5668), .A2(n5254), .B1(n7542), .B2(n5810), .ZN(n5242)
         );
  AOI21_X1 U5930 ( .B1(n7571), .B2(n5808), .A(n5242), .ZN(n5244) );
  NAND2_X1 U5931 ( .A1(n7569), .A2(n5670), .ZN(n5243) );
  OAI211_X1 U5932 ( .C1(n7575), .C2(n5245), .A(n5244), .B(n5243), .ZN(U3027)
         );
  INV_X1 U5933 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5249) );
  OAI22_X1 U5934 ( .A1(n5651), .A2(n5254), .B1(n7542), .B2(n5791), .ZN(n5246)
         );
  AOI21_X1 U5935 ( .B1(n7571), .B2(n5789), .A(n5246), .ZN(n5248) );
  NAND2_X1 U5936 ( .A1(n7569), .A2(n5653), .ZN(n5247) );
  OAI211_X1 U5937 ( .C1(n7575), .C2(n5249), .A(n5248), .B(n5247), .ZN(U3023)
         );
  INV_X1 U5938 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5253) );
  OAI22_X1 U5939 ( .A1(n5657), .A2(n5254), .B1(n7542), .B2(n5803), .ZN(n5250)
         );
  AOI21_X1 U5940 ( .B1(n7571), .B2(n5801), .A(n5250), .ZN(n5252) );
  NAND2_X1 U5941 ( .A1(n7569), .A2(n5659), .ZN(n5251) );
  OAI211_X1 U5942 ( .C1(n7575), .C2(n5253), .A(n5252), .B(n5251), .ZN(U3022)
         );
  INV_X1 U5943 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5258) );
  OAI22_X1 U5944 ( .A1(n5640), .A2(n5254), .B1(n7542), .B2(n5821), .ZN(n5255)
         );
  AOI21_X1 U5945 ( .B1(n7571), .B2(n5819), .A(n5255), .ZN(n5257) );
  NAND2_X1 U5946 ( .A1(n7569), .A2(n5642), .ZN(n5256) );
  OAI211_X1 U5947 ( .C1(n7575), .C2(n5258), .A(n5257), .B(n5256), .ZN(U3026)
         );
  NAND2_X1 U5948 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  XNOR2_X1 U5949 ( .A(n5262), .B(n5261), .ZN(n7133) );
  INV_X1 U5950 ( .A(n7133), .ZN(n5276) );
  OR2_X1 U5951 ( .A1(n6029), .A2(n7197), .ZN(n7175) );
  AOI21_X1 U5952 ( .B1(n5264), .B2(n7175), .A(n5263), .ZN(n7192) );
  OR2_X1 U5953 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5423), .ZN(n7188)
         );
  INV_X1 U5954 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5422) );
  AOI21_X1 U5955 ( .B1(n7192), .B2(n7188), .A(n5422), .ZN(n5274) );
  INV_X1 U5956 ( .A(n5264), .ZN(n5424) );
  NAND2_X1 U5957 ( .A1(n5424), .A2(n7193), .ZN(n7187) );
  OR2_X1 U5958 ( .A1(n4001), .A2(n7187), .ZN(n5421) );
  NOR3_X1 U5959 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5423), .A3(n5421), 
        .ZN(n5273) );
  MUX2_X1 U5960 ( .A(n5947), .B(n5948), .S(EBX_REG_6__SCAN_IN), .Z(n5267) );
  NAND2_X1 U5961 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5962), .ZN(n5265)
         );
  AND2_X1 U5962 ( .A1(n5939), .A2(n5265), .ZN(n5266) );
  NAND2_X1 U5963 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  OR2_X1 U5964 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  NAND2_X1 U5965 ( .A1(n5326), .A2(n5270), .ZN(n7285) );
  INV_X1 U5966 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5271) );
  OAI22_X1 U5967 ( .A1(n7215), .A2(n7285), .B1(n7213), .B2(n5271), .ZN(n5272)
         );
  NOR3_X1 U5968 ( .A1(n5274), .A2(n5273), .A3(n5272), .ZN(n5275) );
  OAI21_X1 U5969 ( .B1(n5276), .B2(n6584), .A(n5275), .ZN(U3012) );
  INV_X1 U5970 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5278) );
  OAI21_X1 U5971 ( .B1(n7132), .B2(n5278), .A(n5277), .ZN(n5280) );
  NOR2_X1 U5972 ( .A1(n7266), .A2(n6489), .ZN(n5279) );
  AOI211_X1 U5973 ( .C1(n7143), .C2(n7263), .A(n5280), .B(n5279), .ZN(n5281)
         );
  OAI21_X1 U5974 ( .B1(n5282), .B2(n7433), .A(n5281), .ZN(U2982) );
  NOR2_X1 U5975 ( .A1(n5283), .A2(n5284), .ZN(n5622) );
  AOI21_X1 U5976 ( .B1(n5284), .B2(n5283), .A(n5622), .ZN(n7290) );
  INV_X1 U5977 ( .A(n7290), .ZN(n5286) );
  INV_X1 U5978 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5285) );
  OAI222_X1 U5979 ( .A1(n5286), .A2(n6357), .B1(n5285), .B2(n7118), .C1(n7105), 
        .C2(n7285), .ZN(U2853) );
  OAI222_X1 U5980 ( .A1(n5287), .A2(n6394), .B1(n6392), .B2(n4699), .C1(n6391), 
        .C2(n5286), .ZN(U2885) );
  INV_X1 U5981 ( .A(n5289), .ZN(n5315) );
  AOI21_X1 U5982 ( .B1(n5291), .B2(n5290), .A(n5315), .ZN(n5297) );
  NAND3_X1 U5983 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4112), .ZN(n5528) );
  AOI22_X1 U5984 ( .A1(n5297), .A2(n5295), .B1(n5379), .B2(n5528), .ZN(n5293)
         );
  NAND2_X1 U5985 ( .A1(n5294), .A2(n5293), .ZN(n5314) );
  INV_X1 U5986 ( .A(n5295), .ZN(n5296) );
  OAI22_X1 U5987 ( .A1(n5297), .A2(n5296), .B1(n5995), .B2(n5528), .ZN(n5313)
         );
  AOI22_X1 U5988 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5314), .B1(n7550), 
        .B2(n5313), .ZN(n5300) );
  NOR2_X2 U5989 ( .A1(n5298), .A2(n6180), .ZN(n5573) );
  AOI22_X1 U5990 ( .A1(n5573), .A2(n7553), .B1(n5315), .B2(n7551), .ZN(n5299)
         );
  OAI211_X1 U5991 ( .C1(n5771), .C2(n5511), .A(n5300), .B(n5299), .ZN(U3077)
         );
  AOI22_X1 U5992 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5314), .B1(n5568), 
        .B2(n5313), .ZN(n5302) );
  AOI22_X1 U5993 ( .A1(n5573), .A2(n5801), .B1(n5315), .B2(n5797), .ZN(n5301)
         );
  OAI211_X1 U5994 ( .C1(n5799), .C2(n5511), .A(n5302), .B(n5301), .ZN(U3078)
         );
  AOI22_X1 U5995 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5314), .B1(n5554), 
        .B2(n5313), .ZN(n5304) );
  AOI22_X1 U5996 ( .A1(n5573), .A2(n5789), .B1(n5315), .B2(n5785), .ZN(n5303)
         );
  OAI211_X1 U5997 ( .C1(n5787), .C2(n5511), .A(n5304), .B(n5303), .ZN(U3079)
         );
  AOI22_X1 U5998 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5314), .B1(n7543), 
        .B2(n5313), .ZN(n5306) );
  AOI22_X1 U5999 ( .A1(n5573), .A2(n7546), .B1(n5315), .B2(n7544), .ZN(n5305)
         );
  OAI211_X1 U6000 ( .C1(n5776), .C2(n5511), .A(n5306), .B(n5305), .ZN(U3076)
         );
  AOI22_X1 U6001 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5314), .B1(n7564), 
        .B2(n5313), .ZN(n5308) );
  AOI22_X1 U6002 ( .A1(n5573), .A2(n7570), .B1(n5315), .B2(n7567), .ZN(n5307)
         );
  OAI211_X1 U6003 ( .C1(n5793), .C2(n5511), .A(n5308), .B(n5307), .ZN(U3081)
         );
  AOI22_X1 U6004 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5314), .B1(n5536), 
        .B2(n5313), .ZN(n5310) );
  AOI22_X1 U6005 ( .A1(n5573), .A2(n5819), .B1(n5315), .B2(n5813), .ZN(n5309)
         );
  OAI211_X1 U6006 ( .C1(n5815), .C2(n5511), .A(n5310), .B(n5309), .ZN(U3082)
         );
  AOI22_X1 U6007 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5314), .B1(n5541), 
        .B2(n5313), .ZN(n5312) );
  AOI22_X1 U6008 ( .A1(n5573), .A2(n5808), .B1(n5315), .B2(n5804), .ZN(n5311)
         );
  OAI211_X1 U6009 ( .C1(n5806), .C2(n5511), .A(n5312), .B(n5311), .ZN(U3083)
         );
  AOI22_X1 U6010 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5314), .B1(n7557), 
        .B2(n5313), .ZN(n5317) );
  AOI22_X1 U6011 ( .A1(n5573), .A2(n7560), .B1(n5315), .B2(n7558), .ZN(n5316)
         );
  OAI211_X1 U6012 ( .C1(n5781), .C2(n5511), .A(n5317), .B(n5316), .ZN(U3080)
         );
  OR2_X1 U6013 ( .A1(n5625), .A2(n5318), .ZN(n5319) );
  AND2_X1 U6014 ( .A1(n5319), .A2(n5578), .ZN(n5618) );
  INV_X1 U6015 ( .A(n5618), .ZN(n5412) );
  INV_X1 U6016 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5328) );
  INV_X1 U6017 ( .A(n4770), .ZN(n5948) );
  MUX2_X1 U6018 ( .A(n5947), .B(n5948), .S(EBX_REG_8__SCAN_IN), .Z(n5321) );
  NAND2_X1 U6019 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n5962), .ZN(n5320)
         );
  AND3_X1 U6020 ( .A1(n5321), .A2(n5939), .A3(n5320), .ZN(n5327) );
  NAND2_X1 U6021 ( .A1(n5322), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5323)
         );
  OAI211_X1 U6022 ( .C1(n5962), .C2(EBX_REG_7__SCAN_IN), .A(n5948), .B(n5323), 
        .ZN(n5324) );
  OAI21_X1 U6023 ( .B1(n5956), .B2(EBX_REG_7__SCAN_IN), .A(n5324), .ZN(n7099)
         );
  OR2_X1 U6024 ( .A1(n5326), .A2(n7099), .ZN(n7101) );
  AOI21_X1 U6025 ( .B1(n5327), .B2(n7101), .A(n5584), .ZN(n5432) );
  INV_X1 U6026 ( .A(n5432), .ZN(n5615) );
  OAI222_X1 U6027 ( .A1(n5412), .A2(n6357), .B1(n7118), .B2(n5328), .C1(n5615), 
        .C2(n7105), .ZN(U2851) );
  INV_X1 U6028 ( .A(n5368), .ZN(n5329) );
  AOI211_X1 U6029 ( .C1(n5527), .C2(n5330), .A(n5365), .B(n5329), .ZN(n5335)
         );
  NOR2_X1 U6030 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5331), .ZN(n5339)
         );
  OAI211_X1 U6031 ( .C1(n4732), .C2(n5339), .A(n5333), .B(n5332), .ZN(n5334)
         );
  NAND2_X1 U6032 ( .A1(n5361), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5342) );
  INV_X1 U6033 ( .A(n5535), .ZN(n5638) );
  NOR3_X1 U6034 ( .A1(n5336), .A2(n5533), .A3(n5529), .ZN(n5337) );
  AOI21_X1 U6035 ( .B1(n5638), .B2(n5338), .A(n5337), .ZN(n5363) );
  INV_X1 U6036 ( .A(n5339), .ZN(n5362) );
  OAI22_X1 U6037 ( .A1(n5363), .A2(n5821), .B1(n5640), .B2(n5362), .ZN(n5340)
         );
  AOI21_X1 U6038 ( .B1(n5642), .B2(n5365), .A(n5340), .ZN(n5341) );
  OAI211_X1 U6039 ( .C1(n5368), .C2(n5645), .A(n5342), .B(n5341), .ZN(U3058)
         );
  NAND2_X1 U6040 ( .A1(n5361), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5345) );
  OAI22_X1 U6041 ( .A1(n5363), .A2(n5784), .B1(n5674), .B2(n5362), .ZN(n5343)
         );
  AOI21_X1 U6042 ( .B1(n7559), .B2(n5365), .A(n5343), .ZN(n5344) );
  OAI211_X1 U6043 ( .C1(n5368), .C2(n5678), .A(n5345), .B(n5344), .ZN(U3056)
         );
  NAND2_X1 U6044 ( .A1(n5361), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5348) );
  OAI22_X1 U6045 ( .A1(n5363), .A2(n5803), .B1(n5657), .B2(n5362), .ZN(n5346)
         );
  AOI21_X1 U6046 ( .B1(n5659), .B2(n5365), .A(n5346), .ZN(n5347) );
  OAI211_X1 U6047 ( .C1(n5368), .C2(n5662), .A(n5348), .B(n5347), .ZN(U3054)
         );
  NAND2_X1 U6048 ( .A1(n5361), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5351) );
  OAI22_X1 U6049 ( .A1(n5363), .A2(n5791), .B1(n5651), .B2(n5362), .ZN(n5349)
         );
  AOI21_X1 U6050 ( .B1(n5653), .B2(n5365), .A(n5349), .ZN(n5350) );
  OAI211_X1 U6051 ( .C1(n5368), .C2(n5656), .A(n5351), .B(n5350), .ZN(U3055)
         );
  NAND2_X1 U6052 ( .A1(n5361), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5354) );
  OAI22_X1 U6053 ( .A1(n5363), .A2(n5779), .B1(n5646), .B2(n5362), .ZN(n5352)
         );
  AOI21_X1 U6054 ( .B1(n7545), .B2(n5365), .A(n5352), .ZN(n5353) );
  OAI211_X1 U6055 ( .C1(n5368), .C2(n5650), .A(n5354), .B(n5353), .ZN(U3052)
         );
  NAND2_X1 U6056 ( .A1(n5361), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5357) );
  OAI22_X1 U6057 ( .A1(n5363), .A2(n5796), .B1(n5681), .B2(n5362), .ZN(n5355)
         );
  AOI21_X1 U6058 ( .B1(n7568), .B2(n5365), .A(n5355), .ZN(n5356) );
  OAI211_X1 U6059 ( .C1(n5368), .C2(n5688), .A(n5357), .B(n5356), .ZN(U3057)
         );
  NAND2_X1 U6060 ( .A1(n5361), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5360) );
  OAI22_X1 U6061 ( .A1(n5363), .A2(n5810), .B1(n5668), .B2(n5362), .ZN(n5358)
         );
  AOI21_X1 U6062 ( .B1(n5670), .B2(n5365), .A(n5358), .ZN(n5359) );
  OAI211_X1 U6063 ( .C1(n5368), .C2(n5673), .A(n5360), .B(n5359), .ZN(U3059)
         );
  NAND2_X1 U6064 ( .A1(n5361), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5367) );
  OAI22_X1 U6065 ( .A1(n5363), .A2(n5774), .B1(n5663), .B2(n5362), .ZN(n5364)
         );
  AOI21_X1 U6066 ( .B1(n7552), .B2(n5365), .A(n5364), .ZN(n5366) );
  OAI211_X1 U6067 ( .C1(n5368), .C2(n5667), .A(n5367), .B(n5366), .ZN(U3053)
         );
  NOR3_X1 U6068 ( .A1(n6175), .A2(n5370), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5378) );
  OR2_X1 U6069 ( .A1(n5371), .A2(n5474), .ZN(n5380) );
  INV_X1 U6070 ( .A(n5380), .ZN(n5372) );
  AOI21_X1 U6071 ( .B1(n5373), .B2(STATEBS16_REG_SCAN_IN), .A(n5372), .ZN(
        n5375) );
  NAND2_X1 U6072 ( .A1(n5382), .A2(n5381), .ZN(n5374) );
  AOI221_X1 U6073 ( .B1(n5375), .B2(n5995), .C1(n5374), .C2(
        STATE2_REG_2__SCAN_IN), .A(STATE2_REG_3__SCAN_IN), .ZN(n5377) );
  OAI21_X1 U6074 ( .B1(n5378), .B2(n5377), .A(n5376), .ZN(n5406) );
  NAND2_X1 U6075 ( .A1(n5406), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5387) );
  INV_X1 U6076 ( .A(n5378), .ZN(n5407) );
  AOI21_X1 U6077 ( .B1(n5380), .B2(n5407), .A(n5379), .ZN(n5384) );
  AND3_X1 U6078 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5382), .A3(n5381), .ZN(
        n5383) );
  NOR2_X1 U6079 ( .A1(n5384), .A2(n5383), .ZN(n5408) );
  OAI22_X1 U6080 ( .A1(n5408), .A2(n5821), .B1(n5407), .B2(n5640), .ZN(n5385)
         );
  AOI21_X1 U6081 ( .B1(n7569), .B2(n5819), .A(n5385), .ZN(n5386) );
  OAI211_X1 U6082 ( .C1(n5687), .C2(n5815), .A(n5387), .B(n5386), .ZN(U3034)
         );
  NAND2_X1 U6083 ( .A1(n5406), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5390) );
  OAI22_X1 U6084 ( .A1(n5408), .A2(n5784), .B1(n5407), .B2(n5674), .ZN(n5388)
         );
  AOI21_X1 U6085 ( .B1(n7569), .B2(n7560), .A(n5388), .ZN(n5389) );
  OAI211_X1 U6086 ( .C1(n5687), .C2(n5781), .A(n5390), .B(n5389), .ZN(U3032)
         );
  NAND2_X1 U6087 ( .A1(n5406), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5393) );
  OAI22_X1 U6088 ( .A1(n5408), .A2(n5791), .B1(n5407), .B2(n5651), .ZN(n5391)
         );
  AOI21_X1 U6089 ( .B1(n7569), .B2(n5789), .A(n5391), .ZN(n5392) );
  OAI211_X1 U6090 ( .C1(n5687), .C2(n5787), .A(n5393), .B(n5392), .ZN(U3031)
         );
  NAND2_X1 U6091 ( .A1(n5406), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5396) );
  OAI22_X1 U6092 ( .A1(n5408), .A2(n5796), .B1(n5407), .B2(n5681), .ZN(n5394)
         );
  AOI21_X1 U6093 ( .B1(n7569), .B2(n7570), .A(n5394), .ZN(n5395) );
  OAI211_X1 U6094 ( .C1(n5687), .C2(n5793), .A(n5396), .B(n5395), .ZN(U3033)
         );
  NAND2_X1 U6095 ( .A1(n5406), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5399) );
  OAI22_X1 U6096 ( .A1(n5408), .A2(n5774), .B1(n5407), .B2(n5663), .ZN(n5397)
         );
  AOI21_X1 U6097 ( .B1(n7569), .B2(n7553), .A(n5397), .ZN(n5398) );
  OAI211_X1 U6098 ( .C1(n5687), .C2(n5771), .A(n5399), .B(n5398), .ZN(U3029)
         );
  NAND2_X1 U6099 ( .A1(n5406), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5402) );
  OAI22_X1 U6100 ( .A1(n5408), .A2(n5779), .B1(n5646), .B2(n5407), .ZN(n5400)
         );
  AOI21_X1 U6101 ( .B1(n7546), .B2(n7569), .A(n5400), .ZN(n5401) );
  OAI211_X1 U6102 ( .C1(n5776), .C2(n5687), .A(n5402), .B(n5401), .ZN(U3028)
         );
  NAND2_X1 U6103 ( .A1(n5406), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5405) );
  OAI22_X1 U6104 ( .A1(n5408), .A2(n5803), .B1(n5407), .B2(n5657), .ZN(n5403)
         );
  AOI21_X1 U6105 ( .B1(n7569), .B2(n5801), .A(n5403), .ZN(n5404) );
  OAI211_X1 U6106 ( .C1(n5687), .C2(n5799), .A(n5405), .B(n5404), .ZN(U3030)
         );
  NAND2_X1 U6107 ( .A1(n5406), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5411) );
  OAI22_X1 U6108 ( .A1(n5408), .A2(n5810), .B1(n5407), .B2(n5668), .ZN(n5409)
         );
  AOI21_X1 U6109 ( .B1(n7569), .B2(n5808), .A(n5409), .ZN(n5410) );
  OAI211_X1 U6110 ( .C1(n5687), .C2(n5806), .A(n5411), .B(n5410), .ZN(U3035)
         );
  INV_X1 U6111 ( .A(DATAI_8_), .ZN(n5413) );
  INV_X1 U6112 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7009) );
  OAI222_X1 U6113 ( .A1(n6394), .A2(n5413), .B1(n6392), .B2(n7009), .C1(n6391), 
        .C2(n5412), .ZN(U2883) );
  OAI21_X1 U6114 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n5434) );
  NAND2_X1 U6115 ( .A1(n7147), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5417)
         );
  NAND2_X1 U6116 ( .A1(n7205), .A2(REIP_REG_8__SCAN_IN), .ZN(n5420) );
  OAI211_X1 U6117 ( .C1(n7152), .C2(n5612), .A(n5417), .B(n5420), .ZN(n5418)
         );
  AOI21_X1 U6118 ( .B1(n5618), .B2(n3628), .A(n5418), .ZN(n5419) );
  OAI21_X1 U6119 ( .B1(n5434), .B2(n7433), .A(n5419), .ZN(U2978) );
  INV_X1 U6120 ( .A(n5420), .ZN(n5431) );
  NOR2_X1 U6121 ( .A1(n5428), .A2(n7209), .ZN(n7220) );
  NOR2_X1 U6122 ( .A1(n5422), .A2(n5421), .ZN(n5426) );
  INV_X1 U6123 ( .A(n5426), .ZN(n5835) );
  NOR2_X1 U6124 ( .A1(n5423), .A2(n5835), .ZN(n7210) );
  OAI21_X1 U6125 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n7210), .ZN(n5429) );
  NAND4_X1 U6126 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n5425), .A4(n5424), .ZN(n5834) );
  NOR2_X1 U6127 ( .A1(n5426), .A2(n6036), .ZN(n5427) );
  AOI211_X1 U6128 ( .C1(n6029), .C2(n5834), .A(n5427), .B(n5839), .ZN(n7218)
         );
  OAI22_X1 U6129 ( .A1(n7220), .A2(n5429), .B1(n7218), .B2(n5428), .ZN(n5430)
         );
  AOI211_X1 U6130 ( .C1(n7238), .C2(n5432), .A(n5431), .B(n5430), .ZN(n5433)
         );
  OAI21_X1 U6131 ( .B1(n5434), .B2(n6584), .A(n5433), .ZN(U3010) );
  NAND3_X1 U6132 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n7495), .ZN(n7488) );
  NAND2_X1 U6133 ( .A1(n6001), .A2(n5435), .ZN(n7485) );
  NAND3_X1 U6134 ( .A1(n7213), .A2(n7488), .A3(n7485), .ZN(n5436) );
  NAND2_X1 U6135 ( .A1(n7390), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5450) );
  INV_X1 U6136 ( .A(n5450), .ZN(n5458) );
  NAND2_X1 U6137 ( .A1(n5458), .A2(n5437), .ZN(n5441) );
  INV_X1 U6138 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6401) );
  INV_X1 U6139 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U6140 ( .A(n5439), .B(n5438), .ZN(n6066) );
  NOR2_X1 U6141 ( .A1(n6066), .A2(n7487), .ZN(n5440) );
  NAND2_X1 U6142 ( .A1(n5441), .A2(n7396), .ZN(n7278) );
  INV_X1 U6143 ( .A(n7278), .ZN(n7265) );
  NAND2_X1 U6144 ( .A1(n5458), .A2(n5442), .ZN(n7261) );
  NOR2_X1 U6145 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5451) );
  INV_X1 U6146 ( .A(n5451), .ZN(n5455) );
  OR2_X1 U6147 ( .A1(n7159), .A2(n5455), .ZN(n7476) );
  AND2_X1 U6148 ( .A1(n3634), .A2(n7476), .ZN(n6013) );
  NOR2_X1 U6149 ( .A1(n5451), .A2(EBX_REG_31__SCAN_IN), .ZN(n5443) );
  AND2_X1 U6150 ( .A1(n5454), .A2(n5443), .ZN(n5444) );
  NOR2_X1 U6151 ( .A1(n6013), .A2(n5444), .ZN(n5445) );
  NOR2_X2 U6152 ( .A1(n5450), .A2(n5445), .ZN(n7403) );
  NAND2_X1 U6153 ( .A1(n7403), .A2(EBX_REG_0__SCAN_IN), .ZN(n5448) );
  AND2_X1 U6154 ( .A1(n6066), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5446) );
  OAI21_X1 U6155 ( .B1(n7424), .B2(n7426), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5447) );
  OAI211_X1 U6156 ( .C1(n7261), .C2(n6184), .A(n5448), .B(n5447), .ZN(n5449)
         );
  INV_X1 U6157 ( .A(n5449), .ZN(n5461) );
  INV_X1 U6158 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5967) );
  NOR2_X1 U6159 ( .A1(n5450), .A2(n5967), .ZN(n6014) );
  NOR2_X1 U6160 ( .A1(n5962), .A2(n5451), .ZN(n5452) );
  NAND2_X1 U6161 ( .A1(n3632), .A2(n5453), .ZN(n5456) );
  AOI21_X1 U6162 ( .B1(n5962), .B2(n5456), .A(n5455), .ZN(n5457) );
  NAND2_X1 U6163 ( .A1(n7415), .A2(n7390), .ZN(n7358) );
  AOI22_X1 U6164 ( .A1(n7409), .A2(n5459), .B1(n7358), .B2(REIP_REG_0__SCAN_IN), .ZN(n5460) );
  OAI211_X1 U6165 ( .C1(n5462), .C2(n7265), .A(n5461), .B(n5460), .ZN(U2827)
         );
  INV_X1 U6166 ( .A(n5463), .ZN(n5464) );
  OAI211_X1 U6167 ( .C1(n5638), .C2(n5464), .A(n5507), .B(n5511), .ZN(n5472)
         );
  NAND2_X1 U6168 ( .A1(n6175), .A2(n5465), .ZN(n5473) );
  INV_X1 U6169 ( .A(n5466), .ZN(n5467) );
  AOI21_X1 U6170 ( .B1(n5473), .B2(STATE2_REG_3__SCAN_IN), .A(n5467), .ZN(
        n5471) );
  NAND2_X1 U6171 ( .A1(n5474), .A2(n5469), .ZN(n5470) );
  NAND4_X1 U6172 ( .A1(n5472), .A2(n5769), .A3(n5471), .A4(n5470), .ZN(n5514)
         );
  NOR2_X1 U6173 ( .A1(n5507), .A2(n5793), .ZN(n5481) );
  INV_X1 U6174 ( .A(n5473), .ZN(n5509) );
  OR2_X1 U6175 ( .A1(n5527), .A2(n5474), .ZN(n5478) );
  OR2_X1 U6176 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  NAND2_X1 U6177 ( .A1(n5478), .A2(n5477), .ZN(n5508) );
  AOI22_X1 U6178 ( .A1(n7567), .A2(n5509), .B1(n7564), .B2(n5508), .ZN(n5479)
         );
  OAI21_X1 U6179 ( .B1(n5511), .B2(n5688), .A(n5479), .ZN(n5480) );
  AOI211_X1 U6180 ( .C1(INSTQUEUE_REG_8__5__SCAN_IN), .C2(n5514), .A(n5481), 
        .B(n5480), .ZN(n5482) );
  INV_X1 U6181 ( .A(n5482), .ZN(U3089) );
  NOR2_X1 U6182 ( .A1(n5507), .A2(n5776), .ZN(n5485) );
  AOI22_X1 U6183 ( .A1(n7544), .A2(n5509), .B1(n7543), .B2(n5508), .ZN(n5483)
         );
  OAI21_X1 U6184 ( .B1(n5511), .B2(n5650), .A(n5483), .ZN(n5484) );
  AOI211_X1 U6185 ( .C1(INSTQUEUE_REG_8__0__SCAN_IN), .C2(n5514), .A(n5485), 
        .B(n5484), .ZN(n5486) );
  INV_X1 U6186 ( .A(n5486), .ZN(U3084) );
  NOR2_X1 U6187 ( .A1(n5507), .A2(n5781), .ZN(n5489) );
  AOI22_X1 U6188 ( .A1(n7558), .A2(n5509), .B1(n7557), .B2(n5508), .ZN(n5487)
         );
  OAI21_X1 U6189 ( .B1(n5511), .B2(n5678), .A(n5487), .ZN(n5488) );
  AOI211_X1 U6190 ( .C1(INSTQUEUE_REG_8__4__SCAN_IN), .C2(n5514), .A(n5489), 
        .B(n5488), .ZN(n5490) );
  INV_X1 U6191 ( .A(n5490), .ZN(U3088) );
  NOR2_X1 U6192 ( .A1(n5507), .A2(n5806), .ZN(n5493) );
  AOI22_X1 U6193 ( .A1(n5804), .A2(n5509), .B1(n5541), .B2(n5508), .ZN(n5491)
         );
  OAI21_X1 U6194 ( .B1(n5511), .B2(n5673), .A(n5491), .ZN(n5492) );
  AOI211_X1 U6195 ( .C1(INSTQUEUE_REG_8__7__SCAN_IN), .C2(n5514), .A(n5493), 
        .B(n5492), .ZN(n5494) );
  INV_X1 U6196 ( .A(n5494), .ZN(U3091) );
  NOR2_X1 U6197 ( .A1(n5507), .A2(n5815), .ZN(n5497) );
  AOI22_X1 U6198 ( .A1(n5813), .A2(n5509), .B1(n5536), .B2(n5508), .ZN(n5495)
         );
  OAI21_X1 U6199 ( .B1(n5511), .B2(n5645), .A(n5495), .ZN(n5496) );
  AOI211_X1 U6200 ( .C1(INSTQUEUE_REG_8__6__SCAN_IN), .C2(n5514), .A(n5497), 
        .B(n5496), .ZN(n5498) );
  INV_X1 U6201 ( .A(n5498), .ZN(U3090) );
  NOR2_X1 U6202 ( .A1(n5507), .A2(n5787), .ZN(n5501) );
  AOI22_X1 U6203 ( .A1(n5785), .A2(n5509), .B1(n5554), .B2(n5508), .ZN(n5499)
         );
  OAI21_X1 U6204 ( .B1(n5511), .B2(n5656), .A(n5499), .ZN(n5500) );
  AOI211_X1 U6205 ( .C1(INSTQUEUE_REG_8__3__SCAN_IN), .C2(n5514), .A(n5501), 
        .B(n5500), .ZN(n5502) );
  INV_X1 U6206 ( .A(n5502), .ZN(U3087) );
  NOR2_X1 U6207 ( .A1(n5507), .A2(n5799), .ZN(n5505) );
  AOI22_X1 U6208 ( .A1(n5797), .A2(n5509), .B1(n5568), .B2(n5508), .ZN(n5503)
         );
  OAI21_X1 U6209 ( .B1(n5511), .B2(n5662), .A(n5503), .ZN(n5504) );
  AOI211_X1 U6210 ( .C1(INSTQUEUE_REG_8__2__SCAN_IN), .C2(n5514), .A(n5505), 
        .B(n5504), .ZN(n5506) );
  INV_X1 U6211 ( .A(n5506), .ZN(U3086) );
  NOR2_X1 U6212 ( .A1(n5507), .A2(n5771), .ZN(n5513) );
  AOI22_X1 U6213 ( .A1(n7551), .A2(n5509), .B1(n7550), .B2(n5508), .ZN(n5510)
         );
  OAI21_X1 U6214 ( .B1(n5511), .B2(n5667), .A(n5510), .ZN(n5512) );
  AOI211_X1 U6215 ( .C1(INSTQUEUE_REG_8__1__SCAN_IN), .C2(n5514), .A(n5513), 
        .B(n5512), .ZN(n5515) );
  INV_X1 U6216 ( .A(n5515), .ZN(U3085) );
  INV_X1 U6217 ( .A(n7390), .ZN(n7360) );
  AOI22_X1 U6218 ( .A1(n7424), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7360), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6219 ( .A1(n7426), .A2(n4796), .ZN(n5516) );
  OAI211_X1 U6220 ( .C1(n7261), .C2(n5518), .A(n5517), .B(n5516), .ZN(n5521)
         );
  INV_X1 U6221 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5519) );
  OAI22_X1 U6222 ( .A1(n7418), .A2(n5519), .B1(REIP_REG_1__SCAN_IN), .B2(n7415), .ZN(n5520) );
  AOI211_X1 U6223 ( .C1(n7409), .C2(n5522), .A(n5521), .B(n5520), .ZN(n5523)
         );
  OAI21_X1 U6224 ( .B1(n7265), .B2(n5524), .A(n5523), .ZN(U2826) );
  INV_X1 U6225 ( .A(n5571), .ZN(n5525) );
  AOI211_X1 U6226 ( .C1(n5527), .C2(n5526), .A(n5525), .B(n5573), .ZN(n5532)
         );
  NOR2_X1 U6227 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5528), .ZN(n5569)
         );
  NAND2_X1 U6228 ( .A1(n5529), .A2(n4112), .ZN(n5635) );
  NAND2_X1 U6229 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5635), .ZN(n5633) );
  OAI211_X1 U6230 ( .C1(n4732), .C2(n5569), .A(n5530), .B(n5633), .ZN(n5531)
         );
  NOR3_X2 U6231 ( .A1(n5532), .A2(n3637), .A3(n5531), .ZN(n5576) );
  INV_X1 U6232 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5540) );
  OAI22_X1 U6233 ( .A1(n5535), .A2(n5534), .B1(n5635), .B2(n5533), .ZN(n5567)
         );
  AOI22_X1 U6234 ( .A1(n5813), .A2(n5569), .B1(n5536), .B2(n5567), .ZN(n5537)
         );
  OAI21_X1 U6235 ( .B1(n5645), .B2(n5571), .A(n5537), .ZN(n5538) );
  AOI21_X1 U6236 ( .B1(n5642), .B2(n5573), .A(n5538), .ZN(n5539) );
  OAI21_X1 U6237 ( .B1(n5576), .B2(n5540), .A(n5539), .ZN(U3074) );
  INV_X1 U6238 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5545) );
  AOI22_X1 U6239 ( .A1(n5804), .A2(n5569), .B1(n5541), .B2(n5567), .ZN(n5542)
         );
  OAI21_X1 U6240 ( .B1(n5673), .B2(n5571), .A(n5542), .ZN(n5543) );
  AOI21_X1 U6241 ( .B1(n5670), .B2(n5573), .A(n5543), .ZN(n5544) );
  OAI21_X1 U6242 ( .B1(n5576), .B2(n5545), .A(n5544), .ZN(U3075) );
  INV_X1 U6243 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5549) );
  AOI22_X1 U6244 ( .A1(n7567), .A2(n5569), .B1(n7564), .B2(n5567), .ZN(n5546)
         );
  OAI21_X1 U6245 ( .B1(n5688), .B2(n5571), .A(n5546), .ZN(n5547) );
  AOI21_X1 U6246 ( .B1(n7568), .B2(n5573), .A(n5547), .ZN(n5548) );
  OAI21_X1 U6247 ( .B1(n5576), .B2(n5549), .A(n5548), .ZN(U3073) );
  INV_X1 U6248 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5553) );
  AOI22_X1 U6249 ( .A1(n7558), .A2(n5569), .B1(n7557), .B2(n5567), .ZN(n5550)
         );
  OAI21_X1 U6250 ( .B1(n5678), .B2(n5571), .A(n5550), .ZN(n5551) );
  AOI21_X1 U6251 ( .B1(n7559), .B2(n5573), .A(n5551), .ZN(n5552) );
  OAI21_X1 U6252 ( .B1(n5576), .B2(n5553), .A(n5552), .ZN(U3072) );
  INV_X1 U6253 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5558) );
  AOI22_X1 U6254 ( .A1(n5785), .A2(n5569), .B1(n5554), .B2(n5567), .ZN(n5555)
         );
  OAI21_X1 U6255 ( .B1(n5656), .B2(n5571), .A(n5555), .ZN(n5556) );
  AOI21_X1 U6256 ( .B1(n5653), .B2(n5573), .A(n5556), .ZN(n5557) );
  OAI21_X1 U6257 ( .B1(n5576), .B2(n5558), .A(n5557), .ZN(U3071) );
  INV_X1 U6258 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5562) );
  AOI22_X1 U6259 ( .A1(n7544), .A2(n5569), .B1(n7543), .B2(n5567), .ZN(n5559)
         );
  OAI21_X1 U6260 ( .B1(n5650), .B2(n5571), .A(n5559), .ZN(n5560) );
  AOI21_X1 U6261 ( .B1(n7545), .B2(n5573), .A(n5560), .ZN(n5561) );
  OAI21_X1 U6262 ( .B1(n5576), .B2(n5562), .A(n5561), .ZN(U3068) );
  INV_X1 U6263 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5566) );
  AOI22_X1 U6264 ( .A1(n7551), .A2(n5569), .B1(n7550), .B2(n5567), .ZN(n5563)
         );
  OAI21_X1 U6265 ( .B1(n5667), .B2(n5571), .A(n5563), .ZN(n5564) );
  AOI21_X1 U6266 ( .B1(n7552), .B2(n5573), .A(n5564), .ZN(n5565) );
  OAI21_X1 U6267 ( .B1(n5576), .B2(n5566), .A(n5565), .ZN(U3069) );
  INV_X1 U6268 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5575) );
  AOI22_X1 U6269 ( .A1(n5797), .A2(n5569), .B1(n5568), .B2(n5567), .ZN(n5570)
         );
  OAI21_X1 U6270 ( .B1(n5662), .B2(n5571), .A(n5570), .ZN(n5572) );
  AOI21_X1 U6271 ( .B1(n5659), .B2(n5573), .A(n5572), .ZN(n5574) );
  OAI21_X1 U6272 ( .B1(n5576), .B2(n5575), .A(n5574), .ZN(U3070) );
  INV_X1 U6273 ( .A(n5699), .ZN(n5577) );
  AOI21_X1 U6274 ( .B1(n5579), .B2(n5578), .A(n5577), .ZN(n5697) );
  INV_X1 U6275 ( .A(n6357), .ZN(n7115) );
  INV_X1 U6276 ( .A(n5956), .ZN(n5934) );
  INV_X1 U6277 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U6278 ( .A1(n5934), .A2(n5586), .ZN(n5582) );
  NAND2_X1 U6279 ( .A1(n5322), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5580)
         );
  OAI211_X1 U6280 ( .C1(n5962), .C2(EBX_REG_9__SCAN_IN), .A(n5948), .B(n5580), 
        .ZN(n5581) );
  AND2_X1 U6281 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  NAND2_X1 U6282 ( .A1(n5584), .A2(n5583), .ZN(n5706) );
  OR2_X1 U6283 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  NAND2_X1 U6284 ( .A1(n5706), .A2(n5585), .ZN(n7225) );
  OAI22_X1 U6285 ( .A1(n7225), .A2(n7105), .B1(n5586), .B2(n7118), .ZN(n5587)
         );
  AOI21_X1 U6286 ( .B1(n5697), .B2(n7115), .A(n5587), .ZN(n5588) );
  INV_X1 U6287 ( .A(n5588), .ZN(U2850) );
  NAND2_X1 U6288 ( .A1(n7409), .A2(n5589), .ZN(n5596) );
  INV_X1 U6289 ( .A(n5590), .ZN(n5591) );
  AOI22_X1 U6290 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n7424), .B1(n7426), 
        .B2(n5591), .ZN(n5595) );
  INV_X1 U6291 ( .A(n7261), .ZN(n7250) );
  NAND2_X1 U6292 ( .A1(n5592), .A2(n7250), .ZN(n5594) );
  NAND2_X1 U6293 ( .A1(n7403), .A2(EBX_REG_3__SCAN_IN), .ZN(n5593) );
  NAND4_X1 U6294 ( .A1(n5596), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(n5599)
         );
  INV_X1 U6295 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7028) );
  NAND3_X1 U6296 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        n7390), .ZN(n5597) );
  OAI21_X1 U6297 ( .B1(n7028), .B2(n5597), .A(n7358), .ZN(n7271) );
  AOI21_X1 U6298 ( .B1(n7028), .B2(n5597), .A(n7271), .ZN(n5598) );
  AOI211_X1 U6299 ( .C1(n5600), .C2(n7278), .A(n5599), .B(n5598), .ZN(n5601)
         );
  INV_X1 U6300 ( .A(n5601), .ZN(U2824) );
  INV_X1 U6301 ( .A(n5697), .ZN(n5689) );
  NAND3_X1 U6302 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .ZN(n5737) );
  NAND4_X1 U6303 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .A4(REIP_REG_4__SCAN_IN), .ZN(n5605) );
  NOR2_X1 U6304 ( .A1(n7415), .A2(n5605), .ZN(n7281) );
  NAND2_X1 U6305 ( .A1(REIP_REG_5__SCAN_IN), .A2(n7281), .ZN(n7298) );
  NOR2_X1 U6306 ( .A1(n5737), .A2(n7298), .ZN(n7307) );
  INV_X1 U6307 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7035) );
  INV_X1 U6308 ( .A(n7424), .ZN(n7405) );
  INV_X1 U6309 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U6310 ( .A1(n7426), .A2(n5693), .ZN(n5603) );
  AND2_X1 U6311 ( .A1(n7390), .A2(n5602), .ZN(n7385) );
  INV_X1 U6312 ( .A(n7385), .ZN(n7274) );
  OAI211_X1 U6313 ( .C1(n7405), .C2(n5695), .A(n5603), .B(n7274), .ZN(n5604)
         );
  AOI21_X1 U6314 ( .B1(n7307), .B2(n7035), .A(n5604), .ZN(n5610) );
  INV_X1 U6315 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7129) );
  NOR2_X1 U6316 ( .A1(n5605), .A2(n7129), .ZN(n6008) );
  NAND2_X1 U6317 ( .A1(n6008), .A2(n7390), .ZN(n5606) );
  NAND2_X1 U6318 ( .A1(n7358), .A2(n5606), .ZN(n7299) );
  INV_X1 U6319 ( .A(n7299), .ZN(n7280) );
  AOI21_X1 U6320 ( .B1(n5737), .B2(n7358), .A(n7280), .ZN(n5621) );
  INV_X1 U6321 ( .A(n5621), .ZN(n5715) );
  AOI22_X1 U6322 ( .A1(EBX_REG_9__SCAN_IN), .A2(n7403), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5715), .ZN(n5607) );
  OAI21_X1 U6323 ( .B1(n7431), .B2(n7225), .A(n5607), .ZN(n5608) );
  INV_X1 U6324 ( .A(n5608), .ZN(n5609) );
  OAI211_X1 U6325 ( .C1(n5689), .C2(n7396), .A(n5610), .B(n5609), .ZN(U2818)
         );
  INV_X1 U6326 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U6327 ( .A1(n7403), .A2(EBX_REG_8__SCAN_IN), .ZN(n5611) );
  OAI21_X1 U6328 ( .B1(n5612), .B2(n7412), .A(n5611), .ZN(n5617) );
  NAND2_X1 U6329 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n7296) );
  NOR3_X1 U6330 ( .A1(REIP_REG_8__SCAN_IN), .A2(n7296), .A3(n7298), .ZN(n5613)
         );
  AOI211_X1 U6331 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n7385), 
        .B(n5613), .ZN(n5614) );
  OAI21_X1 U6332 ( .B1(n7431), .B2(n5615), .A(n5614), .ZN(n5616) );
  AOI211_X1 U6333 ( .C1(n5618), .C2(n7428), .A(n5617), .B(n5616), .ZN(n5619)
         );
  OAI21_X1 U6334 ( .B1(n5621), .B2(n5620), .A(n5619), .ZN(U2819) );
  INV_X1 U6335 ( .A(EAX_REG_7__SCAN_IN), .ZN(n7007) );
  INV_X1 U6336 ( .A(n5622), .ZN(n5624) );
  AND2_X1 U6337 ( .A1(n5624), .A2(n5623), .ZN(n5626) );
  OR2_X1 U6338 ( .A1(n5626), .A2(n5625), .ZN(n7098) );
  OAI222_X1 U6339 ( .A1(n6394), .A2(n6381), .B1(n6392), .B2(n7007), .C1(n6391), 
        .C2(n7098), .ZN(U2884) );
  INV_X1 U6340 ( .A(n5684), .ZN(n5627) );
  NAND2_X1 U6341 ( .A1(n5627), .A2(n5687), .ZN(n5630) );
  AOI22_X1 U6342 ( .A1(n5630), .A2(n5629), .B1(n5628), .B2(n5637), .ZN(n5631)
         );
  NOR2_X1 U6343 ( .A1(n5631), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5634) );
  NOR2_X1 U6344 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5632), .ZN(n5639)
         );
  OAI211_X1 U6345 ( .C1(n5634), .C2(n5639), .A(n5769), .B(n5633), .ZN(n5679)
         );
  NAND2_X1 U6346 ( .A1(n5679), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5644) );
  INV_X1 U6347 ( .A(n5635), .ZN(n5636) );
  AOI22_X1 U6348 ( .A1(n5638), .A2(n5637), .B1(n5760), .B2(n5636), .ZN(n5682)
         );
  INV_X1 U6349 ( .A(n5639), .ZN(n5680) );
  OAI22_X1 U6350 ( .A1(n5682), .A2(n5821), .B1(n5640), .B2(n5680), .ZN(n5641)
         );
  AOI21_X1 U6351 ( .B1(n5684), .B2(n5642), .A(n5641), .ZN(n5643) );
  OAI211_X1 U6352 ( .C1(n5645), .C2(n5687), .A(n5644), .B(n5643), .ZN(U3042)
         );
  NAND2_X1 U6353 ( .A1(n5679), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5649) );
  OAI22_X1 U6354 ( .A1(n5682), .A2(n5779), .B1(n5646), .B2(n5680), .ZN(n5647)
         );
  AOI21_X1 U6355 ( .B1(n5684), .B2(n7545), .A(n5647), .ZN(n5648) );
  OAI211_X1 U6356 ( .C1(n5650), .C2(n5687), .A(n5649), .B(n5648), .ZN(U3036)
         );
  NAND2_X1 U6357 ( .A1(n5679), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5655) );
  OAI22_X1 U6358 ( .A1(n5682), .A2(n5791), .B1(n5651), .B2(n5680), .ZN(n5652)
         );
  AOI21_X1 U6359 ( .B1(n5684), .B2(n5653), .A(n5652), .ZN(n5654) );
  OAI211_X1 U6360 ( .C1(n5656), .C2(n5687), .A(n5655), .B(n5654), .ZN(U3039)
         );
  NAND2_X1 U6361 ( .A1(n5679), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5661) );
  OAI22_X1 U6362 ( .A1(n5682), .A2(n5803), .B1(n5657), .B2(n5680), .ZN(n5658)
         );
  AOI21_X1 U6363 ( .B1(n5684), .B2(n5659), .A(n5658), .ZN(n5660) );
  OAI211_X1 U6364 ( .C1(n5662), .C2(n5687), .A(n5661), .B(n5660), .ZN(U3038)
         );
  NAND2_X1 U6365 ( .A1(n5679), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5666) );
  OAI22_X1 U6366 ( .A1(n5682), .A2(n5774), .B1(n5663), .B2(n5680), .ZN(n5664)
         );
  AOI21_X1 U6367 ( .B1(n5684), .B2(n7552), .A(n5664), .ZN(n5665) );
  OAI211_X1 U6368 ( .C1(n5667), .C2(n5687), .A(n5666), .B(n5665), .ZN(U3037)
         );
  NAND2_X1 U6369 ( .A1(n5679), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5672) );
  OAI22_X1 U6370 ( .A1(n5682), .A2(n5810), .B1(n5668), .B2(n5680), .ZN(n5669)
         );
  AOI21_X1 U6371 ( .B1(n5684), .B2(n5670), .A(n5669), .ZN(n5671) );
  OAI211_X1 U6372 ( .C1(n5673), .C2(n5687), .A(n5672), .B(n5671), .ZN(U3043)
         );
  NAND2_X1 U6373 ( .A1(n5679), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5677) );
  OAI22_X1 U6374 ( .A1(n5682), .A2(n5784), .B1(n5674), .B2(n5680), .ZN(n5675)
         );
  AOI21_X1 U6375 ( .B1(n5684), .B2(n7559), .A(n5675), .ZN(n5676) );
  OAI211_X1 U6376 ( .C1(n5678), .C2(n5687), .A(n5677), .B(n5676), .ZN(U3040)
         );
  NAND2_X1 U6377 ( .A1(n5679), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5686) );
  OAI22_X1 U6378 ( .A1(n5682), .A2(n5796), .B1(n5681), .B2(n5680), .ZN(n5683)
         );
  AOI21_X1 U6379 ( .B1(n5684), .B2(n7568), .A(n5683), .ZN(n5685) );
  OAI211_X1 U6380 ( .C1(n5688), .C2(n5687), .A(n5686), .B(n5685), .ZN(U3041)
         );
  INV_X1 U6381 ( .A(DATAI_9_), .ZN(n5690) );
  INV_X1 U6382 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7011) );
  OAI222_X1 U6383 ( .A1(n6394), .A2(n5690), .B1(n6392), .B2(n7011), .C1(n6391), 
        .C2(n5689), .ZN(U2882) );
  OAI21_X1 U6384 ( .B1(n5692), .B2(n5691), .A(n5748), .ZN(n7229) );
  NAND2_X1 U6385 ( .A1(n7143), .A2(n5693), .ZN(n5694) );
  NAND2_X1 U6386 ( .A1(n7205), .A2(REIP_REG_9__SCAN_IN), .ZN(n7226) );
  OAI211_X1 U6387 ( .C1(n7132), .C2(n5695), .A(n5694), .B(n7226), .ZN(n5696)
         );
  AOI21_X1 U6388 ( .B1(n5697), .B2(n3628), .A(n5696), .ZN(n5698) );
  OAI21_X1 U6389 ( .B1(n7229), .B2(n7433), .A(n5698), .ZN(U2977) );
  AOI21_X1 U6390 ( .B1(n5700), .B2(n5699), .A(n5720), .ZN(n5753) );
  INV_X1 U6391 ( .A(n5947), .ZN(n5954) );
  INV_X1 U6392 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U6393 ( .A1(n5954), .A2(n5708), .ZN(n5704) );
  NAND2_X1 U6394 ( .A1(n5948), .A2(n7212), .ZN(n5702) );
  NAND2_X1 U6395 ( .A1(n5924), .A2(n5708), .ZN(n5701) );
  NAND3_X1 U6396 ( .A1(n5702), .A2(n5322), .A3(n5701), .ZN(n5703) );
  AND2_X1 U6397 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  NOR2_X2 U6398 ( .A1(n5706), .A2(n5705), .ZN(n5733) );
  INV_X1 U6399 ( .A(n5733), .ZN(n5831) );
  NAND2_X1 U6400 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  NAND2_X1 U6401 ( .A1(n5831), .A2(n5707), .ZN(n7216) );
  OAI22_X1 U6402 ( .A1(n7216), .A2(n7105), .B1(n5708), .B2(n7118), .ZN(n5709)
         );
  AOI21_X1 U6403 ( .B1(n5753), .B2(n7115), .A(n5709), .ZN(n5710) );
  INV_X1 U6404 ( .A(n5710), .ZN(U2849) );
  INV_X1 U6405 ( .A(n5753), .ZN(n5717) );
  AOI21_X1 U6406 ( .B1(n7424), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7385), 
        .ZN(n5712) );
  NAND2_X1 U6407 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n7317) );
  OAI211_X1 U6408 ( .C1(REIP_REG_9__SCAN_IN), .C2(REIP_REG_10__SCAN_IN), .A(
        n7307), .B(n7317), .ZN(n5711) );
  OAI211_X1 U6409 ( .C1(n7216), .C2(n7431), .A(n5712), .B(n5711), .ZN(n5714)
         );
  OAI22_X1 U6410 ( .A1(n7418), .A2(n5708), .B1(n5751), .B2(n7412), .ZN(n5713)
         );
  AOI211_X1 U6411 ( .C1(n5715), .C2(REIP_REG_10__SCAN_IN), .A(n5714), .B(n5713), .ZN(n5716) );
  OAI21_X1 U6412 ( .B1(n5717), .B2(n7396), .A(n5716), .ZN(U2817) );
  INV_X1 U6413 ( .A(DATAI_10_), .ZN(n5718) );
  INV_X1 U6414 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7013) );
  OAI222_X1 U6415 ( .A1(n6394), .A2(n5718), .B1(n6392), .B2(n7013), .C1(n6391), 
        .C2(n5717), .ZN(U2881) );
  INV_X1 U6416 ( .A(DATAI_11_), .ZN(n5722) );
  INV_X1 U6417 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7015) );
  NOR2_X1 U6418 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  OR2_X1 U6419 ( .A1(n5725), .A2(n5721), .ZN(n7142) );
  OAI222_X1 U6420 ( .A1(n6394), .A2(n5722), .B1(n6392), .B2(n7015), .C1(n6391), 
        .C2(n7142), .ZN(U2880) );
  OAI21_X1 U6421 ( .B1(n5725), .B2(n5724), .A(n5723), .ZN(n5880) );
  INV_X1 U6422 ( .A(n5876), .ZN(n5744) );
  INV_X1 U6423 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5742) );
  OR2_X1 U6424 ( .A1(n5947), .A2(EBX_REG_12__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6425 ( .A1(n5948), .A2(n6955), .ZN(n5727) );
  NAND2_X1 U6426 ( .A1(n5924), .A2(n5742), .ZN(n5726) );
  NAND3_X1 U6427 ( .A1(n5727), .A2(n5322), .A3(n5726), .ZN(n5728) );
  NAND2_X1 U6428 ( .A1(n5729), .A2(n5728), .ZN(n5734) );
  INV_X1 U6429 ( .A(n5734), .ZN(n5736) );
  NAND2_X1 U6430 ( .A1(n5322), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5730) );
  OAI211_X1 U6431 ( .C1(n5962), .C2(EBX_REG_11__SCAN_IN), .A(n5948), .B(n5730), 
        .ZN(n5731) );
  OAI21_X1 U6432 ( .B1(n5956), .B2(EBX_REG_11__SCAN_IN), .A(n5731), .ZN(n5830)
         );
  AND2_X2 U6433 ( .A1(n5733), .A2(n5732), .ZN(n5833) );
  INV_X1 U6434 ( .A(n5833), .ZN(n5735) );
  AND2_X2 U6435 ( .A1(n5833), .A2(n5734), .ZN(n5853) );
  AOI21_X1 U6436 ( .B1(n5736), .B2(n5735), .A(n5853), .ZN(n6952) );
  INV_X1 U6437 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7306) );
  NOR3_X1 U6438 ( .A1(n5737), .A2(n7317), .A3(n7306), .ZN(n6007) );
  AOI21_X1 U6439 ( .B1(n6007), .B2(n6008), .A(n7415), .ZN(n5738) );
  OR2_X1 U6440 ( .A1(n5738), .A2(n7360), .ZN(n7324) );
  AOI22_X1 U6441 ( .A1(n7409), .A2(n6952), .B1(REIP_REG_12__SCAN_IN), .B2(
        n7324), .ZN(n5741) );
  INV_X1 U6442 ( .A(n6007), .ZN(n5739) );
  NOR3_X1 U6443 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5739), .A3(n7298), .ZN(n7325) );
  AOI211_X1 U6444 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n7385), 
        .B(n7325), .ZN(n5740) );
  OAI211_X1 U6445 ( .C1(n5742), .C2(n7418), .A(n5741), .B(n5740), .ZN(n5743)
         );
  AOI21_X1 U6446 ( .B1(n7426), .B2(n5744), .A(n5743), .ZN(n5745) );
  OAI21_X1 U6447 ( .B1(n5880), .B2(n7396), .A(n5745), .ZN(U2815) );
  AOI22_X1 U6448 ( .A1(n6952), .A2(n7114), .B1(EBX_REG_12__SCAN_IN), .B2(n6338), .ZN(n5746) );
  OAI21_X1 U6449 ( .B1(n5880), .B2(n6357), .A(n5746), .ZN(U2847) );
  NAND2_X1 U6450 ( .A1(n5748), .A2(n5747), .ZN(n5826) );
  NAND2_X1 U6451 ( .A1(n5827), .A2(n5825), .ZN(n5749) );
  XNOR2_X1 U6452 ( .A(n5826), .B(n5749), .ZN(n7221) );
  INV_X1 U6453 ( .A(n7221), .ZN(n5755) );
  AOI22_X1 U6454 ( .A1(n7147), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n7205), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5750) );
  OAI21_X1 U6455 ( .B1(n5751), .B2(n7152), .A(n5750), .ZN(n5752) );
  AOI21_X1 U6456 ( .B1(n5753), .B2(n3628), .A(n5752), .ZN(n5754) );
  OAI21_X1 U6457 ( .B1(n5755), .B2(n7433), .A(n5754), .ZN(U2976) );
  OAI21_X1 U6458 ( .B1(n5818), .B2(n5761), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5757) );
  INV_X1 U6459 ( .A(n5758), .ZN(n5759) );
  AOI22_X1 U6460 ( .A1(n5765), .A2(n5763), .B1(n5760), .B2(n5759), .ZN(n5822)
         );
  NOR2_X1 U6461 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5762), .ZN(n5812)
         );
  INV_X1 U6462 ( .A(n5812), .ZN(n5766) );
  INV_X1 U6463 ( .A(n5763), .ZN(n5764) );
  AOI22_X1 U6464 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5766), .B1(n5765), .B2(
        n5764), .ZN(n5768) );
  NAND3_X1 U6465 ( .A1(n5769), .A2(n5768), .A3(n5767), .ZN(n5811) );
  AOI22_X1 U6466 ( .A1(n7551), .A2(n5812), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5811), .ZN(n5770) );
  OAI21_X1 U6467 ( .B1(n5771), .B2(n5816), .A(n5770), .ZN(n5772) );
  AOI21_X1 U6468 ( .B1(n7553), .B2(n5818), .A(n5772), .ZN(n5773) );
  OAI21_X1 U6469 ( .B1(n5822), .B2(n5774), .A(n5773), .ZN(U3101) );
  AOI22_X1 U6470 ( .A1(n7544), .A2(n5812), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5811), .ZN(n5775) );
  OAI21_X1 U6471 ( .B1(n5816), .B2(n5776), .A(n5775), .ZN(n5777) );
  AOI21_X1 U6472 ( .B1(n7546), .B2(n5818), .A(n5777), .ZN(n5778) );
  OAI21_X1 U6473 ( .B1(n5822), .B2(n5779), .A(n5778), .ZN(U3100) );
  AOI22_X1 U6474 ( .A1(n7558), .A2(n5812), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5811), .ZN(n5780) );
  OAI21_X1 U6475 ( .B1(n5816), .B2(n5781), .A(n5780), .ZN(n5782) );
  AOI21_X1 U6476 ( .B1(n7560), .B2(n5818), .A(n5782), .ZN(n5783) );
  OAI21_X1 U6477 ( .B1(n5822), .B2(n5784), .A(n5783), .ZN(U3104) );
  AOI22_X1 U6478 ( .A1(n5785), .A2(n5812), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5811), .ZN(n5786) );
  OAI21_X1 U6479 ( .B1(n5816), .B2(n5787), .A(n5786), .ZN(n5788) );
  AOI21_X1 U6480 ( .B1(n5789), .B2(n5818), .A(n5788), .ZN(n5790) );
  OAI21_X1 U6481 ( .B1(n5822), .B2(n5791), .A(n5790), .ZN(U3103) );
  AOI22_X1 U6482 ( .A1(n7567), .A2(n5812), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5811), .ZN(n5792) );
  OAI21_X1 U6483 ( .B1(n5816), .B2(n5793), .A(n5792), .ZN(n5794) );
  AOI21_X1 U6484 ( .B1(n7570), .B2(n5818), .A(n5794), .ZN(n5795) );
  OAI21_X1 U6485 ( .B1(n5822), .B2(n5796), .A(n5795), .ZN(U3105) );
  AOI22_X1 U6486 ( .A1(n5797), .A2(n5812), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5811), .ZN(n5798) );
  OAI21_X1 U6487 ( .B1(n5816), .B2(n5799), .A(n5798), .ZN(n5800) );
  AOI21_X1 U6488 ( .B1(n5801), .B2(n5818), .A(n5800), .ZN(n5802) );
  OAI21_X1 U6489 ( .B1(n5822), .B2(n5803), .A(n5802), .ZN(U3102) );
  AOI22_X1 U6490 ( .A1(n5804), .A2(n5812), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5811), .ZN(n5805) );
  OAI21_X1 U6491 ( .B1(n5816), .B2(n5806), .A(n5805), .ZN(n5807) );
  AOI21_X1 U6492 ( .B1(n5808), .B2(n5818), .A(n5807), .ZN(n5809) );
  OAI21_X1 U6493 ( .B1(n5822), .B2(n5810), .A(n5809), .ZN(U3107) );
  AOI22_X1 U6494 ( .A1(n5813), .A2(n5812), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5811), .ZN(n5814) );
  OAI21_X1 U6495 ( .B1(n5816), .B2(n5815), .A(n5814), .ZN(n5817) );
  AOI21_X1 U6496 ( .B1(n5819), .B2(n5818), .A(n5817), .ZN(n5820) );
  OAI21_X1 U6497 ( .B1(n5822), .B2(n5821), .A(n5820), .ZN(U3106) );
  INV_X1 U6498 ( .A(DATAI_12_), .ZN(n5823) );
  INV_X1 U6499 ( .A(EAX_REG_12__SCAN_IN), .ZN(n7017) );
  OAI222_X1 U6500 ( .A1(n6394), .A2(n5823), .B1(n6392), .B2(n7017), .C1(n6391), 
        .C2(n5880), .ZN(U2879) );
  NAND2_X1 U6501 ( .A1(n5824), .A2(n5870), .ZN(n5829) );
  NAND2_X1 U6502 ( .A1(n5826), .A2(n5825), .ZN(n5869) );
  NAND2_X1 U6503 ( .A1(n5869), .A2(n5827), .ZN(n5828) );
  XOR2_X1 U6504 ( .A(n5829), .B(n5828), .Z(n7146) );
  AND2_X1 U6505 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  NOR2_X1 U6506 ( .A1(n5833), .A2(n5832), .ZN(n7308) );
  NAND3_X1 U6507 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n7220), .ZN(n5836) );
  OR2_X1 U6508 ( .A1(n5834), .A2(n5836), .ZN(n6031) );
  OR2_X1 U6509 ( .A1(n6566), .A2(n6031), .ZN(n5838) );
  NOR2_X1 U6510 ( .A1(n5836), .A2(n5835), .ZN(n5841) );
  INV_X1 U6511 ( .A(n5841), .ZN(n5899) );
  OR2_X1 U6512 ( .A1(n6036), .A2(n5899), .ZN(n5837) );
  NAND2_X1 U6513 ( .A1(n5838), .A2(n5837), .ZN(n6578) );
  INV_X1 U6514 ( .A(n6578), .ZN(n6949) );
  INV_X1 U6515 ( .A(n5839), .ZN(n6034) );
  NAND2_X1 U6516 ( .A1(n6029), .A2(n6031), .ZN(n5840) );
  AND2_X1 U6517 ( .A1(n6034), .A2(n5840), .ZN(n6135) );
  OR2_X1 U6518 ( .A1(n6036), .A2(n5841), .ZN(n6134) );
  NAND2_X1 U6519 ( .A1(n6135), .A2(n6134), .ZN(n6945) );
  AOI22_X1 U6520 ( .A1(n7205), .A2(REIP_REG_11__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6945), .ZN(n5842) );
  OAI21_X1 U6521 ( .B1(n6949), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5842), 
        .ZN(n5843) );
  AOI21_X1 U6522 ( .B1(n7308), .B2(n7238), .A(n5843), .ZN(n5844) );
  OAI21_X1 U6523 ( .B1(n7146), .B2(n6584), .A(n5844), .ZN(U3007) );
  NAND2_X1 U6524 ( .A1(n5847), .A2(n5846), .ZN(n6465) );
  OAI21_X1 U6525 ( .B1(n5847), .B2(n5846), .A(n6465), .ZN(n5862) );
  INV_X1 U6526 ( .A(n5862), .ZN(n5858) );
  NOR3_X1 U6527 ( .A1(n5848), .A2(n6955), .A3(n6948), .ZN(n5896) );
  INV_X1 U6528 ( .A(n7175), .ZN(n7219) );
  INV_X1 U6529 ( .A(n6945), .ZN(n6575) );
  OAI21_X1 U6530 ( .B1(n5896), .B2(n7219), .A(n6575), .ZN(n5908) );
  NOR3_X1 U6531 ( .A1(n6949), .A2(n6948), .A3(n6955), .ZN(n5849) );
  AOI22_X1 U6532 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5908), .B1(n5849), .B2(n5848), .ZN(n5857) );
  MUX2_X1 U6533 ( .A(n5956), .B(n5322), .S(EBX_REG_13__SCAN_IN), .Z(n5850) );
  OAI21_X1 U6534 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5963), .A(n5850), 
        .ZN(n5851) );
  INV_X1 U6535 ( .A(n5851), .ZN(n5852) );
  OR2_X1 U6536 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  AND2_X1 U6537 ( .A1(n5913), .A2(n5854), .ZN(n7318) );
  INV_X1 U6538 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5855) );
  NOR2_X1 U6539 ( .A1(n7213), .A2(n5855), .ZN(n5865) );
  AOI21_X1 U6540 ( .B1(n7318), .B2(n7238), .A(n5865), .ZN(n5856) );
  OAI211_X1 U6541 ( .C1(n5858), .C2(n6584), .A(n5857), .B(n5856), .ZN(U3005)
         );
  XNOR2_X1 U6542 ( .A(n5860), .B(n5859), .ZN(n7321) );
  AOI22_X1 U6543 ( .A1(n7318), .A2(n7114), .B1(EBX_REG_13__SCAN_IN), .B2(n6338), .ZN(n5861) );
  OAI21_X1 U6544 ( .B1(n7321), .B2(n6357), .A(n5861), .ZN(U2846) );
  NAND2_X1 U6545 ( .A1(n5862), .A2(n7148), .ZN(n5867) );
  NOR2_X1 U6546 ( .A1(n7132), .A2(n5863), .ZN(n5864) );
  AOI211_X1 U6547 ( .C1(n7143), .C2(n7322), .A(n5865), .B(n5864), .ZN(n5866)
         );
  OAI211_X1 U6548 ( .C1(n7321), .C2(n6489), .A(n5867), .B(n5866), .ZN(U2973)
         );
  NAND2_X1 U6549 ( .A1(n5869), .A2(n5868), .ZN(n5871) );
  AND2_X1 U6550 ( .A1(n5871), .A2(n5870), .ZN(n5875) );
  NAND2_X1 U6551 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  XNOR2_X1 U6552 ( .A(n5875), .B(n5874), .ZN(n6947) );
  NAND2_X1 U6553 ( .A1(n6947), .A2(n7148), .ZN(n5879) );
  INV_X1 U6554 ( .A(REIP_REG_12__SCAN_IN), .ZN(n7039) );
  NOR2_X1 U6555 ( .A1(n7213), .A2(n7039), .ZN(n6951) );
  NOR2_X1 U6556 ( .A1(n7152), .A2(n5876), .ZN(n5877) );
  AOI211_X1 U6557 ( .C1(n7147), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6951), 
        .B(n5877), .ZN(n5878) );
  OAI211_X1 U6558 ( .C1(n6489), .C2(n5880), .A(n5879), .B(n5878), .ZN(U2974)
         );
  OAI21_X1 U6559 ( .B1(n5887), .B2(n6477), .A(n6454), .ZN(n6455) );
  MUX2_X1 U6560 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .B(n5881), .S(n4049), 
        .Z(n5882) );
  XNOR2_X1 U6561 ( .A(n6455), .B(n5882), .ZN(n7149) );
  MUX2_X1 U6562 ( .A(n5947), .B(n5948), .S(EBX_REG_14__SCAN_IN), .Z(n5884) );
  NAND2_X1 U6563 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5962), .ZN(n5883) );
  AND3_X1 U6564 ( .A1(n5884), .A2(n5939), .A3(n5883), .ZN(n5912) );
  NAND2_X1 U6565 ( .A1(n5322), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5885) );
  OAI211_X1 U6566 ( .C1(n5962), .C2(EBX_REG_15__SCAN_IN), .A(n5948), .B(n5885), 
        .ZN(n5886) );
  OAI21_X1 U6567 ( .B1(n5956), .B2(EBX_REG_15__SCAN_IN), .A(n5886), .ZN(n6300)
         );
  OR2_X1 U6568 ( .A1(n5947), .A2(EBX_REG_16__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6569 ( .A1(n5948), .A2(n5887), .ZN(n5889) );
  INV_X1 U6570 ( .A(EBX_REG_16__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U6571 ( .A1(n5924), .A2(n7355), .ZN(n5888) );
  NAND3_X1 U6572 ( .A1(n5889), .A2(n5322), .A3(n5888), .ZN(n5890) );
  NAND2_X1 U6573 ( .A1(n5891), .A2(n5890), .ZN(n6349) );
  MUX2_X1 U6574 ( .A(n5956), .B(n5322), .S(EBX_REG_17__SCAN_IN), .Z(n5892) );
  OAI21_X1 U6575 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5963), .A(n5892), 
        .ZN(n5894) );
  NAND2_X1 U6576 ( .A1(n5893), .A2(n5894), .ZN(n5895) );
  NAND2_X1 U6577 ( .A1(n6336), .A2(n5895), .ZN(n7363) );
  INV_X1 U6578 ( .A(n5896), .ZN(n5916) );
  NOR2_X1 U6579 ( .A1(n5922), .A2(n5916), .ZN(n6579) );
  NAND3_X1 U6580 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6579), .ZN(n6569) );
  NOR2_X1 U6581 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6569), .ZN(n6567)
         );
  AOI22_X1 U6582 ( .A1(n6578), .A2(n6567), .B1(n7205), .B2(
        REIP_REG_17__SCAN_IN), .ZN(n5904) );
  INV_X1 U6583 ( .A(n6569), .ZN(n5897) );
  NAND2_X1 U6584 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5897), .ZN(n5898) );
  OAI21_X1 U6585 ( .B1(n5899), .B2(n5898), .A(n7197), .ZN(n5902) );
  NAND2_X1 U6586 ( .A1(n6029), .A2(n6569), .ZN(n5900) );
  AND2_X1 U6587 ( .A1(n6135), .A2(n5900), .ZN(n5901) );
  NAND2_X1 U6588 ( .A1(n5902), .A2(n5901), .ZN(n6568) );
  NAND2_X1 U6589 ( .A1(n6568), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5903) );
  OAI211_X1 U6590 ( .C1(n7363), .C2(n7215), .A(n5904), .B(n5903), .ZN(n5905)
         );
  AOI21_X1 U6591 ( .B1(n7149), .B2(n7239), .A(n5905), .ZN(n5906) );
  INV_X1 U6592 ( .A(n5906), .ZN(U3001) );
  INV_X1 U6593 ( .A(DATAI_13_), .ZN(n5907) );
  OAI222_X1 U6594 ( .A1(n6394), .A2(n5907), .B1(n6391), .B2(n7321), .C1(n7019), 
        .C2(n6392), .ZN(U2878) );
  INV_X1 U6595 ( .A(n5908), .ZN(n5921) );
  NAND2_X1 U6596 ( .A1(n6465), .A2(n5909), .ZN(n5911) );
  XNOR2_X1 U6597 ( .A(n6477), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5910)
         );
  XNOR2_X1 U6598 ( .A(n5911), .B(n5910), .ZN(n6484) );
  NAND2_X1 U6599 ( .A1(n6484), .A2(n7239), .ZN(n5920) );
  NAND2_X1 U6600 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  NAND2_X1 U6601 ( .A1(n6301), .A2(n5914), .ZN(n7341) );
  INV_X1 U6602 ( .A(n7341), .ZN(n5918) );
  INV_X1 U6603 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U6604 ( .A1(n7213), .A2(n5915), .ZN(n6486) );
  NOR3_X1 U6605 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6949), .A3(n5916), 
        .ZN(n5917) );
  AOI211_X1 U6606 ( .C1(n7238), .C2(n5918), .A(n6486), .B(n5917), .ZN(n5919)
         );
  OAI211_X1 U6607 ( .C1(n5922), .C2(n5921), .A(n5920), .B(n5919), .ZN(U3004)
         );
  INV_X1 U6608 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7378) );
  NAND2_X1 U6609 ( .A1(n5954), .A2(n7378), .ZN(n5928) );
  NAND2_X1 U6610 ( .A1(n5948), .A2(n5923), .ZN(n5926) );
  NAND2_X1 U6611 ( .A1(n5924), .A2(n7378), .ZN(n5925) );
  NAND3_X1 U6612 ( .A1(n5926), .A2(n5322), .A3(n5925), .ZN(n5927) );
  AND2_X1 U6613 ( .A1(n5928), .A2(n5927), .ZN(n6337) );
  OR2_X2 U6614 ( .A1(n6336), .A2(n6337), .ZN(n6334) );
  NAND2_X1 U6615 ( .A1(n5322), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5929) );
  OAI211_X1 U6616 ( .C1(n5962), .C2(EBX_REG_19__SCAN_IN), .A(n5948), .B(n5929), 
        .ZN(n5930) );
  OAI21_X1 U6617 ( .B1(n5956), .B2(EBX_REG_19__SCAN_IN), .A(n5930), .ZN(n6133)
         );
  MUX2_X1 U6618 ( .A(n5947), .B(n5948), .S(EBX_REG_20__SCAN_IN), .Z(n5933) );
  NAND2_X1 U6619 ( .A1(n5962), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5931) );
  AND2_X1 U6620 ( .A1(n5939), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U6621 ( .A1(n5933), .A2(n5932), .ZN(n6124) );
  INV_X1 U6622 ( .A(EBX_REG_21__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U6623 ( .A1(n5934), .A2(n7111), .ZN(n5937) );
  NAND2_X1 U6624 ( .A1(n4768), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5935) );
  OAI211_X1 U6625 ( .C1(n5962), .C2(EBX_REG_21__SCAN_IN), .A(n5948), .B(n5935), 
        .ZN(n5936) );
  AND2_X1 U6626 ( .A1(n5937), .A2(n5936), .ZN(n6544) );
  MUX2_X1 U6627 ( .A(n5947), .B(n5948), .S(EBX_REG_22__SCAN_IN), .Z(n5941) );
  NAND2_X1 U6628 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n5962), .ZN(n5938) );
  AND2_X1 U6629 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  NAND2_X1 U6630 ( .A1(n5941), .A2(n5940), .ZN(n6327) );
  MUX2_X1 U6631 ( .A(n5956), .B(n5322), .S(EBX_REG_23__SCAN_IN), .Z(n5942) );
  OAI21_X1 U6632 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5963), .A(n5942), 
        .ZN(n6290) );
  MUX2_X1 U6633 ( .A(n5947), .B(n5948), .S(EBX_REG_24__SCAN_IN), .Z(n5944) );
  NAND2_X1 U6634 ( .A1(n5962), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5943) );
  AND2_X1 U6635 ( .A1(n5944), .A2(n5943), .ZN(n6090) );
  MUX2_X1 U6636 ( .A(n5956), .B(n5322), .S(EBX_REG_25__SCAN_IN), .Z(n5946) );
  OR2_X1 U6637 ( .A1(n5963), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5945)
         );
  AND2_X1 U6638 ( .A1(n5946), .A2(n5945), .ZN(n6260) );
  OR2_X1 U6639 ( .A1(n5947), .A2(EBX_REG_26__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U6640 ( .A1(n5948), .A2(n6414), .ZN(n5949) );
  OAI211_X1 U6641 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5962), .A(n5949), .B(n5322), 
        .ZN(n5950) );
  NAND2_X1 U6642 ( .A1(n5951), .A2(n5950), .ZN(n6250) );
  AND2_X2 U6643 ( .A1(n6249), .A2(n6250), .ZN(n6024) );
  NOR2_X1 U6644 ( .A1(n5962), .A2(EBX_REG_29__SCAN_IN), .ZN(n5953) );
  AOI21_X1 U6645 ( .B1(n5952), .B2(n6096), .A(n5953), .ZN(n6192) );
  MUX2_X1 U6646 ( .A(n5953), .B(n6192), .S(n5322), .Z(n6095) );
  MUX2_X1 U6647 ( .A(n5954), .B(n4770), .S(EBX_REG_28__SCAN_IN), .Z(n5955) );
  AOI21_X1 U6648 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5962), .A(n5955), 
        .ZN(n6025) );
  MUX2_X1 U6649 ( .A(n5956), .B(n5322), .S(EBX_REG_27__SCAN_IN), .Z(n5957) );
  OAI21_X1 U6650 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5963), .A(n5957), 
        .ZN(n6235) );
  NOR2_X1 U6651 ( .A1(n6025), .A2(n6235), .ZN(n6023) );
  AND2_X1 U6652 ( .A1(n6095), .A2(n6023), .ZN(n5958) );
  AND2_X1 U6654 ( .A1(n5962), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5959)
         );
  AOI21_X1 U6655 ( .B1(n5963), .B2(EBX_REG_30__SCAN_IN), .A(n5959), .ZN(n6194)
         );
  OAI22_X1 U6657 ( .A1(n5963), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5962), .ZN(n5964) );
  INV_X1 U6658 ( .A(n5964), .ZN(n5965) );
  XNOR2_X2 U6659 ( .A(n5966), .B(n5965), .ZN(n6162) );
  OAI22_X1 U6660 ( .A1(n6162), .A2(n7105), .B1(n7118), .B2(n5967), .ZN(U2828)
         );
  AOI22_X1 U6661 ( .A1(n5999), .A2(EAX_REG_31__SCAN_IN), .B1(n5968), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6006) );
  NOR2_X1 U6662 ( .A1(n5970), .A2(n5969), .ZN(n5991) );
  AOI22_X1 U6663 ( .A1(n5971), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5979) );
  AOI22_X1 U6664 ( .A1(n3684), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5972), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5978) );
  AOI22_X1 U6665 ( .A1(n3635), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5973), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5977) );
  AOI22_X1 U6666 ( .A1(n5975), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5974), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5976) );
  NAND4_X1 U6667 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n5989)
         );
  AOI22_X1 U6668 ( .A1(n5980), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5987) );
  AOI22_X1 U6669 ( .A1(n5981), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5986) );
  AOI22_X1 U6670 ( .A1(n3901), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5985) );
  AOI22_X1 U6671 ( .A1(n3800), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5983), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5984) );
  NAND4_X1 U6672 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n5988)
         );
  NOR2_X1 U6673 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  XNOR2_X1 U6674 ( .A(n5991), .B(n5990), .ZN(n5994) );
  INV_X1 U6675 ( .A(n5992), .ZN(n5993) );
  NAND2_X1 U6676 ( .A1(n5994), .A2(n5993), .ZN(n6004) );
  NAND2_X1 U6677 ( .A1(n5995), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5996)
         );
  NAND2_X1 U6678 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  AOI21_X1 U6679 ( .B1(n5999), .B2(EAX_REG_30__SCAN_IN), .A(n5998), .ZN(n6003)
         );
  XNOR2_X1 U6680 ( .A(n6000), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6399)
         );
  AND2_X1 U6681 ( .A1(n6399), .A2(n6001), .ZN(n6002) );
  AOI21_X1 U6682 ( .B1(n6004), .B2(n6003), .A(n6002), .ZN(n6190) );
  NAND2_X1 U6683 ( .A1(n6189), .A2(n6190), .ZN(n6005) );
  XOR2_X1 U6684 ( .A(n6006), .B(n6005), .Z(n6186) );
  NAND2_X1 U6685 ( .A1(n6186), .A2(n7428), .ZN(n6019) );
  INV_X1 U6686 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7070) );
  NOR2_X1 U6687 ( .A1(n7070), .A2(n7065), .ZN(n6011) );
  INV_X1 U6688 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7054) );
  INV_X1 U6689 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7420) );
  INV_X1 U6690 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7391) );
  NAND3_X1 U6691 ( .A1(n6008), .A2(n6007), .A3(REIP_REG_12__SCAN_IN), .ZN(
        n7319) );
  NOR2_X1 U6692 ( .A1(n7319), .A2(n5855), .ZN(n7332) );
  NAND2_X1 U6693 ( .A1(n7332), .A2(REIP_REG_14__SCAN_IN), .ZN(n6304) );
  INV_X1 U6694 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7344) );
  INV_X1 U6695 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7342) );
  NOR3_X1 U6696 ( .A1(n6304), .A2(n7344), .A3(n7342), .ZN(n7356) );
  NAND2_X1 U6697 ( .A1(n7356), .A2(REIP_REG_17__SCAN_IN), .ZN(n7359) );
  NAND2_X1 U6698 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n7393) );
  NOR3_X1 U6699 ( .A1(n7391), .A2(n7359), .A3(n7393), .ZN(n7407) );
  NAND2_X1 U6700 ( .A1(REIP_REG_21__SCAN_IN), .A2(n7407), .ZN(n7414) );
  NOR2_X1 U6701 ( .A1(n7420), .A2(n7414), .ZN(n6291) );
  NAND2_X1 U6702 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6291), .ZN(n6280) );
  NOR2_X1 U6703 ( .A1(n7054), .A2(n6280), .ZN(n6269) );
  AND2_X1 U6704 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6269), .ZN(n6253) );
  AND2_X1 U6705 ( .A1(n6253), .A2(REIP_REG_26__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U6706 ( .A1(n7390), .A2(n6012), .ZN(n6009) );
  AND2_X1 U6707 ( .A1(n7358), .A2(n6009), .ZN(n6238) );
  AOI21_X1 U6708 ( .B1(REIP_REG_28__SCAN_IN), .B2(REIP_REG_27__SCAN_IN), .A(
        n7415), .ZN(n6010) );
  NOR2_X1 U6709 ( .A1(n6238), .A2(n6010), .ZN(n6216) );
  OAI21_X1 U6710 ( .B1(n6011), .B2(n7415), .A(n6216), .ZN(n6213) );
  INV_X1 U6711 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7062) );
  INV_X1 U6712 ( .A(n6012), .ZN(n6240) );
  NOR3_X1 U6713 ( .A1(n7415), .A2(n7062), .A3(n6240), .ZN(n6226) );
  NAND2_X1 U6714 ( .A1(n6226), .A2(REIP_REG_28__SCAN_IN), .ZN(n6221) );
  INV_X1 U6715 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7067) );
  NAND3_X1 U6716 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .A3(
        n7067), .ZN(n6016) );
  AOI22_X1 U6717 ( .A1(n6014), .A2(n6013), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n7424), .ZN(n6015) );
  OAI21_X1 U6718 ( .B1(n6221), .B2(n6016), .A(n6015), .ZN(n6017) );
  AOI21_X1 U6719 ( .B1(REIP_REG_31__SCAN_IN), .B2(n6213), .A(n6017), .ZN(n6018) );
  OAI211_X1 U6720 ( .C1(n6162), .C2(n7431), .A(n6019), .B(n6018), .ZN(U2796)
         );
  OR2_X1 U6721 ( .A1(n4049), .A2(n6414), .ZN(n6405) );
  OAI21_X1 U6722 ( .B1(n6505), .B2(n6477), .A(n6405), .ZN(n6020) );
  XNOR2_X1 U6723 ( .A(n6477), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6021)
         );
  XNOR2_X1 U6724 ( .A(n6022), .B(n6021), .ZN(n6055) );
  OR2_X1 U6725 ( .A1(n6252), .A2(n6235), .ZN(n6237) );
  AOI21_X1 U6726 ( .B1(n6025), .B2(n6237), .A(n6191), .ZN(n6312) );
  NOR2_X1 U6727 ( .A1(n6569), .A2(n6026), .ZN(n6558) );
  AND2_X1 U6728 ( .A1(n6558), .A2(n6080), .ZN(n6028) );
  NAND2_X1 U6729 ( .A1(n6578), .A2(n6028), .ZN(n6039) );
  OR2_X1 U6730 ( .A1(n6039), .A2(n6040), .ZN(n6538) );
  OR2_X1 U6731 ( .A1(n6036), .A2(n6028), .ZN(n6027) );
  AND2_X1 U6732 ( .A1(n6134), .A2(n6027), .ZN(n6033) );
  INV_X1 U6733 ( .A(n6028), .ZN(n6030) );
  OAI21_X1 U6734 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(n6032) );
  AND3_X1 U6735 ( .A1(n6034), .A2(n6033), .A3(n6032), .ZN(n6549) );
  NAND2_X1 U6736 ( .A1(n6538), .A2(n6549), .ZN(n6541) );
  INV_X1 U6737 ( .A(n6035), .ZN(n6041) );
  AOI21_X1 U6738 ( .B1(n6566), .B2(n6036), .A(n6041), .ZN(n6037) );
  NOR2_X1 U6739 ( .A1(n6541), .A2(n6037), .ZN(n6511) );
  NAND2_X1 U6740 ( .A1(n6511), .A2(n7219), .ZN(n6164) );
  NAND2_X1 U6741 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6057) );
  INV_X1 U6742 ( .A(n6057), .ZN(n6038) );
  NAND2_X1 U6743 ( .A1(n6511), .A2(n6038), .ZN(n6500) );
  NAND3_X1 U6744 ( .A1(n6164), .A2(n6500), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6044) );
  INV_X1 U6745 ( .A(n6039), .ZN(n6552) );
  AND2_X1 U6746 ( .A1(n6552), .A2(n6040), .ZN(n6529) );
  NAND2_X1 U6747 ( .A1(n6529), .A2(n6041), .ZN(n6520) );
  OR2_X1 U6748 ( .A1(n6520), .A2(n6057), .ZN(n6168) );
  INV_X1 U6749 ( .A(n6168), .ZN(n6506) );
  AND2_X1 U6750 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6056) );
  INV_X1 U6751 ( .A(n6056), .ZN(n6097) );
  NAND3_X1 U6752 ( .A1(n6506), .A2(n6042), .A3(n6097), .ZN(n6043) );
  NAND2_X1 U6753 ( .A1(n7205), .A2(REIP_REG_28__SCAN_IN), .ZN(n6047) );
  NAND3_X1 U6754 ( .A1(n6044), .A2(n6043), .A3(n6047), .ZN(n6045) );
  AOI21_X1 U6755 ( .B1(n6312), .B2(n7238), .A(n6045), .ZN(n6046) );
  OAI21_X1 U6756 ( .B1(n6055), .B2(n6584), .A(n6046), .ZN(U2990) );
  OAI21_X1 U6757 ( .B1(n7132), .B2(n6048), .A(n6047), .ZN(n6053) );
  OAI21_X1 U6758 ( .B1(n6049), .B2(n6051), .A(n6050), .ZN(n6367) );
  NOR2_X1 U6759 ( .A1(n6367), .A2(n6489), .ZN(n6052) );
  AOI211_X1 U6760 ( .C1(n6227), .C2(n7143), .A(n6053), .B(n6052), .ZN(n6054)
         );
  OAI21_X1 U6761 ( .B1(n6055), .B2(n7433), .A(n6054), .ZN(U2958) );
  AND4_X1 U6762 ( .A1(n4049), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n6062) );
  NAND2_X1 U6763 ( .A1(n6056), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6491) );
  OAI21_X1 U6764 ( .B1(n6057), .B2(n6491), .A(n6395), .ZN(n6059) );
  AOI21_X1 U6765 ( .B1(n6060), .B2(n6059), .A(n6058), .ZN(n6396) );
  NOR3_X1 U6766 ( .A1(n6395), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6061) );
  AOI22_X1 U6767 ( .A1(n6063), .A2(n6062), .B1(n6396), .B2(n6061), .ZN(n6064)
         );
  INV_X1 U6768 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U6769 ( .A(n6064), .B(n6166), .ZN(n6174) );
  NOR2_X1 U6770 ( .A1(n7213), .A2(n7067), .ZN(n6170) );
  AOI21_X1 U6771 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6170), 
        .ZN(n6065) );
  OAI21_X1 U6772 ( .B1(n7152), .B2(n6066), .A(n6065), .ZN(n6067) );
  AOI21_X1 U6773 ( .B1(n6186), .B2(n3628), .A(n6067), .ZN(n6068) );
  OAI21_X1 U6774 ( .B1(n6174), .B2(n7433), .A(n6068), .ZN(U2955) );
  NOR2_X1 U6775 ( .A1(n7487), .A2(n7195), .ZN(n6967) );
  AOI22_X1 U6776 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n3881), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6166), .ZN(n6968) );
  INV_X1 U6777 ( .A(n6968), .ZN(n6072) );
  NOR2_X1 U6778 ( .A1(n6069), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6071)
         );
  AOI222_X1 U6779 ( .A1(n6967), .A2(n6072), .B1(n6960), .B2(n6071), .C1(n6070), 
        .C2(n7481), .ZN(n6077) );
  AOI21_X1 U6780 ( .B1(n7494), .B2(n6073), .A(n6076), .ZN(n6075) );
  OAI22_X1 U6781 ( .A1(n6077), .A2(n6076), .B1(n6075), .B2(n6074), .ZN(U3459)
         );
  INV_X1 U6782 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6551) );
  INV_X1 U6783 ( .A(n6131), .ZN(n6431) );
  INV_X1 U6784 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6140) );
  XNOR2_X1 U6785 ( .A(n6395), .B(n6140), .ZN(n6130) );
  NAND2_X1 U6786 ( .A1(n6431), .A2(n6078), .ZN(n6128) );
  INV_X1 U6787 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6557) );
  NOR2_X1 U6788 ( .A1(n6395), .A2(n6557), .ZN(n6079) );
  INV_X1 U6789 ( .A(n6080), .ZN(n6081) );
  NAND2_X1 U6790 ( .A1(n6477), .A2(n6081), .ZN(n6082) );
  XNOR2_X1 U6791 ( .A(n6395), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6155)
         );
  NAND2_X1 U6792 ( .A1(n6156), .A2(n6155), .ZN(n6157) );
  NAND3_X1 U6793 ( .A1(n6441), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6087) );
  INV_X1 U6794 ( .A(n6083), .ZN(n6085) );
  XNOR2_X1 U6795 ( .A(n6089), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6113)
         );
  AND2_X1 U6796 ( .A1(n6288), .A2(n6090), .ZN(n6091) );
  NOR2_X1 U6797 ( .A1(n6261), .A2(n6091), .ZN(n6317) );
  AOI21_X1 U6798 ( .B1(n6529), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U6799 ( .A1(n7205), .A2(REIP_REG_24__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U6800 ( .B1(n6511), .B2(n6092), .A(n6109), .ZN(n6093) );
  AOI21_X1 U6801 ( .B1(n6317), .B2(n7238), .A(n6093), .ZN(n6094) );
  OAI21_X1 U6802 ( .B1(n6113), .B2(n6584), .A(n6094), .ZN(U2994) );
  OAI21_X1 U6803 ( .B1(n6191), .B2(n6095), .A(n6193), .ZN(n6310) );
  NOR2_X1 U6804 ( .A1(n6310), .A2(n7215), .ZN(n6101) );
  NOR2_X1 U6805 ( .A1(n6500), .A2(n6097), .ZN(n6163) );
  INV_X1 U6806 ( .A(n6164), .ZN(n6502) );
  NOR3_X1 U6807 ( .A1(n6163), .A2(n6502), .A3(n6096), .ZN(n6100) );
  NOR3_X1 U6808 ( .A1(n6168), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n6097), 
        .ZN(n6098) );
  NOR4_X1 U6809 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n6102)
         );
  OAI21_X1 U6810 ( .B1(n6103), .B2(n6584), .A(n6102), .ZN(U2989) );
  NAND2_X1 U6811 ( .A1(n6356), .A2(n6106), .ZN(n6265) );
  INV_X1 U6812 ( .A(n6378), .ZN(n6111) );
  NAND2_X1 U6813 ( .A1(n7147), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6108)
         );
  OAI211_X1 U6814 ( .C1(n7152), .C2(n6279), .A(n6109), .B(n6108), .ZN(n6110)
         );
  AOI21_X1 U6815 ( .B1(n6111), .B2(n3628), .A(n6110), .ZN(n6112) );
  OAI21_X1 U6816 ( .B1(n6113), .B2(n7433), .A(n6112), .ZN(U2962) );
  AND2_X1 U6817 ( .A1(n6356), .A2(n6114), .ZN(n6146) );
  AND2_X1 U6818 ( .A1(n6356), .A2(n6115), .ZN(n6154) );
  INV_X1 U6819 ( .A(n6154), .ZN(n6116) );
  AND2_X1 U6820 ( .A1(n6392), .A2(n6118), .ZN(n7535) );
  INV_X1 U6821 ( .A(n6392), .ZN(n7538) );
  AOI22_X1 U6822 ( .A1(n7535), .A2(DATAI_20_), .B1(n7538), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6123) );
  AND2_X1 U6823 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  NAND2_X1 U6824 ( .A1(n7539), .A2(DATAI_4_), .ZN(n6122) );
  OAI211_X1 U6825 ( .C1(n7397), .C2(n6391), .A(n6123), .B(n6122), .ZN(U2871)
         );
  INV_X1 U6826 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7402) );
  INV_X1 U6827 ( .A(n6124), .ZN(n6127) );
  INV_X1 U6828 ( .A(n6132), .ZN(n6126) );
  AOI21_X1 U6829 ( .B1(n6127), .B2(n6126), .A(n6125), .ZN(n6563) );
  INV_X1 U6830 ( .A(n6563), .ZN(n7395) );
  OAI222_X1 U6831 ( .A1(n7397), .A2(n6357), .B1(n7118), .B2(n7402), .C1(n7395), 
        .C2(n7105), .ZN(U2839) );
  INV_X1 U6832 ( .A(n6446), .ZN(n6129) );
  AOI21_X1 U6833 ( .B1(n6131), .B2(n6130), .A(n6129), .ZN(n6151) );
  AOI21_X1 U6834 ( .B1(n6133), .B2(n6334), .A(n6132), .ZN(n7386) );
  AOI21_X1 U6835 ( .B1(n6558), .B2(n6134), .A(n7219), .ZN(n6137) );
  INV_X1 U6836 ( .A(n6135), .ZN(n6136) );
  NOR2_X1 U6837 ( .A1(n6137), .A2(n6136), .ZN(n6556) );
  AND2_X1 U6838 ( .A1(n6558), .A2(n6140), .ZN(n6138) );
  NAND2_X1 U6839 ( .A1(n6578), .A2(n6138), .ZN(n6555) );
  INV_X1 U6840 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7382) );
  NOR2_X1 U6841 ( .A1(n7213), .A2(n7382), .ZN(n6147) );
  INV_X1 U6842 ( .A(n6147), .ZN(n6139) );
  OAI211_X1 U6843 ( .C1(n6556), .C2(n6140), .A(n6555), .B(n6139), .ZN(n6141)
         );
  AOI21_X1 U6844 ( .B1(n7386), .B2(n7238), .A(n6141), .ZN(n6142) );
  OAI21_X1 U6845 ( .B1(n6151), .B2(n6584), .A(n6142), .ZN(U2999) );
  NAND2_X1 U6846 ( .A1(n6356), .A2(n6143), .ZN(n6331) );
  AND2_X1 U6847 ( .A1(n6331), .A2(n6144), .ZN(n6145) );
  AOI21_X1 U6848 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6147), 
        .ZN(n6148) );
  OAI21_X1 U6849 ( .B1(n7389), .B2(n7152), .A(n6148), .ZN(n6149) );
  AOI21_X1 U6850 ( .B1(n7529), .B2(n3628), .A(n6149), .ZN(n6150) );
  OAI21_X1 U6851 ( .B1(n6151), .B2(n7433), .A(n6150), .ZN(U2967) );
  OAI21_X1 U6852 ( .B1(n6154), .B2(n6153), .A(n6323), .ZN(n7108) );
  NAND3_X1 U6853 ( .A1(n6547), .A2(n6546), .A3(n7148), .ZN(n6161) );
  NAND2_X1 U6854 ( .A1(n7205), .A2(REIP_REG_21__SCAN_IN), .ZN(n6548) );
  INV_X1 U6855 ( .A(n6548), .ZN(n6159) );
  NOR2_X1 U6856 ( .A1(n7152), .A2(n7413), .ZN(n6158) );
  AOI211_X1 U6857 ( .C1(n7147), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n6159), 
        .B(n6158), .ZN(n6160) );
  OAI211_X1 U6858 ( .C1(n6489), .C2(n7108), .A(n6161), .B(n6160), .ZN(U2965)
         );
  NOR2_X1 U6859 ( .A1(n6162), .A2(n7215), .ZN(n6172) );
  NAND2_X1 U6860 ( .A1(n6163), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6165) );
  INV_X1 U6861 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6167) );
  AOI21_X1 U6862 ( .B1(n6165), .B2(n6164), .A(n6167), .ZN(n6495) );
  NOR3_X1 U6863 ( .A1(n6495), .A2(n6502), .A3(n6166), .ZN(n6171) );
  NOR4_X1 U6864 ( .A1(n6168), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6167), 
        .A4(n6491), .ZN(n6169) );
  NOR4_X2 U6865 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n6173)
         );
  OAI21_X1 U6866 ( .B1(n6174), .B2(n6584), .A(n6173), .ZN(U2987) );
  NOR2_X1 U6867 ( .A1(n6990), .A2(n6175), .ZN(n6179) );
  INV_X1 U6868 ( .A(n7484), .ZN(n6176) );
  NOR3_X1 U6869 ( .A1(n6177), .A2(n7490), .A3(n6176), .ZN(n6178) );
  AOI211_X1 U6870 ( .C1(n6181), .C2(n6180), .A(n6179), .B(n6178), .ZN(n6182)
         );
  OAI21_X1 U6871 ( .B1(n6184), .B2(n6183), .A(n6182), .ZN(U3465) );
  NAND3_X1 U6872 ( .A1(n6186), .A2(n6185), .A3(n6392), .ZN(n6188) );
  AOI22_X1 U6873 ( .A1(n7535), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7538), .ZN(n6187) );
  NAND2_X1 U6874 ( .A1(n6188), .A2(n6187), .ZN(U2860) );
  XOR2_X1 U6875 ( .A(n6190), .B(n6189), .Z(n6403) );
  INV_X1 U6876 ( .A(n6403), .ZN(n6361) );
  INV_X1 U6877 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6210) );
  AOI22_X1 U6878 ( .A1(n6193), .A2(n5024), .B1(n6192), .B2(n6191), .ZN(n6195)
         );
  XNOR2_X1 U6879 ( .A(n6195), .B(n6194), .ZN(n6490) );
  OAI222_X1 U6880 ( .A1(n6357), .A2(n6361), .B1(n6210), .B2(n7118), .C1(n6490), 
        .C2(n7105), .ZN(U2829) );
  OR2_X1 U6881 ( .A1(n6196), .A2(n6202), .ZN(n6204) );
  NAND2_X1 U6882 ( .A1(n6198), .A2(n6197), .ZN(n6201) );
  AOI22_X1 U6883 ( .A1(n6202), .A2(n6201), .B1(n6200), .B2(n6199), .ZN(n6203)
         );
  AND2_X1 U6884 ( .A1(n6204), .A2(n6203), .ZN(n7448) );
  INV_X1 U6885 ( .A(n7448), .ZN(n6208) );
  NAND2_X1 U6886 ( .A1(n6205), .A2(n7159), .ZN(n7168) );
  NAND2_X1 U6887 ( .A1(n7168), .A2(n7513), .ZN(n6206) );
  AND2_X1 U6888 ( .A1(n6207), .A2(n6206), .ZN(n7445) );
  NOR2_X1 U6889 ( .A1(n7445), .A2(n7499), .ZN(n7434) );
  MUX2_X1 U6890 ( .A(MORE_REG_SCAN_IN), .B(n6208), .S(n7434), .Z(U3471) );
  NAND2_X1 U6891 ( .A1(n6403), .A2(n7428), .ZN(n6215) );
  OAI21_X1 U6892 ( .B1(n6221), .B2(n7065), .A(n7070), .ZN(n6212) );
  AOI22_X1 U6893 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7424), .B1(n7426), 
        .B2(n6399), .ZN(n6209) );
  OAI21_X1 U6894 ( .B1(n7418), .B2(n6210), .A(n6209), .ZN(n6211) );
  AOI21_X1 U6895 ( .B1(n6213), .B2(n6212), .A(n6211), .ZN(n6214) );
  OAI211_X1 U6896 ( .C1(n7431), .C2(n6490), .A(n6215), .B(n6214), .ZN(U2797)
         );
  NAND2_X1 U6897 ( .A1(n6309), .A2(n7428), .ZN(n6224) );
  INV_X1 U6898 ( .A(n6216), .ZN(n6225) );
  OAI22_X1 U6899 ( .A1(n6218), .A2(n7405), .B1(n7412), .B2(n6217), .ZN(n6219)
         );
  AOI21_X1 U6900 ( .B1(n7403), .B2(EBX_REG_29__SCAN_IN), .A(n6219), .ZN(n6220)
         );
  OAI21_X1 U6901 ( .B1(n6221), .B2(REIP_REG_29__SCAN_IN), .A(n6220), .ZN(n6222) );
  AOI21_X1 U6902 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6225), .A(n6222), .ZN(n6223) );
  OAI211_X1 U6903 ( .C1(n7431), .C2(n6310), .A(n6224), .B(n6223), .ZN(U2798)
         );
  INV_X1 U6904 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U6905 ( .B1(REIP_REG_28__SCAN_IN), .B2(n6226), .A(n6225), .ZN(n6229) );
  AOI22_X1 U6906 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n7424), .B1(n7426), 
        .B2(n6227), .ZN(n6228) );
  OAI211_X1 U6907 ( .C1(n6230), .C2(n7418), .A(n6229), .B(n6228), .ZN(n6231)
         );
  AOI21_X1 U6908 ( .B1(n6312), .B2(n7409), .A(n6231), .ZN(n6232) );
  OAI21_X1 U6909 ( .B1(n6367), .B2(n7396), .A(n6232), .ZN(U2799) );
  NAND2_X1 U6910 ( .A1(n6356), .A2(n6233), .ZN(n6247) );
  AOI21_X1 U6911 ( .B1(n6234), .B2(n6247), .A(n6049), .ZN(n6412) );
  INV_X1 U6912 ( .A(n6412), .ZN(n6370) );
  NAND2_X1 U6913 ( .A1(n6252), .A2(n6235), .ZN(n6236) );
  INV_X1 U6914 ( .A(n6238), .ZN(n6257) );
  OAI22_X1 U6915 ( .A1(n6239), .A2(n7405), .B1(n7412), .B2(n6410), .ZN(n6242)
         );
  NOR3_X1 U6916 ( .A1(n7415), .A2(REIP_REG_27__SCAN_IN), .A3(n6240), .ZN(n6241) );
  AOI211_X1 U6917 ( .C1(EBX_REG_27__SCAN_IN), .C2(n7403), .A(n6242), .B(n6241), 
        .ZN(n6243) );
  OAI21_X1 U6918 ( .B1(n7062), .B2(n6257), .A(n6243), .ZN(n6244) );
  AOI21_X1 U6919 ( .B1(n6507), .B2(n7409), .A(n6244), .ZN(n6245) );
  OAI21_X1 U6920 ( .B1(n6370), .B2(n7396), .A(n6245), .ZN(U2800) );
  AND2_X1 U6921 ( .A1(n6356), .A2(n6246), .ZN(n6263) );
  OAI21_X1 U6922 ( .B1(n6263), .B2(n6248), .A(n6247), .ZN(n6418) );
  OR2_X1 U6923 ( .A1(n6249), .A2(n6250), .ZN(n6251) );
  AND2_X1 U6924 ( .A1(n6252), .A2(n6251), .ZN(n6515) );
  INV_X1 U6925 ( .A(n7415), .ZN(n7357) );
  AOI21_X1 U6926 ( .B1(n7357), .B2(n6253), .A(REIP_REG_26__SCAN_IN), .ZN(n6256) );
  AOI22_X1 U6927 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n7424), .B1(n7426), 
        .B2(n6421), .ZN(n6255) );
  NAND2_X1 U6928 ( .A1(n7403), .A2(EBX_REG_26__SCAN_IN), .ZN(n6254) );
  OAI211_X1 U6929 ( .C1(n6257), .C2(n6256), .A(n6255), .B(n6254), .ZN(n6258)
         );
  AOI21_X1 U6930 ( .B1(n6515), .B2(n7409), .A(n6258), .ZN(n6259) );
  OAI21_X1 U6931 ( .B1(n6418), .B2(n7396), .A(n6259), .ZN(U2801) );
  NOR2_X1 U6932 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  OR2_X1 U6933 ( .A1(n6249), .A2(n6262), .ZN(n6523) );
  AOI21_X1 U6934 ( .B1(n6265), .B2(n6264), .A(n6263), .ZN(n6428) );
  NAND2_X1 U6935 ( .A1(n6428), .A2(n7428), .ZN(n6277) );
  INV_X1 U6936 ( .A(n6280), .ZN(n6266) );
  NAND2_X1 U6937 ( .A1(n7390), .A2(n6266), .ZN(n6267) );
  NAND2_X1 U6938 ( .A1(n7358), .A2(n6267), .ZN(n6292) );
  INV_X1 U6939 ( .A(n6292), .ZN(n6275) );
  NAND2_X1 U6940 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6268) );
  OAI21_X1 U6941 ( .B1(REIP_REG_25__SCAN_IN), .B2(n6269), .A(n6268), .ZN(n6273) );
  INV_X1 U6942 ( .A(n6426), .ZN(n6270) );
  AOI22_X1 U6943 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n7424), .B1(n7426), 
        .B2(n6270), .ZN(n6272) );
  NAND2_X1 U6944 ( .A1(n7403), .A2(EBX_REG_25__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U6945 ( .C1(n7415), .C2(n6273), .A(n6272), .B(n6271), .ZN(n6274)
         );
  AOI21_X1 U6946 ( .B1(n6275), .B2(REIP_REG_25__SCAN_IN), .A(n6274), .ZN(n6276) );
  OAI211_X1 U6947 ( .C1(n6523), .C2(n7431), .A(n6277), .B(n6276), .ZN(U2802)
         );
  INV_X1 U6948 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6278) );
  OAI22_X1 U6949 ( .A1(n6279), .A2(n7412), .B1(n7405), .B2(n6278), .ZN(n6282)
         );
  NOR3_X1 U6950 ( .A1(n7415), .A2(REIP_REG_24__SCAN_IN), .A3(n6280), .ZN(n6281) );
  AOI211_X1 U6951 ( .C1(EBX_REG_24__SCAN_IN), .C2(n7403), .A(n6282), .B(n6281), 
        .ZN(n6283) );
  OAI21_X1 U6952 ( .B1(n7054), .B2(n6292), .A(n6283), .ZN(n6284) );
  AOI21_X1 U6953 ( .B1(n6317), .B2(n7409), .A(n6284), .ZN(n6285) );
  OAI21_X1 U6954 ( .B1(n6378), .B2(n7396), .A(n6285), .ZN(U2803) );
  AOI21_X1 U6955 ( .B1(n6287), .B2(n6325), .A(n6286), .ZN(n6438) );
  INV_X1 U6956 ( .A(n6438), .ZN(n6321) );
  INV_X1 U6957 ( .A(n6288), .ZN(n6289) );
  AOI21_X1 U6958 ( .B1(n6290), .B2(n6329), .A(n6289), .ZN(n6534) );
  AOI21_X1 U6959 ( .B1(n7357), .B2(n6291), .A(REIP_REG_23__SCAN_IN), .ZN(n6293) );
  OAI22_X1 U6960 ( .A1(n6293), .A2(n6292), .B1(n4405), .B2(n7405), .ZN(n6295)
         );
  INV_X1 U6961 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6320) );
  OAI22_X1 U6962 ( .A1(n7418), .A2(n6320), .B1(n6436), .B2(n7412), .ZN(n6294)
         );
  AOI211_X1 U6963 ( .C1(n6534), .C2(n7409), .A(n6295), .B(n6294), .ZN(n6296)
         );
  OAI21_X1 U6964 ( .B1(n6321), .B2(n7396), .A(n6296), .ZN(U2804) );
  NAND2_X1 U6965 ( .A1(n6356), .A2(n6297), .ZN(n6347) );
  NAND2_X1 U6966 ( .A1(n6356), .A2(n6355), .ZN(n6354) );
  NAND2_X1 U6967 ( .A1(n6354), .A2(n6298), .ZN(n6299) );
  INV_X1 U6968 ( .A(n7116), .ZN(n6389) );
  AND2_X1 U6969 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NOR2_X1 U6970 ( .A1(n6350), .A2(n6302), .ZN(n7237) );
  INV_X1 U6971 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6303) );
  OAI22_X1 U6972 ( .A1(n7418), .A2(n6303), .B1(n7412), .B2(n6481), .ZN(n6307)
         );
  INV_X1 U6973 ( .A(n6304), .ZN(n7330) );
  NAND2_X1 U6974 ( .A1(n7357), .A2(n7330), .ZN(n7346) );
  OAI21_X1 U6975 ( .B1(n7360), .B2(n6304), .A(n7358), .ZN(n7343) );
  AOI21_X1 U6976 ( .B1(n7424), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7385), 
        .ZN(n6305) );
  OAI221_X1 U6977 ( .B1(REIP_REG_15__SCAN_IN), .B2(n7346), .C1(n7342), .C2(
        n7343), .A(n6305), .ZN(n6306) );
  AOI211_X1 U6978 ( .C1(n7237), .C2(n7409), .A(n6307), .B(n6306), .ZN(n6308)
         );
  OAI21_X1 U6979 ( .B1(n6389), .B2(n7396), .A(n6308), .ZN(U2812) );
  INV_X1 U6980 ( .A(n6309), .ZN(n6364) );
  INV_X1 U6981 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6311) );
  OAI222_X1 U6982 ( .A1(n6357), .A2(n6364), .B1(n6311), .B2(n7118), .C1(n6310), 
        .C2(n7105), .ZN(U2830) );
  AOI22_X1 U6983 ( .A1(n6312), .A2(n7114), .B1(EBX_REG_28__SCAN_IN), .B2(n6338), .ZN(n6313) );
  OAI21_X1 U6984 ( .B1(n6367), .B2(n6357), .A(n6313), .ZN(U2831) );
  AOI22_X1 U6985 ( .A1(n6507), .A2(n7114), .B1(EBX_REG_27__SCAN_IN), .B2(n6338), .ZN(n6314) );
  OAI21_X1 U6986 ( .B1(n6370), .B2(n6357), .A(n6314), .ZN(U2832) );
  AOI22_X1 U6987 ( .A1(n6515), .A2(n7114), .B1(EBX_REG_26__SCAN_IN), .B2(n6338), .ZN(n6315) );
  OAI21_X1 U6988 ( .B1(n6418), .B2(n6357), .A(n6315), .ZN(U2833) );
  INV_X1 U6989 ( .A(n6428), .ZN(n6375) );
  INV_X1 U6990 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6316) );
  OAI222_X1 U6991 ( .A1(n6375), .A2(n6357), .B1(n6316), .B2(n7118), .C1(n6523), 
        .C2(n7105), .ZN(U2834) );
  AOI22_X1 U6992 ( .A1(n6317), .A2(n7114), .B1(EBX_REG_24__SCAN_IN), .B2(n6338), .ZN(n6318) );
  OAI21_X1 U6993 ( .B1(n6378), .B2(n6357), .A(n6318), .ZN(U2835) );
  INV_X1 U6994 ( .A(n6534), .ZN(n6319) );
  OAI222_X1 U6995 ( .A1(n6357), .A2(n6321), .B1(n6320), .B2(n7118), .C1(n6319), 
        .C2(n7105), .ZN(U2836) );
  NAND2_X1 U6996 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U6997 ( .A1(n6325), .A2(n6324), .ZN(n7425) );
  INV_X1 U6998 ( .A(EBX_REG_22__SCAN_IN), .ZN(n7419) );
  OR2_X1 U6999 ( .A1(n6326), .A2(n6327), .ZN(n6328) );
  NAND2_X1 U7000 ( .A1(n6329), .A2(n6328), .ZN(n7432) );
  OAI222_X1 U7001 ( .A1(n6357), .A2(n7425), .B1(n7118), .B2(n7419), .C1(n7432), 
        .C2(n7105), .ZN(U2837) );
  NAND2_X1 U7002 ( .A1(n6356), .A2(n6330), .ZN(n6343) );
  INV_X1 U7003 ( .A(n6331), .ZN(n6332) );
  AOI21_X1 U7004 ( .B1(n6333), .B2(n6343), .A(n6332), .ZN(n6461) );
  INV_X1 U7005 ( .A(n6461), .ZN(n7373) );
  INV_X1 U7006 ( .A(n6334), .ZN(n6335) );
  AOI21_X1 U7007 ( .B1(n6337), .B2(n6336), .A(n6335), .ZN(n7371) );
  AOI22_X1 U7008 ( .A1(n7371), .A2(n7114), .B1(EBX_REG_18__SCAN_IN), .B2(n6338), .ZN(n6339) );
  OAI21_X1 U7009 ( .B1(n7373), .B2(n6357), .A(n6339), .ZN(U2841) );
  AND2_X1 U7010 ( .A1(n6356), .A2(n6340), .ZN(n6346) );
  OR2_X1 U7011 ( .A1(n6346), .A2(n6341), .ZN(n6342) );
  INV_X1 U7012 ( .A(n7526), .ZN(n6345) );
  INV_X1 U7013 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6344) );
  OAI222_X1 U7014 ( .A1(n6345), .A2(n6357), .B1(n6344), .B2(n7118), .C1(n7105), 
        .C2(n7363), .ZN(U2842) );
  OR2_X1 U7015 ( .A1(n6350), .A2(n6349), .ZN(n6351) );
  NAND2_X1 U7016 ( .A1(n5893), .A2(n6351), .ZN(n7349) );
  OAI22_X1 U7017 ( .A1(n7349), .A2(n7105), .B1(n7355), .B2(n7118), .ZN(n6352)
         );
  AOI21_X1 U7018 ( .B1(n7348), .B2(n7115), .A(n6352), .ZN(n6353) );
  INV_X1 U7019 ( .A(n6353), .ZN(U2843) );
  INV_X1 U7020 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U7021 ( .B1(n6356), .B2(n6355), .A(n6354), .ZN(n7335) );
  OAI222_X1 U7022 ( .A1(n7341), .A2(n7105), .B1(n7118), .B2(n6358), .C1(n7335), 
        .C2(n6357), .ZN(U2845) );
  AOI22_X1 U7023 ( .A1(n7535), .A2(DATAI_30_), .B1(n7538), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7024 ( .A1(n7539), .A2(DATAI_14_), .ZN(n6359) );
  OAI211_X1 U7025 ( .C1(n6361), .C2(n6391), .A(n6360), .B(n6359), .ZN(U2861)
         );
  AOI22_X1 U7026 ( .A1(n7535), .A2(DATAI_29_), .B1(n7538), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U7027 ( .A1(n7539), .A2(DATAI_13_), .ZN(n6362) );
  OAI211_X1 U7028 ( .C1(n6364), .C2(n6391), .A(n6363), .B(n6362), .ZN(U2862)
         );
  AOI22_X1 U7029 ( .A1(n7535), .A2(DATAI_28_), .B1(n7538), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U7030 ( .A1(n7539), .A2(DATAI_12_), .ZN(n6365) );
  OAI211_X1 U7031 ( .C1(n6367), .C2(n6391), .A(n6366), .B(n6365), .ZN(U2863)
         );
  AOI22_X1 U7032 ( .A1(n7535), .A2(DATAI_27_), .B1(n7538), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U7033 ( .A1(n7539), .A2(DATAI_11_), .ZN(n6368) );
  OAI211_X1 U7034 ( .C1(n6370), .C2(n6391), .A(n6369), .B(n6368), .ZN(U2864)
         );
  AOI22_X1 U7035 ( .A1(n7535), .A2(DATAI_26_), .B1(n7538), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7036 ( .A1(n7539), .A2(DATAI_10_), .ZN(n6371) );
  OAI211_X1 U7037 ( .C1(n6418), .C2(n6391), .A(n6372), .B(n6371), .ZN(U2865)
         );
  AOI22_X1 U7038 ( .A1(n7535), .A2(DATAI_25_), .B1(n7538), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7039 ( .A1(n7539), .A2(DATAI_9_), .ZN(n6373) );
  OAI211_X1 U7040 ( .C1(n6375), .C2(n6391), .A(n6374), .B(n6373), .ZN(U2866)
         );
  AOI22_X1 U7041 ( .A1(n7535), .A2(DATAI_24_), .B1(n7538), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U7042 ( .A1(n7539), .A2(DATAI_8_), .ZN(n6376) );
  OAI211_X1 U7043 ( .C1(n6378), .C2(n6391), .A(n6377), .B(n6376), .ZN(U2867)
         );
  INV_X1 U7044 ( .A(n7539), .ZN(n6388) );
  INV_X1 U7045 ( .A(n6391), .ZN(n7536) );
  NAND2_X1 U7046 ( .A1(n6438), .A2(n7536), .ZN(n6380) );
  AOI22_X1 U7047 ( .A1(n7535), .A2(DATAI_23_), .B1(n7538), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6379) );
  OAI211_X1 U7048 ( .C1(n6388), .C2(n6381), .A(n6380), .B(n6379), .ZN(U2868)
         );
  NAND2_X1 U7049 ( .A1(n6461), .A2(n7536), .ZN(n6383) );
  AOI22_X1 U7050 ( .A1(n7535), .A2(DATAI_18_), .B1(n7538), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6382) );
  OAI211_X1 U7051 ( .C1(n6388), .C2(n6384), .A(n6383), .B(n6382), .ZN(U2873)
         );
  NAND2_X1 U7052 ( .A1(n7348), .A2(n7536), .ZN(n6386) );
  AOI22_X1 U7053 ( .A1(n7535), .A2(DATAI_16_), .B1(n7538), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6385) );
  OAI211_X1 U7054 ( .C1(n6388), .C2(n6387), .A(n6386), .B(n6385), .ZN(U2875)
         );
  INV_X1 U7055 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7025) );
  OAI222_X1 U7056 ( .A1(n6390), .A2(n6394), .B1(n6392), .B2(n7025), .C1(n6391), 
        .C2(n6389), .ZN(U2876) );
  INV_X1 U7057 ( .A(DATAI_14_), .ZN(n6393) );
  INV_X1 U7058 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7021) );
  OAI222_X1 U7059 ( .A1(n6394), .A2(n6393), .B1(n6392), .B2(n7021), .C1(n6391), 
        .C2(n7335), .ZN(U2877) );
  NOR2_X1 U7060 ( .A1(n6395), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6397)
         );
  MUX2_X1 U7061 ( .A(n4049), .B(n6397), .S(n6396), .Z(n6398) );
  XNOR2_X1 U7062 ( .A(n6398), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6499)
         );
  NAND2_X1 U7063 ( .A1(n7143), .A2(n6399), .ZN(n6400) );
  NAND2_X1 U7064 ( .A1(n7205), .A2(REIP_REG_30__SCAN_IN), .ZN(n6493) );
  OAI211_X1 U7065 ( .C1(n7132), .C2(n6401), .A(n6400), .B(n6493), .ZN(n6402)
         );
  AOI21_X1 U7066 ( .B1(n6403), .B2(n3628), .A(n6402), .ZN(n6404) );
  OAI21_X1 U7067 ( .B1(n6499), .B2(n7433), .A(n6404), .ZN(U2956) );
  NAND2_X1 U7068 ( .A1(n6406), .A2(n6405), .ZN(n6408) );
  XNOR2_X1 U7069 ( .A(n6395), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6407)
         );
  XNOR2_X1 U7070 ( .A(n6408), .B(n6407), .ZN(n6510) );
  NOR2_X1 U7071 ( .A1(n7213), .A2(n7062), .ZN(n6504) );
  AOI21_X1 U7072 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6504), 
        .ZN(n6409) );
  OAI21_X1 U7073 ( .B1(n7152), .B2(n6410), .A(n6409), .ZN(n6411) );
  AOI21_X1 U7074 ( .B1(n6412), .B2(n3628), .A(n6411), .ZN(n6413) );
  OAI21_X1 U7075 ( .B1(n6510), .B2(n7433), .A(n6413), .ZN(U2959) );
  XNOR2_X1 U7076 ( .A(n6395), .B(n6414), .ZN(n6415) );
  XNOR2_X1 U7077 ( .A(n6416), .B(n6415), .ZN(n6518) );
  NAND2_X1 U7078 ( .A1(n7205), .A2(REIP_REG_26__SCAN_IN), .ZN(n6512) );
  OAI21_X1 U7079 ( .B1(n7132), .B2(n6417), .A(n6512), .ZN(n6420) );
  NOR2_X1 U7080 ( .A1(n6418), .A2(n6489), .ZN(n6419) );
  AOI211_X1 U7081 ( .C1(n6421), .C2(n7143), .A(n6420), .B(n6419), .ZN(n6422)
         );
  OAI21_X1 U7082 ( .B1(n7433), .B2(n6518), .A(n6422), .ZN(U2960) );
  XNOR2_X1 U7083 ( .A(n6477), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6423)
         );
  XNOR2_X1 U7084 ( .A(n6424), .B(n6423), .ZN(n6527) );
  NAND2_X1 U7085 ( .A1(n7205), .A2(REIP_REG_25__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U7086 ( .A1(n7147), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6425)
         );
  OAI211_X1 U7087 ( .C1(n7152), .C2(n6426), .A(n6519), .B(n6425), .ZN(n6427)
         );
  AOI21_X1 U7088 ( .B1(n6428), .B2(n3628), .A(n6427), .ZN(n6429) );
  OAI21_X1 U7089 ( .B1(n6527), .B2(n7433), .A(n6429), .ZN(U2961) );
  NOR2_X1 U7090 ( .A1(n6431), .A2(n6430), .ZN(n6433) );
  MUX2_X1 U7091 ( .A(n6433), .B(n6432), .S(n6447), .Z(n6434) );
  XNOR2_X1 U7092 ( .A(n6434), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6536)
         );
  INV_X1 U7093 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7053) );
  NOR2_X1 U7094 ( .A1(n7213), .A2(n7053), .ZN(n6528) );
  AOI21_X1 U7095 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6528), 
        .ZN(n6435) );
  OAI21_X1 U7096 ( .B1(n6436), .B2(n7152), .A(n6435), .ZN(n6437) );
  AOI21_X1 U7097 ( .B1(n6438), .B2(n3628), .A(n6437), .ZN(n6439) );
  OAI21_X1 U7098 ( .B1(n6536), .B2(n7433), .A(n6439), .ZN(U2963) );
  XNOR2_X1 U7099 ( .A(n6395), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6440)
         );
  XNOR2_X1 U7100 ( .A(n6441), .B(n6440), .ZN(n6543) );
  INV_X1 U7101 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U7102 ( .A1(n7205), .A2(REIP_REG_22__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U7103 ( .B1(n7132), .B2(n6442), .A(n6537), .ZN(n6444) );
  NOR2_X1 U7104 ( .A1(n7425), .A2(n6489), .ZN(n6443) );
  AOI211_X1 U7105 ( .C1(n7143), .C2(n7427), .A(n6444), .B(n6443), .ZN(n6445)
         );
  OAI21_X1 U7106 ( .B1(n6543), .B2(n7433), .A(n6445), .ZN(U2964) );
  OAI21_X1 U7107 ( .B1(n6447), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6446), 
        .ZN(n6449) );
  XNOR2_X1 U7108 ( .A(n6447), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6448)
         );
  XNOR2_X1 U7109 ( .A(n6449), .B(n6448), .ZN(n6565) );
  NAND2_X1 U7110 ( .A1(n7205), .A2(REIP_REG_20__SCAN_IN), .ZN(n6559) );
  OAI21_X1 U7111 ( .B1(n7132), .B2(n6450), .A(n6559), .ZN(n6452) );
  NOR2_X1 U7112 ( .A1(n7397), .A2(n6489), .ZN(n6451) );
  AOI211_X1 U7113 ( .C1(n7143), .C2(n7399), .A(n6452), .B(n6451), .ZN(n6453)
         );
  OAI21_X1 U7114 ( .B1(n7433), .B2(n6565), .A(n6453), .ZN(U2966) );
  NOR2_X1 U7115 ( .A1(n6454), .A2(n5881), .ZN(n6457) );
  NOR2_X1 U7116 ( .A1(n6455), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6456)
         );
  MUX2_X1 U7117 ( .A(n6457), .B(n6456), .S(n6447), .Z(n6458) );
  XNOR2_X1 U7118 ( .A(n6458), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6574)
         );
  INV_X1 U7119 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7379) );
  NOR2_X1 U7120 ( .A1(n7213), .A2(n7379), .ZN(n6571) );
  NOR2_X1 U7121 ( .A1(n7132), .A2(n6459), .ZN(n6460) );
  AOI211_X1 U7122 ( .C1(n7143), .C2(n7375), .A(n6571), .B(n6460), .ZN(n6463)
         );
  NAND2_X1 U7123 ( .A1(n6461), .A2(n3628), .ZN(n6462) );
  OAI211_X1 U7124 ( .C1(n6574), .C2(n7433), .A(n6463), .B(n6462), .ZN(U2968)
         );
  NAND2_X1 U7125 ( .A1(n6465), .A2(n6464), .ZN(n6476) );
  AND2_X1 U7126 ( .A1(n6476), .A2(n6466), .ZN(n6468) );
  NOR2_X1 U7127 ( .A1(n6468), .A2(n6467), .ZN(n6470) );
  MUX2_X1 U7128 ( .A(n5887), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .S(n4049), 
        .Z(n6469) );
  XNOR2_X1 U7129 ( .A(n6470), .B(n6469), .ZN(n6585) );
  NOR2_X1 U7130 ( .A1(n7213), .A2(n7344), .ZN(n6576) );
  AOI21_X1 U7131 ( .B1(n7147), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6576), 
        .ZN(n6471) );
  OAI21_X1 U7132 ( .B1(n6472), .B2(n7152), .A(n6471), .ZN(n6473) );
  AOI21_X1 U7133 ( .B1(n7348), .B2(n3628), .A(n6473), .ZN(n6474) );
  OAI21_X1 U7134 ( .B1(n6585), .B2(n7433), .A(n6474), .ZN(U2970) );
  AND2_X1 U7135 ( .A1(n6476), .A2(n6475), .ZN(n6479) );
  XNOR2_X1 U7136 ( .A(n6477), .B(n6580), .ZN(n6478) );
  XNOR2_X1 U7137 ( .A(n6479), .B(n6478), .ZN(n7236) );
  AOI22_X1 U7138 ( .A1(n7147), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n7205), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n6480) );
  OAI21_X1 U7139 ( .B1(n7152), .B2(n6481), .A(n6480), .ZN(n6482) );
  AOI21_X1 U7140 ( .B1(n7116), .B2(n3628), .A(n6482), .ZN(n6483) );
  OAI21_X1 U7141 ( .B1(n7236), .B2(n7433), .A(n6483), .ZN(U2971) );
  NAND2_X1 U7142 ( .A1(n6484), .A2(n7148), .ZN(n6488) );
  NOR2_X1 U7143 ( .A1(n7152), .A2(n7336), .ZN(n6485) );
  AOI211_X1 U7144 ( .C1(n7147), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6486), 
        .B(n6485), .ZN(n6487) );
  OAI211_X1 U7145 ( .C1(n6489), .C2(n7335), .A(n6488), .B(n6487), .ZN(U2972)
         );
  INV_X1 U7146 ( .A(n6490), .ZN(n6497) );
  INV_X1 U7147 ( .A(n6491), .ZN(n6492) );
  AOI21_X1 U7148 ( .B1(n6506), .B2(n6492), .A(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n6494) );
  OAI21_X1 U7149 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(n6496) );
  AOI21_X1 U7150 ( .B1(n6497), .B2(n7238), .A(n6496), .ZN(n6498) );
  OAI21_X1 U7151 ( .B1(n6499), .B2(n6584), .A(n6498), .ZN(U2988) );
  INV_X1 U7152 ( .A(n6500), .ZN(n6501) );
  NOR3_X1 U7153 ( .A1(n6502), .A2(n6501), .A3(n6505), .ZN(n6503) );
  AOI211_X1 U7154 ( .C1(n6506), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6509)
         );
  NAND2_X1 U7155 ( .A1(n6507), .A2(n7238), .ZN(n6508) );
  OAI211_X1 U7156 ( .C1(n6510), .C2(n6584), .A(n6509), .B(n6508), .ZN(U2991)
         );
  INV_X1 U7157 ( .A(n6511), .ZN(n6522) );
  XNOR2_X1 U7158 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6513) );
  OAI21_X1 U7159 ( .B1(n6520), .B2(n6513), .A(n6512), .ZN(n6514) );
  AOI21_X1 U7160 ( .B1(n6522), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6514), 
        .ZN(n6517) );
  NAND2_X1 U7161 ( .A1(n6515), .A2(n7238), .ZN(n6516) );
  OAI211_X1 U7162 ( .C1(n6518), .C2(n6584), .A(n6517), .B(n6516), .ZN(U2992)
         );
  OAI21_X1 U7163 ( .B1(n6520), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6519), 
        .ZN(n6521) );
  AOI21_X1 U7164 ( .B1(n6522), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6521), 
        .ZN(n6526) );
  INV_X1 U7165 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U7166 ( .A1(n6524), .A2(n7238), .ZN(n6525) );
  OAI211_X1 U7167 ( .C1(n6527), .C2(n6584), .A(n6526), .B(n6525), .ZN(U2993)
         );
  INV_X1 U7168 ( .A(n6541), .ZN(n6532) );
  AOI21_X1 U7169 ( .B1(n6529), .B2(n6531), .A(n6528), .ZN(n6530) );
  OAI21_X1 U7170 ( .B1(n6532), .B2(n6531), .A(n6530), .ZN(n6533) );
  AOI21_X1 U7171 ( .B1(n6534), .B2(n7238), .A(n6533), .ZN(n6535) );
  OAI21_X1 U7172 ( .B1(n6536), .B2(n6584), .A(n6535), .ZN(U2995) );
  OAI21_X1 U7173 ( .B1(n6538), .B2(n6551), .A(n6537), .ZN(n6540) );
  NOR2_X1 U7174 ( .A1(n7432), .A2(n7215), .ZN(n6539) );
  AOI211_X1 U7175 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n6541), .A(n6540), .B(n6539), .ZN(n6542) );
  OAI21_X1 U7176 ( .B1(n6543), .B2(n6584), .A(n6542), .ZN(U2996) );
  NOR2_X1 U7177 ( .A1(n6125), .A2(n6544), .ZN(n6545) );
  OR2_X1 U7178 ( .A1(n6326), .A2(n6545), .ZN(n7109) );
  NAND3_X1 U7179 ( .A1(n6547), .A2(n6546), .A3(n7239), .ZN(n6554) );
  OAI21_X1 U7180 ( .B1(n6549), .B2(n6551), .A(n6548), .ZN(n6550) );
  AOI21_X1 U7181 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(n6553) );
  OAI211_X1 U7182 ( .C1(n7215), .C2(n7109), .A(n6554), .B(n6553), .ZN(U2997)
         );
  AOI21_X1 U7183 ( .B1(n6556), .B2(n6555), .A(n6557), .ZN(n6562) );
  NAND4_X1 U7184 ( .A1(n6578), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n6558), .A4(n6557), .ZN(n6560) );
  NAND2_X1 U7185 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  AOI211_X1 U7186 ( .C1(n6563), .C2(n7238), .A(n6562), .B(n6561), .ZN(n6564)
         );
  OAI21_X1 U7187 ( .B1(n6565), .B2(n6584), .A(n6564), .ZN(U2998) );
  INV_X1 U7188 ( .A(n6566), .ZN(n6946) );
  OAI221_X1 U7189 ( .B1(n6568), .B2(n6946), .C1(n6568), .C2(n6567), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6573) );
  NOR4_X1 U7190 ( .A1(n6949), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5881), 
        .A4(n6569), .ZN(n6570) );
  AOI211_X1 U7191 ( .C1(n7371), .C2(n7238), .A(n6571), .B(n6570), .ZN(n6572)
         );
  OAI211_X1 U7192 ( .C1(n6574), .C2(n6584), .A(n6573), .B(n6572), .ZN(U3000)
         );
  OAI21_X1 U7193 ( .B1(n6579), .B2(n7219), .A(n6575), .ZN(n7235) );
  INV_X1 U7194 ( .A(n6576), .ZN(n6577) );
  OAI21_X1 U7195 ( .B1(n7349), .B2(n7215), .A(n6577), .ZN(n6582) );
  NAND2_X1 U7196 ( .A1(n6579), .A2(n6578), .ZN(n7243) );
  AOI221_X1 U7197 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n5887), .C2(n6580), .A(n7243), 
        .ZN(n6581) );
  AOI211_X1 U7198 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n7235), .A(n6582), .B(n6581), .ZN(n6583) );
  OAI21_X1 U7199 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(U3002) );
  XNOR2_X1 U7200 ( .A(DATAI_30_), .B(keyinput_129), .ZN(n6588) );
  XNOR2_X1 U7201 ( .A(DATAI_29_), .B(keyinput_130), .ZN(n6587) );
  XNOR2_X1 U7202 ( .A(DATAI_31_), .B(keyinput_128), .ZN(n6586) );
  NOR3_X1 U7203 ( .A1(n6588), .A2(n6587), .A3(n6586), .ZN(n6592) );
  XOR2_X1 U7204 ( .A(DATAI_28_), .B(keyinput_131), .Z(n6591) );
  XNOR2_X1 U7205 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n6590) );
  XNOR2_X1 U7206 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n6589) );
  OAI211_X1 U7207 ( .C1(n6592), .C2(n6591), .A(n6590), .B(n6589), .ZN(n6595)
         );
  XOR2_X1 U7208 ( .A(DATAI_25_), .B(keyinput_134), .Z(n6594) );
  XNOR2_X1 U7209 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n6593) );
  AOI21_X1 U7210 ( .B1(n6595), .B2(n6594), .A(n6593), .ZN(n6598) );
  XOR2_X1 U7211 ( .A(DATAI_22_), .B(keyinput_137), .Z(n6597) );
  XOR2_X1 U7212 ( .A(DATAI_23_), .B(keyinput_136), .Z(n6596) );
  NOR3_X1 U7213 ( .A1(n6598), .A2(n6597), .A3(n6596), .ZN(n6607) );
  XOR2_X1 U7214 ( .A(DATAI_21_), .B(keyinput_138), .Z(n6606) );
  XOR2_X1 U7215 ( .A(DATAI_20_), .B(keyinput_139), .Z(n6601) );
  XNOR2_X1 U7216 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n6600) );
  XNOR2_X1 U7217 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n6599) );
  NAND3_X1 U7218 ( .A1(n6601), .A2(n6600), .A3(n6599), .ZN(n6604) );
  XOR2_X1 U7219 ( .A(DATAI_18_), .B(keyinput_141), .Z(n6603) );
  XNOR2_X1 U7220 ( .A(DATAI_17_), .B(keyinput_142), .ZN(n6602) );
  NOR3_X1 U7221 ( .A1(n6604), .A2(n6603), .A3(n6602), .ZN(n6605) );
  OAI21_X1 U7222 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6610) );
  XNOR2_X1 U7223 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n6609) );
  XNOR2_X1 U7224 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n6608) );
  AOI21_X1 U7225 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(n6613) );
  XOR2_X1 U7226 ( .A(DATAI_13_), .B(keyinput_146), .Z(n6612) );
  XOR2_X1 U7227 ( .A(DATAI_12_), .B(keyinput_147), .Z(n6611) );
  OAI21_X1 U7228 ( .B1(n6613), .B2(n6612), .A(n6611), .ZN(n6617) );
  XNOR2_X1 U7229 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n6616) );
  XOR2_X1 U7230 ( .A(DATAI_9_), .B(keyinput_150), .Z(n6615) );
  XNOR2_X1 U7231 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n6614) );
  AOI211_X1 U7232 ( .C1(n6617), .C2(n6616), .A(n6615), .B(n6614), .ZN(n6620)
         );
  XOR2_X1 U7233 ( .A(DATAI_8_), .B(keyinput_151), .Z(n6619) );
  XOR2_X1 U7234 ( .A(DATAI_7_), .B(keyinput_152), .Z(n6618) );
  NOR3_X1 U7235 ( .A1(n6620), .A2(n6619), .A3(n6618), .ZN(n6623) );
  XNOR2_X1 U7236 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n6622) );
  XNOR2_X1 U7237 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n6621) );
  NOR3_X1 U7238 ( .A1(n6623), .A2(n6622), .A3(n6621), .ZN(n6626) );
  XOR2_X1 U7239 ( .A(DATAI_4_), .B(keyinput_155), .Z(n6625) );
  XOR2_X1 U7240 ( .A(DATAI_3_), .B(keyinput_156), .Z(n6624) );
  OAI21_X1 U7241 ( .B1(n6626), .B2(n6625), .A(n6624), .ZN(n6630) );
  XOR2_X1 U7242 ( .A(DATAI_2_), .B(keyinput_157), .Z(n6629) );
  XNOR2_X1 U7243 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n6628) );
  XNOR2_X1 U7244 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n6627) );
  AOI211_X1 U7245 ( .C1(n6630), .C2(n6629), .A(n6628), .B(n6627), .ZN(n6634)
         );
  XOR2_X1 U7246 ( .A(NA_N), .B(keyinput_161), .Z(n6633) );
  XOR2_X1 U7247 ( .A(BS16_N), .B(keyinput_162), .Z(n6632) );
  XNOR2_X1 U7248 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_160), .ZN(n6631)
         );
  NOR4_X1 U7249 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6638)
         );
  XNOR2_X1 U7250 ( .A(n7513), .B(keyinput_163), .ZN(n6637) );
  XOR2_X1 U7251 ( .A(HOLD), .B(keyinput_164), .Z(n6636) );
  XNOR2_X1 U7252 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_165), .ZN(n6635)
         );
  OAI211_X1 U7253 ( .C1(n6638), .C2(n6637), .A(n6636), .B(n6635), .ZN(n6641)
         );
  XOR2_X1 U7254 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_167), .Z(n6640) );
  XNOR2_X1 U7255 ( .A(ADS_N_REG_SCAN_IN), .B(keyinput_166), .ZN(n6639) );
  NAND3_X1 U7256 ( .A1(n6641), .A2(n6640), .A3(n6639), .ZN(n6644) );
  INV_X1 U7257 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7523) );
  XNOR2_X1 U7258 ( .A(n7523), .B(keyinput_168), .ZN(n6643) );
  XNOR2_X1 U7259 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_169), .ZN(n6642) );
  AOI21_X1 U7260 ( .B1(n6644), .B2(n6643), .A(n6642), .ZN(n6650) );
  XNOR2_X1 U7261 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_170), .ZN(n6649) );
  XOR2_X1 U7262 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_173), .Z(n6647) );
  XNOR2_X1 U7263 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_171), .ZN(n6646) );
  XNOR2_X1 U7264 ( .A(MORE_REG_SCAN_IN), .B(keyinput_172), .ZN(n6645) );
  NOR3_X1 U7265 ( .A1(n6647), .A2(n6646), .A3(n6645), .ZN(n6648) );
  OAI21_X1 U7266 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(n6654) );
  XOR2_X1 U7267 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_175), .Z(n6653)
         );
  INV_X1 U7268 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7093) );
  XNOR2_X1 U7269 ( .A(n7093), .B(keyinput_176), .ZN(n6652) );
  XNOR2_X1 U7270 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_174), .ZN(n6651) );
  NAND4_X1 U7271 ( .A1(n6654), .A2(n6653), .A3(n6652), .A4(n6651), .ZN(n6658)
         );
  XOR2_X1 U7272 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .Z(n6657) );
  INV_X1 U7273 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7089) );
  XNOR2_X1 U7274 ( .A(n7089), .B(keyinput_177), .ZN(n6656) );
  XNOR2_X1 U7275 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_178), .ZN(n6655)
         );
  NAND4_X1 U7276 ( .A1(n6658), .A2(n6657), .A3(n6656), .A4(n6655), .ZN(n6664)
         );
  INV_X1 U7277 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7060) );
  OAI22_X1 U7278 ( .A1(n7060), .A2(keyinput_184), .B1(REIP_REG_28__SCAN_IN), 
        .B2(keyinput_182), .ZN(n6659) );
  AOI221_X1 U7279 ( .B1(n7060), .B2(keyinput_184), .C1(keyinput_182), .C2(
        REIP_REG_28__SCAN_IN), .A(n6659), .ZN(n6663) );
  XOR2_X1 U7280 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_181), .Z(n6662) );
  OAI22_X1 U7281 ( .A1(n7070), .A2(keyinput_180), .B1(n7062), .B2(keyinput_183), .ZN(n6660) );
  AOI221_X1 U7282 ( .B1(n7070), .B2(keyinput_180), .C1(keyinput_183), .C2(
        n7062), .A(n6660), .ZN(n6661) );
  NAND4_X1 U7283 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6668)
         );
  XNOR2_X1 U7284 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .ZN(n6667) );
  XOR2_X1 U7285 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .Z(n6666) );
  XNOR2_X1 U7286 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n6665) );
  AOI211_X1 U7287 ( .C1(n6668), .C2(n6667), .A(n6666), .B(n6665), .ZN(n6672)
         );
  XNOR2_X1 U7288 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .ZN(n6671) );
  XNOR2_X1 U7289 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .ZN(n6670) );
  XNOR2_X1 U7290 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .ZN(n6669) );
  NOR4_X1 U7291 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6675)
         );
  XNOR2_X1 U7292 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .ZN(n6674) );
  XOR2_X1 U7293 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .Z(n6673) );
  OAI21_X1 U7294 ( .B1(n6675), .B2(n6674), .A(n6673), .ZN(n6679) );
  XOR2_X1 U7295 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .Z(n6678) );
  XNOR2_X1 U7296 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_195), .ZN(n6677) );
  XNOR2_X1 U7297 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .ZN(n6676) );
  NAND4_X1 U7298 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6681)
         );
  XNOR2_X1 U7299 ( .A(BE_N_REG_2__SCAN_IN), .B(keyinput_196), .ZN(n6680) );
  NAND2_X1 U7300 ( .A1(n6681), .A2(n6680), .ZN(n6685) );
  XOR2_X1 U7301 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_197), .Z(n6684) );
  XOR2_X1 U7302 ( .A(ADDRESS_REG_29__SCAN_IN), .B(keyinput_199), .Z(n6683) );
  XNOR2_X1 U7303 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_198), .ZN(n6682) );
  NAND4_X1 U7304 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6695)
         );
  INV_X1 U7305 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7063) );
  XNOR2_X1 U7306 ( .A(n7063), .B(keyinput_201), .ZN(n6689) );
  INV_X1 U7307 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7066) );
  XNOR2_X1 U7308 ( .A(n7066), .B(keyinput_200), .ZN(n6688) );
  INV_X1 U7309 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7061) );
  XNOR2_X1 U7310 ( .A(n7061), .B(keyinput_202), .ZN(n6687) );
  XNOR2_X1 U7311 ( .A(ADDRESS_REG_25__SCAN_IN), .B(keyinput_203), .ZN(n6686)
         );
  NOR4_X1 U7312 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6694)
         );
  XNOR2_X1 U7313 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_204), .ZN(n6693)
         );
  XNOR2_X1 U7314 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_205), .ZN(n6691)
         );
  XNOR2_X1 U7315 ( .A(ADDRESS_REG_22__SCAN_IN), .B(keyinput_206), .ZN(n6690)
         );
  NAND2_X1 U7316 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  AOI211_X1 U7317 ( .C1(n6695), .C2(n6694), .A(n6693), .B(n6692), .ZN(n6701)
         );
  XNOR2_X1 U7318 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_207), .ZN(n6700)
         );
  INV_X1 U7319 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7048) );
  XNOR2_X1 U7320 ( .A(n7048), .B(keyinput_209), .ZN(n6698) );
  INV_X1 U7321 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7047) );
  XNOR2_X1 U7322 ( .A(n7047), .B(keyinput_210), .ZN(n6697) );
  XNOR2_X1 U7323 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_208), .ZN(n6696)
         );
  NOR3_X1 U7324 ( .A1(n6698), .A2(n6697), .A3(n6696), .ZN(n6699) );
  OAI21_X1 U7325 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(n6704) );
  INV_X1 U7326 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7046) );
  XNOR2_X1 U7327 ( .A(n7046), .B(keyinput_211), .ZN(n6703) );
  XNOR2_X1 U7328 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_212), .ZN(n6702)
         );
  NAND3_X1 U7329 ( .A1(n6704), .A2(n6703), .A3(n6702), .ZN(n6707) );
  XOR2_X1 U7330 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_213), .Z(n6706) );
  XNOR2_X1 U7331 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_214), .ZN(n6705)
         );
  NAND3_X1 U7332 ( .A1(n6707), .A2(n6706), .A3(n6705), .ZN(n6710) );
  INV_X1 U7333 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7042) );
  XNOR2_X1 U7334 ( .A(n7042), .B(keyinput_215), .ZN(n6709) );
  XNOR2_X1 U7335 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_216), .ZN(n6708)
         );
  AOI21_X1 U7336 ( .B1(n6710), .B2(n6709), .A(n6708), .ZN(n6716) );
  INV_X1 U7337 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7034) );
  INV_X1 U7338 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7339 ( .A1(n7034), .A2(keyinput_221), .B1(keyinput_220), .B2(n7036), .ZN(n6711) );
  OAI221_X1 U7340 ( .B1(n7034), .B2(keyinput_221), .C1(n7036), .C2(
        keyinput_220), .A(n6711), .ZN(n6715) );
  INV_X1 U7341 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7040) );
  AOI22_X1 U7342 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(keyinput_218), .B1(n7040), 
        .B2(keyinput_217), .ZN(n6712) );
  OAI221_X1 U7343 ( .B1(ADDRESS_REG_10__SCAN_IN), .B2(keyinput_218), .C1(n7040), .C2(keyinput_217), .A(n6712), .ZN(n6714) );
  XNOR2_X1 U7344 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_219), .ZN(n6713) );
  NOR4_X1 U7345 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6719)
         );
  INV_X1 U7346 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7033) );
  XNOR2_X1 U7347 ( .A(n7033), .B(keyinput_222), .ZN(n6718) );
  INV_X1 U7348 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7032) );
  XNOR2_X1 U7349 ( .A(n7032), .B(keyinput_223), .ZN(n6717) );
  OAI21_X1 U7350 ( .B1(n6719), .B2(n6718), .A(n6717), .ZN(n6722) );
  XNOR2_X1 U7351 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_224), .ZN(n6721) );
  XNOR2_X1 U7352 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_225), .ZN(n6720) );
  NAND3_X1 U7353 ( .A1(n6722), .A2(n6721), .A3(n6720), .ZN(n6725) );
  INV_X1 U7354 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7029) );
  XNOR2_X1 U7355 ( .A(n7029), .B(keyinput_226), .ZN(n6724) );
  XNOR2_X1 U7356 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_227), .ZN(n6723) );
  AOI21_X1 U7357 ( .B1(n6725), .B2(n6724), .A(n6723), .ZN(n6733) );
  XNOR2_X1 U7358 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_229), .ZN(n6732) );
  XNOR2_X1 U7359 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_230), .ZN(n6731) );
  XOR2_X1 U7360 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_228), .Z(n6729) );
  XOR2_X1 U7361 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_233), .Z(n6728) );
  XNOR2_X1 U7362 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_231), .ZN(n6727) );
  XNOR2_X1 U7363 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_232), .ZN(n6726)
         );
  NAND4_X1 U7364 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6730)
         );
  NOR4_X1 U7365 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6739)
         );
  INV_X1 U7366 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6978) );
  INV_X1 U7367 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6976) );
  AOI22_X1 U7368 ( .A1(n6978), .A2(keyinput_238), .B1(keyinput_234), .B2(n6976), .ZN(n6734) );
  OAI221_X1 U7369 ( .B1(n6978), .B2(keyinput_238), .C1(n6976), .C2(
        keyinput_234), .A(n6734), .ZN(n6738) );
  INV_X1 U7370 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6977) );
  AOI22_X1 U7371 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput_235), .B1(n6977), .B2(keyinput_236), .ZN(n6735) );
  OAI221_X1 U7372 ( .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput_235), .C1(
        n6977), .C2(keyinput_236), .A(n6735), .ZN(n6737) );
  XNOR2_X1 U7373 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_237), .ZN(n6736)
         );
  NOR4_X1 U7374 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6742)
         );
  INV_X1 U7375 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6979) );
  XNOR2_X1 U7376 ( .A(n6979), .B(keyinput_239), .ZN(n6741) );
  XNOR2_X1 U7377 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_240), .ZN(n6740)
         );
  OAI21_X1 U7378 ( .B1(n6742), .B2(n6741), .A(n6740), .ZN(n6748) );
  INV_X1 U7379 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6983) );
  INV_X1 U7380 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6981) );
  OAI22_X1 U7381 ( .A1(n6983), .A2(keyinput_243), .B1(n6981), .B2(keyinput_241), .ZN(n6743) );
  AOI221_X1 U7382 ( .B1(n6983), .B2(keyinput_243), .C1(keyinput_241), .C2(
        n6981), .A(n6743), .ZN(n6747) );
  XOR2_X1 U7383 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_245), .Z(n6746)
         );
  INV_X1 U7384 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6982) );
  OAI22_X1 U7385 ( .A1(n6982), .A2(keyinput_242), .B1(
        DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_244), .ZN(n6744) );
  AOI221_X1 U7386 ( .B1(n6982), .B2(keyinput_242), .C1(keyinput_244), .C2(
        DATAWIDTH_REG_12__SCAN_IN), .A(n6744), .ZN(n6745) );
  NAND4_X1 U7387 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6752)
         );
  XNOR2_X1 U7388 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_247), .ZN(n6751)
         );
  XNOR2_X1 U7389 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_246), .ZN(n6750)
         );
  XNOR2_X1 U7390 ( .A(DATAWIDTH_REG_16__SCAN_IN), .B(keyinput_248), .ZN(n6749)
         );
  AND4_X1 U7391 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6759)
         );
  XOR2_X1 U7392 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_249), .Z(n6758)
         );
  INV_X1 U7393 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6987) );
  XNOR2_X1 U7394 ( .A(n6987), .B(keyinput_251), .ZN(n6756) );
  XNOR2_X1 U7395 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_253), .ZN(n6755)
         );
  XNOR2_X1 U7396 ( .A(DATAWIDTH_REG_18__SCAN_IN), .B(keyinput_250), .ZN(n6754)
         );
  XNOR2_X1 U7397 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_252), .ZN(n6753)
         );
  NOR4_X1 U7398 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6757)
         );
  OAI21_X1 U7399 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n6944) );
  XOR2_X1 U7400 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .Z(n6943)
         );
  XOR2_X1 U7401 ( .A(DATAI_29_), .B(keyinput_2), .Z(n6762) );
  XNOR2_X1 U7402 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n6761) );
  XNOR2_X1 U7403 ( .A(DATAI_31_), .B(keyinput_0), .ZN(n6760) );
  NOR3_X1 U7404 ( .A1(n6762), .A2(n6761), .A3(n6760), .ZN(n6766) );
  XNOR2_X1 U7405 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n6765) );
  XOR2_X1 U7406 ( .A(DATAI_27_), .B(keyinput_4), .Z(n6764) );
  XNOR2_X1 U7407 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n6763) );
  OAI211_X1 U7408 ( .C1(n6766), .C2(n6765), .A(n6764), .B(n6763), .ZN(n6769)
         );
  XNOR2_X1 U7409 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n6768) );
  XNOR2_X1 U7410 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n6767) );
  AOI21_X1 U7411 ( .B1(n6769), .B2(n6768), .A(n6767), .ZN(n6772) );
  XOR2_X1 U7412 ( .A(DATAI_23_), .B(keyinput_8), .Z(n6771) );
  XNOR2_X1 U7413 ( .A(keyinput_9), .B(DATAI_22_), .ZN(n6770) );
  NOR3_X1 U7414 ( .A1(n6772), .A2(n6771), .A3(n6770), .ZN(n6781) );
  XNOR2_X1 U7415 ( .A(keyinput_10), .B(DATAI_21_), .ZN(n6780) );
  XOR2_X1 U7416 ( .A(keyinput_13), .B(DATAI_18_), .Z(n6778) );
  XOR2_X1 U7417 ( .A(keyinput_15), .B(DATAI_16_), .Z(n6777) );
  XNOR2_X1 U7418 ( .A(keyinput_12), .B(DATAI_19_), .ZN(n6776) );
  XNOR2_X1 U7419 ( .A(keyinput_11), .B(DATAI_20_), .ZN(n6774) );
  XNOR2_X1 U7420 ( .A(keyinput_14), .B(DATAI_17_), .ZN(n6773) );
  NAND2_X1 U7421 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  NOR4_X1 U7422 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6779)
         );
  OAI21_X1 U7423 ( .B1(n6781), .B2(n6780), .A(n6779), .ZN(n6784) );
  XNOR2_X1 U7424 ( .A(keyinput_16), .B(DATAI_15_), .ZN(n6783) );
  XOR2_X1 U7425 ( .A(DATAI_14_), .B(keyinput_17), .Z(n6782) );
  AOI21_X1 U7426 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(n6787) );
  XOR2_X1 U7427 ( .A(DATAI_13_), .B(keyinput_18), .Z(n6786) );
  XNOR2_X1 U7428 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n6785) );
  OAI21_X1 U7429 ( .B1(n6787), .B2(n6786), .A(n6785), .ZN(n6791) );
  XOR2_X1 U7430 ( .A(DATAI_11_), .B(keyinput_20), .Z(n6790) );
  XOR2_X1 U7431 ( .A(DATAI_10_), .B(keyinput_21), .Z(n6789) );
  XOR2_X1 U7432 ( .A(DATAI_9_), .B(keyinput_22), .Z(n6788) );
  AOI211_X1 U7433 ( .C1(n6791), .C2(n6790), .A(n6789), .B(n6788), .ZN(n6794)
         );
  XOR2_X1 U7434 ( .A(DATAI_8_), .B(keyinput_23), .Z(n6793) );
  XOR2_X1 U7435 ( .A(DATAI_7_), .B(keyinput_24), .Z(n6792) );
  NOR3_X1 U7436 ( .A1(n6794), .A2(n6793), .A3(n6792), .ZN(n6797) );
  XOR2_X1 U7437 ( .A(keyinput_25), .B(DATAI_6_), .Z(n6796) );
  XNOR2_X1 U7438 ( .A(keyinput_26), .B(DATAI_5_), .ZN(n6795) );
  NOR3_X1 U7439 ( .A1(n6797), .A2(n6796), .A3(n6795), .ZN(n6800) );
  XOR2_X1 U7440 ( .A(keyinput_27), .B(DATAI_4_), .Z(n6799) );
  XNOR2_X1 U7441 ( .A(keyinput_28), .B(DATAI_3_), .ZN(n6798) );
  OAI21_X1 U7442 ( .B1(n6800), .B2(n6799), .A(n6798), .ZN(n6804) );
  XOR2_X1 U7443 ( .A(keyinput_29), .B(DATAI_2_), .Z(n6803) );
  XOR2_X1 U7444 ( .A(keyinput_30), .B(DATAI_1_), .Z(n6802) );
  XOR2_X1 U7445 ( .A(keyinput_31), .B(DATAI_0_), .Z(n6801) );
  AOI211_X1 U7446 ( .C1(n6804), .C2(n6803), .A(n6802), .B(n6801), .ZN(n6808)
         );
  XOR2_X1 U7447 ( .A(keyinput_33), .B(NA_N), .Z(n6807) );
  XOR2_X1 U7448 ( .A(keyinput_34), .B(BS16_N), .Z(n6806) );
  XNOR2_X1 U7449 ( .A(keyinput_32), .B(MEMORYFETCH_REG_SCAN_IN), .ZN(n6805) );
  NOR4_X1 U7450 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6812)
         );
  XNOR2_X1 U7451 ( .A(n7513), .B(keyinput_35), .ZN(n6811) );
  XOR2_X1 U7452 ( .A(keyinput_36), .B(HOLD), .Z(n6810) );
  XNOR2_X1 U7453 ( .A(keyinput_37), .B(READREQUEST_REG_SCAN_IN), .ZN(n6809) );
  OAI211_X1 U7454 ( .C1(n6812), .C2(n6811), .A(n6810), .B(n6809), .ZN(n6815)
         );
  XNOR2_X1 U7455 ( .A(keyinput_38), .B(ADS_N_REG_SCAN_IN), .ZN(n6814) );
  XNOR2_X1 U7456 ( .A(keyinput_39), .B(CODEFETCH_REG_SCAN_IN), .ZN(n6813) );
  NAND3_X1 U7457 ( .A1(n6815), .A2(n6814), .A3(n6813), .ZN(n6818) );
  XNOR2_X1 U7458 ( .A(keyinput_40), .B(M_IO_N_REG_SCAN_IN), .ZN(n6817) );
  INV_X1 U7459 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7154) );
  XNOR2_X1 U7460 ( .A(n7154), .B(keyinput_41), .ZN(n6816) );
  AOI21_X1 U7461 ( .B1(n6818), .B2(n6817), .A(n6816), .ZN(n6824) );
  XNOR2_X1 U7462 ( .A(keyinput_42), .B(REQUESTPENDING_REG_SCAN_IN), .ZN(n6823)
         );
  XOR2_X1 U7463 ( .A(keyinput_45), .B(FLUSH_REG_SCAN_IN), .Z(n6821) );
  XNOR2_X1 U7464 ( .A(n7502), .B(keyinput_43), .ZN(n6820) );
  XNOR2_X1 U7465 ( .A(keyinput_44), .B(MORE_REG_SCAN_IN), .ZN(n6819) );
  NOR3_X1 U7466 ( .A1(n6821), .A2(n6820), .A3(n6819), .ZN(n6822) );
  OAI21_X1 U7467 ( .B1(n6824), .B2(n6823), .A(n6822), .ZN(n6828) );
  INV_X1 U7468 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7156) );
  XNOR2_X1 U7469 ( .A(n7156), .B(keyinput_46), .ZN(n6827) );
  XOR2_X1 U7470 ( .A(keyinput_47), .B(BYTEENABLE_REG_0__SCAN_IN), .Z(n6826) );
  XNOR2_X1 U7471 ( .A(keyinput_48), .B(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6825)
         );
  NAND4_X1 U7472 ( .A1(n6828), .A2(n6827), .A3(n6826), .A4(n6825), .ZN(n6833)
         );
  INV_X1 U7473 ( .A(keyinput_51), .ZN(n6829) );
  XNOR2_X1 U7474 ( .A(n6829), .B(REIP_REG_31__SCAN_IN), .ZN(n6832) );
  XNOR2_X1 U7475 ( .A(keyinput_50), .B(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6831)
         );
  XNOR2_X1 U7476 ( .A(keyinput_49), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6830)
         );
  NAND4_X1 U7477 ( .A1(n6833), .A2(n6832), .A3(n6831), .A4(n6830), .ZN(n6839)
         );
  OAI22_X1 U7478 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_53), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput_56), .ZN(n6834) );
  AOI221_X1 U7479 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_53), .C1(
        keyinput_56), .C2(REIP_REG_26__SCAN_IN), .A(n6834), .ZN(n6838) );
  XNOR2_X1 U7480 ( .A(n7070), .B(keyinput_52), .ZN(n6837) );
  INV_X1 U7481 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7064) );
  OAI22_X1 U7482 ( .A1(n7064), .A2(keyinput_54), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_55), .ZN(n6835) );
  AOI221_X1 U7483 ( .B1(n7064), .B2(keyinput_54), .C1(keyinput_55), .C2(
        REIP_REG_27__SCAN_IN), .A(n6835), .ZN(n6836) );
  NAND4_X1 U7484 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6843)
         );
  XOR2_X1 U7485 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .Z(n6842) );
  XNOR2_X1 U7486 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_59), .ZN(n6841) );
  XNOR2_X1 U7487 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .ZN(n6840) );
  AOI211_X1 U7488 ( .C1(n6843), .C2(n6842), .A(n6841), .B(n6840), .ZN(n6847)
         );
  XNOR2_X1 U7489 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n6846) );
  XNOR2_X1 U7490 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n6845) );
  XNOR2_X1 U7491 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .ZN(n6844) );
  OR4_X1 U7492 ( .A1(n6847), .A2(n6846), .A3(n6845), .A4(n6844), .ZN(n6850) );
  XNOR2_X1 U7493 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .ZN(n6849) );
  XNOR2_X1 U7494 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .ZN(n6848) );
  AOI21_X1 U7495 ( .B1(n6850), .B2(n6849), .A(n6848), .ZN(n6857) );
  INV_X1 U7496 ( .A(keyinput_67), .ZN(n6854) );
  INV_X1 U7497 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7072) );
  XOR2_X1 U7498 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .Z(n6853) );
  INV_X1 U7499 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7368) );
  OAI22_X1 U7500 ( .A1(n7368), .A2(keyinput_65), .B1(keyinput_67), .B2(
        BE_N_REG_3__SCAN_IN), .ZN(n6851) );
  AOI21_X1 U7501 ( .B1(n7368), .B2(keyinput_65), .A(n6851), .ZN(n6852) );
  OAI211_X1 U7502 ( .C1(n6854), .C2(n7072), .A(n6853), .B(n6852), .ZN(n6856)
         );
  XOR2_X1 U7503 ( .A(keyinput_68), .B(BE_N_REG_2__SCAN_IN), .Z(n6855) );
  OAI21_X1 U7504 ( .B1(n6857), .B2(n6856), .A(n6855), .ZN(n6861) );
  XOR2_X1 U7505 ( .A(keyinput_71), .B(ADDRESS_REG_29__SCAN_IN), .Z(n6860) );
  XOR2_X1 U7506 ( .A(keyinput_69), .B(BE_N_REG_1__SCAN_IN), .Z(n6859) );
  XNOR2_X1 U7507 ( .A(keyinput_70), .B(BE_N_REG_0__SCAN_IN), .ZN(n6858) );
  NAND4_X1 U7508 ( .A1(n6861), .A2(n6860), .A3(n6859), .A4(n6858), .ZN(n6871)
         );
  INV_X1 U7509 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7059) );
  XNOR2_X1 U7510 ( .A(n7059), .B(keyinput_75), .ZN(n6865) );
  XNOR2_X1 U7511 ( .A(keyinput_73), .B(ADDRESS_REG_27__SCAN_IN), .ZN(n6864) );
  XNOR2_X1 U7512 ( .A(n7066), .B(keyinput_72), .ZN(n6863) );
  XNOR2_X1 U7513 ( .A(keyinput_74), .B(ADDRESS_REG_26__SCAN_IN), .ZN(n6862) );
  NOR4_X1 U7514 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6870)
         );
  XOR2_X1 U7515 ( .A(keyinput_76), .B(ADDRESS_REG_24__SCAN_IN), .Z(n6868) );
  INV_X1 U7516 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7055) );
  XNOR2_X1 U7517 ( .A(n7055), .B(keyinput_77), .ZN(n6867) );
  INV_X1 U7518 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7052) );
  XNOR2_X1 U7519 ( .A(n7052), .B(keyinput_78), .ZN(n6866) );
  NAND3_X1 U7520 ( .A1(n6868), .A2(n6867), .A3(n6866), .ZN(n6869) );
  AOI21_X1 U7521 ( .B1(n6871), .B2(n6870), .A(n6869), .ZN(n6877) );
  INV_X1 U7522 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7051) );
  XNOR2_X1 U7523 ( .A(n7051), .B(keyinput_79), .ZN(n6876) );
  XNOR2_X1 U7524 ( .A(keyinput_80), .B(ADDRESS_REG_20__SCAN_IN), .ZN(n6874) );
  XNOR2_X1 U7525 ( .A(keyinput_81), .B(ADDRESS_REG_19__SCAN_IN), .ZN(n6873) );
  XNOR2_X1 U7526 ( .A(keyinput_82), .B(ADDRESS_REG_18__SCAN_IN), .ZN(n6872) );
  NOR3_X1 U7527 ( .A1(n6874), .A2(n6873), .A3(n6872), .ZN(n6875) );
  OAI21_X1 U7528 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n6880) );
  INV_X1 U7529 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7045) );
  XNOR2_X1 U7530 ( .A(n7045), .B(keyinput_84), .ZN(n6879) );
  XNOR2_X1 U7531 ( .A(keyinput_83), .B(ADDRESS_REG_17__SCAN_IN), .ZN(n6878) );
  NAND3_X1 U7532 ( .A1(n6880), .A2(n6879), .A3(n6878), .ZN(n6883) );
  XOR2_X1 U7533 ( .A(keyinput_85), .B(ADDRESS_REG_15__SCAN_IN), .Z(n6882) );
  INV_X1 U7534 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7043) );
  XNOR2_X1 U7535 ( .A(n7043), .B(keyinput_86), .ZN(n6881) );
  NAND3_X1 U7536 ( .A1(n6883), .A2(n6882), .A3(n6881), .ZN(n6886) );
  XNOR2_X1 U7537 ( .A(n7042), .B(keyinput_87), .ZN(n6885) );
  XNOR2_X1 U7538 ( .A(keyinput_88), .B(ADDRESS_REG_12__SCAN_IN), .ZN(n6884) );
  AOI21_X1 U7539 ( .B1(n6886), .B2(n6885), .A(n6884), .ZN(n6892) );
  AOI22_X1 U7540 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput_93), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(keyinput_91), .ZN(n6887) );
  OAI221_X1 U7541 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput_93), .C1(
        ADDRESS_REG_9__SCAN_IN), .C2(keyinput_91), .A(n6887), .ZN(n6891) );
  AOI22_X1 U7542 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput_89), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(keyinput_92), .ZN(n6888) );
  OAI221_X1 U7543 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput_89), .C1(
        ADDRESS_REG_8__SCAN_IN), .C2(keyinput_92), .A(n6888), .ZN(n6890) );
  XNOR2_X1 U7544 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_90), .ZN(n6889) );
  OR4_X1 U7545 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6895) );
  XNOR2_X1 U7546 ( .A(n7033), .B(keyinput_94), .ZN(n6894) );
  XNOR2_X1 U7547 ( .A(keyinput_95), .B(ADDRESS_REG_5__SCAN_IN), .ZN(n6893) );
  AOI21_X1 U7548 ( .B1(n6895), .B2(n6894), .A(n6893), .ZN(n6898) );
  INV_X1 U7549 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7031) );
  XNOR2_X1 U7550 ( .A(n7031), .B(keyinput_96), .ZN(n6897) );
  INV_X1 U7551 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7030) );
  XNOR2_X1 U7552 ( .A(n7030), .B(keyinput_97), .ZN(n6896) );
  NOR3_X1 U7553 ( .A1(n6898), .A2(n6897), .A3(n6896), .ZN(n6901) );
  XNOR2_X1 U7554 ( .A(n7029), .B(keyinput_98), .ZN(n6900) );
  XNOR2_X1 U7555 ( .A(keyinput_99), .B(ADDRESS_REG_1__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U7556 ( .B1(n6901), .B2(n6900), .A(n6899), .ZN(n6909) );
  XOR2_X1 U7557 ( .A(keyinput_100), .B(ADDRESS_REG_0__SCAN_IN), .Z(n6908) );
  XOR2_X1 U7558 ( .A(keyinput_105), .B(DATAWIDTH_REG_1__SCAN_IN), .Z(n6907) );
  XNOR2_X1 U7559 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_103), .ZN(n6905) );
  XNOR2_X1 U7560 ( .A(keyinput_104), .B(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6904)
         );
  XNOR2_X1 U7561 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .ZN(n6903) );
  XNOR2_X1 U7562 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .ZN(n6902) );
  NOR4_X1 U7563 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6906)
         );
  NAND4_X1 U7564 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n6916)
         );
  XOR2_X1 U7565 ( .A(keyinput_109), .B(DATAWIDTH_REG_5__SCAN_IN), .Z(n6912) );
  XOR2_X1 U7566 ( .A(keyinput_110), .B(DATAWIDTH_REG_6__SCAN_IN), .Z(n6911) );
  XNOR2_X1 U7567 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_107), .ZN(n6910)
         );
  NOR3_X1 U7568 ( .A1(n6912), .A2(n6911), .A3(n6910), .ZN(n6915) );
  XNOR2_X1 U7569 ( .A(keyinput_106), .B(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6914)
         );
  XNOR2_X1 U7570 ( .A(keyinput_108), .B(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6913)
         );
  NAND4_X1 U7571 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), .ZN(n6919)
         );
  XNOR2_X1 U7572 ( .A(keyinput_111), .B(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6918)
         );
  XNOR2_X1 U7573 ( .A(keyinput_112), .B(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6917)
         );
  AOI21_X1 U7574 ( .B1(n6919), .B2(n6918), .A(n6917), .ZN(n6925) );
  AOI22_X1 U7575 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput_117), .B1(
        n6983), .B2(keyinput_115), .ZN(n6920) );
  OAI221_X1 U7576 ( .B1(DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_117), .C1(
        n6983), .C2(keyinput_115), .A(n6920), .ZN(n6924) );
  AOI22_X1 U7577 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput_114), .B1(
        n6981), .B2(keyinput_113), .ZN(n6921) );
  OAI221_X1 U7578 ( .B1(DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_114), .C1(
        n6981), .C2(keyinput_113), .A(n6921), .ZN(n6923) );
  XNOR2_X1 U7579 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_116), .ZN(n6922)
         );
  NOR4_X1 U7580 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6930)
         );
  INV_X1 U7581 ( .A(keyinput_118), .ZN(n6926) );
  XNOR2_X1 U7582 ( .A(n6926), .B(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6929) );
  XNOR2_X1 U7583 ( .A(keyinput_120), .B(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6928)
         );
  XNOR2_X1 U7584 ( .A(keyinput_119), .B(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6927)
         );
  NOR4_X1 U7585 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n6937)
         );
  XNOR2_X1 U7586 ( .A(keyinput_121), .B(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6936)
         );
  INV_X1 U7587 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6986) );
  XNOR2_X1 U7588 ( .A(n6986), .B(keyinput_122), .ZN(n6934) );
  XNOR2_X1 U7589 ( .A(keyinput_124), .B(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6933)
         );
  INV_X1 U7590 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6988) );
  XNOR2_X1 U7591 ( .A(n6988), .B(keyinput_125), .ZN(n6932) );
  XNOR2_X1 U7592 ( .A(keyinput_123), .B(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6931)
         );
  NOR4_X1 U7593 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n6935)
         );
  OAI21_X1 U7594 ( .B1(n6937), .B2(n6936), .A(n6935), .ZN(n6940) );
  INV_X1 U7595 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6989) );
  XNOR2_X1 U7596 ( .A(n6989), .B(keyinput_126), .ZN(n6939) );
  XOR2_X1 U7597 ( .A(keyinput_127), .B(DATAWIDTH_REG_23__SCAN_IN), .Z(n6938)
         );
  NAND3_X1 U7598 ( .A1(n6940), .A2(n6939), .A3(n6938), .ZN(n6942) );
  XNOR2_X1 U7599 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_254), .ZN(n6941)
         );
  NAND4_X1 U7600 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6958)
         );
  AOI221_X1 U7601 ( .B1(n7197), .B2(n6948), .C1(n6946), .C2(n6948), .A(n6945), 
        .ZN(n6956) );
  NAND2_X1 U7602 ( .A1(n6947), .A2(n7239), .ZN(n6954) );
  NOR3_X1 U7603 ( .A1(n6949), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n6948), 
        .ZN(n6950) );
  AOI211_X1 U7604 ( .C1(n6952), .C2(n7238), .A(n6951), .B(n6950), .ZN(n6953)
         );
  OAI211_X1 U7605 ( .C1(n6956), .C2(n6955), .A(n6954), .B(n6953), .ZN(n6957)
         );
  XNOR2_X1 U7606 ( .A(n6958), .B(n6957), .ZN(U3006) );
  NAND2_X1 U7607 ( .A1(n4892), .A2(n6959), .ZN(n6966) );
  NOR2_X1 U7608 ( .A1(n6961), .A2(n6960), .ZN(n6969) );
  AOI22_X1 U7609 ( .A1(n6964), .A2(n6963), .B1(n6969), .B2(n6962), .ZN(n6965)
         );
  NAND2_X1 U7610 ( .A1(n6966), .A2(n6965), .ZN(n7457) );
  INV_X1 U7611 ( .A(n7457), .ZN(n6972) );
  AOI22_X1 U7612 ( .A1(n7494), .A2(n6969), .B1(n6968), .B2(n6967), .ZN(n6970)
         );
  OAI21_X1 U7613 ( .B1(n6972), .B2(n6971), .A(n6970), .ZN(n6973) );
  MUX2_X1 U7614 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n6973), .S(n7441), 
        .Z(U3460) );
  INV_X1 U7615 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6975) );
  INV_X1 U7616 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6974) );
  NOR2_X1 U7617 ( .A1(n6974), .A2(STATE_REG_2__SCAN_IN), .ZN(n7512) );
  NOR2_X1 U7618 ( .A1(n6974), .A2(STATE_REG_0__SCAN_IN), .ZN(n7068) );
  INV_X1 U7619 ( .A(n7068), .ZN(n7522) );
  OAI21_X2 U7620 ( .B1(n7512), .B2(n7158), .A(n7522), .ZN(n7505) );
  NOR2_X1 U7621 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n7153) );
  INV_X1 U7622 ( .A(n7505), .ZN(n7503) );
  OAI21_X1 U7623 ( .B1(BS16_N), .B2(n7153), .A(n7503), .ZN(n7501) );
  INV_X1 U7624 ( .A(n7501), .ZN(n7504) );
  AOI21_X1 U7625 ( .B1(n6975), .B2(n7505), .A(n7504), .ZN(U3451) );
  NOR2_X1 U7626 ( .A1(n7503), .A2(n6976), .ZN(U3180) );
  AND2_X1 U7627 ( .A1(n7505), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  NOR2_X1 U7628 ( .A1(n7503), .A2(n6977), .ZN(U3178) );
  AND2_X1 U7629 ( .A1(n7505), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  NOR2_X1 U7630 ( .A1(n7503), .A2(n6978), .ZN(U3176) );
  NOR2_X1 U7631 ( .A1(n7503), .A2(n6979), .ZN(U3175) );
  INV_X1 U7632 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U7633 ( .A1(n7503), .A2(n6980), .ZN(U3174) );
  NOR2_X1 U7634 ( .A1(n7503), .A2(n6981), .ZN(U3173) );
  NOR2_X1 U7635 ( .A1(n7503), .A2(n6982), .ZN(U3172) );
  NOR2_X1 U7636 ( .A1(n7503), .A2(n6983), .ZN(U3171) );
  AND2_X1 U7637 ( .A1(n7505), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7638 ( .A1(n7505), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  INV_X1 U7639 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6984) );
  NOR2_X1 U7640 ( .A1(n7503), .A2(n6984), .ZN(U3168) );
  INV_X1 U7641 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6985) );
  NOR2_X1 U7642 ( .A1(n7503), .A2(n6985), .ZN(U3167) );
  AND2_X1 U7643 ( .A1(n7505), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U7644 ( .A1(n7505), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  NOR2_X1 U7645 ( .A1(n7503), .A2(n6986), .ZN(U3164) );
  NOR2_X1 U7646 ( .A1(n7503), .A2(n6987), .ZN(U3163) );
  AND2_X1 U7647 ( .A1(n7505), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  NOR2_X1 U7648 ( .A1(n7503), .A2(n6988), .ZN(U3161) );
  NOR2_X1 U7649 ( .A1(n7503), .A2(n6989), .ZN(U3160) );
  AND2_X1 U7650 ( .A1(n7505), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7651 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7505), .ZN(U3158) );
  AND2_X1 U7652 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7505), .ZN(U3157) );
  AND2_X1 U7653 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7505), .ZN(U3156) );
  AND2_X1 U7654 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7505), .ZN(U3155) );
  AND2_X1 U7655 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7505), .ZN(U3154) );
  AND2_X1 U7656 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7505), .ZN(U3153) );
  AND2_X1 U7657 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7505), .ZN(U3152) );
  AND2_X1 U7658 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7505), .ZN(U3151) );
  NOR2_X1 U7659 ( .A1(n6991), .A2(n6990), .ZN(U3019) );
  AND2_X1 U7660 ( .A1(n6992), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7661 ( .A(n7522), .ZN(n7525) );
  INV_X1 U7662 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6993) );
  OAI21_X1 U7663 ( .B1(n7525), .B2(n6993), .A(n7505), .ZN(U2789) );
  AOI22_X1 U7664 ( .A1(n7167), .A2(LWORD_REG_0__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6994) );
  OAI21_X1 U7665 ( .B1(n6995), .B2(n7024), .A(n6994), .ZN(U2923) );
  AOI22_X1 U7666 ( .A1(n7167), .A2(LWORD_REG_1__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6996) );
  OAI21_X1 U7667 ( .B1(n6997), .B2(n7024), .A(n6996), .ZN(U2922) );
  AOI22_X1 U7668 ( .A1(n7167), .A2(LWORD_REG_2__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6998) );
  OAI21_X1 U7669 ( .B1(n6999), .B2(n7024), .A(n6998), .ZN(U2921) );
  AOI22_X1 U7670 ( .A1(n7167), .A2(LWORD_REG_3__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7000) );
  OAI21_X1 U7671 ( .B1(n7001), .B2(n7024), .A(n7000), .ZN(U2920) );
  AOI22_X1 U7672 ( .A1(n7167), .A2(LWORD_REG_4__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7002) );
  OAI21_X1 U7673 ( .B1(n7003), .B2(n7024), .A(n7002), .ZN(U2919) );
  AOI22_X1 U7674 ( .A1(n7167), .A2(LWORD_REG_5__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7004) );
  OAI21_X1 U7675 ( .B1(n4697), .B2(n7024), .A(n7004), .ZN(U2918) );
  AOI22_X1 U7676 ( .A1(n7167), .A2(LWORD_REG_6__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7005) );
  OAI21_X1 U7677 ( .B1(n4699), .B2(n7024), .A(n7005), .ZN(U2917) );
  AOI22_X1 U7678 ( .A1(n7167), .A2(LWORD_REG_7__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7006) );
  OAI21_X1 U7679 ( .B1(n7007), .B2(n7024), .A(n7006), .ZN(U2916) );
  AOI22_X1 U7680 ( .A1(n7167), .A2(LWORD_REG_8__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7008) );
  OAI21_X1 U7681 ( .B1(n7009), .B2(n7024), .A(n7008), .ZN(U2915) );
  AOI22_X1 U7682 ( .A1(n7167), .A2(LWORD_REG_9__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7010) );
  OAI21_X1 U7683 ( .B1(n7011), .B2(n7024), .A(n7010), .ZN(U2914) );
  AOI22_X1 U7684 ( .A1(n7167), .A2(LWORD_REG_10__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7012) );
  OAI21_X1 U7685 ( .B1(n7013), .B2(n7024), .A(n7012), .ZN(U2913) );
  AOI22_X1 U7686 ( .A1(n7167), .A2(LWORD_REG_11__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7014) );
  OAI21_X1 U7687 ( .B1(n7015), .B2(n7024), .A(n7014), .ZN(U2912) );
  AOI22_X1 U7688 ( .A1(n7167), .A2(LWORD_REG_12__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7016) );
  OAI21_X1 U7689 ( .B1(n7017), .B2(n7024), .A(n7016), .ZN(U2911) );
  AOI22_X1 U7690 ( .A1(n7167), .A2(LWORD_REG_13__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7018) );
  OAI21_X1 U7691 ( .B1(n7019), .B2(n7024), .A(n7018), .ZN(U2910) );
  AOI22_X1 U7692 ( .A1(n7167), .A2(LWORD_REG_14__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7020) );
  OAI21_X1 U7693 ( .B1(n7021), .B2(n7024), .A(n7020), .ZN(U2909) );
  AOI22_X1 U7694 ( .A1(n7167), .A2(LWORD_REG_15__SCAN_IN), .B1(n7022), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U7695 ( .B1(n7025), .B2(n7024), .A(n7023), .ZN(U2908) );
  INV_X1 U7696 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7198) );
  INV_X1 U7697 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7026) );
  INV_X1 U7698 ( .A(n7522), .ZN(n7157) );
  INV_X1 U7699 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7086) );
  OAI222_X1 U7700 ( .A1(n7056), .A2(n7198), .B1(n7026), .B2(n7157), .C1(n7086), 
        .C2(n7071), .ZN(U3184) );
  INV_X1 U7701 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7027) );
  OAI222_X1 U7702 ( .A1(n7056), .A2(n7028), .B1(n7027), .B2(n7068), .C1(n7198), 
        .C2(n7071), .ZN(U3185) );
  OAI222_X1 U7703 ( .A1(n7056), .A2(n7272), .B1(n7029), .B2(n7157), .C1(n7028), 
        .C2(n7071), .ZN(U3186) );
  OAI222_X1 U7704 ( .A1(n7056), .A2(n7129), .B1(n7030), .B2(n7068), .C1(n7272), 
        .C2(n7071), .ZN(U3187) );
  OAI222_X1 U7705 ( .A1(n7056), .A2(n5271), .B1(n7031), .B2(n7157), .C1(n7129), 
        .C2(n7071), .ZN(U3188) );
  INV_X1 U7706 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7300) );
  OAI222_X1 U7707 ( .A1(n7056), .A2(n7300), .B1(n7032), .B2(n7068), .C1(n5271), 
        .C2(n7071), .ZN(U3189) );
  OAI222_X1 U7708 ( .A1(n7056), .A2(n5620), .B1(n7033), .B2(n7157), .C1(n7300), 
        .C2(n7071), .ZN(U3190) );
  OAI222_X1 U7709 ( .A1(n7056), .A2(n7035), .B1(n7034), .B2(n7157), .C1(n5620), 
        .C2(n7071), .ZN(U3191) );
  INV_X1 U7710 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7214) );
  OAI222_X1 U7711 ( .A1(n7056), .A2(n7214), .B1(n7036), .B2(n7157), .C1(n7035), 
        .C2(n7071), .ZN(U3192) );
  INV_X1 U7712 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7037) );
  OAI222_X1 U7713 ( .A1(n7056), .A2(n7306), .B1(n7037), .B2(n7157), .C1(n7214), 
        .C2(n7071), .ZN(U3193) );
  INV_X1 U7714 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7038) );
  OAI222_X1 U7715 ( .A1(n7056), .A2(n7039), .B1(n7038), .B2(n7157), .C1(n7306), 
        .C2(n7071), .ZN(U3194) );
  OAI222_X1 U7716 ( .A1(n7056), .A2(n5855), .B1(n7040), .B2(n7157), .C1(n7039), 
        .C2(n7071), .ZN(U3195) );
  INV_X1 U7717 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7041) );
  OAI222_X1 U7718 ( .A1(n7056), .A2(n5915), .B1(n7041), .B2(n7157), .C1(n5855), 
        .C2(n7071), .ZN(U3196) );
  OAI222_X1 U7719 ( .A1(n7056), .A2(n7342), .B1(n7042), .B2(n7157), .C1(n5915), 
        .C2(n7071), .ZN(U3197) );
  OAI222_X1 U7720 ( .A1(n7071), .A2(n7342), .B1(n7043), .B2(n7157), .C1(n7344), 
        .C2(n7056), .ZN(U3198) );
  INV_X1 U7721 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7044) );
  OAI222_X1 U7722 ( .A1(n7056), .A2(n7368), .B1(n7044), .B2(n7157), .C1(n7344), 
        .C2(n7071), .ZN(U3199) );
  OAI222_X1 U7723 ( .A1(n7071), .A2(n7368), .B1(n7045), .B2(n7157), .C1(n7379), 
        .C2(n7056), .ZN(U3200) );
  OAI222_X1 U7724 ( .A1(n7056), .A2(n7382), .B1(n7046), .B2(n7157), .C1(n7379), 
        .C2(n7071), .ZN(U3201) );
  OAI222_X1 U7725 ( .A1(n7071), .A2(n7382), .B1(n7047), .B2(n7157), .C1(n7391), 
        .C2(n7056), .ZN(U3202) );
  INV_X1 U7726 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7050) );
  OAI222_X1 U7727 ( .A1(n7071), .A2(n7391), .B1(n7048), .B2(n7157), .C1(n7050), 
        .C2(n7056), .ZN(U3203) );
  INV_X1 U7728 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7049) );
  OAI222_X1 U7729 ( .A1(n7071), .A2(n7050), .B1(n7049), .B2(n7157), .C1(n7420), 
        .C2(n7056), .ZN(U3204) );
  OAI222_X1 U7730 ( .A1(n7056), .A2(n7053), .B1(n7051), .B2(n7157), .C1(n7420), 
        .C2(n7071), .ZN(U3205) );
  OAI222_X1 U7731 ( .A1(n7071), .A2(n7053), .B1(n7052), .B2(n7157), .C1(n7054), 
        .C2(n7056), .ZN(U3206) );
  INV_X1 U7732 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7058) );
  OAI222_X1 U7733 ( .A1(n7056), .A2(n7058), .B1(n7055), .B2(n7068), .C1(n7054), 
        .C2(n7071), .ZN(U3207) );
  INV_X1 U7734 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7057) );
  OAI222_X1 U7735 ( .A1(n7071), .A2(n7058), .B1(n7057), .B2(n7068), .C1(n7060), 
        .C2(n7056), .ZN(U3208) );
  OAI222_X1 U7736 ( .A1(n7071), .A2(n7060), .B1(n7059), .B2(n7068), .C1(n7062), 
        .C2(n7056), .ZN(U3209) );
  OAI222_X1 U7737 ( .A1(n7071), .A2(n7062), .B1(n7061), .B2(n7068), .C1(n7064), 
        .C2(n7056), .ZN(U3210) );
  OAI222_X1 U7738 ( .A1(n7071), .A2(n7064), .B1(n7063), .B2(n7068), .C1(n7065), 
        .C2(n7056), .ZN(U3211) );
  OAI222_X1 U7739 ( .A1(n7056), .A2(n7070), .B1(n7066), .B2(n7068), .C1(n7065), 
        .C2(n7071), .ZN(U3212) );
  INV_X1 U7740 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7069) );
  OAI222_X1 U7741 ( .A1(n7071), .A2(n7070), .B1(n7069), .B2(n7068), .C1(n7067), 
        .C2(n7056), .ZN(U3213) );
  INV_X1 U7742 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7073) );
  AOI22_X1 U7743 ( .A1(n7525), .A2(n7073), .B1(n7072), .B2(n7522), .ZN(U3445)
         );
  AOI221_X1 U7744 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7084) );
  NOR4_X1 U7745 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7077) );
  NOR4_X1 U7746 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n7076) );
  NOR4_X1 U7747 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7075) );
  NOR4_X1 U7748 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n7074) );
  NAND4_X1 U7749 ( .A1(n7077), .A2(n7076), .A3(n7075), .A4(n7074), .ZN(n7083)
         );
  NOR4_X1 U7750 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7081) );
  AOI211_X1 U7751 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_11__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n7080) );
  NOR4_X1 U7752 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n7079) );
  NOR4_X1 U7753 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7078) );
  NAND4_X1 U7754 ( .A1(n7081), .A2(n7080), .A3(n7079), .A4(n7078), .ZN(n7082)
         );
  NOR2_X1 U7755 ( .A1(n7083), .A2(n7082), .ZN(n7097) );
  MUX2_X1 U7756 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n7084), .S(n7097), .Z(
        U2795) );
  OAI22_X1 U7757 ( .A1(n7522), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n7157), .ZN(n7085) );
  INV_X1 U7758 ( .A(n7085), .ZN(U3446) );
  AOI21_X1 U7759 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7087) );
  OAI221_X1 U7760 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7087), .C1(n7086), .C2(
        REIP_REG_0__SCAN_IN), .A(n7097), .ZN(n7088) );
  OAI21_X1 U7761 ( .B1(n7097), .B2(n7089), .A(n7088), .ZN(U3468) );
  OAI22_X1 U7762 ( .A1(n7522), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n7157), .ZN(n7090) );
  INV_X1 U7763 ( .A(n7090), .ZN(U3447) );
  NOR3_X1 U7764 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7091) );
  OAI21_X1 U7765 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7091), .A(n7097), .ZN(n7092)
         );
  OAI21_X1 U7766 ( .B1(n7097), .B2(n7093), .A(n7092), .ZN(U2794) );
  INV_X1 U7767 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7096) );
  INV_X1 U7768 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U7769 ( .A1(n7157), .A2(n7096), .B1(n7094), .B2(n7522), .ZN(U3448)
         );
  OAI21_X1 U7770 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n7097), .ZN(n7095) );
  OAI21_X1 U7771 ( .B1(n7097), .B2(n7096), .A(n7095), .ZN(U3469) );
  INV_X1 U7772 ( .A(EBX_REG_7__SCAN_IN), .ZN(n7103) );
  INV_X1 U7773 ( .A(n7098), .ZN(n7302) );
  NAND2_X1 U7774 ( .A1(n5326), .A2(n7099), .ZN(n7100) );
  AND2_X1 U7775 ( .A1(n7101), .A2(n7100), .ZN(n7295) );
  AOI22_X1 U7776 ( .A1(n7302), .A2(n7115), .B1(n7114), .B2(n7295), .ZN(n7102)
         );
  OAI21_X1 U7777 ( .B1(n7118), .B2(n7103), .A(n7102), .ZN(U2852) );
  INV_X1 U7778 ( .A(EBX_REG_11__SCAN_IN), .ZN(n7310) );
  INV_X1 U7779 ( .A(n7308), .ZN(n7104) );
  OAI22_X1 U7780 ( .A1(n7142), .A2(n6357), .B1(n7105), .B2(n7104), .ZN(n7106)
         );
  INV_X1 U7781 ( .A(n7106), .ZN(n7107) );
  OAI21_X1 U7782 ( .B1(n7118), .B2(n7310), .A(n7107), .ZN(U2848) );
  INV_X1 U7783 ( .A(n7108), .ZN(n7532) );
  INV_X1 U7784 ( .A(n7109), .ZN(n7408) );
  AOI22_X1 U7785 ( .A1(n7532), .A2(n7115), .B1(n7114), .B2(n7408), .ZN(n7110)
         );
  OAI21_X1 U7786 ( .B1(n7118), .B2(n7111), .A(n7110), .ZN(U2838) );
  INV_X1 U7787 ( .A(EBX_REG_19__SCAN_IN), .ZN(n7113) );
  AOI22_X1 U7788 ( .A1(n7529), .A2(n7115), .B1(n7114), .B2(n7386), .ZN(n7112)
         );
  OAI21_X1 U7789 ( .B1(n7118), .B2(n7113), .A(n7112), .ZN(U2840) );
  AOI22_X1 U7790 ( .A1(n7116), .A2(n7115), .B1(n7114), .B2(n7237), .ZN(n7117)
         );
  OAI21_X1 U7791 ( .B1(n7118), .B2(n6303), .A(n7117), .ZN(U2844) );
  AOI22_X1 U7792 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7147), .B1(n7205), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U7793 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  XOR2_X1 U7794 ( .A(n7122), .B(n7121), .Z(n7201) );
  AOI22_X1 U7795 ( .A1(n7148), .A2(n7201), .B1(n7255), .B2(n3628), .ZN(n7123)
         );
  OAI211_X1 U7796 ( .C1(n7152), .C2(n7247), .A(n7124), .B(n7123), .ZN(U2984)
         );
  INV_X1 U7797 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7276) );
  CLKBUF_X1 U7798 ( .A(n7125), .Z(n7126) );
  XOR2_X1 U7799 ( .A(n7127), .B(n7126), .Z(n7190) );
  INV_X1 U7800 ( .A(n7284), .ZN(n7128) );
  AOI222_X1 U7801 ( .A1(n7190), .A2(n7148), .B1(n3628), .B2(n7279), .C1(n7128), 
        .C2(n7143), .ZN(n7131) );
  NOR2_X1 U7802 ( .A1(n7213), .A2(n7129), .ZN(n7185) );
  INV_X1 U7803 ( .A(n7185), .ZN(n7130) );
  OAI211_X1 U7804 ( .C1(n7132), .C2(n7276), .A(n7131), .B(n7130), .ZN(U2981)
         );
  AOI22_X1 U7805 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n7147), .B1(n7205), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n7135) );
  AOI22_X1 U7806 ( .A1(n7133), .A2(n7148), .B1(n3628), .B2(n7290), .ZN(n7134)
         );
  OAI211_X1 U7807 ( .C1(n7152), .C2(n7292), .A(n7135), .B(n7134), .ZN(U2980)
         );
  AOI22_X1 U7808 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n7147), .B1(n7205), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U7809 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n7139) );
  INV_X1 U7810 ( .A(n7139), .ZN(n7206) );
  AOI22_X1 U7811 ( .A1(n7206), .A2(n7148), .B1(n3628), .B2(n7302), .ZN(n7140)
         );
  OAI211_X1 U7812 ( .C1(n7152), .C2(n7305), .A(n7141), .B(n7140), .ZN(U2979)
         );
  AOI22_X1 U7813 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7147), .B1(n7205), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n7145) );
  INV_X1 U7814 ( .A(n7142), .ZN(n7313) );
  AOI22_X1 U7815 ( .A1(n7313), .A2(n3628), .B1(n7143), .B2(n7312), .ZN(n7144)
         );
  OAI211_X1 U7816 ( .C1(n7146), .C2(n7433), .A(n7145), .B(n7144), .ZN(U2975)
         );
  AOI22_X1 U7817 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7147), .B1(n7205), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n7151) );
  AOI22_X1 U7818 ( .A1(n7149), .A2(n7148), .B1(n3628), .B2(n7526), .ZN(n7150)
         );
  OAI211_X1 U7819 ( .C1(n7152), .C2(n7362), .A(n7151), .B(n7150), .ZN(U2969)
         );
  INV_X1 U7820 ( .A(n7153), .ZN(n7155) );
  OAI222_X1 U7821 ( .A1(n7525), .A2(n7155), .B1(n7525), .B2(n7154), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(n7522), .ZN(U2791) );
  AOI22_X1 U7822 ( .A1(n7157), .A2(READREQUEST_REG_SCAN_IN), .B1(n7156), .B2(
        n7522), .ZN(U3470) );
  AND2_X1 U7823 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7508) );
  INV_X1 U7824 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7515) );
  NOR2_X1 U7825 ( .A1(n7158), .A2(n7515), .ZN(n7518) );
  AOI21_X1 U7826 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7518), .ZN(n7160)
         );
  NAND2_X1 U7827 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7507) );
  OAI211_X1 U7828 ( .C1(n7508), .C2(n7160), .A(n7159), .B(n7507), .ZN(U3182)
         );
  NOR2_X1 U7829 ( .A1(READY_N), .A2(n7161), .ZN(n7162) );
  OAI21_X1 U7830 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7162), .A(n7491), .ZN(
        n7164) );
  OAI21_X1 U7831 ( .B1(n7495), .B2(n7164), .A(n7163), .ZN(U3150) );
  AOI211_X1 U7832 ( .C1(n7167), .C2(n7513), .A(n7166), .B(n7165), .ZN(n7174)
         );
  INV_X1 U7833 ( .A(n7168), .ZN(n7171) );
  OAI211_X1 U7834 ( .C1(n7169), .C2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .B(n7513), .ZN(n7170) );
  OAI21_X1 U7835 ( .B1(n7171), .B2(n7170), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n7173) );
  NOR2_X1 U7836 ( .A1(n7174), .A2(n7495), .ZN(n7172) );
  AOI22_X1 U7837 ( .A1(n7515), .A2(n7174), .B1(n7173), .B2(n7172), .ZN(U3472)
         );
  NAND3_X1 U7838 ( .A1(n3881), .A2(n7176), .A3(n7175), .ZN(n7178) );
  OAI211_X1 U7839 ( .C1(n7215), .C2(n7179), .A(n7178), .B(n7177), .ZN(n7180)
         );
  AOI21_X1 U7840 ( .B1(n7239), .B2(n7181), .A(n7180), .ZN(n7182) );
  OAI221_X1 U7841 ( .B1(n3881), .B2(n7184), .C1(n3881), .C2(n7183), .A(n7182), 
        .ZN(U3017) );
  AOI21_X1 U7842 ( .B1(n7273), .B2(n7238), .A(n7185), .ZN(n7186) );
  OAI21_X1 U7843 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7189) );
  AOI21_X1 U7844 ( .B1(n7190), .B2(n7239), .A(n7189), .ZN(n7191) );
  OAI21_X1 U7845 ( .B1(n7192), .B2(n4001), .A(n7191), .ZN(U3013) );
  NAND2_X1 U7846 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6946), .ZN(n7204)
         );
  OAI21_X1 U7847 ( .B1(n7195), .B2(n7194), .A(n7193), .ZN(n7196) );
  AND2_X1 U7848 ( .A1(n7197), .A2(n7196), .ZN(n7200) );
  OAI22_X1 U7849 ( .A1(n7215), .A2(n7258), .B1(n7198), .B2(n7213), .ZN(n7199)
         );
  AOI211_X1 U7850 ( .C1(n7201), .C2(n7239), .A(n7200), .B(n7199), .ZN(n7202)
         );
  OAI221_X1 U7851 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n7204), .C1(n4849), .C2(n7203), .A(n7202), .ZN(U3016) );
  AOI22_X1 U7852 ( .A1(n7295), .A2(n7238), .B1(n7205), .B2(REIP_REG_7__SCAN_IN), .ZN(n7208) );
  AOI22_X1 U7853 ( .A1(n7206), .A2(n7239), .B1(n7210), .B2(n7209), .ZN(n7207)
         );
  OAI211_X1 U7854 ( .C1(n7218), .C2(n7209), .A(n7208), .B(n7207), .ZN(U3011)
         );
  NAND2_X1 U7855 ( .A1(n7220), .A2(n7210), .ZN(n7234) );
  INV_X1 U7856 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7211) );
  AOI22_X1 U7857 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n7212), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n7211), .ZN(n7224) );
  OAI22_X1 U7858 ( .A1(n7216), .A2(n7215), .B1(n7214), .B2(n7213), .ZN(n7217)
         );
  INV_X1 U7859 ( .A(n7217), .ZN(n7223) );
  OAI21_X1 U7860 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7230) );
  AOI22_X1 U7861 ( .A1(n7221), .A2(n7239), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n7230), .ZN(n7222) );
  OAI211_X1 U7862 ( .C1(n7234), .C2(n7224), .A(n7223), .B(n7222), .ZN(U3008)
         );
  INV_X1 U7863 ( .A(n7225), .ZN(n7228) );
  INV_X1 U7864 ( .A(n7226), .ZN(n7227) );
  AOI21_X1 U7865 ( .B1(n7228), .B2(n7238), .A(n7227), .ZN(n7233) );
  INV_X1 U7866 ( .A(n7229), .ZN(n7231) );
  AOI22_X1 U7867 ( .A1(n7231), .A2(n7239), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n7230), .ZN(n7232) );
  OAI211_X1 U7868 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n7234), .A(n7233), 
        .B(n7232), .ZN(U3009) );
  AOI22_X1 U7869 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n7235), .B1(n7205), .B2(REIP_REG_15__SCAN_IN), .ZN(n7242) );
  INV_X1 U7870 ( .A(n7236), .ZN(n7240) );
  AOI22_X1 U7871 ( .A1(n7240), .A2(n7239), .B1(n7238), .B2(n7237), .ZN(n7241)
         );
  OAI211_X1 U7872 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n7243), .A(n7242), .B(n7241), .ZN(U3003) );
  NOR2_X1 U7873 ( .A1(n7415), .A2(REIP_REG_2__SCAN_IN), .ZN(n7244) );
  AOI22_X1 U7874 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7424), .B1(
        REIP_REG_1__SCAN_IN), .B2(n7244), .ZN(n7257) );
  INV_X1 U7875 ( .A(n7358), .ZN(n7245) );
  AOI211_X1 U7876 ( .C1(REIP_REG_1__SCAN_IN), .C2(n7390), .A(n7198), .B(n7245), 
        .ZN(n7254) );
  INV_X1 U7877 ( .A(n7246), .ZN(n7249) );
  INV_X1 U7878 ( .A(n7247), .ZN(n7248) );
  AOI22_X1 U7879 ( .A1(n7250), .A2(n7249), .B1(n7426), .B2(n7248), .ZN(n7251)
         );
  OAI21_X1 U7880 ( .B1(n7252), .B2(n7418), .A(n7251), .ZN(n7253) );
  AOI211_X1 U7881 ( .C1(n7255), .C2(n7278), .A(n7254), .B(n7253), .ZN(n7256)
         );
  OAI211_X1 U7882 ( .C1(n7431), .C2(n7258), .A(n7257), .B(n7256), .ZN(U2825)
         );
  NAND3_X1 U7883 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n7259) );
  NOR3_X1 U7884 ( .A1(n7415), .A2(REIP_REG_4__SCAN_IN), .A3(n7259), .ZN(n7260)
         );
  AOI211_X1 U7885 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7385), 
        .B(n7260), .ZN(n7270) );
  OAI22_X1 U7886 ( .A1(n7431), .A2(n7262), .B1(n7435), .B2(n7261), .ZN(n7268)
         );
  INV_X1 U7887 ( .A(n7263), .ZN(n7264) );
  OAI22_X1 U7888 ( .A1(n7266), .A2(n7265), .B1(n7264), .B2(n7412), .ZN(n7267)
         );
  AOI211_X1 U7889 ( .C1(EBX_REG_4__SCAN_IN), .C2(n7403), .A(n7268), .B(n7267), 
        .ZN(n7269) );
  OAI211_X1 U7890 ( .C1(n7272), .C2(n7271), .A(n7270), .B(n7269), .ZN(U2823)
         );
  AOI22_X1 U7891 ( .A1(EBX_REG_5__SCAN_IN), .A2(n7403), .B1(n7409), .B2(n7273), 
        .ZN(n7275) );
  OAI211_X1 U7892 ( .C1(n7405), .C2(n7276), .A(n7275), .B(n7274), .ZN(n7277)
         );
  AOI21_X1 U7893 ( .B1(n7279), .B2(n7278), .A(n7277), .ZN(n7283) );
  OAI21_X1 U7894 ( .B1(REIP_REG_5__SCAN_IN), .B2(n7281), .A(n7280), .ZN(n7282)
         );
  OAI211_X1 U7895 ( .C1(n7412), .C2(n7284), .A(n7283), .B(n7282), .ZN(U2822)
         );
  OAI22_X1 U7896 ( .A1(n7286), .A2(n7405), .B1(n7431), .B2(n7285), .ZN(n7287)
         );
  AOI211_X1 U7897 ( .C1(n7403), .C2(EBX_REG_6__SCAN_IN), .A(n7385), .B(n7287), 
        .ZN(n7288) );
  OAI221_X1 U7898 ( .B1(REIP_REG_6__SCAN_IN), .B2(n7298), .C1(n5271), .C2(
        n7299), .A(n7288), .ZN(n7289) );
  AOI21_X1 U7899 ( .B1(n7290), .B2(n7428), .A(n7289), .ZN(n7291) );
  OAI21_X1 U7900 ( .B1(n7292), .B2(n7412), .A(n7291), .ZN(U2821) );
  AOI22_X1 U7901 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n7424), .B1(
        EBX_REG_7__SCAN_IN), .B2(n7403), .ZN(n7293) );
  INV_X1 U7902 ( .A(n7293), .ZN(n7294) );
  AOI211_X1 U7903 ( .C1(n7409), .C2(n7295), .A(n7385), .B(n7294), .ZN(n7304)
         );
  OAI21_X1 U7904 ( .B1(REIP_REG_6__SCAN_IN), .B2(REIP_REG_7__SCAN_IN), .A(
        n7296), .ZN(n7297) );
  OAI22_X1 U7905 ( .A1(n7300), .A2(n7299), .B1(n7298), .B2(n7297), .ZN(n7301)
         );
  AOI21_X1 U7906 ( .B1(n7302), .B2(n7428), .A(n7301), .ZN(n7303) );
  OAI211_X1 U7907 ( .C1(n7305), .C2(n7412), .A(n7304), .B(n7303), .ZN(U2820)
         );
  NAND2_X1 U7908 ( .A1(n7307), .A2(n7306), .ZN(n7316) );
  AOI22_X1 U7909 ( .A1(n7409), .A2(n7308), .B1(REIP_REG_11__SCAN_IN), .B2(
        n7324), .ZN(n7309) );
  OAI21_X1 U7910 ( .B1(n7310), .B2(n7418), .A(n7309), .ZN(n7311) );
  AOI211_X1 U7911 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n7385), 
        .B(n7311), .ZN(n7315) );
  AOI22_X1 U7912 ( .A1(n7313), .A2(n7428), .B1(n7426), .B2(n7312), .ZN(n7314)
         );
  OAI211_X1 U7913 ( .C1(n7317), .C2(n7316), .A(n7315), .B(n7314), .ZN(U2816)
         );
  AOI22_X1 U7914 ( .A1(EBX_REG_13__SCAN_IN), .A2(n7403), .B1(n7409), .B2(n7318), .ZN(n7329) );
  NOR3_X1 U7915 ( .A1(n7415), .A2(REIP_REG_13__SCAN_IN), .A3(n7319), .ZN(n7320) );
  AOI211_X1 U7916 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n7385), 
        .B(n7320), .ZN(n7328) );
  INV_X1 U7917 ( .A(n7321), .ZN(n7323) );
  AOI22_X1 U7918 ( .A1(n7323), .A2(n7428), .B1(n7426), .B2(n7322), .ZN(n7327)
         );
  OAI21_X1 U7919 ( .B1(n7325), .B2(n7324), .A(REIP_REG_13__SCAN_IN), .ZN(n7326) );
  NAND4_X1 U7920 ( .A1(n7329), .A2(n7328), .A3(n7327), .A4(n7326), .ZN(U2814)
         );
  NOR2_X1 U7921 ( .A1(n7415), .A2(n7330), .ZN(n7331) );
  AOI22_X1 U7922 ( .A1(EBX_REG_14__SCAN_IN), .A2(n7403), .B1(n7332), .B2(n7331), .ZN(n7333) );
  OAI21_X1 U7923 ( .B1(n7343), .B2(n5915), .A(n7333), .ZN(n7334) );
  AOI211_X1 U7924 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n7385), 
        .B(n7334), .ZN(n7340) );
  INV_X1 U7925 ( .A(n7335), .ZN(n7338) );
  INV_X1 U7926 ( .A(n7336), .ZN(n7337) );
  AOI22_X1 U7927 ( .A1(n7338), .A2(n7428), .B1(n7337), .B2(n7426), .ZN(n7339)
         );
  OAI211_X1 U7928 ( .C1(n7431), .C2(n7341), .A(n7340), .B(n7339), .ZN(U2813)
         );
  XOR2_X1 U7929 ( .A(REIP_REG_16__SCAN_IN), .B(n7342), .Z(n7345) );
  OAI22_X1 U7930 ( .A1(n7346), .A2(n7345), .B1(n7344), .B2(n7343), .ZN(n7347)
         );
  AOI211_X1 U7931 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7385), 
        .B(n7347), .ZN(n7354) );
  INV_X1 U7932 ( .A(n7348), .ZN(n7350) );
  OAI22_X1 U7933 ( .A1(n7350), .A2(n7396), .B1(n7431), .B2(n7349), .ZN(n7351)
         );
  AOI21_X1 U7934 ( .B1(n7352), .B2(n7426), .A(n7351), .ZN(n7353) );
  OAI211_X1 U7935 ( .C1(n7355), .C2(n7418), .A(n7354), .B(n7353), .ZN(U2811)
         );
  INV_X1 U7936 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7367) );
  NAND2_X1 U7937 ( .A1(n7357), .A2(n7356), .ZN(n7369) );
  OAI21_X1 U7938 ( .B1(n7360), .B2(n7359), .A(n7358), .ZN(n7383) );
  AOI21_X1 U7939 ( .B1(n7368), .B2(n7369), .A(n7383), .ZN(n7361) );
  AOI211_X1 U7940 ( .C1(n7403), .C2(EBX_REG_17__SCAN_IN), .A(n7385), .B(n7361), 
        .ZN(n7366) );
  OAI22_X1 U7941 ( .A1(n7363), .A2(n7431), .B1(n7362), .B2(n7412), .ZN(n7364)
         );
  AOI21_X1 U7942 ( .B1(n7526), .B2(n7428), .A(n7364), .ZN(n7365) );
  OAI211_X1 U7943 ( .C1(n7367), .C2(n7405), .A(n7366), .B(n7365), .ZN(U2810)
         );
  OR2_X1 U7944 ( .A1(n7369), .A2(n7368), .ZN(n7392) );
  AOI22_X1 U7945 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7383), .B1(n7392), .B2(
        n7379), .ZN(n7370) );
  AOI211_X1 U7946 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n7385), 
        .B(n7370), .ZN(n7377) );
  INV_X1 U7947 ( .A(n7371), .ZN(n7372) );
  OAI22_X1 U7948 ( .A1(n7373), .A2(n7396), .B1(n7431), .B2(n7372), .ZN(n7374)
         );
  AOI21_X1 U7949 ( .B1(n7375), .B2(n7426), .A(n7374), .ZN(n7376) );
  OAI211_X1 U7950 ( .C1(n7378), .C2(n7418), .A(n7377), .B(n7376), .ZN(U2809)
         );
  AOI21_X1 U7951 ( .B1(n7379), .B2(n7382), .A(n7392), .ZN(n7380) );
  AOI22_X1 U7952 ( .A1(EBX_REG_19__SCAN_IN), .A2(n7403), .B1(n7380), .B2(n7393), .ZN(n7381) );
  OAI21_X1 U7953 ( .B1(n7383), .B2(n7382), .A(n7381), .ZN(n7384) );
  AOI211_X1 U7954 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7385), 
        .B(n7384), .ZN(n7388) );
  AOI22_X1 U7955 ( .A1(n7529), .A2(n7428), .B1(n7409), .B2(n7386), .ZN(n7387)
         );
  OAI211_X1 U7956 ( .C1(n7389), .C2(n7412), .A(n7388), .B(n7387), .ZN(U2808)
         );
  OAI21_X1 U7957 ( .B1(n7415), .B2(n7407), .A(n7390), .ZN(n7417) );
  OAI21_X1 U7958 ( .B1(n7393), .B2(n7392), .A(n7391), .ZN(n7394) );
  AOI22_X1 U7959 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n7424), .B1(n7417), 
        .B2(n7394), .ZN(n7401) );
  OAI22_X1 U7960 ( .A1(n7397), .A2(n7396), .B1(n7431), .B2(n7395), .ZN(n7398)
         );
  AOI21_X1 U7961 ( .B1(n7399), .B2(n7426), .A(n7398), .ZN(n7400) );
  OAI211_X1 U7962 ( .C1(n7402), .C2(n7418), .A(n7401), .B(n7400), .ZN(U2807)
         );
  NOR2_X1 U7963 ( .A1(n7415), .A2(REIP_REG_21__SCAN_IN), .ZN(n7416) );
  AOI22_X1 U7964 ( .A1(EBX_REG_21__SCAN_IN), .A2(n7403), .B1(
        REIP_REG_21__SCAN_IN), .B2(n7417), .ZN(n7404) );
  OAI21_X1 U7965 ( .B1(n4447), .B2(n7405), .A(n7404), .ZN(n7406) );
  AOI21_X1 U7966 ( .B1(n7407), .B2(n7416), .A(n7406), .ZN(n7411) );
  AOI22_X1 U7967 ( .A1(n7532), .A2(n7428), .B1(n7409), .B2(n7408), .ZN(n7410)
         );
  OAI211_X1 U7968 ( .C1(n7413), .C2(n7412), .A(n7411), .B(n7410), .ZN(U2806)
         );
  NOR3_X1 U7969 ( .A1(n7415), .A2(REIP_REG_22__SCAN_IN), .A3(n7414), .ZN(n7423) );
  NOR2_X1 U7970 ( .A1(n7417), .A2(n7416), .ZN(n7421) );
  OAI22_X1 U7971 ( .A1(n7421), .A2(n7420), .B1(n7419), .B2(n7418), .ZN(n7422)
         );
  AOI211_X1 U7972 ( .C1(n7424), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n7423), 
        .B(n7422), .ZN(n7430) );
  INV_X1 U7973 ( .A(n7425), .ZN(n7537) );
  AOI22_X1 U7974 ( .A1(n7537), .A2(n7428), .B1(n7427), .B2(n7426), .ZN(n7429)
         );
  OAI211_X1 U7975 ( .C1(n7432), .C2(n7431), .A(n7430), .B(n7429), .ZN(U2805)
         );
  OAI21_X1 U7976 ( .B1(n7434), .B2(n7443), .A(n7433), .ZN(U2793) );
  INV_X1 U7977 ( .A(n7435), .ZN(n7439) );
  NOR3_X1 U7978 ( .A1(n7436), .A2(STATE2_REG_1__SCAN_IN), .A3(
        STATE2_REG_3__SCAN_IN), .ZN(n7438) );
  NAND3_X1 U7979 ( .A1(n7439), .A2(n7438), .A3(n7437), .ZN(n7440) );
  OAI21_X1 U7980 ( .B1(n7441), .B2(n5171), .A(n7440), .ZN(U3455) );
  INV_X1 U7981 ( .A(MORE_REG_SCAN_IN), .ZN(n7442) );
  NAND2_X1 U7982 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  NAND2_X1 U7983 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  NAND3_X1 U7984 ( .A1(n7448), .A2(n7447), .A3(n7446), .ZN(n7449) );
  NOR2_X1 U7985 ( .A1(n7450), .A2(n7449), .ZN(n7451) );
  AND2_X1 U7986 ( .A1(n7452), .A2(n7451), .ZN(n7472) );
  INV_X1 U7987 ( .A(n7463), .ZN(n7465) );
  NAND2_X1 U7988 ( .A1(n7453), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7454) );
  NOR2_X1 U7989 ( .A1(n7455), .A2(n7454), .ZN(n7459) );
  NAND2_X1 U7990 ( .A1(n7459), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U7991 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  OAI21_X1 U7992 ( .B1(n7459), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n7458), 
        .ZN(n7460) );
  OAI211_X1 U7993 ( .C1(n7463), .C2(n7462), .A(n7461), .B(n7460), .ZN(n7464)
         );
  OAI21_X1 U7994 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7465), .A(n7464), 
        .ZN(n7466) );
  OAI21_X1 U7995 ( .B1(n7467), .B2(n4112), .A(n7466), .ZN(n7469) );
  NAND2_X1 U7996 ( .A1(n7467), .A2(n4112), .ZN(n7468) );
  NAND2_X1 U7997 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  NAND2_X1 U7998 ( .A1(n7470), .A2(n6991), .ZN(n7471) );
  AND2_X1 U7999 ( .A1(n7472), .A2(n7471), .ZN(n7500) );
  NAND2_X1 U8000 ( .A1(n7500), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U8001 ( .A1(READY_N), .A2(n7167), .ZN(n7474) );
  NAND2_X1 U8002 ( .A1(n7475), .A2(n7474), .ZN(n7479) );
  OR2_X1 U8003 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  NAND2_X1 U8004 ( .A1(n7479), .A2(n7478), .ZN(n7492) );
  OAI21_X1 U8005 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7513), .A(n7492), .ZN(
        n7480) );
  NAND2_X1 U8006 ( .A1(n7480), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7489) );
  NAND3_X1 U8007 ( .A1(n7481), .A2(STATE2_REG_0__SCAN_IN), .A3(n7513), .ZN(
        n7482) );
  NAND3_X1 U8008 ( .A1(n7482), .A2(n7499), .A3(n7492), .ZN(n7483) );
  OAI21_X1 U8009 ( .B1(n7484), .B2(n7492), .A(n7483), .ZN(n7486) );
  OAI211_X1 U8010 ( .C1(n7487), .C2(n7489), .A(n7486), .B(n7485), .ZN(U3149)
         );
  OAI221_X1 U8011 ( .B1(n4732), .B2(STATE2_REG_0__SCAN_IN), .C1(n4732), .C2(
        n7492), .A(n7491), .ZN(U3453) );
  OAI211_X1 U8012 ( .C1(n7491), .C2(n7490), .A(n7489), .B(n7488), .ZN(n7497)
         );
  INV_X1 U8013 ( .A(n7492), .ZN(n7493) );
  AOI211_X1 U8014 ( .C1(n7495), .C2(n7494), .A(STATE2_REG_0__SCAN_IN), .B(
        n7493), .ZN(n7496) );
  NOR2_X1 U8015 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  OAI21_X1 U8016 ( .B1(n7500), .B2(n7499), .A(n7498), .ZN(U3148) );
  OAI21_X1 U8017 ( .B1(n7503), .B2(n7502), .A(n7501), .ZN(U2792) );
  AOI21_X1 U8018 ( .B1(n7505), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n7504), .ZN(
        n7506) );
  INV_X1 U8019 ( .A(n7506), .ZN(U3452) );
  NAND2_X1 U8020 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7511) );
  INV_X1 U8021 ( .A(n7507), .ZN(n7516) );
  INV_X1 U8022 ( .A(NA_N), .ZN(n7517) );
  AOI221_X1 U8023 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7517), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7521) );
  AOI221_X1 U8024 ( .B1(n7516), .B2(n7509), .C1(n7508), .C2(n7509), .A(n7521), 
        .ZN(n7510) );
  OAI221_X1 U8025 ( .B1(n7525), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7525), 
        .C2(n7511), .A(n7510), .ZN(U3181) );
  OAI21_X1 U8026 ( .B1(NA_N), .B2(n7513), .A(n7512), .ZN(n7514) );
  OAI211_X1 U8027 ( .C1(STATE_REG_2__SCAN_IN), .C2(n7515), .A(HOLD), .B(n7514), 
        .ZN(n7520) );
  OAI221_X1 U8028 ( .B1(STATE_REG_2__SCAN_IN), .B2(n7518), .C1(
        STATE_REG_2__SCAN_IN), .C2(n7517), .A(n7516), .ZN(n7519) );
  OAI221_X1 U8029 ( .B1(n7521), .B2(STATE_REG_0__SCAN_IN), .C1(n7521), .C2(
        n7520), .A(n7519), .ZN(U3183) );
  AOI22_X1 U8030 ( .A1(n7525), .A2(n7524), .B1(n7523), .B2(n7522), .ZN(U3473)
         );
  AOI22_X1 U8031 ( .A1(n7526), .A2(n7536), .B1(n7535), .B2(DATAI_17_), .ZN(
        n7528) );
  AOI22_X1 U8032 ( .A1(n7539), .A2(DATAI_1_), .B1(n7538), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U8033 ( .A1(n7528), .A2(n7527), .ZN(U2874) );
  AOI22_X1 U8034 ( .A1(n7529), .A2(n7536), .B1(n7535), .B2(DATAI_19_), .ZN(
        n7531) );
  AOI22_X1 U8035 ( .A1(n7539), .A2(DATAI_3_), .B1(n7538), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U8036 ( .A1(n7531), .A2(n7530), .ZN(U2872) );
  AOI22_X1 U8037 ( .A1(n7532), .A2(n7536), .B1(n7535), .B2(DATAI_21_), .ZN(
        n7534) );
  AOI22_X1 U8038 ( .A1(n7539), .A2(DATAI_5_), .B1(n7538), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U8039 ( .A1(n7534), .A2(n7533), .ZN(U2870) );
  AOI22_X1 U8040 ( .A1(n7537), .A2(n7536), .B1(n7535), .B2(DATAI_22_), .ZN(
        n7541) );
  AOI22_X1 U8041 ( .A1(n7539), .A2(DATAI_6_), .B1(n7538), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n7540) );
  NAND2_X1 U8042 ( .A1(n7541), .A2(n7540), .ZN(U2869) );
  INV_X1 U8043 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n7549) );
  INV_X1 U8044 ( .A(n7542), .ZN(n7565) );
  AOI22_X1 U8045 ( .A1(n7544), .A2(n7566), .B1(n7565), .B2(n7543), .ZN(n7548)
         );
  AOI22_X1 U8046 ( .A1(n7571), .A2(n7546), .B1(n7569), .B2(n7545), .ZN(n7547)
         );
  OAI211_X1 U8047 ( .C1(n7575), .C2(n7549), .A(n7548), .B(n7547), .ZN(U3020)
         );
  AOI22_X1 U8048 ( .A1(n7551), .A2(n7566), .B1(n7565), .B2(n7550), .ZN(n7555)
         );
  AOI22_X1 U8049 ( .A1(n7571), .A2(n7553), .B1(n7569), .B2(n7552), .ZN(n7554)
         );
  OAI211_X1 U8050 ( .C1(n7575), .C2(n7556), .A(n7555), .B(n7554), .ZN(U3021)
         );
  INV_X1 U8051 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n7563) );
  AOI22_X1 U8052 ( .A1(n7558), .A2(n7566), .B1(n7565), .B2(n7557), .ZN(n7562)
         );
  AOI22_X1 U8053 ( .A1(n7571), .A2(n7560), .B1(n7569), .B2(n7559), .ZN(n7561)
         );
  OAI211_X1 U8054 ( .C1(n7575), .C2(n7563), .A(n7562), .B(n7561), .ZN(U3024)
         );
  INV_X1 U8055 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n7574) );
  AOI22_X1 U8056 ( .A1(n7567), .A2(n7566), .B1(n7565), .B2(n7564), .ZN(n7573)
         );
  AOI22_X1 U8057 ( .A1(n7571), .A2(n7570), .B1(n7569), .B2(n7568), .ZN(n7572)
         );
  OAI211_X1 U8058 ( .C1(n7575), .C2(n7574), .A(n7573), .B(n7572), .ZN(U3025)
         );
  NOR2_X1 U6656 ( .A1(n6193), .A2(n5960), .ZN(n5961) );
  CLKBUF_X1 U3698 ( .A(n3836), .Z(n3683) );
  CLKBUF_X1 U3739 ( .A(n3838), .Z(n5974) );
  CLKBUF_X1 U3751 ( .A(n3760), .Z(n4753) );
  CLKBUF_X1 U3993 ( .A(n4618), .Z(n4736) );
  NAND2_X1 U4152 ( .A1(n6024), .A2(n5958), .ZN(n6193) );
  CLKBUF_X1 U6653 ( .A(n6992), .Z(n7022) );
endmodule

