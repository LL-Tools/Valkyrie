

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859;

  AND2_X1 U4994 ( .A1(n9850), .A2(n9853), .ZN(n9935) );
  OR2_X1 U4995 ( .A1(n10590), .A2(n10591), .ZN(n10588) );
  XNOR2_X1 U4996 ( .A(n6879), .B(n10563), .ZN(n10573) );
  INV_X2 U4997 ( .A(n7350), .ZN(n8722) );
  AND2_X1 U4998 ( .A1(n8649), .A2(n8659), .ZN(n8590) );
  CLKBUF_X2 U4999 ( .A(n5713), .Z(n8596) );
  INV_X2 U5000 ( .A(n7785), .ZN(n9425) );
  MUX2_X1 U5001 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6217), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n6219) );
  OR2_X1 U5002 ( .A1(n6873), .A2(n6875), .ZN(n5354) );
  OAI21_X1 U5003 ( .B1(n10506), .B2(n5354), .A(n5353), .ZN(n6876) );
  NAND2_X1 U5004 ( .A1(n5365), .A2(n5363), .ZN(n6887) );
  INV_X1 U5005 ( .A(n8590), .ZN(n8576) );
  INV_X1 U5006 ( .A(n7349), .ZN(n7453) );
  NOR2_X1 U5007 ( .A1(n8376), .A2(n8268), .ZN(n5341) );
  NAND2_X1 U5008 ( .A1(n6410), .A2(n6409), .ZN(n7684) );
  NOR2_X1 U5009 ( .A1(n8946), .A2(n5351), .ZN(n10491) );
  NOR2_X1 U5010 ( .A1(n10573), .A2(n10572), .ZN(n10571) );
  XNOR2_X1 U5011 ( .A(n6882), .B(n7309), .ZN(n10607) );
  NOR2_X1 U5012 ( .A1(n10639), .A2(n10638), .ZN(n10637) );
  XNOR2_X1 U5013 ( .A(n8803), .B(n8966), .ZN(n8795) );
  AND2_X1 U5014 ( .A1(n5779), .A2(n5778), .ZN(n7669) );
  AND3_X1 U5015 ( .A1(n5748), .A2(n5747), .A3(n5746), .ZN(n7544) );
  NAND2_X1 U5016 ( .A1(n6810), .A2(n6747), .ZN(n8197) );
  NAND2_X1 U5017 ( .A1(n6514), .A2(n6513), .ZN(n8268) );
  OR2_X1 U5018 ( .A1(n6395), .A2(n6394), .ZN(n7834) );
  NAND2_X1 U5019 ( .A1(n6451), .A2(n6450), .ZN(n8142) );
  AND4_X1 U5020 ( .A1(n6406), .A2(n6405), .A3(n6404), .A4(n6403), .ZN(n7785)
         );
  NAND2_X1 U5021 ( .A1(n5843), .A2(n5610), .ZN(n5846) );
  INV_X1 U5022 ( .A(n9412), .ZN(n5338) );
  NOR2_X1 U5023 ( .A1(n8284), .A2(n8928), .ZN(n4930) );
  XOR2_X1 U5024 ( .A(n8454), .B(n8801), .Z(n4931) );
  NAND2_X2 U5025 ( .A1(n5437), .A2(n5438), .ZN(n9645) );
  XNOR2_X2 U5026 ( .A(n6229), .B(n6228), .ZN(n6239) );
  NAND2_X2 U5027 ( .A1(n9987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  NAND2_X4 U5028 ( .A1(n5062), .A2(n5061), .ZN(n5586) );
  NAND2_X2 U5029 ( .A1(n6063), .A2(n6062), .ZN(n9195) );
  INV_X2 U5030 ( .A(n6238), .ZN(n5034) );
  XNOR2_X2 U5031 ( .A(n6223), .B(n6225), .ZN(n6238) );
  XNOR2_X2 U5032 ( .A(n6158), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8281) );
  NOR2_X2 U5033 ( .A1(n10507), .A2(n10508), .ZN(n10506) );
  XNOR2_X2 U5034 ( .A(n6254), .B(n6255), .ZN(n6253) );
  NAND2_X2 U5035 ( .A1(n6200), .A2(n6199), .ZN(n6254) );
  XNOR2_X2 U5036 ( .A(n5317), .B(n5678), .ZN(n6967) );
  AOI21_X2 U5037 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7247), .A(n10555), .ZN(
        n6879) );
  NAND2_X2 U5038 ( .A1(n6428), .A2(n6427), .ZN(n9841) );
  AND2_X1 U5039 ( .A1(n9784), .A2(n9580), .ZN(n5545) );
  NAND2_X2 U5040 ( .A1(n9425), .A2(n7784), .ZN(n6795) );
  NAND2_X1 U5041 ( .A1(n7836), .A2(n6716), .ZN(n7809) );
  INV_X1 U5042 ( .A(n7820), .ZN(n10744) );
  INV_X1 U5043 ( .A(n7590), .ZN(n7585) );
  XNOR2_X1 U5044 ( .A(n6363), .B(n10735), .ZN(n7557) );
  INV_X1 U5045 ( .A(n7554), .ZN(n7774) );
  CLKBUF_X2 U5047 ( .A(n5376), .Z(n4935) );
  INV_X1 U5048 ( .A(n7553), .ZN(n4933) );
  NAND2_X1 U5049 ( .A1(n8109), .A2(n10222), .ZN(n7553) );
  INV_X1 U5050 ( .A(n6357), .ZN(n5376) );
  INV_X1 U5052 ( .A(n6673), .ZN(n6340) );
  AND2_X1 U5053 ( .A1(n5217), .A2(n5216), .ZN(n6336) );
  OAI21_X1 U5054 ( .B1(n6781), .B2(n6780), .A(n7563), .ZN(n6782) );
  NOR2_X1 U5055 ( .A1(n9858), .A2(n5247), .ZN(n5032) );
  AND2_X1 U5056 ( .A1(n9626), .A2(n9625), .ZN(n9864) );
  NAND2_X1 U5057 ( .A1(n5547), .A2(n7173), .ZN(n7186) );
  OR2_X1 U5058 ( .A1(n6150), .A2(n9165), .ZN(n5562) );
  NOR4_X1 U5059 ( .A1(n6731), .A2(n6730), .A3(n6832), .A4(n6770), .ZN(n6774)
         );
  NAND2_X1 U5060 ( .A1(n7157), .A2(n7156), .ZN(n8608) );
  OR2_X1 U5061 ( .A1(n6729), .A2(n9567), .ZN(n6768) );
  OR2_X1 U5062 ( .A1(n8586), .A2(n8587), .ZN(n8592) );
  AND2_X1 U5063 ( .A1(n8595), .A2(n8594), .ZN(n9178) );
  NAND2_X1 U5064 ( .A1(n8453), .A2(n8452), .ZN(n8586) );
  NAND2_X1 U5065 ( .A1(n6264), .A2(n6263), .ZN(n9557) );
  CLKBUF_X1 U5066 ( .A(n9726), .Z(n5031) );
  OAI21_X1 U5067 ( .B1(n9726), .B2(n5447), .A(n5446), .ZN(n9589) );
  NAND2_X1 U5068 ( .A1(n9653), .A2(n9944), .ZN(n9640) );
  AOI21_X1 U5069 ( .B1(n4944), .B2(n8568), .A(n5038), .ZN(n5037) );
  AOI21_X1 U5070 ( .B1(n5233), .B2(n5236), .A(n5232), .ZN(n5231) );
  XNOR2_X1 U5071 ( .A(n6691), .B(n6690), .ZN(n9257) );
  INV_X1 U5072 ( .A(n9637), .ZN(n9653) );
  NAND2_X1 U5073 ( .A1(n6221), .A2(n6220), .ZN(n9560) );
  NAND2_X1 U5074 ( .A1(n6144), .A2(n6143), .ZN(n8993) );
  AND2_X1 U5075 ( .A1(n8567), .A2(n8566), .ZN(n8978) );
  NAND2_X1 U5076 ( .A1(n9607), .A2(n9606), .ZN(n9714) );
  AND2_X1 U5077 ( .A1(n8613), .A2(n8612), .ZN(n8994) );
  NAND2_X1 U5078 ( .A1(n6643), .A2(n6642), .ZN(n9672) );
  NAND2_X1 U5079 ( .A1(n5444), .A2(n5442), .ZN(n9784) );
  NAND2_X1 U5080 ( .A1(n6074), .A2(n6073), .ZN(n8678) );
  NAND2_X1 U5081 ( .A1(n9605), .A2(n9604), .ZN(n9727) );
  NAND2_X1 U5082 ( .A1(n5681), .A2(n5680), .ZN(n9185) );
  NOR2_X1 U5083 ( .A1(n10675), .A2(n10674), .ZN(n10673) );
  AOI21_X1 U5084 ( .B1(n5270), .B2(n4943), .A(n8559), .ZN(n5269) );
  NAND2_X1 U5085 ( .A1(n6050), .A2(n6049), .ZN(n9201) );
  NAND2_X1 U5086 ( .A1(n6612), .A2(n6611), .ZN(n9885) );
  NAND2_X1 U5087 ( .A1(n6280), .A2(n6279), .ZN(n9736) );
  NAND2_X1 U5088 ( .A1(n6018), .A2(n6017), .ZN(n9053) );
  NAND2_X1 U5089 ( .A1(n6290), .A2(n6289), .ZN(n9754) );
  NAND2_X1 U5090 ( .A1(n6272), .A2(n6271), .ZN(n9889) );
  AOI21_X1 U5091 ( .B1(n5243), .B2(n9575), .A(n5242), .ZN(n5241) );
  AOI21_X1 U5092 ( .B1(n8308), .B2(n5245), .A(n5244), .ZN(n5243) );
  NAND2_X1 U5093 ( .A1(n6580), .A2(n6579), .ZN(n9919) );
  AND2_X1 U5094 ( .A1(n6710), .A2(n6748), .ZN(n8173) );
  OAI211_X1 U5095 ( .C1(n5043), .C2(n5046), .A(n5045), .B(n8504), .ZN(n8224)
         );
  OR2_X1 U5096 ( .A1(n5047), .A2(n5043), .ZN(n5045) );
  NAND2_X1 U5097 ( .A1(n6566), .A2(n6565), .ZN(n9577) );
  INV_X1 U5098 ( .A(n10815), .ZN(n8376) );
  AND2_X1 U5099 ( .A1(n7975), .A2(n8090), .ZN(n8018) );
  AOI21_X1 U5100 ( .B1(n8096), .B2(n5532), .A(n4999), .ZN(n5531) );
  NAND2_X1 U5101 ( .A1(n6484), .A2(n6483), .ZN(n8390) );
  OR2_X1 U5102 ( .A1(n8165), .A2(n8289), .ZN(n8509) );
  OAI21_X2 U5103 ( .B1(n7248), .B2(n5741), .A(n5849), .ZN(n5856) );
  NAND2_X2 U5104 ( .A1(n7628), .A2(n10829), .ZN(n10837) );
  OAI21_X1 U5105 ( .B1(n6365), .B2(n7557), .A(n6364), .ZN(n7811) );
  NAND2_X1 U5106 ( .A1(n5597), .A2(n5596), .ZN(n5812) );
  INV_X2 U5107 ( .A(n10712), .ZN(n4932) );
  AND2_X1 U5108 ( .A1(n5352), .A2(n7207), .ZN(n8946) );
  OAI211_X2 U5109 ( .C1(n6625), .C2(n7205), .A(n6377), .B(n6376), .ZN(n7820)
         );
  INV_X1 U5110 ( .A(n7517), .ZN(n7538) );
  OAI211_X1 U5111 ( .C1(P1_DATAO_REG_1__SCAN_IN), .C2(n5774), .A(n5727), .B(
        n4995), .ZN(n7590) );
  AND3_X1 U5112 ( .A1(n5289), .A2(n5736), .A3(n5288), .ZN(n7517) );
  NAND2_X1 U5113 ( .A1(n4968), .A2(n5357), .ZN(n7396) );
  NAND2_X1 U5114 ( .A1(n7763), .A2(n5117), .ZN(n7349) );
  INV_X1 U5115 ( .A(n7560), .ZN(n10226) );
  AND4_X1 U5116 ( .A1(n5842), .A2(n5841), .A3(n5840), .A4(n5839), .ZN(n8289)
         );
  INV_X1 U5117 ( .A(n7661), .ZN(n7527) );
  XNOR2_X1 U5118 ( .A(n6105), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8649) );
  AND2_X1 U5119 ( .A1(n5358), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5357) );
  NAND4_X2 U5120 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .ZN(n6363)
         );
  NAND2_X1 U5121 ( .A1(n6104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U5122 ( .A1(n6157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6158) );
  INV_X1 U5123 ( .A(n5774), .ZN(n5994) );
  CLKBUF_X3 U5124 ( .A(n6666), .Z(n4938) );
  AND2_X2 U5126 ( .A1(n8690), .A2(n9265), .ZN(n5764) );
  AND2_X1 U5127 ( .A1(n5595), .A2(n5593), .ZN(n5490) );
  NAND2_X1 U5128 ( .A1(n6102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6106) );
  AND2_X1 U5129 ( .A1(n6161), .A2(n6160), .ZN(n6166) );
  CLKBUF_X3 U5130 ( .A(n6350), .Z(n6670) );
  INV_X2 U5131 ( .A(n6962), .ZN(n8788) );
  OR2_X1 U5132 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  AND2_X2 U5133 ( .A1(n6357), .A2(n7195), .ZN(n6666) );
  OAI21_X1 U5134 ( .B1(n5464), .B2(n5462), .A(n4997), .ZN(n5461) );
  NAND2_X4 U5135 ( .A1(n7002), .A2(n6967), .ZN(n5726) );
  XNOR2_X1 U5136 ( .A(n5684), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5691) );
  NOR2_X1 U5137 ( .A1(n7329), .A2(n6866), .ZN(n7316) );
  OR2_X1 U5138 ( .A1(n5889), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5905) );
  NOR2_X1 U5139 ( .A1(n4985), .A2(n5055), .ZN(n5054) );
  AND2_X1 U5140 ( .A1(n5569), .A2(n5570), .ZN(n5718) );
  OAI21_X1 U5141 ( .B1(n5993), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6101) );
  XNOR2_X1 U5142 ( .A(n5677), .B(n5285), .ZN(n7002) );
  NAND2_X1 U5143 ( .A1(n6160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U5144 ( .A1(n5682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5677) );
  AND2_X1 U5145 ( .A1(n4971), .A2(n5541), .ZN(n5686) );
  AND2_X1 U5146 ( .A1(n5725), .A2(n6904), .ZN(n6864) );
  NAND2_X1 U5147 ( .A1(n5745), .A2(n5744), .ZN(n8449) );
  AND2_X1 U5148 ( .A1(n5977), .A2(n5006), .ZN(n5286) );
  AND3_X1 U5149 ( .A1(n5672), .A2(n5671), .A3(n5707), .ZN(n5977) );
  INV_X1 U5150 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6250) );
  INV_X1 U5151 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6103) );
  NOR2_X1 U5152 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5666) );
  INV_X1 U5153 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6850) );
  INV_X1 U5154 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5707) );
  NOR2_X1 U5155 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5373) );
  NOR2_X1 U5156 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5374) );
  INV_X1 U5157 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6153) );
  INV_X1 U5158 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5981) );
  INV_X1 U5159 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6100) );
  CLKBUF_X1 U5160 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10302) );
  INV_X1 U5161 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5667) );
  NOR2_X2 U5162 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6386) );
  INV_X1 U5163 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7656) );
  OR2_X1 U5164 ( .A1(n9861), .A2(n10810), .ZN(n5033) );
  INV_X2 U5165 ( .A(n7050), .ZN(n7474) );
  NAND2_X2 U5166 ( .A1(n7069), .A2(n8351), .ZN(n8284) );
  NOR4_X2 U5167 ( .A1(n8646), .A2(n8645), .A3(n8605), .A4(n8644), .ZN(n8650)
         );
  NAND2_X1 U5168 ( .A1(n5845), .A2(n5846), .ZN(n7248) );
  INV_X1 U5169 ( .A(n8966), .ZN(n4936) );
  INV_X1 U5170 ( .A(n4936), .ZN(n4937) );
  NOR2_X2 U5171 ( .A1(n9789), .A2(n9906), .ZN(n9774) );
  OAI21_X2 U5172 ( .B1(n6165), .B2(P2_D_REG_0__SCAN_IN), .A(n6163), .ZN(n6164)
         );
  NAND4_X2 U5173 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5099), .ZN(n5668)
         );
  XNOR2_X2 U5174 ( .A(n7111), .B(n7112), .ZN(n8815) );
  NAND2_X2 U5175 ( .A1(n8875), .A2(n7110), .ZN(n7111) );
  NAND2_X2 U5176 ( .A1(n6309), .A2(n6308), .ZN(n9412) );
  AOI21_X2 U5177 ( .B1(n8670), .B2(n7125), .A(n5546), .ZN(n8793) );
  INV_X1 U5178 ( .A(n7474), .ZN(n4940) );
  INV_X4 U5179 ( .A(n7474), .ZN(n8794) );
  BUF_X4 U5180 ( .A(n6348), .Z(n6669) );
  AOI21_X1 U5181 ( .B1(n5298), .B2(n5301), .A(n5003), .ZN(n5296) );
  INV_X1 U5182 ( .A(n5561), .ZN(n5301) );
  AND2_X1 U5183 ( .A1(n5542), .A2(n5678), .ZN(n5541) );
  AOI21_X1 U5184 ( .B1(n5448), .B2(n5450), .A(n4982), .ZN(n5446) );
  INV_X1 U5185 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6202) );
  INV_X1 U5186 ( .A(n6372), .ZN(n6393) );
  NAND2_X1 U5187 ( .A1(n5086), .A2(n5084), .ZN(n6606) );
  NOR2_X1 U5188 ( .A1(n9575), .A2(n5085), .ZN(n5084) );
  NAND2_X1 U5189 ( .A1(n6562), .A2(n5087), .ZN(n5086) );
  NAND2_X1 U5190 ( .A1(n5083), .A2(n5082), .ZN(n5085) );
  NAND2_X1 U5191 ( .A1(n4963), .A2(n5208), .ZN(n5207) );
  INV_X1 U5192 ( .A(n8560), .ZN(n5208) );
  NOR2_X1 U5193 ( .A1(n5543), .A2(n5676), .ZN(n5542) );
  NAND2_X1 U5194 ( .A1(n5544), .A2(n5674), .ZN(n5543) );
  INV_X1 U5195 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5544) );
  AND2_X1 U5196 ( .A1(n9630), .A2(n5234), .ZN(n5233) );
  NAND2_X1 U5197 ( .A1(n5235), .A2(n9612), .ZN(n5234) );
  INV_X1 U5198 ( .A(n5943), .ZN(n5482) );
  INV_X1 U5199 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U5200 ( .A1(n7406), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U5201 ( .A1(n8941), .A2(n5102), .ZN(n6909) );
  OR2_X1 U5202 ( .A1(n8944), .A2(n6908), .ZN(n5102) );
  INV_X1 U5203 ( .A(n8514), .ZN(n8504) );
  NAND2_X1 U5204 ( .A1(n7942), .A2(n6125), .ZN(n5046) );
  INV_X1 U5205 ( .A(n8490), .ZN(n5260) );
  INV_X1 U5206 ( .A(n8495), .ZN(n5259) );
  OR2_X1 U5207 ( .A1(n9226), .A2(n9063), .ZN(n8547) );
  NAND2_X1 U5208 ( .A1(n5405), .A2(n5130), .ZN(n5129) );
  INV_X1 U5209 ( .A(n5131), .ZN(n5130) );
  AOI21_X1 U5210 ( .B1(n5425), .B2(n5426), .A(n5424), .ZN(n5423) );
  INV_X1 U5211 ( .A(n8365), .ZN(n5424) );
  BUF_X1 U5212 ( .A(n7451), .Z(n8767) );
  NAND2_X1 U5213 ( .A1(n9597), .A2(n5228), .ZN(n5227) );
  NAND2_X1 U5214 ( .A1(n5231), .A2(n5229), .ZN(n5228) );
  INV_X1 U5215 ( .A(n5233), .ZN(n5229) );
  NAND2_X1 U5216 ( .A1(n9614), .A2(n5231), .ZN(n5226) );
  NAND2_X1 U5217 ( .A1(n9767), .A2(n5246), .ZN(n9605) );
  AND2_X1 U5218 ( .A1(n6822), .A2(n6823), .ZN(n5246) );
  INV_X1 U5219 ( .A(n6059), .ZN(n5661) );
  AOI21_X1 U5220 ( .B1(n5466), .B2(n5813), .A(n4998), .ZN(n5464) );
  NAND2_X1 U5221 ( .A1(n5491), .A2(n5490), .ZN(n5597) );
  INV_X1 U5222 ( .A(n8857), .ZN(n7103) );
  OAI21_X1 U5223 ( .B1(n5511), .B2(n4947), .A(n8864), .ZN(n5510) );
  AOI21_X1 U5224 ( .B1(n7897), .B2(n5527), .A(n5526), .ZN(n7068) );
  INV_X1 U5225 ( .A(n5531), .ZN(n5526) );
  NOR2_X1 U5226 ( .A1(n5533), .A2(n5528), .ZN(n5527) );
  OAI21_X1 U5227 ( .B1(n5523), .B2(n4987), .A(n5520), .ZN(n5519) );
  NAND2_X1 U5228 ( .A1(n5523), .A2(n8671), .ZN(n5520) );
  INV_X1 U5229 ( .A(n8671), .ZN(n5521) );
  NAND2_X1 U5230 ( .A1(n7083), .A2(n7082), .ZN(n8807) );
  NAND2_X1 U5232 ( .A1(n6884), .A2(n5368), .ZN(n5364) );
  NAND2_X1 U5233 ( .A1(n5297), .A2(n5561), .ZN(n7162) );
  INV_X1 U5234 ( .A(n8509), .ZN(n5279) );
  OR2_X1 U5235 ( .A1(n9016), .A2(n9026), .ZN(n5316) );
  OR2_X1 U5236 ( .A1(n9141), .A2(n9048), .ZN(n9039) );
  AOI21_X1 U5237 ( .B1(n5332), .B2(n5334), .A(n5001), .ZN(n5331) );
  NAND2_X1 U5238 ( .A1(n9097), .A2(n5018), .ZN(n9079) );
  INV_X1 U5239 ( .A(n9106), .ZN(n9082) );
  AND2_X1 U5240 ( .A1(n5777), .A2(n5550), .ZN(n5778) );
  NOR2_X1 U5241 ( .A1(n9255), .A2(n8344), .ZN(n7187) );
  NAND2_X1 U5242 ( .A1(n8606), .A2(n7127), .ZN(n9103) );
  NAND2_X1 U5243 ( .A1(n9258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5684) );
  OR2_X1 U5244 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  AND2_X1 U5245 ( .A1(n8762), .A2(n5418), .ZN(n5417) );
  NAND2_X1 U5246 ( .A1(n5420), .A2(n5422), .ZN(n5418) );
  NAND2_X1 U5247 ( .A1(n5070), .A2(n6705), .ZN(n6781) );
  OAI211_X1 U5248 ( .C1(n6700), .C2(n6701), .A(n6699), .B(n6698), .ZN(n5070)
         );
  INV_X1 U5249 ( .A(n6673), .ZN(n6590) );
  NAND2_X1 U5250 ( .A1(n6239), .A2(n5034), .ZN(n6350) );
  AND2_X1 U5251 ( .A1(n6238), .A2(n9991), .ZN(n6348) );
  OR2_X1 U5252 ( .A1(n9624), .A2(n9630), .ZN(n9626) );
  NAND2_X1 U5253 ( .A1(n5239), .A2(n5237), .ZN(n9704) );
  NOR2_X1 U5254 ( .A1(n9700), .A2(n5238), .ZN(n5237) );
  INV_X1 U5255 ( .A(n9608), .ZN(n5238) );
  AOI21_X1 U5256 ( .B1(n5451), .B2(n5449), .A(n4988), .ZN(n5448) );
  INV_X1 U5257 ( .A(n4961), .ZN(n5449) );
  NAND2_X1 U5258 ( .A1(n9578), .A2(n4962), .ZN(n5444) );
  AND2_X1 U5259 ( .A1(n7569), .A2(n9440), .ZN(n10225) );
  NAND2_X1 U5260 ( .A1(n6694), .A2(n6693), .ZN(n9568) );
  NOR2_X1 U5261 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n6209), .ZN(n5336) );
  NAND2_X1 U5262 ( .A1(n6850), .A2(n6208), .ZN(n6209) );
  INV_X1 U5263 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U5264 ( .A1(n5705), .A2(n5627), .ZN(n5944) );
  NOR2_X1 U5265 ( .A1(n5897), .A2(n5473), .ZN(n5468) );
  INV_X1 U5266 ( .A(n5726), .ZN(n6862) );
  NAND2_X1 U5267 ( .A1(n6091), .A2(n6090), .ZN(n8803) );
  OAI21_X1 U5268 ( .B1(n8489), .B2(n5251), .A(n4989), .ZN(n5210) );
  OAI21_X1 U5269 ( .B1(n8489), .B2(n8485), .A(n4972), .ZN(n5212) );
  NAND2_X1 U5270 ( .A1(n8505), .A2(n8504), .ZN(n5172) );
  NAND2_X1 U5271 ( .A1(n8516), .A2(n8515), .ZN(n5175) );
  NAND2_X1 U5272 ( .A1(n6606), .A2(n4980), .ZN(n6594) );
  NAND2_X1 U5273 ( .A1(n8557), .A2(n8556), .ZN(n5201) );
  OAI21_X1 U5274 ( .B1(n5191), .B2(n5189), .A(n5185), .ZN(n8545) );
  INV_X1 U5275 ( .A(n5207), .ZN(n5199) );
  NOR2_X1 U5276 ( .A1(n5207), .A2(n4994), .ZN(n5202) );
  NAND2_X1 U5277 ( .A1(n5206), .A2(n5204), .ZN(n5203) );
  NAND2_X1 U5278 ( .A1(n6610), .A2(n9606), .ZN(n5090) );
  AND2_X1 U5279 ( .A1(n8625), .A2(n8626), .ZN(n5875) );
  NAND2_X1 U5280 ( .A1(n7040), .A2(n7590), .ZN(n8473) );
  AND2_X1 U5281 ( .A1(n7451), .A2(n7349), .ZN(n7448) );
  NOR2_X1 U5282 ( .A1(n9597), .A2(n6681), .ZN(n6682) );
  AOI21_X1 U5283 ( .B1(n6656), .B2(n6655), .A(n5235), .ZN(n5066) );
  INV_X1 U5284 ( .A(SI_17_), .ZN(n10137) );
  NAND3_X1 U5285 ( .A1(n5060), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5061) );
  INV_X1 U5286 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5063) );
  NAND2_X1 U5287 ( .A1(n8608), .A2(n8607), .ZN(n5051) );
  NOR2_X1 U5288 ( .A1(n5267), .A2(n4983), .ZN(n5050) );
  OR2_X1 U5289 ( .A1(n8605), .A2(n8606), .ZN(n5267) );
  NAND2_X1 U5290 ( .A1(n6906), .A2(n5105), .ZN(n5104) );
  OR2_X1 U5291 ( .A1(n5359), .A2(n7206), .ZN(n5105) );
  AND2_X1 U5292 ( .A1(n6906), .A2(n7206), .ZN(n5111) );
  OR2_X1 U5293 ( .A1(n7408), .A2(n4970), .ZN(n5352) );
  NAND2_X1 U5294 ( .A1(n10515), .A2(n6911), .ZN(n6912) );
  NAND2_X1 U5295 ( .A1(n10547), .A2(n6914), .ZN(n6915) );
  NAND2_X1 U5296 ( .A1(n5669), .A2(n5505), .ZN(n5504) );
  INV_X1 U5297 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U5298 ( .A1(n10580), .A2(n6917), .ZN(n6918) );
  NAND2_X1 U5299 ( .A1(n10614), .A2(n6920), .ZN(n6921) );
  NAND2_X1 U5300 ( .A1(n10654), .A2(n5362), .ZN(n5361) );
  NOR2_X1 U5301 ( .A1(n5276), .A2(n5048), .ZN(n5047) );
  INV_X1 U5302 ( .A(n8498), .ZN(n5048) );
  NAND2_X1 U5303 ( .A1(n7041), .A2(n7585), .ZN(n8475) );
  OR2_X1 U5304 ( .A1(n9185), .A2(n8976), .ZN(n8572) );
  AND2_X1 U5305 ( .A1(n8459), .A2(n8458), .ZN(n8614) );
  NOR2_X1 U5306 ( .A1(n9071), .A2(n5333), .ZN(n5332) );
  NOR2_X1 U5307 ( .A1(n5990), .A2(n5334), .ZN(n5333) );
  NOR2_X1 U5308 ( .A1(n9061), .A2(n5329), .ZN(n5328) );
  INV_X1 U5309 ( .A(n5331), .ZN(n5329) );
  OR2_X1 U5310 ( .A1(n9243), .A2(n9095), .ZN(n8534) );
  NAND2_X1 U5311 ( .A1(n5926), .A2(n5319), .ZN(n5318) );
  NOR2_X1 U5312 ( .A1(n5942), .A2(n5320), .ZN(n5319) );
  INV_X1 U5313 ( .A(n5925), .ZN(n5320) );
  INV_X1 U5314 ( .A(n5504), .ZN(n5500) );
  NAND2_X1 U5315 ( .A1(n6107), .A2(n5542), .ZN(n6160) );
  NAND2_X1 U5316 ( .A1(n5980), .A2(n5979), .ZN(n5993) );
  OAI21_X1 U5317 ( .B1(n7680), .B2(n5153), .A(n5155), .ZN(n8049) );
  NOR2_X1 U5318 ( .A1(n5391), .A2(n5154), .ZN(n5153) );
  NOR2_X1 U5319 ( .A1(n4993), .A2(n5156), .ZN(n5155) );
  NOR2_X1 U5320 ( .A1(n5158), .A2(n7679), .ZN(n5154) );
  NOR2_X1 U5321 ( .A1(n8711), .A2(n8709), .ZN(n5131) );
  INV_X1 U5322 ( .A(n9612), .ZN(n5236) );
  INV_X1 U5323 ( .A(n9613), .ZN(n5232) );
  NOR2_X1 U5324 ( .A1(n9732), .A2(n9736), .ZN(n9719) );
  INV_X1 U5325 ( .A(n5434), .ZN(n5433) );
  OAI21_X1 U5326 ( .B1(n9815), .B2(n5435), .A(n9575), .ZN(n5434) );
  INV_X1 U5327 ( .A(n8307), .ZN(n5435) );
  OR2_X1 U5328 ( .A1(n8331), .A2(n8250), .ZN(n6801) );
  NAND2_X1 U5329 ( .A1(n6848), .A2(n7961), .ZN(n7346) );
  NAND2_X1 U5330 ( .A1(n5454), .A2(n4961), .ZN(n5453) );
  INV_X1 U5331 ( .A(n5031), .ZN(n5454) );
  AND2_X1 U5332 ( .A1(n7774), .A2(n10725), .ZN(n10221) );
  INV_X1 U5333 ( .A(n5495), .ZN(n5494) );
  OAI22_X1 U5334 ( .A1(n5661), .A2(n5496), .B1(n5663), .B2(SI_26_), .ZN(n5495)
         );
  NAND2_X1 U5335 ( .A1(n5488), .A2(n5647), .ZN(n5487) );
  INV_X1 U5336 ( .A(n6026), .ZN(n5488) );
  INV_X1 U5337 ( .A(n5487), .ZN(n5484) );
  OAI21_X1 U5338 ( .B1(n5163), .B2(n9985), .A(n6778), .ZN(n5161) );
  OR2_X1 U5339 ( .A1(n6575), .A2(n9985), .ZN(n5162) );
  INV_X1 U5340 ( .A(n6015), .ZN(n5646) );
  AND2_X1 U5341 ( .A1(n6246), .A2(n6250), .ZN(n5163) );
  INV_X1 U5342 ( .A(n5960), .ZN(n5476) );
  AND2_X1 U5343 ( .A1(n5479), .A2(n5630), .ZN(n5478) );
  NAND2_X1 U5344 ( .A1(n5482), .A2(n5627), .ZN(n5481) );
  NAND2_X1 U5345 ( .A1(n5812), .A2(n5602), .ZN(n5816) );
  XNOR2_X1 U5346 ( .A(n7050), .B(n7585), .ZN(n7042) );
  NAND2_X1 U5347 ( .A1(n5540), .A2(n5538), .ZN(n5537) );
  INV_X1 U5348 ( .A(n7053), .ZN(n5538) );
  INV_X1 U5349 ( .A(n8394), .ZN(n5513) );
  OR3_X1 U5350 ( .A1(n8649), .A2(n7958), .A3(n7127), .ZN(n7178) );
  NAND2_X1 U5351 ( .A1(n7095), .A2(n9107), .ZN(n7096) );
  AND4_X1 U5352 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n8832)
         );
  NOR2_X1 U5353 ( .A1(n7410), .A2(n7409), .ZN(n7408) );
  OR2_X1 U5354 ( .A1(n7406), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U5355 ( .A1(n5103), .A2(n8937), .ZN(n8941) );
  NAND2_X1 U5356 ( .A1(n10481), .A2(n5026), .ZN(n5103) );
  XNOR2_X1 U5357 ( .A(n6909), .B(n10500), .ZN(n10499) );
  NAND2_X1 U5358 ( .A1(n10516), .A2(n10517), .ZN(n10515) );
  XNOR2_X1 U5359 ( .A(n6912), .B(n10530), .ZN(n10532) );
  NAND2_X1 U5360 ( .A1(n10548), .A2(n10549), .ZN(n10547) );
  XNOR2_X1 U5361 ( .A(n6915), .B(n10563), .ZN(n10565) );
  NAND2_X1 U5362 ( .A1(n10582), .A2(n10581), .ZN(n10580) );
  XNOR2_X1 U5363 ( .A(n6918), .B(n10597), .ZN(n10599) );
  NAND2_X1 U5364 ( .A1(n10615), .A2(n10616), .ZN(n10614) );
  NAND2_X1 U5365 ( .A1(n5367), .A2(n5366), .ZN(n5365) );
  AND2_X1 U5366 ( .A1(n5368), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5366) );
  NOR2_X1 U5367 ( .A1(n10597), .A2(n6883), .ZN(n6884) );
  NOR2_X1 U5368 ( .A1(n10607), .A2(n10606), .ZN(n10605) );
  XNOR2_X1 U5369 ( .A(n6887), .B(n6886), .ZN(n10639) );
  XNOR2_X1 U5370 ( .A(n6921), .B(n10629), .ZN(n10631) );
  OR2_X1 U5371 ( .A1(n7138), .A2(n8217), .ZN(n7008) );
  OAI21_X1 U5372 ( .B1(n4931), .B2(n5294), .A(n5293), .ZN(n5292) );
  OR2_X1 U5373 ( .A1(n8965), .A2(n5008), .ZN(n5291) );
  NAND2_X1 U5374 ( .A1(n5309), .A2(n5308), .ZN(n8973) );
  NAND2_X1 U5375 ( .A1(n5005), .A2(n4950), .ZN(n5308) );
  OAI21_X1 U5376 ( .B1(n8222), .B2(n5911), .A(n8220), .ZN(n8235) );
  INV_X1 U5377 ( .A(n8628), .ZN(n5274) );
  NAND2_X1 U5378 ( .A1(n8511), .A2(n8512), .ZN(n8626) );
  NAND2_X1 U5379 ( .A1(n5879), .A2(n5878), .ZN(n8112) );
  NAND2_X1 U5380 ( .A1(n5046), .A2(n8498), .ZN(n8125) );
  NAND2_X1 U5381 ( .A1(n5256), .A2(n5255), .ZN(n6124) );
  OR2_X1 U5382 ( .A1(n5259), .A2(n8622), .ZN(n5255) );
  NAND2_X1 U5383 ( .A1(n7916), .A2(n5257), .ZN(n5256) );
  AOI21_X1 U5384 ( .B1(n8622), .B2(n5260), .A(n5259), .ZN(n5253) );
  OAI21_X1 U5385 ( .B1(n7606), .B2(n5252), .A(n5041), .ZN(n7716) );
  AOI21_X1 U5386 ( .B1(n8479), .B2(n5251), .A(n5250), .ZN(n5041) );
  AND2_X1 U5387 ( .A1(n8490), .A2(n8488), .ZN(n8617) );
  NAND2_X1 U5388 ( .A1(n7716), .A2(n8617), .ZN(n7916) );
  NAND2_X1 U5389 ( .A1(n5165), .A2(n5762), .ZN(n7530) );
  AND2_X1 U5390 ( .A1(n5760), .A2(n5761), .ZN(n5165) );
  OAI21_X1 U5391 ( .B1(n8462), .B2(n7536), .A(n5733), .ZN(n7545) );
  OR2_X1 U5392 ( .A1(n8576), .A2(n6188), .ZN(n7179) );
  NAND2_X1 U5393 ( .A1(n8567), .A2(n5040), .ZN(n5039) );
  INV_X1 U5394 ( .A(n8612), .ZN(n5040) );
  NAND2_X1 U5395 ( .A1(n5311), .A2(n8641), .ZN(n5310) );
  INV_X1 U5396 ( .A(n5314), .ZN(n5311) );
  AOI21_X1 U5397 ( .B1(n6046), .B2(n5316), .A(n5315), .ZN(n5314) );
  INV_X1 U5398 ( .A(n8640), .ZN(n5315) );
  OR2_X1 U5399 ( .A1(n9036), .A2(n5017), .ZN(n6138) );
  INV_X1 U5400 ( .A(n5271), .ZN(n5270) );
  OAI21_X1 U5401 ( .B1(n6137), .B2(n4943), .A(n6140), .ZN(n5271) );
  NAND2_X1 U5402 ( .A1(n6138), .A2(n6137), .ZN(n9042) );
  NAND2_X1 U5403 ( .A1(n9079), .A2(n5332), .ZN(n5330) );
  NAND2_X1 U5404 ( .A1(n5042), .A2(n5261), .ZN(n9036) );
  AOI21_X1 U5405 ( .B1(n5264), .B2(n5266), .A(n5262), .ZN(n5261) );
  NAND2_X1 U5406 ( .A1(n9090), .A2(n5264), .ZN(n5042) );
  INV_X1 U5407 ( .A(n5265), .ZN(n5264) );
  AND2_X1 U5408 ( .A1(n8547), .A2(n9056), .ZN(n9071) );
  AND2_X1 U5409 ( .A1(n8541), .A2(n8537), .ZN(n9078) );
  AND2_X1 U5410 ( .A1(n5964), .A2(n5963), .ZN(n8536) );
  AND4_X1 U5411 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n9094)
         );
  NAND2_X1 U5412 ( .A1(n9091), .A2(n9089), .ZN(n9097) );
  OR2_X1 U5413 ( .A1(n7148), .A2(n8576), .ZN(n9170) );
  INV_X1 U5414 ( .A(n9170), .ZN(n9080) );
  INV_X1 U5415 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U5416 ( .A1(n6107), .A2(n5541), .ZN(n5682) );
  INV_X1 U5417 ( .A(n6967), .ZN(n6962) );
  NAND2_X1 U5418 ( .A1(n5100), .A2(n5099), .ZN(n5789) );
  INV_X1 U5419 ( .A(n5744), .ZN(n5100) );
  NOR2_X1 U5420 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5724) );
  NOR2_X1 U5421 ( .A1(n5397), .A2(n5396), .ZN(n5395) );
  INV_X1 U5422 ( .A(n7730), .ZN(n5396) );
  INV_X1 U5423 ( .A(n5417), .ZN(n5414) );
  NOR2_X1 U5424 ( .A1(n5122), .A2(n5121), .ZN(n5120) );
  NOR2_X1 U5425 ( .A1(n5126), .A2(n5125), .ZN(n5124) );
  NAND2_X1 U5426 ( .A1(n9352), .A2(n5408), .ZN(n5407) );
  INV_X1 U5427 ( .A(n5410), .ZN(n5408) );
  INV_X1 U5428 ( .A(n8257), .ZN(n5426) );
  AOI21_X1 U5429 ( .B1(n8257), .B2(n4952), .A(n5024), .ZN(n5425) );
  INV_X1 U5430 ( .A(n8245), .ZN(n5427) );
  NOR2_X1 U5431 ( .A1(n9400), .A2(n9399), .ZN(n5150) );
  NAND2_X1 U5432 ( .A1(n9400), .A2(n9399), .ZN(n5151) );
  INV_X1 U5433 ( .A(n5150), .ZN(n5147) );
  OR2_X1 U5434 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  OR2_X1 U5435 ( .A1(n6440), .A2(n6439), .ZN(n6452) );
  NAND2_X1 U5436 ( .A1(n8733), .A2(n8732), .ZN(n5144) );
  NAND2_X1 U5437 ( .A1(n7680), .A2(n7679), .ZN(n7729) );
  NAND2_X1 U5438 ( .A1(n8752), .A2(n8751), .ZN(n5421) );
  OAI21_X1 U5439 ( .B1(n8420), .B2(n5380), .A(n5378), .ZN(n5382) );
  INV_X1 U5440 ( .A(n5379), .ZN(n5378) );
  OAI21_X1 U5441 ( .B1(n8419), .B2(n5380), .A(n8692), .ZN(n5379) );
  NAND2_X1 U5442 ( .A1(n8424), .A2(n5381), .ZN(n5380) );
  INV_X1 U5443 ( .A(n7961), .ZN(n7563) );
  NAND2_X1 U5444 ( .A1(n5069), .A2(n10222), .ZN(n5068) );
  NAND2_X1 U5445 ( .A1(n6781), .A2(n4986), .ZN(n5069) );
  NAND2_X1 U5446 ( .A1(n6776), .A2(n9552), .ZN(n5067) );
  AND2_X1 U5447 ( .A1(n7961), .A2(n9552), .ZN(n7548) );
  INV_X1 U5448 ( .A(n6842), .ZN(n6844) );
  AND4_X1 U5449 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n9281)
         );
  AND4_X1 U5450 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n7752)
         );
  NOR2_X1 U5451 ( .A1(n5096), .A2(n4978), .ZN(n7466) );
  NAND2_X1 U5452 ( .A1(n6341), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U5453 ( .A1(n9646), .A2(n9612), .ZN(n9631) );
  NAND2_X1 U5454 ( .A1(n9652), .A2(n9948), .ZN(n9637) );
  AOI21_X1 U5455 ( .B1(n5439), .B2(n5441), .A(n4973), .ZN(n5438) );
  AND2_X1 U5456 ( .A1(n6760), .A2(n9611), .ZN(n9665) );
  INV_X1 U5457 ( .A(n9690), .ZN(n9591) );
  AND4_X1 U5458 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n9702)
         );
  NAND2_X1 U5459 ( .A1(n9714), .A2(n9715), .ZN(n5239) );
  INV_X1 U5460 ( .A(n9586), .ZN(n5452) );
  AND2_X1 U5461 ( .A1(n6706), .A2(n9608), .ZN(n9715) );
  NAND2_X1 U5462 ( .A1(n9719), .A2(n9559), .ZN(n9720) );
  INV_X1 U5463 ( .A(n9719), .ZN(n9733) );
  AND4_X1 U5464 ( .A1(n6278), .A2(n6277), .A3(n6276), .A4(n6275), .ZN(n9729)
         );
  NOR2_X1 U5465 ( .A1(n9787), .A2(n5443), .ZN(n5442) );
  INV_X1 U5466 ( .A(n9579), .ZN(n5443) );
  NAND2_X1 U5467 ( .A1(n9788), .A2(n9558), .ZN(n9789) );
  NAND2_X1 U5468 ( .A1(n8306), .A2(n8305), .ZN(n9814) );
  NAND2_X1 U5469 ( .A1(n8072), .A2(n8071), .ZN(n8074) );
  AND4_X1 U5470 ( .A1(n6422), .A2(n6421), .A3(n6420), .A4(n6419), .ZN(n7800)
         );
  INV_X1 U5471 ( .A(n6736), .ZN(n5223) );
  NAND2_X1 U5472 ( .A1(n7837), .A2(n6791), .ZN(n6737) );
  INV_X1 U5473 ( .A(n7788), .ZN(n5220) );
  AND2_X1 U5474 ( .A1(n9998), .A2(n7569), .ZN(n10227) );
  NOR2_X1 U5475 ( .A1(n7827), .A2(n7834), .ZN(n7830) );
  OR2_X1 U5476 ( .A1(n9819), .A2(n9552), .ZN(n7575) );
  NAND2_X1 U5477 ( .A1(n8028), .A2(n8109), .ZN(n10702) );
  INV_X1 U5478 ( .A(n10225), .ZN(n10704) );
  NAND2_X1 U5479 ( .A1(n6627), .A2(n6626), .ZN(n9879) );
  OR2_X1 U5480 ( .A1(n8447), .A2(n6625), .ZN(n6627) );
  INV_X1 U5481 ( .A(n9984), .ZN(n7694) );
  INV_X1 U5482 ( .A(n10806), .ZN(n10810) );
  NAND2_X1 U5483 ( .A1(n7359), .A2(n8417), .ZN(n9980) );
  INV_X1 U5484 ( .A(n9980), .ZN(n7372) );
  NOR2_X1 U5485 ( .A1(n8448), .A2(n8273), .ZN(n6855) );
  INV_X1 U5486 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U5487 ( .A1(n6222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6223) );
  NOR2_X1 U5488 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6213) );
  NAND2_X1 U5489 ( .A1(n5498), .A2(n5661), .ZN(n6061) );
  NAND2_X1 U5490 ( .A1(n6849), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6851) );
  XNOR2_X1 U5491 ( .A(n6852), .B(P1_IR_REG_24__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U5492 ( .A1(n4960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6852) );
  AND2_X1 U5493 ( .A1(n6300), .A2(n5335), .ZN(n6575) );
  NAND2_X1 U5494 ( .A1(n5928), .A2(n5927), .ZN(n5930) );
  NAND2_X1 U5495 ( .A1(n5846), .A2(n5470), .ZN(n5469) );
  NAND2_X1 U5496 ( .A1(n5466), .A2(n5830), .ZN(n5463) );
  INV_X1 U5497 ( .A(n5461), .ZN(n5460) );
  INV_X1 U5498 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U5499 ( .A1(n5491), .A2(n5593), .ZN(n5807) );
  NAND2_X1 U5500 ( .A1(n7080), .A2(n7079), .ZN(n7081) );
  NAND2_X1 U5501 ( .A1(n5530), .A2(n5529), .ZN(n7069) );
  AOI21_X1 U5502 ( .B1(n5533), .B2(n5531), .A(n7067), .ZN(n5529) );
  AND4_X1 U5503 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n9048)
         );
  NAND2_X1 U5504 ( .A1(n5904), .A2(n5903), .ZN(n8402) );
  NAND2_X1 U5505 ( .A1(n7093), .A2(n7092), .ZN(n10851) );
  AND4_X1 U5506 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n8868)
         );
  AND4_X1 U5507 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n8359)
         );
  AND4_X1 U5508 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n9063)
         );
  NOR2_X1 U5509 ( .A1(n5517), .A2(n8907), .ZN(n5515) );
  AND2_X1 U5510 ( .A1(n5519), .A2(n5015), .ZN(n5517) );
  NAND2_X1 U5511 ( .A1(n5519), .A2(n5522), .ZN(n5518) );
  NAND2_X1 U5512 ( .A1(n8674), .A2(n8671), .ZN(n5522) );
  NAND2_X1 U5513 ( .A1(n7136), .A2(n10829), .ZN(n10853) );
  INV_X1 U5514 ( .A(n5180), .ZN(n5176) );
  OAI21_X1 U5515 ( .B1(n5183), .B2(n4941), .A(n5181), .ZN(n5180) );
  NAND2_X1 U5516 ( .A1(n5183), .A2(n5182), .ZN(n5181) );
  NAND2_X1 U5517 ( .A1(n8646), .A2(n8655), .ZN(n5182) );
  NAND2_X1 U5518 ( .A1(n5002), .A2(n5184), .ZN(n5179) );
  INV_X1 U5519 ( .A(n8878), .ZN(n9026) );
  AND4_X1 U5520 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n9171)
         );
  XNOR2_X1 U5521 ( .A(n5809), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U5522 ( .A1(n10664), .A2(n6924), .ZN(n7022) );
  NAND2_X1 U5523 ( .A1(n7031), .A2(n4979), .ZN(n5115) );
  AND2_X1 U5524 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  AOI21_X1 U5525 ( .B1(n7012), .B2(n10670), .A(n7011), .ZN(n7013) );
  NAND2_X1 U5526 ( .A1(n5371), .A2(n5369), .ZN(n6897) );
  NOR2_X1 U5527 ( .A1(n6895), .A2(n5370), .ZN(n5369) );
  NAND2_X1 U5528 ( .A1(n10673), .A2(n5372), .ZN(n5371) );
  NOR2_X1 U5529 ( .A1(n7018), .A2(n9085), .ZN(n5370) );
  NAND2_X1 U5530 ( .A1(n7255), .A2(n6962), .ZN(n10677) );
  AOI21_X1 U5531 ( .B1(n6119), .B2(n9103), .A(n6118), .ZN(n8786) );
  NAND2_X1 U5532 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  NAND2_X1 U5533 ( .A1(n5248), .A2(n8612), .ZN(n8977) );
  NAND2_X1 U5534 ( .A1(n6039), .A2(n6038), .ZN(n9016) );
  NAND2_X1 U5535 ( .A1(n7171), .A2(n8156), .ZN(n7173) );
  INV_X1 U5536 ( .A(n8803), .ZN(n8782) );
  INV_X1 U5537 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U5538 ( .A1(n5135), .A2(n5133), .ZN(n5377) );
  AOI21_X1 U5539 ( .B1(n5136), .B2(n5138), .A(n5134), .ZN(n5133) );
  NAND2_X1 U5540 ( .A1(n8736), .A2(n9361), .ZN(n5142) );
  NAND2_X1 U5541 ( .A1(n8733), .A2(n4975), .ZN(n5139) );
  NAND2_X1 U5542 ( .A1(n6551), .A2(n6550), .ZN(n9930) );
  INV_X1 U5543 ( .A(n7752), .ZN(n9423) );
  INV_X1 U5544 ( .A(n7466), .ZN(n9426) );
  XNOR2_X1 U5545 ( .A(n9571), .B(n9561), .ZN(n9563) );
  NAND2_X1 U5546 ( .A1(n9626), .A2(n9596), .ZN(n9598) );
  NAND2_X1 U5547 ( .A1(n9638), .A2(n9595), .ZN(n9596) );
  AND2_X2 U5548 ( .A1(n7580), .A2(n9984), .ZN(n10819) );
  NAND2_X1 U5549 ( .A1(n8467), .A2(n8486), .ZN(n8470) );
  AOI21_X1 U5550 ( .B1(n5078), .B2(n4933), .A(n5077), .ZN(n5076) );
  INV_X1 U5551 ( .A(n7794), .ZN(n5078) );
  NOR2_X1 U5552 ( .A1(n6738), .A2(n4933), .ZN(n5077) );
  OR2_X1 U5553 ( .A1(n6400), .A2(n6399), .ZN(n5075) );
  INV_X1 U5554 ( .A(n5080), .ZN(n5079) );
  OAI22_X1 U5555 ( .A1(n6460), .A2(n4933), .B1(n5222), .B2(n7553), .ZN(n5080)
         );
  NAND2_X1 U5556 ( .A1(n5074), .A2(n5076), .ZN(n6463) );
  OR2_X1 U5557 ( .A1(n5081), .A2(n5079), .ZN(n5074) );
  NAND2_X1 U5558 ( .A1(n5073), .A2(n5071), .ZN(n6446) );
  AOI21_X1 U5559 ( .B1(n4948), .B2(n5079), .A(n5072), .ZN(n5071) );
  NAND2_X1 U5560 ( .A1(n5081), .A2(n4948), .ZN(n5073) );
  NAND2_X1 U5561 ( .A1(n7858), .A2(n7789), .ZN(n5072) );
  AND2_X1 U5562 ( .A1(n8497), .A2(n8620), .ZN(n5213) );
  NAND2_X1 U5563 ( .A1(n5175), .A2(n5174), .ZN(n5173) );
  NAND2_X1 U5564 ( .A1(n5172), .A2(n8590), .ZN(n5171) );
  NOR2_X1 U5565 ( .A1(n8514), .A2(n8590), .ZN(n5174) );
  NAND2_X1 U5566 ( .A1(n6560), .A2(n7553), .ZN(n5082) );
  NAND2_X1 U5567 ( .A1(n5245), .A2(n4933), .ZN(n5083) );
  NAND2_X1 U5568 ( .A1(n5004), .A2(n5088), .ZN(n5087) );
  NAND2_X1 U5569 ( .A1(n6561), .A2(n7553), .ZN(n5088) );
  NAND2_X1 U5570 ( .A1(n8543), .A2(n5195), .ZN(n5194) );
  NOR2_X1 U5571 ( .A1(n5197), .A2(n5196), .ZN(n5195) );
  INV_X1 U5572 ( .A(n8542), .ZN(n5196) );
  INV_X1 U5573 ( .A(n8535), .ZN(n5197) );
  NAND2_X1 U5574 ( .A1(n5169), .A2(n5166), .ZN(n8529) );
  NOR2_X1 U5575 ( .A1(n5168), .A2(n5167), .ZN(n5166) );
  NAND2_X1 U5576 ( .A1(n5170), .A2(n8521), .ZN(n5169) );
  INV_X1 U5577 ( .A(n8524), .ZN(n5167) );
  OAI21_X1 U5578 ( .B1(n5188), .B2(n5187), .A(n5186), .ZN(n5185) );
  NAND2_X1 U5579 ( .A1(n8537), .A2(n8536), .ZN(n5187) );
  NOR3_X1 U5580 ( .A1(n4951), .A2(n8576), .A3(n5262), .ZN(n5186) );
  INV_X1 U5581 ( .A(n5194), .ZN(n5188) );
  NOR2_X1 U5582 ( .A1(n5192), .A2(n5262), .ZN(n5191) );
  AOI21_X1 U5583 ( .B1(n5194), .B2(n9107), .A(n5193), .ZN(n5192) );
  INV_X1 U5584 ( .A(n8537), .ZN(n5193) );
  NAND2_X1 U5585 ( .A1(n5190), .A2(n8576), .ZN(n5189) );
  NAND2_X1 U5586 ( .A1(n8540), .A2(n9078), .ZN(n5190) );
  INV_X1 U5587 ( .A(n8557), .ZN(n5206) );
  NAND2_X1 U5588 ( .A1(n5205), .A2(n9049), .ZN(n5204) );
  AOI21_X1 U5589 ( .B1(n6609), .B2(n5092), .A(n9751), .ZN(n5091) );
  AND2_X1 U5590 ( .A1(n6823), .A2(n7553), .ZN(n5092) );
  NAND2_X1 U5591 ( .A1(n6605), .A2(n5094), .ZN(n5093) );
  NOR2_X1 U5592 ( .A1(n7553), .A2(n5095), .ZN(n5094) );
  INV_X1 U5593 ( .A(n9743), .ZN(n5095) );
  NAND2_X1 U5594 ( .A1(n8614), .A2(n5201), .ZN(n5200) );
  INV_X1 U5595 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5064) );
  INV_X1 U5596 ( .A(n5296), .ZN(n5295) );
  AND2_X1 U5597 ( .A1(n7161), .A2(n5299), .ZN(n5298) );
  NAND2_X1 U5598 ( .A1(n5300), .A2(n5561), .ZN(n5299) );
  INV_X1 U5599 ( .A(n5302), .ZN(n5300) );
  NAND2_X1 U5600 ( .A1(n5875), .A2(n5872), .ZN(n5874) );
  INV_X1 U5601 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U5602 ( .A1(n5401), .A2(n5029), .ZN(n5158) );
  AND2_X1 U5603 ( .A1(n5391), .A2(n5157), .ZN(n5156) );
  INV_X1 U5604 ( .A(n7679), .ZN(n5157) );
  OR2_X1 U5605 ( .A1(n8043), .A2(n5402), .ZN(n5400) );
  OR3_X1 U5606 ( .A1(n5393), .A2(n7750), .A3(n5397), .ZN(n5390) );
  NOR2_X1 U5607 ( .A1(n5393), .A2(n5392), .ZN(n5391) );
  INV_X1 U5608 ( .A(n5395), .ZN(n5392) );
  NAND2_X1 U5609 ( .A1(n5497), .A2(n5662), .ZN(n5496) );
  INV_X1 U5610 ( .A(n6070), .ZN(n5497) );
  INV_X1 U5611 ( .A(n5496), .ZN(n5493) );
  INV_X1 U5612 ( .A(n5702), .ZN(n5480) );
  INV_X1 U5613 ( .A(SI_16_), .ZN(n10143) );
  INV_X1 U5614 ( .A(SI_9_), .ZN(n10047) );
  INV_X1 U5615 ( .A(SI_8_), .ZN(n10040) );
  INV_X1 U5616 ( .A(n7062), .ZN(n5528) );
  AND2_X1 U5617 ( .A1(n5112), .A2(n5114), .ZN(n6907) );
  NAND2_X1 U5618 ( .A1(n10524), .A2(n6874), .ZN(n5353) );
  INV_X1 U5619 ( .A(n10623), .ZN(n5368) );
  AND2_X1 U5620 ( .A1(n5364), .A2(n6885), .ZN(n5363) );
  NAND2_X1 U5621 ( .A1(n4931), .A2(n5296), .ZN(n5293) );
  NOR2_X1 U5622 ( .A1(n5295), .A2(n5298), .ZN(n5294) );
  INV_X1 U5623 ( .A(n8572), .ZN(n5038) );
  NAND2_X1 U5624 ( .A1(n5303), .A2(n8976), .ZN(n5302) );
  OR2_X1 U5625 ( .A1(n5303), .A2(n8976), .ZN(n5561) );
  NOR2_X1 U5626 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n6052), .ZN(n6051) );
  INV_X1 U5627 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10179) );
  NOR2_X1 U5628 ( .A1(n5259), .A2(n5260), .ZN(n5257) );
  OR2_X1 U5629 ( .A1(n6165), .A2(n6179), .ZN(n7129) );
  AOI21_X1 U5630 ( .B1(n5328), .B2(n5326), .A(n9043), .ZN(n5325) );
  INV_X1 U5631 ( .A(n5332), .ZN(n5326) );
  INV_X1 U5632 ( .A(n6133), .ZN(n5266) );
  OAI21_X1 U5633 ( .B1(n9092), .B2(n5266), .A(n9078), .ZN(n5265) );
  AND2_X1 U5634 ( .A1(n8534), .A2(n8538), .ZN(n8633) );
  INV_X1 U5635 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6415) );
  INV_X1 U5636 ( .A(n5129), .ZN(n5121) );
  INV_X1 U5637 ( .A(n8701), .ZN(n5122) );
  NOR2_X1 U5638 ( .A1(n5409), .A2(n9279), .ZN(n5405) );
  INV_X1 U5639 ( .A(n9352), .ZN(n5409) );
  OR2_X1 U5640 ( .A1(n5552), .A2(n8714), .ZN(n5126) );
  OAI21_X1 U5641 ( .B1(n5066), .B2(n5065), .A(n6682), .ZN(n6683) );
  NAND2_X1 U5642 ( .A1(n9630), .A2(n6678), .ZN(n5065) );
  NAND2_X1 U5643 ( .A1(n5089), .A2(n5098), .ZN(n5097) );
  INV_X1 U5644 ( .A(n7831), .ZN(n5098) );
  INV_X1 U5645 ( .A(n5440), .ZN(n5439) );
  OAI21_X1 U5646 ( .B1(n9590), .B2(n5441), .A(n9594), .ZN(n5440) );
  INV_X1 U5647 ( .A(n9593), .ZN(n5441) );
  NOR2_X1 U5648 ( .A1(n9682), .A2(n9672), .ZN(n9652) );
  INV_X1 U5649 ( .A(n9806), .ZN(n5244) );
  INV_X1 U5650 ( .A(n5341), .ZN(n5340) );
  AND2_X1 U5651 ( .A1(n7889), .A2(n10793), .ZN(n7975) );
  OR2_X1 U5652 ( .A1(n5223), .A2(n5222), .ZN(n5221) );
  NOR2_X1 U5653 ( .A1(n7850), .A2(n9841), .ZN(n5343) );
  NAND2_X1 U5654 ( .A1(n5545), .A2(n9581), .ZN(n9762) );
  NOR2_X1 U5655 ( .A1(n7987), .A2(n8142), .ZN(n7889) );
  NOR2_X1 U5656 ( .A1(n5215), .A2(n5214), .ZN(n5337) );
  INV_X1 U5657 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6212) );
  NOR2_X1 U5658 ( .A1(n6211), .A2(n9985), .ZN(n6210) );
  INV_X1 U5659 ( .A(SI_27_), .ZN(n10122) );
  INV_X1 U5660 ( .A(SI_28_), .ZN(n10017) );
  INV_X1 U5661 ( .A(SI_24_), .ZN(n10012) );
  NAND2_X1 U5662 ( .A1(n5387), .A2(n5386), .ZN(n5385) );
  INV_X1 U5663 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5386) );
  INV_X1 U5664 ( .A(SI_23_), .ZN(n10132) );
  INV_X1 U5665 ( .A(SI_20_), .ZN(n10116) );
  INV_X1 U5666 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6246) );
  INV_X1 U5667 ( .A(SI_15_), .ZN(n10147) );
  INV_X1 U5668 ( .A(n5830), .ZN(n5462) );
  INV_X1 U5669 ( .A(SI_10_), .ZN(n10043) );
  INV_X1 U5670 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6447) );
  INV_X1 U5671 ( .A(n5603), .ZN(n5467) );
  INV_X1 U5672 ( .A(n5591), .ZN(n5055) );
  OAI21_X1 U5673 ( .B1(n7195), .B2(n5580), .A(n5579), .ZN(n5581) );
  NAND2_X1 U5674 ( .A1(n5458), .A2(n5457), .ZN(n5570) );
  AND2_X1 U5675 ( .A1(n5567), .A2(SI_1_), .ZN(n5457) );
  OR2_X1 U5676 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  NAND2_X1 U5677 ( .A1(n8096), .A2(n5534), .ZN(n5533) );
  INV_X1 U5678 ( .A(n7064), .ZN(n5534) );
  INV_X1 U5679 ( .A(n7063), .ZN(n5532) );
  NAND2_X1 U5680 ( .A1(n7503), .A2(n7055), .ZN(n7619) );
  NOR2_X1 U5681 ( .A1(n5905), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5919) );
  OR2_X1 U5682 ( .A1(n5850), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5889) );
  INV_X1 U5683 ( .A(n7056), .ZN(n5539) );
  OR2_X1 U5684 ( .A1(n5800), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U5685 ( .A1(n5051), .A2(n4976), .ZN(n5049) );
  AND4_X1 U5686 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n7252)
         );
  NAND2_X1 U5687 ( .A1(n5348), .A2(n6865), .ZN(n7330) );
  NAND2_X1 U5688 ( .A1(n6864), .A2(n5349), .ZN(n5348) );
  NAND2_X1 U5689 ( .A1(n5350), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U5690 ( .A(n6906), .B(n5359), .ZN(n7395) );
  OAI211_X1 U5691 ( .C1(n5111), .C2(P2_REG1_REG_3__SCAN_IN), .A(n5110), .B(
        n5109), .ZN(n5112) );
  INV_X1 U5692 ( .A(n7413), .ZN(n5110) );
  NAND2_X1 U5693 ( .A1(n5106), .A2(n5104), .ZN(n5109) );
  OR2_X1 U5694 ( .A1(n5359), .A2(n6906), .ZN(n5106) );
  AND2_X1 U5695 ( .A1(n7396), .A2(n4968), .ZN(n7410) );
  AND2_X1 U5696 ( .A1(n5108), .A2(n5107), .ZN(n7412) );
  INV_X1 U5697 ( .A(n5111), .ZN(n5107) );
  NAND2_X1 U5698 ( .A1(n7395), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5108) );
  NOR2_X1 U5699 ( .A1(n5352), .A2(n7207), .ZN(n5351) );
  NOR2_X1 U5700 ( .A1(n5808), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U5701 ( .A1(n10498), .A2(n6910), .ZN(n10516) );
  INV_X1 U5702 ( .A(n10524), .ZN(n5355) );
  NAND2_X1 U5703 ( .A1(n10531), .A2(n6913), .ZN(n10548) );
  NOR2_X1 U5704 ( .A1(n5744), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U5705 ( .A1(n10564), .A2(n6916), .ZN(n10582) );
  NAND2_X1 U5706 ( .A1(n5501), .A2(n5287), .ZN(n5706) );
  NAND2_X1 U5707 ( .A1(n10598), .A2(n6919), .ZN(n10615) );
  NAND2_X1 U5708 ( .A1(n10630), .A2(n6922), .ZN(n10647) );
  NAND2_X1 U5709 ( .A1(n10647), .A2(n10648), .ZN(n10646) );
  XNOR2_X1 U5710 ( .A(n6923), .B(n10663), .ZN(n10665) );
  OAI21_X1 U5711 ( .B1(n7635), .B2(n6892), .A(n7018), .ZN(n10675) );
  NAND2_X1 U5712 ( .A1(n10646), .A2(n5101), .ZN(n6923) );
  NAND2_X1 U5713 ( .A1(n7512), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5101) );
  INV_X1 U5714 ( .A(n7020), .ZN(n5372) );
  OR2_X1 U5715 ( .A1(n6075), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6077) );
  OR2_X1 U5716 ( .A1(n6040), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U5717 ( .A1(n5689), .A2(n10179), .ZN(n6007) );
  INV_X1 U5718 ( .A(n5997), .ZN(n5689) );
  AND2_X1 U5719 ( .A1(n5966), .A2(n5965), .ZN(n5984) );
  INV_X1 U5720 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10081) );
  AND2_X1 U5721 ( .A1(n5953), .A2(n10081), .ZN(n5966) );
  NAND2_X1 U5722 ( .A1(n8409), .A2(n5321), .ZN(n9105) );
  NAND2_X1 U5723 ( .A1(n8413), .A2(n5322), .ZN(n5321) );
  INV_X1 U5724 ( .A(n9171), .ZN(n5322) );
  NAND2_X1 U5725 ( .A1(n9105), .A2(n9113), .ZN(n9104) );
  OR2_X1 U5726 ( .A1(n5934), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5936) );
  NOR2_X1 U5727 ( .A1(n5936), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5953) );
  OR3_X1 U5728 ( .A1(n7629), .A2(n4941), .A3(n6148), .ZN(n7529) );
  AOI21_X1 U5729 ( .B1(n8234), .B2(n8629), .A(n6129), .ZN(n9164) );
  NAND2_X1 U5730 ( .A1(n5304), .A2(n5305), .ZN(n8222) );
  INV_X1 U5731 ( .A(n5306), .ZN(n5305) );
  NAND2_X1 U5732 ( .A1(n5879), .A2(n4946), .ZN(n5304) );
  OAI21_X1 U5733 ( .B1(n5881), .B2(n5307), .A(n5896), .ZN(n5306) );
  NAND2_X1 U5734 ( .A1(n5867), .A2(n5837), .ZN(n5850) );
  NOR2_X1 U5735 ( .A1(n5821), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5865) );
  INV_X1 U5736 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10187) );
  AND2_X1 U5737 ( .A1(n8491), .A2(n8498), .ZN(n8621) );
  INV_X1 U5738 ( .A(n7669), .ZN(n7610) );
  NAND2_X1 U5739 ( .A1(n5764), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5736) );
  AND2_X1 U5740 ( .A1(n8486), .A2(n8483), .ZN(n8618) );
  AND3_X1 U5741 ( .A1(n5752), .A2(n5753), .A3(n5164), .ZN(n7605) );
  NAND2_X1 U5742 ( .A1(n5764), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5752) );
  NOR2_X1 U5743 ( .A1(n4953), .A2(n4984), .ZN(n5164) );
  NOR2_X1 U5744 ( .A1(n7252), .A2(n7432), .ZN(n7536) );
  INV_X1 U5745 ( .A(n6120), .ZN(n8462) );
  NAND2_X1 U5746 ( .A1(n7252), .A2(n7631), .ZN(n7044) );
  NAND2_X1 U5747 ( .A1(n6083), .A2(n5553), .ZN(n8965) );
  OR2_X1 U5748 ( .A1(n9192), .A2(n8832), .ZN(n5553) );
  OR2_X1 U5749 ( .A1(n8678), .A2(n8988), .ZN(n6082) );
  OR2_X1 U5750 ( .A1(n9053), .A2(n9025), .ZN(n9024) );
  NAND2_X1 U5751 ( .A1(n5324), .A2(n5323), .ZN(n9022) );
  AOI21_X1 U5752 ( .B1(n5325), .B2(n5327), .A(n8637), .ZN(n5323) );
  NAND2_X1 U5753 ( .A1(n9079), .A2(n5325), .ZN(n5324) );
  INV_X1 U5754 ( .A(n5328), .ZN(n5327) );
  AND4_X1 U5755 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n9095)
         );
  NAND2_X1 U5756 ( .A1(n9104), .A2(n5556), .ZN(n9091) );
  OR2_X1 U5757 ( .A1(n8846), .A2(n9095), .ZN(n5556) );
  INV_X1 U5758 ( .A(n8633), .ZN(n9113) );
  NAND2_X1 U5759 ( .A1(n5318), .A2(n5941), .ZN(n8407) );
  OAI22_X1 U5760 ( .A1(n7184), .A2(n7183), .B1(n7182), .B2(n7181), .ZN(n7188)
         );
  INV_X1 U5761 ( .A(n7631), .ZN(n7432) );
  OR2_X1 U5762 ( .A1(n8649), .A2(n8659), .ZN(n8344) );
  AND2_X1 U5763 ( .A1(n5500), .A2(n5284), .ZN(n5283) );
  AND2_X1 U5764 ( .A1(n5670), .A2(n5285), .ZN(n5284) );
  NAND2_X1 U5765 ( .A1(n6152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U5766 ( .A1(n6154), .A2(n6153), .ZN(n6157) );
  OR2_X1 U5767 ( .A1(n5789), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5808) );
  INV_X1 U5768 ( .A(n8419), .ZN(n5134) );
  NOR2_X1 U5769 ( .A1(n8736), .A2(n9361), .ZN(n5143) );
  INV_X1 U5770 ( .A(n8732), .ZN(n5140) );
  NAND2_X1 U5771 ( .A1(n8246), .A2(n8245), .ZN(n8321) );
  INV_X1 U5772 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U5773 ( .A1(n8047), .A2(n8046), .ZN(n8050) );
  INV_X1 U5774 ( .A(n8049), .ZN(n8047) );
  INV_X1 U5775 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6515) );
  OR2_X1 U5776 ( .A1(n6554), .A2(n6553), .ZN(n6568) );
  AND2_X1 U5777 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6401) );
  AND2_X1 U5778 ( .A1(n5118), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7347) );
  INV_X1 U5779 ( .A(n6588), .ZN(n6598) );
  NAND2_X1 U5780 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n6598), .ZN(n6597) );
  NAND2_X1 U5781 ( .A1(n8718), .A2(n8717), .ZN(n5410) );
  NAND2_X1 U5782 ( .A1(n9377), .A2(n9380), .ZN(n8715) );
  INV_X1 U5783 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6504) );
  INV_X1 U5784 ( .A(n5423), .ZN(n5138) );
  AOI21_X1 U5785 ( .B1(n5423), .B2(n5137), .A(n5020), .ZN(n5136) );
  INV_X1 U5786 ( .A(n5425), .ZN(n5137) );
  NOR2_X1 U5787 ( .A1(n6568), .A2(n6567), .ZN(n6581) );
  NAND2_X1 U5788 ( .A1(n5127), .A2(n5126), .ZN(n9377) );
  NAND2_X1 U5789 ( .A1(n8702), .A2(n4949), .ZN(n5127) );
  NAND2_X1 U5790 ( .A1(n5128), .A2(n5131), .ZN(n9378) );
  AOI21_X1 U5791 ( .B1(n8109), .B2(n7548), .A(n5118), .ZN(n5117) );
  OR2_X1 U5792 ( .A1(n6599), .A2(n9392), .ZN(n6648) );
  NAND2_X1 U5793 ( .A1(n6669), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6334) );
  NOR2_X1 U5794 ( .A1(n5027), .A2(n4934), .ZN(n9430) );
  NAND2_X1 U5795 ( .A1(n9597), .A2(n5231), .ZN(n5230) );
  NAND2_X1 U5796 ( .A1(n5227), .A2(n5226), .ZN(n5225) );
  NAND2_X1 U5797 ( .A1(n9695), .A2(n9685), .ZN(n9682) );
  INV_X1 U5798 ( .A(n9652), .ZN(n9669) );
  INV_X1 U5799 ( .A(n5448), .ZN(n5447) );
  NAND2_X1 U5800 ( .A1(n9767), .A2(n6823), .ZN(n9744) );
  AND2_X1 U5801 ( .A1(n6823), .A2(n9743), .ZN(n9766) );
  AOI21_X1 U5802 ( .B1(n5433), .B2(n5435), .A(n4965), .ZN(n5431) );
  NAND2_X1 U5803 ( .A1(n8309), .A2(n8308), .ZN(n9805) );
  NAND2_X1 U5804 ( .A1(n9826), .A2(n6749), .ZN(n8309) );
  AND4_X1 U5805 ( .A1(n6559), .A2(n6558), .A3(n6557), .A4(n6556), .ZN(n9403)
         );
  OR2_X1 U5806 ( .A1(n6518), .A2(n6504), .ZN(n6506) );
  NAND2_X1 U5807 ( .A1(n8018), .A2(n5339), .ZN(n8208) );
  NOR2_X1 U5808 ( .A1(n8076), .A2(n5456), .ZN(n5455) );
  INV_X1 U5809 ( .A(n8073), .ZN(n5456) );
  NAND2_X1 U5810 ( .A1(n8018), .A2(n10803), .ZN(n8080) );
  AND2_X1 U5811 ( .A1(n6745), .A2(n6804), .ZN(n7967) );
  AND4_X1 U5812 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n8250)
         );
  AND2_X1 U5813 ( .A1(n6475), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6485) );
  AND4_X1 U5814 ( .A1(n6458), .A2(n6457), .A3(n6456), .A4(n6455), .ZN(n8138)
         );
  NAND2_X1 U5815 ( .A1(n7887), .A2(n7886), .ZN(n7963) );
  NAND2_X1 U5816 ( .A1(n5343), .A2(n5342), .ZN(n7987) );
  NAND2_X1 U5817 ( .A1(n7985), .A2(n7984), .ZN(n7983) );
  AND4_X1 U5818 ( .A1(n6445), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(n8151)
         );
  INV_X1 U5819 ( .A(n5343), .ZN(n7986) );
  OAI21_X1 U5820 ( .B1(n7787), .B2(n7788), .A(n7786), .ZN(n7849) );
  NAND2_X1 U5821 ( .A1(n7849), .A2(n7848), .ZN(n7847) );
  NAND2_X1 U5822 ( .A1(n10221), .A2(n10735), .ZN(n10220) );
  OR2_X1 U5823 ( .A1(n10220), .A2(n7820), .ZN(n7827) );
  INV_X1 U5824 ( .A(n6363), .ZN(n7767) );
  OR2_X1 U5825 ( .A1(n7346), .A2(n9552), .ZN(n7763) );
  NAND2_X1 U5826 ( .A1(n6658), .A2(n6657), .ZN(n9654) );
  NAND2_X1 U5827 ( .A1(n5453), .A2(n5451), .ZN(n9709) );
  INV_X1 U5828 ( .A(n10814), .ZN(n9931) );
  OR2_X1 U5829 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  NOR2_X1 U5830 ( .A1(n7693), .A2(n7577), .ZN(n7580) );
  AND2_X1 U5831 ( .A1(n6856), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7572) );
  AND2_X1 U5832 ( .A1(n6212), .A2(n6211), .ZN(n6224) );
  INV_X1 U5833 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6225) );
  XNOR2_X1 U5834 ( .A(n6253), .B(n6201), .ZN(n9262) );
  NAND2_X1 U5835 ( .A1(n6061), .A2(n5662), .ZN(n6071) );
  INV_X1 U5836 ( .A(n5486), .ZN(n5485) );
  OAI21_X1 U5837 ( .B1(n5646), .B2(n5487), .A(n5651), .ZN(n5486) );
  NAND2_X1 U5838 ( .A1(n6013), .A2(n5647), .ZN(n6027) );
  NAND2_X1 U5839 ( .A1(n6703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U5840 ( .A1(n5162), .A2(n5160), .ZN(n6703) );
  INV_X1 U5841 ( .A(n5161), .ZN(n5160) );
  INV_X1 U5842 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6778) );
  AOI21_X1 U5843 ( .B1(n5477), .B2(n5475), .A(n5474), .ZN(n5972) );
  NOR2_X1 U5844 ( .A1(n5481), .A2(n5476), .ZN(n5475) );
  OAI21_X1 U5845 ( .B1(n5478), .B2(n5476), .A(n5021), .ZN(n5474) );
  OAI21_X1 U5846 ( .B1(n5703), .B2(n5481), .A(n5478), .ZN(n5959) );
  AND2_X1 U5847 ( .A1(n5623), .A2(n5622), .ZN(n5927) );
  AND2_X1 U5848 ( .A1(n5618), .A2(n5617), .ZN(n5912) );
  NAND2_X1 U5849 ( .A1(n5816), .A2(n5603), .ZN(n5858) );
  AND2_X1 U5850 ( .A1(n5388), .A2(n5387), .ZN(n6300) );
  INV_X1 U5851 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5217) );
  NOR2_X2 U5852 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5436) );
  NAND2_X1 U5853 ( .A1(n5723), .A2(n5570), .ZN(n5739) );
  NAND2_X1 U5854 ( .A1(n5933), .A2(n5932), .ZN(n10827) );
  AND4_X1 U5855 ( .A1(n8600), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n8801)
         );
  OR2_X1 U5856 ( .A1(n8790), .A2(n8976), .ZN(n8791) );
  AND4_X1 U5857 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8400)
         );
  OR2_X1 U5858 ( .A1(n7087), .A2(n9171), .ZN(n7088) );
  NAND2_X1 U5859 ( .A1(n5537), .A2(n5536), .ZN(n7621) );
  AND4_X1 U5860 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n8133)
         );
  OAI21_X1 U5861 ( .B1(n7999), .B2(n7064), .A(n7063), .ZN(n8097) );
  INV_X1 U5862 ( .A(n8898), .ZN(n10847) );
  NAND2_X1 U5863 ( .A1(n8821), .A2(n7102), .ZN(n8856) );
  INV_X1 U5864 ( .A(n5510), .ZN(n5509) );
  NAND2_X1 U5865 ( .A1(n5508), .A2(n5512), .ZN(n8865) );
  NAND2_X1 U5866 ( .A1(n8354), .A2(n4947), .ZN(n5508) );
  AND2_X1 U5867 ( .A1(n7106), .A2(n9064), .ZN(n7107) );
  NOR2_X1 U5868 ( .A1(n7475), .A2(n7047), .ZN(n7481) );
  NAND2_X1 U5869 ( .A1(n10851), .A2(n7096), .ZN(n8883) );
  AND2_X1 U5870 ( .A1(n5535), .A2(n5536), .ZN(n8894) );
  INV_X1 U5871 ( .A(n10845), .ZN(n8914) );
  NAND2_X1 U5872 ( .A1(n7145), .A2(n7144), .ZN(n10856) );
  NAND2_X1 U5873 ( .A1(n8807), .A2(n7085), .ZN(n8909) );
  NOR2_X1 U5874 ( .A1(n8661), .A2(n8655), .ZN(n5178) );
  INV_X1 U5875 ( .A(n8133), .ZN(n8000) );
  INV_X1 U5876 ( .A(n7605), .ZN(n8932) );
  NAND2_X1 U5877 ( .A1(n5764), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U5878 ( .A1(n4968), .A2(n5358), .ZN(n7398) );
  OR2_X1 U5879 ( .A1(n10506), .A2(n6873), .ZN(n5356) );
  NAND2_X1 U5880 ( .A1(n5365), .A2(n5364), .ZN(n10622) );
  NOR2_X1 U5881 ( .A1(n6889), .A2(n10637), .ZN(n10655) );
  NAND2_X1 U5882 ( .A1(n7007), .A2(n7006), .ZN(n10662) );
  NAND2_X1 U5883 ( .A1(n6006), .A2(n6005), .ZN(n9141) );
  NAND2_X1 U5884 ( .A1(n5926), .A2(n5925), .ZN(n9166) );
  NAND2_X1 U5885 ( .A1(n8112), .A2(n5881), .ZN(n8184) );
  NAND2_X1 U5886 ( .A1(n5272), .A2(n5275), .ZN(n8187) );
  NAND2_X1 U5887 ( .A1(n5044), .A2(n5273), .ZN(n8186) );
  NAND2_X1 U5888 ( .A1(n8125), .A2(n5278), .ZN(n5272) );
  NAND2_X1 U5889 ( .A1(n5282), .A2(n5281), .ZN(n5280) );
  INV_X1 U5890 ( .A(n8125), .ZN(n5282) );
  OAI21_X1 U5891 ( .B1(n7916), .B2(n5254), .A(n5253), .ZN(n7932) );
  OR2_X1 U5892 ( .A1(n7628), .A2(n10831), .ZN(n8981) );
  AND2_X1 U5893 ( .A1(n5811), .A2(n5810), .ZN(n8036) );
  NAND2_X1 U5894 ( .A1(n5258), .A2(n8622), .ZN(n7918) );
  NAND2_X1 U5895 ( .A1(n7916), .A2(n8490), .ZN(n5258) );
  OR2_X1 U5896 ( .A1(n7135), .A2(n7661), .ZN(n10829) );
  AND2_X1 U5897 ( .A1(n10837), .A2(n10835), .ZN(n9115) );
  INV_X1 U5898 ( .A(n8981), .ZN(n9112) );
  INV_X1 U5899 ( .A(n10829), .ZN(n9111) );
  NAND2_X1 U5900 ( .A1(n5036), .A2(n4944), .ZN(n8963) );
  OR2_X1 U5901 ( .A1(n5248), .A2(n8568), .ZN(n5036) );
  INV_X1 U5902 ( .A(n8678), .ZN(n9192) );
  OR2_X1 U5903 ( .A1(n8447), .A2(n5741), .ZN(n6063) );
  NAND2_X1 U5904 ( .A1(n5312), .A2(n5310), .ZN(n8986) );
  NAND2_X1 U5905 ( .A1(n9010), .A2(n4942), .ZN(n5312) );
  NAND2_X1 U5906 ( .A1(n5313), .A2(n5316), .ZN(n8998) );
  OAI21_X1 U5907 ( .B1(n6138), .B2(n4943), .A(n5270), .ZN(n9008) );
  NAND2_X1 U5908 ( .A1(n9042), .A2(n6139), .ZN(n9020) );
  NAND2_X1 U5909 ( .A1(n5330), .A2(n5331), .ZN(n9060) );
  NAND2_X1 U5910 ( .A1(n5996), .A2(n5995), .ZN(n9226) );
  AOI21_X1 U5911 ( .B1(n9079), .B2(n5990), .A(n5334), .ZN(n9070) );
  NAND2_X1 U5912 ( .A1(n5983), .A2(n5982), .ZN(n9232) );
  OR2_X1 U5913 ( .A1(n7666), .A2(n5741), .ZN(n5983) );
  NAND2_X1 U5914 ( .A1(n5263), .A2(n6133), .ZN(n9077) );
  NAND2_X1 U5915 ( .A1(n9090), .A2(n9092), .ZN(n5263) );
  INV_X1 U5916 ( .A(n8536), .ZN(n10852) );
  NAND2_X1 U5917 ( .A1(n5952), .A2(n5951), .ZN(n9243) );
  INV_X1 U5918 ( .A(n10843), .ZN(n10840) );
  NAND2_X1 U5919 ( .A1(n5726), .A2(n5499), .ZN(n5727) );
  NOR2_X1 U5920 ( .A1(n7196), .A2(n7195), .ZN(n5499) );
  AND2_X1 U5921 ( .A1(n6168), .A2(n6167), .ZN(n9256) );
  NAND2_X1 U5922 ( .A1(n7138), .A2(n6183), .ZN(n9255) );
  XNOR2_X1 U5923 ( .A(n6181), .B(n6182), .ZN(n7239) );
  INV_X1 U5924 ( .A(n6166), .ZN(n8437) );
  AND2_X1 U5925 ( .A1(n5679), .A2(P2_U3151), .ZN(n9267) );
  INV_X1 U5926 ( .A(n10546), .ZN(n7247) );
  INV_X1 U5927 ( .A(n10514), .ZN(n7225) );
  INV_X1 U5928 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7209) );
  XNOR2_X1 U5929 ( .A(n5776), .B(n5775), .ZN(n7406) );
  INV_X1 U5930 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U5931 ( .A1(n5744), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5758) );
  OAI21_X1 U5932 ( .B1(n5743), .B2(n5667), .A(n5742), .ZN(n5745) );
  NAND2_X1 U5933 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5667), .ZN(n5742) );
  INV_X1 U5934 ( .A(n6864), .ZN(n7334) );
  NAND2_X1 U5935 ( .A1(n5398), .A2(n5394), .ZN(n8042) );
  NAND2_X1 U5936 ( .A1(n7729), .A2(n5395), .ZN(n5394) );
  OAI21_X1 U5937 ( .B1(n7728), .B2(n5399), .A(n5029), .ZN(n5398) );
  NAND2_X1 U5938 ( .A1(n8715), .A2(n9378), .ZN(n9278) );
  NAND2_X1 U5939 ( .A1(n6586), .A2(n6585), .ZN(n9791) );
  NAND2_X1 U5940 ( .A1(n8774), .A2(n5420), .ZN(n5415) );
  NAND2_X1 U5941 ( .A1(n5414), .A2(n8774), .ZN(n5413) );
  NAND2_X1 U5942 ( .A1(n8050), .A2(n8143), .ZN(n8053) );
  AND2_X1 U5943 ( .A1(n5407), .A2(n8726), .ZN(n5406) );
  OR2_X1 U5944 ( .A1(n8026), .A2(n6625), .ZN(n6290) );
  NAND2_X1 U5945 ( .A1(n8694), .A2(n5149), .ZN(n5148) );
  NOR2_X1 U5946 ( .A1(n5150), .A2(n5381), .ZN(n5149) );
  OR2_X1 U5947 ( .A1(n6670), .A2(n9463), .ZN(n6369) );
  OAI22_X1 U5948 ( .A1(n6393), .A2(n7203), .B1(n6357), .B2(n9489), .ZN(n6394)
         );
  NAND2_X1 U5949 ( .A1(n6357), .A2(n10002), .ZN(n6347) );
  NAND2_X1 U5950 ( .A1(n5376), .A2(n10302), .ZN(n5375) );
  NAND2_X1 U5951 ( .A1(n5141), .A2(n8736), .ZN(n9359) );
  INV_X1 U5952 ( .A(n5144), .ZN(n5141) );
  OAI22_X1 U5953 ( .A1(n9961), .A2(n7350), .B1(n9717), .B2(n7349), .ZN(n9361)
         );
  NAND2_X1 U5954 ( .A1(n7729), .A2(n7730), .ZN(n5403) );
  AND4_X1 U5955 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n9666)
         );
  NAND2_X1 U5956 ( .A1(n7444), .A2(n8195), .ZN(n9395) );
  NAND2_X1 U5957 ( .A1(n5152), .A2(n5382), .ZN(n9402) );
  NAND2_X1 U5958 ( .A1(n8694), .A2(n8693), .ZN(n5152) );
  INV_X1 U5959 ( .A(n9398), .ZN(n9411) );
  INV_X1 U5960 ( .A(n9395), .ZN(n9409) );
  XNOR2_X1 U5961 ( .A(n6249), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7564) );
  OAI21_X1 U5962 ( .B1(n6702), .B2(n6248), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6249) );
  INV_X1 U5963 ( .A(n6782), .ZN(n6783) );
  NAND2_X1 U5964 ( .A1(n5068), .A2(n5067), .ZN(n6784) );
  NAND2_X1 U5965 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  INV_X1 U5966 ( .A(n9729), .ZN(n9587) );
  INV_X1 U5967 ( .A(n9769), .ZN(n9809) );
  NAND2_X1 U5968 ( .A1(n5089), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6343) );
  INV_X1 U5969 ( .A(n10470), .ZN(n10685) );
  NAND2_X1 U5970 ( .A1(n6668), .A2(n6667), .ZN(n9638) );
  NAND2_X1 U5971 ( .A1(n9688), .A2(n9593), .ZN(n9662) );
  NAND2_X1 U5972 ( .A1(n5239), .A2(n9608), .ZN(n9701) );
  NAND2_X1 U5973 ( .A1(n5445), .A2(n5448), .ZN(n9693) );
  NAND2_X1 U5974 ( .A1(n5031), .A2(n5451), .ZN(n5445) );
  AND2_X1 U5975 ( .A1(n9721), .A2(n9720), .ZN(n9891) );
  NAND2_X1 U5976 ( .A1(n6596), .A2(n6595), .ZN(n9906) );
  NAND2_X1 U5977 ( .A1(n5444), .A2(n9579), .ZN(n9786) );
  NAND2_X1 U5978 ( .A1(n9814), .A2(n9815), .ZN(n5432) );
  NAND2_X1 U5979 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  CLKBUF_X1 U5980 ( .A(n8169), .Z(n8077) );
  OAI211_X1 U5981 ( .C1(n6737), .C2(n5220), .A(n6738), .B(n5219), .ZN(n7844)
         );
  NAND2_X1 U5982 ( .A1(n5223), .A2(n7788), .ZN(n5219) );
  NAND2_X1 U5983 ( .A1(n6787), .A2(n7788), .ZN(n7567) );
  INV_X1 U5984 ( .A(n9835), .ZN(n9842) );
  INV_X1 U5985 ( .A(n9844), .ZN(n9739) );
  INV_X1 U5986 ( .A(n4932), .ZN(n10235) );
  INV_X1 U5987 ( .A(n9557), .ZN(n9940) );
  NAND2_X1 U5988 ( .A1(n9859), .A2(n4966), .ZN(n5247) );
  INV_X1 U5989 ( .A(n9654), .ZN(n9948) );
  INV_X1 U5990 ( .A(n9672), .ZN(n9952) );
  INV_X1 U5991 ( .A(n9736), .ZN(n9961) );
  INV_X1 U5992 ( .A(n9791), .ZN(n9558) );
  AND2_X1 U5993 ( .A1(n7363), .A2(n7362), .ZN(n9984) );
  NAND2_X1 U5994 ( .A1(n7383), .A2(n7572), .ZN(n9983) );
  XNOR2_X1 U5995 ( .A(n6196), .B(n6195), .ZN(n9996) );
  XNOR2_X1 U5996 ( .A(n6854), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8417) );
  INV_X1 U5997 ( .A(n7357), .ZN(n8273) );
  INV_X1 U5998 ( .A(n7564), .ZN(n8109) );
  XNOR2_X1 U5999 ( .A(n6779), .B(n6778), .ZN(n7961) );
  NAND2_X1 U6000 ( .A1(n6702), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6779) );
  AND2_X1 U6001 ( .A1(n6317), .A2(n6316), .ZN(n10364) );
  NAND2_X1 U6002 ( .A1(n5469), .A2(n5472), .ZN(n5898) );
  NAND2_X1 U6003 ( .A1(n5459), .A2(n5844), .ZN(n5845) );
  AND2_X1 U6004 ( .A1(n6481), .A2(n6473), .ZN(n10476) );
  INV_X1 U6005 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U6006 ( .A1(n5518), .A2(n10854), .ZN(n5516) );
  NAND2_X1 U6007 ( .A1(n5176), .A2(n5184), .ZN(n5053) );
  AOI21_X1 U6008 ( .B1(n5116), .B2(n10671), .A(n5115), .ZN(n7034) );
  XNOR2_X1 U6009 ( .A(n7022), .B(n7023), .ZN(n5116) );
  OAI21_X1 U6010 ( .B1(n7014), .B2(n8939), .A(n7013), .ZN(n7015) );
  NAND2_X1 U6011 ( .A1(n7186), .A2(n8349), .ZN(n7177) );
  NAND2_X1 U6012 ( .A1(n8686), .A2(n8349), .ZN(n6194) );
  OAI21_X1 U6013 ( .B1(n8782), .B2(n9158), .A(n6191), .ZN(n6192) );
  AOI21_X1 U6014 ( .B1(n8454), .B2(n7191), .A(n7190), .ZN(n7192) );
  OAI21_X1 U6015 ( .B1(n9935), .B2(n10820), .A(n5345), .ZN(P1_U3521) );
  INV_X1 U6016 ( .A(n5346), .ZN(n5345) );
  OR2_X1 U6017 ( .A1(n10823), .A2(n9936), .ZN(n5347) );
  OAI21_X1 U6018 ( .B1(n9942), .B2(n10820), .A(n5056), .ZN(P1_U3518) );
  INV_X1 U6019 ( .A(n5057), .ZN(n5056) );
  OAI22_X1 U6020 ( .A1(n9944), .A2(n9977), .B1(n10823), .B2(n9943), .ZN(n5057)
         );
  NAND2_X1 U6021 ( .A1(n8467), .A2(n8464), .ZN(n6121) );
  AND2_X1 U6022 ( .A1(n8641), .A2(n5316), .ZN(n4942) );
  INV_X1 U6023 ( .A(n8693), .ZN(n5381) );
  NAND2_X1 U6024 ( .A1(n6347), .A2(n5375), .ZN(n7554) );
  INV_X1 U6025 ( .A(n7040), .ZN(n7041) );
  NAND2_X1 U6026 ( .A1(n4996), .A2(n6139), .ZN(n4943) );
  AND2_X1 U6027 ( .A1(n8566), .A2(n5039), .ZN(n4944) );
  INV_X1 U6028 ( .A(n9163), .ZN(n5168) );
  AND2_X1 U6029 ( .A1(n5389), .A2(n7354), .ZN(n4945) );
  AND2_X1 U6030 ( .A1(n5878), .A2(n5895), .ZN(n4946) );
  AND2_X1 U6031 ( .A1(n5023), .A2(n7075), .ZN(n4947) );
  AND2_X1 U6032 ( .A1(n5076), .A2(n6795), .ZN(n4948) );
  AND2_X1 U6033 ( .A1(n5132), .A2(n8701), .ZN(n4949) );
  NAND2_X1 U6034 ( .A1(n7530), .A2(n7605), .ZN(n8486) );
  NAND2_X2 U6035 ( .A1(n9565), .A2(n9440), .ZN(n6357) );
  INV_X1 U6036 ( .A(n5029), .ZN(n5397) );
  OR2_X1 U6037 ( .A1(n9195), .A2(n8999), .ZN(n4950) );
  NOR3_X1 U6038 ( .A1(n8635), .A2(n9107), .A3(n8534), .ZN(n4951) );
  OR2_X1 U6039 ( .A1(n5427), .A2(n8258), .ZN(n4952) );
  AND2_X1 U6040 ( .A1(n5713), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U6041 ( .A1(n7049), .A2(n7517), .ZN(n4954) );
  INV_X1 U6042 ( .A(n5401), .ZN(n5393) );
  NAND2_X1 U6043 ( .A1(n8043), .A2(n5402), .ZN(n5401) );
  AND2_X1 U6044 ( .A1(n4949), .A2(n9380), .ZN(n4955) );
  AND2_X1 U6045 ( .A1(n5339), .A2(n5338), .ZN(n4956) );
  AND2_X1 U6046 ( .A1(n5540), .A2(n7055), .ZN(n4957) );
  AND2_X1 U6047 ( .A1(n7086), .A2(n7085), .ZN(n4958) );
  AND2_X1 U6048 ( .A1(n7097), .A2(n7096), .ZN(n4959) );
  AND2_X1 U6049 ( .A1(n5403), .A2(n5159), .ZN(n7751) );
  INV_X1 U6050 ( .A(n5356), .ZN(n10523) );
  AND2_X1 U6051 ( .A1(n5961), .A2(n5950), .ZN(n10645) );
  INV_X1 U6052 ( .A(n8661), .ZN(n5184) );
  AND2_X1 U6053 ( .A1(n5691), .A2(n5688), .ZN(n5734) );
  AND3_X1 U6054 ( .A1(n5287), .A2(n5501), .A3(n5286), .ZN(n6107) );
  NAND3_X1 U6055 ( .A1(n5335), .A2(n5388), .A3(n5384), .ZN(n4960) );
  AND2_X1 U6056 ( .A1(n6679), .A2(n6833), .ZN(n9614) );
  INV_X1 U6057 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U6058 ( .A1(n5139), .A2(n5142), .ZN(n9272) );
  XNOR2_X1 U6059 ( .A(n6704), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6848) );
  XNOR2_X1 U6060 ( .A(n6106), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6149) );
  OR2_X1 U6061 ( .A1(n9736), .A2(n9747), .ZN(n4961) );
  NAND2_X1 U6062 ( .A1(n9919), .A2(n9781), .ZN(n4962) );
  INV_X1 U6063 ( .A(n5276), .ZN(n5275) );
  OAI21_X1 U6064 ( .B1(n5281), .B2(n5277), .A(n8512), .ZN(n5276) );
  INV_X1 U6065 ( .A(n9614), .ZN(n9597) );
  OR2_X1 U6066 ( .A1(n8562), .A2(n8639), .ZN(n4963) );
  INV_X1 U6067 ( .A(n5459), .ZN(n5843) );
  OAI21_X1 U6068 ( .B1(n5812), .B2(n5463), .A(n5460), .ZN(n5459) );
  NAND2_X1 U6069 ( .A1(n6575), .A2(n6246), .ZN(n4964) );
  NAND2_X1 U6070 ( .A1(n5411), .A2(n5410), .ZN(n9351) );
  INV_X1 U6071 ( .A(n7206), .ZN(n5359) );
  OAI21_X1 U6072 ( .B1(n5992), .B2(n5991), .A(n5640), .ZN(n6003) );
  NAND2_X1 U6073 ( .A1(n5492), .A2(n5494), .ZN(n6085) );
  NAND2_X1 U6074 ( .A1(n5483), .A2(n5485), .ZN(n6036) );
  INV_X1 U6075 ( .A(n6749), .ZN(n5245) );
  AND2_X1 U6076 ( .A1(n9577), .A2(n9830), .ZN(n4965) );
  AOI21_X1 U6077 ( .B1(n5275), .B2(n5277), .A(n5274), .ZN(n5273) );
  INV_X1 U6078 ( .A(n5273), .ZN(n5043) );
  NAND4_X1 U6079 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n7040)
         );
  OR2_X1 U6080 ( .A1(n9860), .A2(n10814), .ZN(n4966) );
  NAND2_X1 U6081 ( .A1(n6855), .A2(n8417), .ZN(n7383) );
  INV_X1 U6082 ( .A(n7383), .ZN(n5118) );
  AND2_X1 U6083 ( .A1(n5330), .A2(n5328), .ZN(n4967) );
  XNOR2_X1 U6084 ( .A(n5687), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5688) );
  OAI21_X1 U6085 ( .B1(n9272), .B2(n5419), .A(n5417), .ZN(n9389) );
  OR2_X1 U6086 ( .A1(n6868), .A2(n5359), .ZN(n4968) );
  OR2_X1 U6087 ( .A1(n6151), .A2(n5676), .ZN(n4969) );
  AND2_X1 U6088 ( .A1(n7406), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6089 ( .A1(n5144), .A2(n8735), .ZN(n9358) );
  XNOR2_X1 U6090 ( .A(n9598), .B(n9597), .ZN(n9861) );
  INV_X1 U6091 ( .A(n7899), .ZN(n7930) );
  AND3_X1 U6092 ( .A1(n5286), .A2(n5501), .A3(n5283), .ZN(n4971) );
  AND2_X1 U6093 ( .A1(n8490), .A2(n8484), .ZN(n4972) );
  AND4_X1 U6094 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n8976)
         );
  INV_X1 U6095 ( .A(n5451), .ZN(n5450) );
  NOR2_X1 U6096 ( .A1(n9715), .A2(n5452), .ZN(n5451) );
  INV_X1 U6097 ( .A(n5512), .ZN(n5511) );
  NAND2_X1 U6098 ( .A1(n5023), .A2(n5513), .ZN(n5512) );
  INV_X1 U6099 ( .A(n5388), .ZN(n6423) );
  AND2_X1 U6100 ( .A1(n9672), .A2(n9680), .ZN(n4973) );
  AND4_X1 U6101 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n7915)
         );
  NOR2_X1 U6102 ( .A1(n10605), .A2(n6884), .ZN(n4974) );
  INV_X1 U6103 ( .A(n9279), .ZN(n5412) );
  INV_X1 U6104 ( .A(n7717), .ZN(n8930) );
  AND4_X1 U6105 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n7717)
         );
  NOR2_X1 U6106 ( .A1(n5143), .A2(n5140), .ZN(n4975) );
  AND2_X1 U6107 ( .A1(n8610), .A2(n5050), .ZN(n4976) );
  AND2_X1 U6108 ( .A1(n5453), .A2(n9586), .ZN(n4977) );
  NAND2_X1 U6109 ( .A1(n6319), .A2(n6318), .ZN(n8433) );
  NOR2_X1 U6110 ( .A1(n6670), .A2(n6383), .ZN(n4978) );
  AND2_X1 U6111 ( .A1(n7033), .A2(n8886), .ZN(n4979) );
  AND2_X1 U6112 ( .A1(n6708), .A2(n6815), .ZN(n4980) );
  NOR2_X1 U6113 ( .A1(n10655), .A2(n10654), .ZN(n4981) );
  AND2_X1 U6114 ( .A1(n9885), .A2(n9679), .ZN(n4982) );
  AND2_X1 U6115 ( .A1(n9178), .A2(n8586), .ZN(n4983) );
  AND2_X1 U6116 ( .A1(n5734), .A2(n10178), .ZN(n4984) );
  AND2_X1 U6117 ( .A1(n6809), .A2(n6805), .ZN(n8076) );
  INV_X1 U6118 ( .A(n7750), .ZN(n5399) );
  INV_X1 U6119 ( .A(n5420), .ZN(n5419) );
  AND2_X1 U6120 ( .A1(n5421), .A2(n9314), .ZN(n5420) );
  INV_X1 U6121 ( .A(n5473), .ZN(n5472) );
  NOR2_X1 U6122 ( .A1(n5792), .A2(n5793), .ZN(n4985) );
  AND2_X1 U6123 ( .A1(n6732), .A2(n5551), .ZN(n4986) );
  AND2_X1 U6124 ( .A1(n6755), .A2(n9610), .ZN(n9689) );
  AND2_X1 U6125 ( .A1(n6707), .A2(n6821), .ZN(n9787) );
  INV_X1 U6126 ( .A(n5895), .ZN(n5307) );
  OR2_X1 U6127 ( .A1(n9232), .A2(n9094), .ZN(n8541) );
  INV_X1 U6128 ( .A(n8541), .ZN(n5262) );
  NOR2_X1 U6129 ( .A1(n8831), .A2(n5521), .ZN(n4987) );
  NOR2_X1 U6130 ( .A1(n9889), .A2(n9587), .ZN(n4988) );
  AND2_X1 U6131 ( .A1(n8488), .A2(n8487), .ZN(n4989) );
  OR2_X1 U6132 ( .A1(n9426), .A2(n7834), .ZN(n4990) );
  OR2_X1 U6133 ( .A1(n7042), .A2(n7041), .ZN(n4991) );
  NAND2_X1 U6134 ( .A1(n9195), .A2(n8999), .ZN(n4992) );
  INV_X1 U6135 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U6136 ( .A1(n5390), .A2(n5400), .ZN(n4993) );
  NAND2_X1 U6137 ( .A1(n8554), .A2(n5203), .ZN(n4994) );
  OR2_X1 U6138 ( .A1(n5726), .A2(n6864), .ZN(n4995) );
  AND2_X1 U6139 ( .A1(n6761), .A2(n9612), .ZN(n9648) );
  INV_X1 U6140 ( .A(n9648), .ZN(n5235) );
  OR2_X1 U6141 ( .A1(n9033), .A2(n9049), .ZN(n4996) );
  OR2_X1 U6142 ( .A1(n5606), .A2(SI_9_), .ZN(n4997) );
  INV_X1 U6143 ( .A(n5466), .ZN(n5465) );
  NOR2_X1 U6144 ( .A1(n5857), .A2(n5467), .ZN(n5466) );
  AND2_X1 U6145 ( .A1(n5605), .A2(n10040), .ZN(n4998) );
  AND2_X1 U6146 ( .A1(n7066), .A2(n8005), .ZN(n4999) );
  NAND2_X1 U6147 ( .A1(n5416), .A2(n5420), .ZN(n9312) );
  NAND2_X1 U6148 ( .A1(n5405), .A2(n9331), .ZN(n5000) );
  NOR2_X1 U6149 ( .A1(n8829), .A2(n9063), .ZN(n5001) );
  AND2_X1 U6150 ( .A1(n5183), .A2(n8655), .ZN(n5002) );
  INV_X1 U6151 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5350) );
  AND2_X1 U6152 ( .A1(n8803), .A2(n4937), .ZN(n5003) );
  NAND2_X1 U6153 ( .A1(n6811), .A2(n4933), .ZN(n5004) );
  NAND2_X1 U6154 ( .A1(n9591), .A2(n9590), .ZN(n9688) );
  INV_X1 U6155 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U6156 ( .A1(n5310), .A2(n4992), .ZN(n5005) );
  AND3_X1 U6157 ( .A1(n5673), .A2(n5981), .A3(n6100), .ZN(n5006) );
  AND2_X1 U6158 ( .A1(n4931), .A2(n5298), .ZN(n5007) );
  OR2_X1 U6159 ( .A1(n4931), .A2(n5295), .ZN(n5008) );
  INV_X1 U6160 ( .A(n5552), .ZN(n5132) );
  NAND2_X1 U6161 ( .A1(n5489), .A2(n5646), .ZN(n6013) );
  NAND2_X1 U6162 ( .A1(n8221), .A2(n8220), .ZN(n5009) );
  AND2_X1 U6163 ( .A1(n7103), .A2(n7102), .ZN(n5010) );
  AND2_X1 U6164 ( .A1(n9614), .A2(n5233), .ZN(n5011) );
  AOI21_X1 U6165 ( .B1(n5000), .B2(n5129), .A(n5124), .ZN(n5123) );
  AND2_X1 U6166 ( .A1(n8631), .A2(n5941), .ZN(n5012) );
  AND2_X1 U6167 ( .A1(n4950), .A2(n4942), .ZN(n5013) );
  INV_X1 U6168 ( .A(n8751), .ZN(n5422) );
  AND2_X1 U6169 ( .A1(n8750), .A2(n9343), .ZN(n8751) );
  OR2_X1 U6170 ( .A1(n5120), .A2(n4955), .ZN(n5014) );
  NAND2_X1 U6171 ( .A1(n5523), .A2(n8831), .ZN(n5015) );
  INV_X1 U6172 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5387) );
  OR2_X1 U6173 ( .A1(n5539), .A2(n8895), .ZN(n5016) );
  OR2_X1 U6174 ( .A1(n9037), .A2(n6135), .ZN(n5017) );
  INV_X1 U6175 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6176 ( .A1(n7159), .A2(n7158), .ZN(n8454) );
  INV_X1 U6177 ( .A(n8041), .ZN(n5402) );
  NAND2_X1 U6178 ( .A1(n5706), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5980) );
  INV_X1 U6179 ( .A(n8735), .ZN(n8736) );
  INV_X1 U6180 ( .A(n8060), .ZN(n5342) );
  NAND2_X1 U6181 ( .A1(n6737), .A2(n6736), .ZN(n6787) );
  OR2_X1 U6182 ( .A1(n8536), .A2(n9107), .ZN(n5018) );
  OR2_X1 U6183 ( .A1(n7912), .A2(n5828), .ZN(n7924) );
  INV_X1 U6184 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6301) );
  INV_X1 U6185 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5572) );
  OAI21_X1 U6186 ( .B1(n8246), .B2(n5138), .A(n5136), .ZN(n8420) );
  NAND2_X1 U6187 ( .A1(n5280), .A2(n8509), .ZN(n8110) );
  NAND2_X1 U6188 ( .A1(n5377), .A2(n8424), .ZN(n8694) );
  NAND2_X1 U6189 ( .A1(n5432), .A2(n8307), .ZN(n9576) );
  NAND2_X1 U6190 ( .A1(n8354), .A2(n7075), .ZN(n8393) );
  NAND2_X1 U6191 ( .A1(n8702), .A2(n8701), .ZN(n9330) );
  INV_X1 U6192 ( .A(n9380), .ZN(n5125) );
  INV_X1 U6193 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5285) );
  OR3_X1 U6194 ( .A1(n5504), .A2(n5668), .A3(n5744), .ZN(n5019) );
  CLKBUF_X3 U6195 ( .A(n6367), .Z(n6599) );
  INV_X1 U6196 ( .A(n6367), .ZN(n5089) );
  NAND2_X1 U6197 ( .A1(n5503), .A2(n5502), .ZN(n5884) );
  NAND2_X1 U6198 ( .A1(n5335), .A2(n5383), .ZN(n6839) );
  NOR2_X1 U6199 ( .A1(n9799), .A2(n9919), .ZN(n9788) );
  INV_X1 U6200 ( .A(n5344), .ZN(n9799) );
  NOR2_X1 U6201 ( .A1(n9817), .A2(n9577), .ZN(n5344) );
  INV_X1 U6202 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5216) );
  AND2_X1 U6203 ( .A1(n6708), .A2(n6750), .ZN(n9804) );
  INV_X1 U6204 ( .A(n9804), .ZN(n5242) );
  NOR2_X1 U6205 ( .A1(n8368), .A2(n8367), .ZN(n5020) );
  OR2_X1 U6206 ( .A1(n5631), .A2(SI_17_), .ZN(n5021) );
  NOR2_X1 U6207 ( .A1(n7073), .A2(n7072), .ZN(n8354) );
  INV_X1 U6208 ( .A(n8674), .ZN(n5523) );
  AND2_X1 U6209 ( .A1(n7525), .A2(n6190), .ZN(n8349) );
  INV_X1 U6210 ( .A(n8907), .ZN(n10854) );
  NAND2_X1 U6211 ( .A1(n6029), .A2(n6028), .ZN(n9033) );
  INV_X1 U6212 ( .A(n9033), .ZN(n5205) );
  NAND2_X1 U6213 ( .A1(n8018), .A2(n5341), .ZN(n5022) );
  INV_X1 U6214 ( .A(n9390), .ZN(n9414) );
  AND2_X1 U6215 ( .A1(n7377), .A2(n7375), .ZN(n9390) );
  OR2_X1 U6216 ( .A1(n6149), .A2(n8655), .ZN(n7661) );
  INV_X1 U6217 ( .A(n8625), .ZN(n5281) );
  OR2_X1 U6218 ( .A1(n7077), .A2(n8926), .ZN(n5023) );
  AND2_X1 U6219 ( .A1(n8260), .A2(n8259), .ZN(n5024) );
  AND2_X1 U6220 ( .A1(n8495), .A2(n8496), .ZN(n8622) );
  INV_X1 U6221 ( .A(n8622), .ZN(n5254) );
  INV_X1 U6222 ( .A(n5278), .ZN(n5277) );
  NOR2_X1 U6223 ( .A1(n6126), .A2(n5279), .ZN(n5278) );
  INV_X1 U6224 ( .A(n6738), .ZN(n5222) );
  AND2_X1 U6225 ( .A1(n5356), .A2(n5355), .ZN(n5025) );
  INV_X1 U6226 ( .A(n5159), .ZN(n7728) );
  OR2_X1 U6227 ( .A1(n7680), .A2(n7679), .ZN(n5159) );
  INV_X1 U6228 ( .A(n5557), .ZN(n5362) );
  AND2_X2 U6229 ( .A1(n7580), .A2(n7694), .ZN(n10823) );
  INV_X1 U6230 ( .A(n8939), .ZN(n10671) );
  INV_X1 U6231 ( .A(n10230), .ZN(n10716) );
  NAND2_X1 U6232 ( .A1(n7566), .A2(n7565), .ZN(n10230) );
  NAND2_X1 U6233 ( .A1(n5429), .A2(n7561), .ZN(n7826) );
  OR2_X1 U6234 ( .A1(n6907), .A2(n10483), .ZN(n5026) );
  NOR2_X1 U6235 ( .A1(n7568), .A2(n7222), .ZN(n5027) );
  NOR2_X1 U6236 ( .A1(n7481), .A2(n7482), .ZN(n5028) );
  NAND2_X1 U6237 ( .A1(n7736), .A2(n7737), .ZN(n5029) );
  XNOR2_X1 U6238 ( .A(n6251), .B(n6250), .ZN(n9552) );
  INV_X1 U6239 ( .A(n9552), .ZN(n10222) );
  INV_X1 U6240 ( .A(n6147), .ZN(n8655) );
  NAND2_X1 U6241 ( .A1(n5033), .A2(n5032), .ZN(n9941) );
  NAND2_X1 U6242 ( .A1(n9585), .A2(n9584), .ZN(n9726) );
  OAI22_X1 U6243 ( .A1(n9645), .A2(n9648), .B1(n9654), .B2(n9633), .ZN(n9624)
         );
  AND2_X1 U6244 ( .A1(n7053), .A2(n7052), .ZN(n7594) );
  NAND2_X1 U6245 ( .A1(n5030), .A2(n7717), .ZN(n7053) );
  INV_X1 U6246 ( .A(n7051), .ZN(n5030) );
  AOI21_X2 U6247 ( .B1(n8662), .B2(n8663), .A(n7107), .ZN(n8874) );
  NAND2_X1 U6248 ( .A1(n4957), .A2(n7503), .ZN(n5536) );
  NOR2_X1 U6249 ( .A1(n8284), .A2(n7070), .ZN(n7073) );
  NAND2_X2 U6250 ( .A1(n7039), .A2(n7038), .ZN(n7050) );
  NAND2_X2 U6251 ( .A1(n9663), .A2(n9611), .ZN(n9647) );
  NAND2_X1 U6252 ( .A1(n5560), .A2(n9689), .ZN(n9678) );
  NAND2_X1 U6253 ( .A1(n9780), .A2(n9787), .ZN(n9779) );
  AOI21_X1 U6254 ( .B1(n9864), .B2(n10806), .A(n9863), .ZN(n5058) );
  INV_X1 U6255 ( .A(n9862), .ZN(n5059) );
  NAND2_X2 U6256 ( .A1(n6155), .A2(n6157), .ZN(n8335) );
  NAND2_X1 U6257 ( .A1(n8821), .A2(n5010), .ZN(n8854) );
  NAND2_X1 U6258 ( .A1(n5428), .A2(n7562), .ZN(n7787) );
  NAND2_X2 U6259 ( .A1(n6219), .A2(n6218), .ZN(n9565) );
  NAND2_X1 U6260 ( .A1(n5035), .A2(n5037), .ZN(n6145) );
  NAND2_X1 U6261 ( .A1(n5248), .A2(n4944), .ZN(n5035) );
  NOR2_X2 U6262 ( .A1(n5744), .A2(n5668), .ZN(n5501) );
  NAND2_X1 U6263 ( .A1(n7526), .A2(n8618), .ZN(n7606) );
  NAND2_X1 U6264 ( .A1(n5046), .A2(n5047), .ZN(n5044) );
  NOR2_X4 U6265 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6902) );
  AND2_X2 U6266 ( .A1(n5049), .A2(n8654), .ZN(n5183) );
  NAND4_X1 U6267 ( .A1(n5053), .A2(n8660), .A3(n5177), .A4(n5052), .ZN(
        P2_U3296) );
  OR2_X2 U6268 ( .A1(n5179), .A2(n8611), .ZN(n5052) );
  NAND2_X2 U6269 ( .A1(n5726), .A2(n7195), .ZN(n5774) );
  NAND2_X2 U6270 ( .A1(n9779), .A2(n6821), .ZN(n9767) );
  AND2_X2 U6271 ( .A1(n9704), .A2(n9609), .ZN(n5560) );
  NAND2_X1 U6272 ( .A1(n5773), .A2(n5591), .ZN(n5796) );
  NAND2_X1 U6273 ( .A1(n5773), .A2(n5054), .ZN(n5491) );
  AND2_X2 U6274 ( .A1(n5059), .A2(n5058), .ZN(n9942) );
  OAI21_X2 U6275 ( .B1(n7248), .B2(n6625), .A(n6474), .ZN(n8331) );
  INV_X2 U6276 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5060) );
  NAND3_X1 U6277 ( .A1(n7656), .A2(n5064), .A3(n5063), .ZN(n5062) );
  NAND2_X1 U6278 ( .A1(n6398), .A2(n5075), .ZN(n5081) );
  NAND2_X1 U6279 ( .A1(n5089), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6352) );
  NAND2_X2 U6280 ( .A1(n5034), .A2(n9991), .ZN(n6367) );
  AOI21_X1 U6281 ( .B1(n5093), .B2(n5091), .A(n5090), .ZN(n6623) );
  NAND2_X1 U6282 ( .A1(n7834), .A2(n7466), .ZN(n6736) );
  NAND3_X1 U6283 ( .A1(n6385), .A2(n6384), .A3(n5097), .ZN(n5096) );
  INV_X1 U6284 ( .A(n5112), .ZN(n7411) );
  NAND2_X1 U6285 ( .A1(n5114), .A2(n5113), .ZN(n7413) );
  NAND2_X1 U6286 ( .A1(n5119), .A2(n5123), .ZN(n5404) );
  NAND2_X1 U6287 ( .A1(n8702), .A2(n5014), .ZN(n5119) );
  NAND2_X1 U6288 ( .A1(n9330), .A2(n9331), .ZN(n5128) );
  NAND2_X1 U6289 ( .A1(n8246), .A2(n5136), .ZN(n5135) );
  NAND2_X1 U6290 ( .A1(n5145), .A2(n5147), .ZN(n5146) );
  NAND2_X1 U6291 ( .A1(n5382), .A2(n5151), .ZN(n5145) );
  NAND2_X1 U6292 ( .A1(n5148), .A2(n5146), .ZN(n9322) );
  NAND2_X1 U6293 ( .A1(n6575), .A2(n5163), .ZN(n6702) );
  AND4_X2 U6294 ( .A1(n6336), .A2(n6386), .A3(n6202), .A4(n5436), .ZN(n5388)
         );
  NAND2_X2 U6295 ( .A1(n6902), .A2(n5667), .ZN(n5744) );
  INV_X1 U6296 ( .A(n7530), .ZN(n7709) );
  NAND3_X1 U6297 ( .A1(n5173), .A2(n5171), .A3(n5009), .ZN(n5170) );
  NAND3_X1 U6298 ( .A1(n8611), .A2(n8610), .A3(n5178), .ZN(n5177) );
  AOI22_X1 U6299 ( .A1(n8555), .A2(n5202), .B1(n5200), .B2(n5199), .ZN(n5198)
         );
  INV_X1 U6300 ( .A(n5198), .ZN(n8561) );
  NAND4_X1 U6301 ( .A1(n8507), .A2(n5213), .A3(n5211), .A4(n5209), .ZN(n8510)
         );
  NAND4_X1 U6302 ( .A1(n5210), .A2(n8590), .A3(n8490), .A4(n8495), .ZN(n5209)
         );
  NAND4_X1 U6303 ( .A1(n5212), .A2(n8488), .A3(n8496), .A4(n8576), .ZN(n5211)
         );
  NAND3_X1 U6304 ( .A1(n6204), .A2(n5374), .A3(n5373), .ZN(n5214) );
  NAND2_X1 U6305 ( .A1(n6203), .A2(n6547), .ZN(n5215) );
  AND4_X2 U6306 ( .A1(n5384), .A2(n5336), .A3(n5388), .A4(n5337), .ZN(n6227)
         );
  NOR2_X2 U6307 ( .A1(n6206), .A2(n5385), .ZN(n5384) );
  NAND3_X1 U6308 ( .A1(n6205), .A2(n6247), .A3(n6250), .ZN(n6206) );
  INV_X1 U6309 ( .A(n6737), .ZN(n5218) );
  OAI22_X1 U6310 ( .A1(n5221), .A2(n5218), .B1(n5222), .B2(n7788), .ZN(n6739)
         );
  NAND2_X1 U6311 ( .A1(n9647), .A2(n9648), .ZN(n9646) );
  OAI211_X1 U6312 ( .C1(n9647), .C2(n5230), .A(n5225), .B(n5224), .ZN(n9615)
         );
  NAND2_X1 U6313 ( .A1(n9647), .A2(n5011), .ZN(n5224) );
  NAND2_X1 U6314 ( .A1(n9826), .A2(n5243), .ZN(n5240) );
  NAND2_X1 U6315 ( .A1(n5240), .A2(n5241), .ZN(n9807) );
  NAND2_X1 U6316 ( .A1(n8993), .A2(n8613), .ZN(n5248) );
  NAND2_X1 U6317 ( .A1(n5249), .A2(n8479), .ZN(n7608) );
  NAND2_X1 U6318 ( .A1(n7606), .A2(n8486), .ZN(n5249) );
  INV_X1 U6319 ( .A(n8484), .ZN(n5250) );
  INV_X1 U6320 ( .A(n8486), .ZN(n5251) );
  INV_X1 U6321 ( .A(n8479), .ZN(n5252) );
  NAND2_X1 U6322 ( .A1(n5268), .A2(n5269), .ZN(n6141) );
  NAND2_X1 U6323 ( .A1(n6138), .A2(n5270), .ZN(n5268) );
  AND2_X1 U6324 ( .A1(n5500), .A2(n5670), .ZN(n5287) );
  NAND2_X1 U6325 ( .A1(n5713), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6326 ( .A1(n5749), .A2(n7517), .ZN(n8467) );
  AND2_X1 U6327 ( .A1(n5737), .A2(n5738), .ZN(n5288) );
  NAND2_X1 U6328 ( .A1(n6124), .A2(n8620), .ZN(n7942) );
  NAND2_X1 U6329 ( .A1(n6146), .A2(n8795), .ZN(n7157) );
  AOI21_X1 U6330 ( .B1(n9162), .B2(n6131), .A(n6130), .ZN(n9114) );
  NAND2_X1 U6331 ( .A1(n5458), .A2(n5567), .ZN(n5568) );
  NOR2_X1 U6332 ( .A1(n6713), .A2(n6712), .ZN(n6786) );
  NAND2_X2 U6333 ( .A1(n6437), .A2(n6436), .ZN(n8060) );
  NAND3_X1 U6334 ( .A1(n5291), .A2(n5290), .A3(n5292), .ZN(n7163) );
  NAND2_X1 U6335 ( .A1(n8965), .A2(n5007), .ZN(n5290) );
  NAND2_X1 U6336 ( .A1(n8965), .A2(n5302), .ZN(n5297) );
  INV_X1 U6337 ( .A(n9185), .ZN(n5303) );
  NAND2_X1 U6338 ( .A1(n9010), .A2(n5013), .ZN(n5309) );
  OR2_X1 U6339 ( .A1(n9010), .A2(n6046), .ZN(n5313) );
  NAND2_X1 U6340 ( .A1(n5318), .A2(n5012), .ZN(n8409) );
  AND2_X1 U6341 ( .A1(n9232), .A2(n10846), .ZN(n5334) );
  CLKBUF_X1 U6342 ( .A(n5337), .Z(n5335) );
  NAND4_X1 U6343 ( .A1(n5384), .A2(n5388), .A3(n6207), .A4(n5335), .ZN(n6849)
         );
  AND2_X2 U6344 ( .A1(n8018), .A2(n4956), .ZN(n9816) );
  NOR2_X2 U6345 ( .A1(n5340), .A2(n8433), .ZN(n5339) );
  INV_X1 U6346 ( .A(n10725), .ZN(n7777) );
  NOR2_X2 U6347 ( .A1(n9720), .A2(n9885), .ZN(n9695) );
  OAI21_X1 U6348 ( .B1(n9561), .B2(n9977), .A(n5347), .ZN(n5346) );
  NAND2_X1 U6349 ( .A1(n9563), .A2(n9562), .ZN(n9850) );
  XNOR2_X1 U6350 ( .A(n6876), .B(n10530), .ZN(n10540) );
  NAND2_X1 U6351 ( .A1(n6868), .A2(n5359), .ZN(n5358) );
  OR2_X1 U6352 ( .A1(n6889), .A2(n5557), .ZN(n5360) );
  OAI21_X1 U6353 ( .B1(n10637), .B2(n5360), .A(n5361), .ZN(n6891) );
  INV_X1 U6354 ( .A(n10607), .ZN(n5367) );
  NOR3_X1 U6355 ( .A1(n6423), .A2(n6206), .A3(P1_IR_REG_7__SCAN_IN), .ZN(n5383) );
  XNOR2_X1 U6356 ( .A(n5389), .B(n7354), .ZN(n7355) );
  NOR2_X1 U6357 ( .A1(n8680), .A2(n7352), .ZN(n5389) );
  NOR2_X1 U6358 ( .A1(n7355), .A2(n7356), .ZN(n7461) );
  NAND2_X1 U6359 ( .A1(n5404), .A2(n5406), .ZN(n9305) );
  NAND3_X1 U6360 ( .A1(n8715), .A2(n9378), .A3(n5412), .ZN(n5411) );
  OAI21_X1 U6361 ( .B1(n9272), .B2(n5415), .A(n5413), .ZN(n9295) );
  NAND2_X1 U6362 ( .A1(n9272), .A2(n8751), .ZN(n5416) );
  OAI21_X1 U6363 ( .B1(n9272), .B2(n8752), .A(n8751), .ZN(n9313) );
  OAI21_X1 U6364 ( .B1(n8246), .B2(n5426), .A(n5425), .ZN(n8366) );
  NAND3_X1 U6365 ( .A1(n8050), .A2(n8143), .A3(n8051), .ZN(n8144) );
  NAND2_X1 U6366 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  NAND2_X1 U6367 ( .A1(n7808), .A2(n7809), .ZN(n5429) );
  NAND3_X1 U6368 ( .A1(n4990), .A2(n7561), .A3(n5429), .ZN(n5428) );
  NAND2_X1 U6369 ( .A1(n9814), .A2(n5433), .ZN(n5430) );
  NAND2_X1 U6370 ( .A1(n5430), .A2(n5431), .ZN(n9797) );
  NAND3_X1 U6371 ( .A1(n5436), .A2(n6386), .A3(n6336), .ZN(n6411) );
  NAND2_X1 U6372 ( .A1(n9591), .A2(n5439), .ZN(n5437) );
  NAND2_X1 U6373 ( .A1(n8074), .A2(n5455), .ZN(n8169) );
  NAND2_X1 U6374 ( .A1(n8169), .A2(n8168), .ZN(n8198) );
  INV_X1 U6375 ( .A(n5565), .ZN(n5458) );
  OAI21_X1 U6376 ( .B1(n5812), .B2(n5465), .A(n5464), .ZN(n5829) );
  NAND2_X1 U6377 ( .A1(n5469), .A2(n5468), .ZN(n5900) );
  NAND2_X1 U6378 ( .A1(n5846), .A2(n5611), .ZN(n5883) );
  NOR2_X1 U6379 ( .A1(n5882), .A2(n5471), .ZN(n5470) );
  INV_X1 U6380 ( .A(n5611), .ZN(n5471) );
  NOR2_X1 U6381 ( .A1(n5612), .A2(SI_11_), .ZN(n5473) );
  INV_X1 U6382 ( .A(n5703), .ZN(n5477) );
  NAND2_X1 U6383 ( .A1(n5703), .A2(n5702), .ZN(n5705) );
  NAND3_X1 U6384 ( .A1(n5480), .A2(n5627), .A3(n5482), .ZN(n5479) );
  INV_X1 U6385 ( .A(n6014), .ZN(n5489) );
  NAND2_X1 U6386 ( .A1(n6014), .A2(n5484), .ZN(n5483) );
  INV_X1 U6387 ( .A(n6058), .ZN(n5498) );
  NAND2_X1 U6388 ( .A1(n6058), .A2(n5493), .ZN(n5492) );
  NAND2_X2 U6389 ( .A1(n5726), .A2(n5679), .ZN(n5741) );
  INV_X1 U6390 ( .A(n5668), .ZN(n5503) );
  NOR2_X1 U6391 ( .A1(n5668), .A2(n5744), .ZN(n5847) );
  NAND2_X1 U6392 ( .A1(n7072), .A2(n5512), .ZN(n5506) );
  NAND2_X1 U6393 ( .A1(n7073), .A2(n5512), .ZN(n5507) );
  NAND3_X1 U6394 ( .A1(n5507), .A2(n5509), .A3(n5506), .ZN(n8863) );
  NAND2_X1 U6395 ( .A1(n8830), .A2(n5515), .ZN(n5514) );
  OAI211_X1 U6396 ( .C1(n8830), .C2(n5516), .A(n5514), .B(n8679), .ZN(P2_U3180) );
  NAND2_X1 U6397 ( .A1(n4954), .A2(n7482), .ZN(n5524) );
  NAND2_X1 U6398 ( .A1(n4954), .A2(n7046), .ZN(n5525) );
  OAI21_X2 U6399 ( .B1(n5525), .B2(n7475), .A(n5524), .ZN(n7505) );
  NOR2_X2 U6400 ( .A1(n7472), .A2(n7045), .ZN(n7475) );
  NAND2_X1 U6401 ( .A1(n10851), .A2(n4959), .ZN(n8884) );
  NAND2_X1 U6402 ( .A1(n8807), .A2(n4958), .ZN(n8910) );
  NAND2_X1 U6403 ( .A1(n7897), .A2(n7062), .ZN(n7999) );
  NAND2_X1 U6404 ( .A1(n7999), .A2(n5531), .ZN(n5530) );
  NAND2_X1 U6405 ( .A1(n8854), .A2(n7105), .ZN(n8662) );
  NAND3_X1 U6406 ( .A1(n5536), .A2(n5535), .A3(n8893), .ZN(n8892) );
  AND2_X1 U6407 ( .A1(n5537), .A2(n5016), .ZN(n5535) );
  INV_X1 U6408 ( .A(n7618), .ZN(n5540) );
  NAND2_X1 U6409 ( .A1(n6107), .A2(n5674), .ZN(n6151) );
  OAI21_X1 U6410 ( .B1(n7603), .B2(n5781), .A(n5780), .ZN(n7715) );
  INV_X1 U6411 ( .A(n6222), .ZN(n6214) );
  OR2_X1 U6412 ( .A1(n6227), .A2(n9985), .ZN(n6217) );
  NAND2_X1 U6413 ( .A1(n6227), .A2(n6224), .ZN(n6222) );
  NAND4_X2 U6414 ( .A1(n6345), .A2(n6344), .A3(n6343), .A4(n6342), .ZN(n7351)
         );
  NAND4_X4 U6415 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n10228)
         );
  OAI21_X1 U6416 ( .B1(n5586), .B2(n5572), .A(n5571), .ZN(n5573) );
  NAND2_X1 U6417 ( .A1(n5586), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5571) );
  INV_X1 U6418 ( .A(n8586), .ZN(n9181) );
  NAND2_X1 U6419 ( .A1(n5586), .A2(n5566), .ZN(n5567) );
  NAND2_X2 U6420 ( .A1(n6239), .A2(n6238), .ZN(n6673) );
  INV_X1 U6421 ( .A(n9158), .ZN(n7174) );
  INV_X1 U6422 ( .A(n9107), .ZN(n9081) );
  AND4_X1 U6423 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n9107)
         );
  NOR2_X1 U6424 ( .A1(n7124), .A2(n7123), .ZN(n5546) );
  AND3_X1 U6425 ( .A1(n7170), .A2(n7169), .A3(n7168), .ZN(n5547) );
  AND2_X1 U6426 ( .A1(n8689), .A2(n8688), .ZN(n5548) );
  AND2_X1 U6427 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5549) );
  OR2_X1 U6428 ( .A1(n5726), .A2(n7406), .ZN(n5550) );
  OR2_X1 U6429 ( .A1(n8028), .A2(n7564), .ZN(n5551) );
  INV_X1 U6430 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U6431 ( .A1(n8713), .A2(n8712), .ZN(n5552) );
  AND2_X1 U6432 ( .A1(n7176), .A2(n7175), .ZN(n5554) );
  OR2_X1 U6433 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6007), .ZN(n5555) );
  AND2_X1 U6434 ( .A1(n7512), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5557) );
  OR2_X1 U6435 ( .A1(n10702), .A2(n7563), .ZN(n9819) );
  INV_X1 U6436 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5783) );
  INV_X1 U6437 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5918) );
  INV_X1 U6438 ( .A(n10629), .ZN(n6886) );
  AND2_X1 U6439 ( .A1(n6846), .A2(n6845), .ZN(n5558) );
  AND2_X1 U6440 ( .A1(n6506), .A2(n6320), .ZN(n5559) );
  INV_X1 U6441 ( .A(n9766), .ZN(n9581) );
  AND4_X1 U6442 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n8975)
         );
  INV_X1 U6443 ( .A(n8975), .ZN(n8999) );
  INV_X1 U6444 ( .A(n8454), .ZN(n8588) );
  INV_X1 U6445 ( .A(n9568), .ZN(n9561) );
  NOR3_X1 U6446 ( .A1(n9009), .A2(n9058), .A3(n8638), .ZN(n5563) );
  INV_X1 U6447 ( .A(n9249), .ZN(n7191) );
  AND2_X1 U6448 ( .A1(n9185), .A2(n10853), .ZN(n5564) );
  OAI21_X1 U6449 ( .B1(n7461), .B2(n4945), .A(n9368), .ZN(n9367) );
  NAND2_X1 U6450 ( .A1(n7697), .A2(n10709), .ZN(n10712) );
  NAND2_X1 U6451 ( .A1(n8803), .A2(n8590), .ZN(n8456) );
  INV_X1 U6452 ( .A(n6680), .ZN(n6681) );
  NOR2_X1 U6453 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5673) );
  NAND2_X1 U6454 ( .A1(n8589), .A2(n8455), .ZN(n8605) );
  INV_X1 U6455 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5675) );
  INV_X1 U6456 ( .A(n9169), .ZN(n7079) );
  AND2_X1 U6457 ( .A1(n7944), .A2(n5874), .ZN(n5873) );
  INV_X1 U6458 ( .A(n6809), .ZN(n6746) );
  INV_X1 U6459 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6211) );
  INV_X1 U6460 ( .A(SI_19_), .ZN(n10030) );
  OR2_X1 U6461 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  XNOR2_X1 U6462 ( .A(n7050), .B(n7669), .ZN(n7051) );
  NOR2_X1 U6463 ( .A1(n6872), .A2(n10500), .ZN(n6873) );
  INV_X1 U6464 ( .A(n6887), .ZN(n6888) );
  OR2_X1 U6465 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  INV_X1 U6466 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5670) );
  INV_X1 U6467 ( .A(n8712), .ZN(n8709) );
  INV_X1 U6468 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6320) );
  INV_X1 U6469 ( .A(n9618), .ZN(n9595) );
  NOR2_X1 U6470 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6547) );
  INV_X1 U6471 ( .A(SI_13_), .ZN(n10114) );
  NAND2_X1 U6472 ( .A1(n7057), .A2(n7899), .ZN(n7058) );
  INV_X1 U6473 ( .A(n8882), .ZN(n7097) );
  INV_X1 U6474 ( .A(n8908), .ZN(n7086) );
  NAND2_X1 U6475 ( .A1(n7051), .A2(n8930), .ZN(n7052) );
  OR2_X1 U6476 ( .A1(n7074), .A2(n8927), .ZN(n7075) );
  NAND2_X1 U6477 ( .A1(n7084), .A2(n8915), .ZN(n7085) );
  NAND2_X1 U6478 ( .A1(n10661), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U6479 ( .A1(n5555), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6019) );
  INV_X1 U6480 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10096) );
  OAI21_X1 U6481 ( .B1(n6120), .B2(n7044), .A(n8475), .ZN(n7543) );
  NAND2_X1 U6482 ( .A1(n8421), .A2(n8423), .ZN(n8424) );
  INV_X1 U6483 ( .A(n9420), .ZN(n8385) );
  NOR2_X1 U6484 ( .A1(n6452), .A2(n8149), .ZN(n6475) );
  OR2_X1 U6485 ( .A1(n6516), .A2(n6515), .ZN(n6518) );
  OAI22_X1 U6486 ( .A1(n9618), .A2(n9770), .B1(n9617), .B2(n9616), .ZN(n9619)
         );
  AND2_X1 U6487 ( .A1(n6758), .A2(n9613), .ZN(n9630) );
  INV_X1 U6488 ( .A(n9689), .ZN(n9590) );
  INV_X1 U6489 ( .A(n9889), .ZN(n9559) );
  NOR2_X1 U6490 ( .A1(n6506), .A2(n6320), .ZN(n6321) );
  NAND2_X1 U6491 ( .A1(n6485), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U6492 ( .A1(n10226), .A2(n10744), .ZN(n7836) );
  INV_X1 U6493 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U6494 ( .A1(n6218), .A2(n6210), .ZN(n6216) );
  AND2_X1 U6495 ( .A1(n6511), .A2(n6304), .ZN(n6497) );
  INV_X1 U6496 ( .A(n7894), .ZN(n7059) );
  OR2_X1 U6497 ( .A1(n7149), .A2(n7147), .ZN(n8898) );
  NOR2_X1 U6498 ( .A1(n10538), .A2(n6877), .ZN(n10557) );
  NOR2_X1 U6499 ( .A1(n10571), .A2(n6880), .ZN(n10590) );
  NAND2_X1 U6500 ( .A1(n8922), .A2(n9082), .ZN(n6116) );
  AND2_X1 U6501 ( .A1(n6136), .A2(n8637), .ZN(n6137) );
  NAND2_X1 U6502 ( .A1(n10096), .A2(n5984), .ZN(n5997) );
  AND2_X1 U6503 ( .A1(n5865), .A2(n10187), .ZN(n5867) );
  OR2_X1 U6504 ( .A1(n8590), .A2(n6186), .ZN(n7520) );
  INV_X1 U6505 ( .A(n8987), .ZN(n9012) );
  AND2_X1 U6506 ( .A1(n8515), .A2(n8504), .ZN(n8628) );
  INV_X1 U6507 ( .A(n9103), .ZN(n9168) );
  AND2_X1 U6508 ( .A1(n7498), .A2(n7495), .ZN(n7496) );
  AND3_X1 U6509 ( .A1(n7695), .A2(n9984), .A3(n7574), .ZN(n7377) );
  AND2_X1 U6510 ( .A1(n6581), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6587) );
  INV_X1 U6511 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8149) );
  OR2_X1 U6512 ( .A1(n10304), .A2(n9998), .ZN(n10461) );
  AND3_X1 U6513 ( .A1(n6593), .A2(n6592), .A3(n6591), .ZN(n9769) );
  NAND2_X1 U6514 ( .A1(n10235), .A2(n7702), .ZN(n10237) );
  OR2_X1 U6515 ( .A1(n9567), .A2(n9617), .ZN(n9853) );
  INV_X1 U6516 ( .A(n8268), .ZN(n10803) );
  INV_X1 U6517 ( .A(n10227), .ZN(n9770) );
  OR2_X1 U6518 ( .A1(n10702), .A2(n7548), .ZN(n10814) );
  XNOR2_X1 U6519 ( .A(n5631), .B(n10137), .ZN(n5960) );
  AND2_X1 U6520 ( .A1(n5627), .A2(n5626), .ZN(n5702) );
  INV_X1 U6521 ( .A(SI_5_), .ZN(n5793) );
  INV_X1 U6522 ( .A(n7152), .ZN(n7153) );
  AND4_X1 U6523 ( .A1(n8600), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(n8587)
         );
  AND4_X1 U6524 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n8878)
         );
  AND4_X1 U6525 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n9169)
         );
  INV_X1 U6526 ( .A(n7207), .ZN(n10483) );
  OR2_X1 U6527 ( .A1(n8344), .A2(n7527), .ZN(n10831) );
  INV_X1 U6528 ( .A(n8614), .ZN(n9009) );
  AND2_X1 U6529 ( .A1(n8530), .A2(n8531), .ZN(n8615) );
  NAND2_X1 U6530 ( .A1(n7148), .A2(n8590), .ZN(n9106) );
  AND2_X1 U6531 ( .A1(n7529), .A2(n7172), .ZN(n9165) );
  NOR2_X1 U6532 ( .A1(n7126), .A2(n6184), .ZN(n7525) );
  INV_X1 U6533 ( .A(n9165), .ZN(n9182) );
  AND2_X1 U6534 ( .A1(n7239), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6183) );
  NAND2_X1 U6535 ( .A1(n8281), .A2(n6180), .ZN(n7138) );
  XNOR2_X1 U6536 ( .A(n6109), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8659) );
  INV_X1 U6537 ( .A(n9404), .ZN(n9372) );
  AND4_X1 U6538 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n9618)
         );
  AND4_X1 U6539 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(n9771)
         );
  AND4_X1 U6540 ( .A1(n6325), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n8371)
         );
  INV_X1 U6541 ( .A(n8138), .ZN(n8327) );
  INV_X1 U6542 ( .A(n10466), .ZN(n10689) );
  INV_X1 U6543 ( .A(n9819), .ZN(n9562) );
  INV_X1 U6544 ( .A(n9700), .ZN(n9694) );
  AND2_X1 U6545 ( .A1(n6711), .A2(n7968), .ZN(n8014) );
  AND2_X1 U6546 ( .A1(n10712), .A2(n9552), .ZN(n9844) );
  INV_X1 U6547 ( .A(n10237), .ZN(n9840) );
  OR2_X1 U6548 ( .A1(n7575), .A2(n9983), .ZN(n10709) );
  NAND2_X1 U6549 ( .A1(n8207), .A2(n10731), .ZN(n10806) );
  INV_X1 U6550 ( .A(n6239), .ZN(n9991) );
  AND2_X1 U6551 ( .A1(n6563), .A2(n6549), .ZN(n9546) );
  AND2_X1 U6552 ( .A1(n6501), .A2(n6500), .ZN(n10433) );
  AND2_X1 U6553 ( .A1(n6426), .A2(n6425), .ZN(n10325) );
  NOR2_X1 U6554 ( .A1(n5564), .A2(n7153), .ZN(n7154) );
  INV_X1 U6555 ( .A(n10856), .ZN(n7626) );
  NAND2_X1 U6556 ( .A1(n7133), .A2(n7132), .ZN(n8907) );
  INV_X1 U6557 ( .A(n8832), .ZN(n8988) );
  INV_X1 U6558 ( .A(n9094), .ZN(n10846) );
  INV_X1 U6559 ( .A(n8868), .ZN(n8926) );
  OR2_X1 U6560 ( .A1(n7008), .A2(P2_U3151), .ZN(n8931) );
  OR2_X1 U6561 ( .A1(n9175), .A2(n9165), .ZN(n9159) );
  OR2_X1 U6562 ( .A1(n9175), .A2(n8344), .ZN(n9158) );
  INV_X2 U6563 ( .A(n8349), .ZN(n9175) );
  AND3_X1 U6564 ( .A1(n8033), .A2(n8032), .A3(n8031), .ZN(n10781) );
  AND2_X2 U6565 ( .A1(n7188), .A2(n7185), .ZN(n10843) );
  NOR2_X1 U6566 ( .A1(n7226), .A2(n9255), .ZN(n7279) );
  INV_X1 U6567 ( .A(n5688), .ZN(n9265) );
  INV_X1 U6568 ( .A(n6149), .ZN(n7958) );
  INV_X1 U6569 ( .A(n10597), .ZN(n7309) );
  AND2_X1 U6570 ( .A1(n7223), .A2(n9429), .ZN(n10683) );
  OR3_X1 U6571 ( .A1(n9295), .A2(n9299), .A3(n9294), .ZN(n9304) );
  INV_X1 U6572 ( .A(n9879), .ZN(n9685) );
  AND2_X1 U6573 ( .A1(n7378), .A2(n10709), .ZN(n9398) );
  INV_X1 U6574 ( .A(n9666), .ZN(n9633) );
  INV_X1 U6575 ( .A(n9281), .ZN(n9782) );
  INV_X1 U6576 ( .A(n8371), .ZN(n9418) );
  OR2_X1 U6577 ( .A1(n7383), .A2(n7194), .ZN(n9427) );
  AND3_X1 U6578 ( .A1(n10416), .A2(n10415), .A3(n10414), .ZN(n10418) );
  NAND2_X1 U6579 ( .A1(n10235), .A2(n10233), .ZN(n9835) );
  NAND2_X1 U6580 ( .A1(n10819), .A2(n9931), .ZN(n9928) );
  INV_X1 U6581 ( .A(n10819), .ZN(n10818) );
  INV_X1 U6582 ( .A(n9638), .ZN(n9944) );
  INV_X1 U6583 ( .A(n9754), .ZN(n9965) );
  INV_X1 U6584 ( .A(n8433), .ZN(n8302) );
  INV_X1 U6585 ( .A(n10823), .ZN(n10820) );
  NAND2_X1 U6586 ( .A1(n9981), .A2(n9980), .ZN(n10003) );
  OAI21_X1 U6587 ( .B1(n6851), .B2(n6850), .A(n6853), .ZN(n8448) );
  INV_X1 U6588 ( .A(n6848), .ZN(n8028) );
  CLKBUF_X1 U6589 ( .A(n8027), .Z(n10000) );
  INV_X1 U6590 ( .A(n9997), .ZN(n8445) );
  INV_X2 U6591 ( .A(n8931), .ZN(P2_U3893) );
  OAI21_X1 U6592 ( .B1(n7035), .B2(n10677), .A(n7034), .ZN(P2_U3200) );
  NAND2_X1 U6593 ( .A1(n6194), .A2(n6193), .ZN(P2_U3487) );
  INV_X2 U6594 ( .A(n9427), .ZN(P1_U3973) );
  OAI21_X1 U6595 ( .B1(n5586), .B2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .ZN(
        n5565) );
  INV_X1 U6596 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5566) );
  INV_X1 U6597 ( .A(SI_1_), .ZN(n10164) );
  NAND2_X1 U6598 ( .A1(n5568), .A2(n10164), .ZN(n5569) );
  MUX2_X1 U6599 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5586), .Z(n5719) );
  NAND2_X1 U6600 ( .A1(n5718), .A2(n5719), .ZN(n5723) );
  OR2_X1 U6601 ( .A1(n5573), .A2(SI_2_), .ZN(n5574) );
  NAND2_X1 U6602 ( .A1(n5573), .A2(SI_2_), .ZN(n5575) );
  AND2_X1 U6603 ( .A1(n5574), .A2(n5575), .ZN(n5740) );
  NAND2_X1 U6604 ( .A1(n5739), .A2(n5740), .ZN(n5576) );
  NAND2_X1 U6605 ( .A1(n5576), .A2(n5575), .ZN(n5755) );
  INV_X2 U6606 ( .A(n5586), .ZN(n5578) );
  INV_X8 U6607 ( .A(n5578), .ZN(n7195) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U6609 ( .A1(n5581), .A2(SI_3_), .ZN(n5585) );
  INV_X1 U6610 ( .A(n5581), .ZN(n5583) );
  INV_X1 U6611 ( .A(SI_3_), .ZN(n5582) );
  NAND2_X1 U6612 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  AND2_X2 U6613 ( .A1(n5585), .A2(n5584), .ZN(n5754) );
  NAND2_X1 U6614 ( .A1(n5755), .A2(n5754), .ZN(n5757) );
  NAND2_X1 U6615 ( .A1(n5757), .A2(n5585), .ZN(n5771) );
  MUX2_X1 U6616 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5586), .Z(n5587) );
  NAND2_X1 U6617 ( .A1(n5587), .A2(SI_4_), .ZN(n5591) );
  INV_X1 U6618 ( .A(n5587), .ZN(n5589) );
  INV_X1 U6619 ( .A(SI_4_), .ZN(n5588) );
  NAND2_X1 U6620 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  AND2_X1 U6621 ( .A1(n5591), .A2(n5590), .ZN(n5770) );
  NAND2_X1 U6622 ( .A1(n5771), .A2(n5770), .ZN(n5773) );
  MUX2_X1 U6623 ( .A(n7209), .B(n5592), .S(n7195), .Z(n5792) );
  NAND2_X1 U6624 ( .A1(n5792), .A2(n5793), .ZN(n5593) );
  MUX2_X1 U6625 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7195), .Z(n5594) );
  NAND2_X1 U6626 ( .A1(n5594), .A2(SI_6_), .ZN(n5596) );
  OAI21_X1 U6627 ( .B1(n5594), .B2(SI_6_), .A(n5596), .ZN(n5806) );
  INV_X1 U6628 ( .A(n5806), .ZN(n5595) );
  MUX2_X1 U6629 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5586), .Z(n5598) );
  NAND2_X1 U6630 ( .A1(n5598), .A2(SI_7_), .ZN(n5603) );
  INV_X1 U6631 ( .A(n5598), .ZN(n5600) );
  INV_X1 U6632 ( .A(SI_7_), .ZN(n5599) );
  NAND2_X1 U6633 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  NAND2_X1 U6634 ( .A1(n5603), .A2(n5601), .ZN(n5813) );
  INV_X1 U6635 ( .A(n5813), .ZN(n5602) );
  MUX2_X1 U6636 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5586), .Z(n5604) );
  XNOR2_X1 U6637 ( .A(n5604), .B(SI_8_), .ZN(n5857) );
  INV_X1 U6638 ( .A(n5604), .ZN(n5605) );
  MUX2_X1 U6639 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7195), .Z(n5606) );
  XNOR2_X1 U6640 ( .A(n5606), .B(n10047), .ZN(n5830) );
  MUX2_X1 U6641 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7195), .Z(n5607) );
  NAND2_X1 U6642 ( .A1(n5607), .A2(SI_10_), .ZN(n5611) );
  INV_X1 U6643 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U6644 ( .A1(n5608), .A2(n10043), .ZN(n5609) );
  NAND2_X1 U6645 ( .A1(n5611), .A2(n5609), .ZN(n5844) );
  INV_X1 U6646 ( .A(n5844), .ZN(n5610) );
  MUX2_X1 U6647 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7195), .Z(n5612) );
  XNOR2_X1 U6648 ( .A(n5612), .B(SI_11_), .ZN(n5882) );
  MUX2_X1 U6649 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7195), .Z(n5613) );
  NAND2_X1 U6650 ( .A1(n5613), .A2(SI_12_), .ZN(n5614) );
  OAI21_X1 U6651 ( .B1(n5613), .B2(SI_12_), .A(n5614), .ZN(n5897) );
  NAND2_X1 U6652 ( .A1(n5900), .A2(n5614), .ZN(n5913) );
  MUX2_X1 U6653 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7195), .Z(n5615) );
  NAND2_X1 U6654 ( .A1(n5615), .A2(SI_13_), .ZN(n5618) );
  INV_X1 U6655 ( .A(n5615), .ZN(n5616) );
  NAND2_X1 U6656 ( .A1(n5616), .A2(n10114), .ZN(n5617) );
  NAND2_X1 U6657 ( .A1(n5913), .A2(n5912), .ZN(n5915) );
  NAND2_X1 U6658 ( .A1(n5915), .A2(n5618), .ZN(n5928) );
  MUX2_X1 U6659 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7195), .Z(n5619) );
  NAND2_X1 U6660 ( .A1(n5619), .A2(SI_14_), .ZN(n5623) );
  INV_X1 U6661 ( .A(n5619), .ZN(n5621) );
  INV_X1 U6662 ( .A(SI_14_), .ZN(n5620) );
  NAND2_X1 U6663 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U6664 ( .A1(n5930), .A2(n5623), .ZN(n5703) );
  MUX2_X1 U6665 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7195), .Z(n5624) );
  NAND2_X1 U6666 ( .A1(n5624), .A2(SI_15_), .ZN(n5627) );
  INV_X1 U6667 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U6668 ( .A1(n5625), .A2(n10147), .ZN(n5626) );
  MUX2_X1 U6669 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7195), .Z(n5628) );
  XNOR2_X1 U6670 ( .A(n5628), .B(SI_16_), .ZN(n5943) );
  INV_X1 U6671 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U6672 ( .A1(n5629), .A2(n10143), .ZN(n5630) );
  MUX2_X1 U6673 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7195), .Z(n5631) );
  MUX2_X1 U6674 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7195), .Z(n5632) );
  NAND2_X1 U6675 ( .A1(n5632), .A2(SI_18_), .ZN(n5637) );
  INV_X1 U6676 ( .A(n5632), .ZN(n5634) );
  INV_X1 U6677 ( .A(SI_18_), .ZN(n5633) );
  NAND2_X1 U6678 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  NAND2_X1 U6679 ( .A1(n5637), .A2(n5635), .ZN(n5973) );
  INV_X1 U6680 ( .A(n5973), .ZN(n5636) );
  NAND2_X1 U6681 ( .A1(n5972), .A2(n5636), .ZN(n5976) );
  NAND2_X1 U6682 ( .A1(n5976), .A2(n5637), .ZN(n5992) );
  MUX2_X1 U6683 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7195), .Z(n5638) );
  XNOR2_X1 U6684 ( .A(n5638), .B(SI_19_), .ZN(n5991) );
  INV_X1 U6685 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U6686 ( .A1(n5639), .A2(n10030), .ZN(n5640) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7195), .Z(n5641) );
  XNOR2_X1 U6688 ( .A(n5641), .B(n10116), .ZN(n6004) );
  NAND2_X1 U6689 ( .A1(n6003), .A2(n6004), .ZN(n5644) );
  INV_X1 U6690 ( .A(n5641), .ZN(n5642) );
  NAND2_X1 U6691 ( .A1(n5642), .A2(n10116), .ZN(n5643) );
  NAND2_X1 U6692 ( .A1(n5644), .A2(n5643), .ZN(n6014) );
  MUX2_X1 U6693 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7195), .Z(n5645) );
  NAND2_X1 U6694 ( .A1(n5645), .A2(SI_21_), .ZN(n5647) );
  OAI21_X1 U6695 ( .B1(n5645), .B2(SI_21_), .A(n5647), .ZN(n6015) );
  MUX2_X1 U6696 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7195), .Z(n5648) );
  XNOR2_X1 U6697 ( .A(n5648), .B(SI_22_), .ZN(n6026) );
  INV_X1 U6698 ( .A(n5648), .ZN(n5650) );
  INV_X1 U6699 ( .A(SI_22_), .ZN(n5649) );
  NAND2_X1 U6700 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  MUX2_X1 U6701 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7195), .Z(n5652) );
  XNOR2_X1 U6702 ( .A(n5652), .B(n10132), .ZN(n6037) );
  NAND2_X1 U6703 ( .A1(n6036), .A2(n6037), .ZN(n5655) );
  INV_X1 U6704 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U6705 ( .A1(n5653), .A2(n10132), .ZN(n5654) );
  NAND2_X1 U6706 ( .A1(n5655), .A2(n5654), .ZN(n6047) );
  MUX2_X1 U6707 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7195), .Z(n5656) );
  XNOR2_X1 U6708 ( .A(n5656), .B(n10012), .ZN(n6048) );
  NAND2_X1 U6709 ( .A1(n6047), .A2(n6048), .ZN(n5659) );
  INV_X1 U6710 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U6711 ( .A1(n5657), .A2(n10012), .ZN(n5658) );
  NAND2_X1 U6712 ( .A1(n5659), .A2(n5658), .ZN(n6058) );
  MUX2_X1 U6713 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7195), .Z(n5660) );
  NAND2_X1 U6714 ( .A1(n5660), .A2(SI_25_), .ZN(n5662) );
  OAI21_X1 U6715 ( .B1(n5660), .B2(SI_25_), .A(n5662), .ZN(n6059) );
  MUX2_X1 U6716 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7195), .Z(n5663) );
  XNOR2_X1 U6717 ( .A(n5663), .B(SI_26_), .ZN(n6070) );
  MUX2_X1 U6718 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7195), .Z(n6086) );
  XNOR2_X1 U6719 ( .A(n6086), .B(n10122), .ZN(n6084) );
  XNOR2_X1 U6720 ( .A(n6085), .B(n6084), .ZN(n8438) );
  NOR2_X2 U6721 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5665) );
  NOR2_X2 U6722 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5664) );
  NOR2_X1 U6723 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5672) );
  NOR2_X1 U6724 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5671) );
  NAND3_X1 U6725 ( .A1(n6153), .A2(n6182), .A3(n5675), .ZN(n5676) );
  INV_X1 U6726 ( .A(n7195), .ZN(n5679) );
  INV_X2 U6727 ( .A(n5741), .ZN(n8593) );
  NAND2_X1 U6728 ( .A1(n8438), .A2(n8593), .ZN(n5681) );
  INV_X1 U6729 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8787) );
  OR2_X1 U6730 ( .A1(n5774), .A2(n8787), .ZN(n5680) );
  INV_X1 U6731 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6732 ( .A1(n5686), .A2(n5683), .ZN(n9258) );
  INV_X1 U6733 ( .A(n5691), .ZN(n8690) );
  NAND2_X1 U6734 ( .A1(n5764), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5695) );
  NOR2_X1 U6735 ( .A1(n5691), .A2(n9265), .ZN(n5713) );
  NAND2_X1 U6736 ( .A1(n8596), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5694) );
  NOR2_X1 U6737 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5782) );
  NAND2_X1 U6738 ( .A1(n5782), .A2(n5783), .ZN(n5800) );
  NAND2_X1 U6739 ( .A1(n5919), .A2(n5918), .ZN(n5934) );
  INV_X1 U6740 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U6741 ( .A1(n10206), .A2(n6019), .ZN(n6040) );
  INV_X1 U6742 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U6743 ( .A1(n6051), .A2(n10192), .ZN(n6075) );
  NOR2_X1 U6744 ( .A1(n6077), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6093) );
  INV_X1 U6745 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U6746 ( .A1(n6077), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U6747 ( .A1(n6094), .A2(n5690), .ZN(n8969) );
  NAND2_X1 U6748 ( .A1(n6112), .A2(n8969), .ZN(n5693) );
  AND2_X2 U6749 ( .A1(n5691), .A2(n9265), .ZN(n5735) );
  NAND2_X1 U6750 ( .A1(n5735), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5692) );
  INV_X1 U6751 ( .A(n8976), .ZN(n8923) );
  NAND2_X1 U6752 ( .A1(n5764), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U6753 ( .A1(n8596), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5700) );
  INV_X1 U6754 ( .A(n5953), .ZN(n5697) );
  NAND2_X1 U6755 ( .A1(n5936), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6756 ( .A1(n5697), .A2(n5696), .ZN(n8917) );
  NAND2_X1 U6757 ( .A1(n6112), .A2(n8917), .ZN(n5699) );
  NAND2_X1 U6758 ( .A1(n5735), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5698) );
  OR2_X1 U6759 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U6760 ( .A1(n5705), .A2(n5704), .ZN(n7442) );
  OR2_X1 U6761 ( .A1(n7442), .A2(n5741), .ZN(n5712) );
  NAND2_X1 U6762 ( .A1(n5980), .A2(n5707), .ZN(n5708) );
  NAND2_X1 U6763 ( .A1(n5708), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5931) );
  INV_X1 U6764 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6765 ( .A1(n5931), .A2(n5709), .ZN(n5710) );
  NAND2_X1 U6766 ( .A1(n5710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U6767 ( .A(n5946), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U6768 ( .A1(n5994), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6862), .B2(
        n10629), .ZN(n5711) );
  NAND2_X1 U6769 ( .A1(n5712), .A2(n5711), .ZN(n8413) );
  INV_X1 U6770 ( .A(n8413), .ZN(n9250) );
  NAND2_X1 U6771 ( .A1(n5713), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U6772 ( .A1(n5735), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U6773 ( .A1(n5734), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5714) );
  INV_X1 U6774 ( .A(n5718), .ZN(n5721) );
  INV_X1 U6775 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U6776 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  AND2_X1 U6777 ( .A1(n5723), .A2(n5722), .ZN(n7196) );
  AOI21_X1 U6778 ( .B1(n5549), .B2(P2_IR_REG_1__SCAN_IN), .A(n5724), .ZN(n5725) );
  INV_X1 U6779 ( .A(n6902), .ZN(n6904) );
  NAND2_X1 U6780 ( .A1(n8473), .A2(n8475), .ZN(n6120) );
  NAND2_X1 U6781 ( .A1(n5734), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6782 ( .A1(n5713), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6783 ( .A1(n5735), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6784 ( .A1(n5764), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U6785 ( .A1(n5679), .A2(SI_0_), .ZN(n5732) );
  XNOR2_X1 U6786 ( .A(n5732), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9271) );
  MUX2_X1 U6787 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9271), .S(n5726), .Z(n7631) );
  NAND2_X1 U6788 ( .A1(n7041), .A2(n7590), .ZN(n5733) );
  NAND2_X1 U6789 ( .A1(n5734), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U6790 ( .A1(n5735), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5737) );
  XNOR2_X1 U6791 ( .A(n5739), .B(n5740), .ZN(n8450) );
  OR2_X1 U6792 ( .A1(n5741), .A2(n8450), .ZN(n5748) );
  OR2_X1 U6793 ( .A1(n5774), .A2(n5572), .ZN(n5747) );
  NOR2_X1 U6794 ( .A1(n6902), .A2(n5685), .ZN(n5743) );
  OR2_X1 U6795 ( .A1(n5726), .A2(n8449), .ZN(n5746) );
  INV_X1 U6796 ( .A(n7544), .ZN(n5749) );
  NAND2_X1 U6797 ( .A1(n7538), .A2(n7544), .ZN(n8464) );
  NAND2_X1 U6798 ( .A1(n7545), .A2(n6121), .ZN(n5751) );
  NAND2_X1 U6799 ( .A1(n7517), .A2(n7544), .ZN(n5750) );
  NAND2_X1 U6800 ( .A1(n5751), .A2(n5750), .ZN(n7515) );
  INV_X1 U6801 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U6802 ( .A1(n5735), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5753) );
  OR2_X1 U6803 ( .A1(n5774), .A2(n5580), .ZN(n5762) );
  OR2_X1 U6804 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  NAND2_X1 U6805 ( .A1(n5757), .A2(n5756), .ZN(n7205) );
  OR2_X1 U6806 ( .A1(n5741), .A2(n7205), .ZN(n5761) );
  MUX2_X1 U6807 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5758), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5759) );
  NAND2_X1 U6808 ( .A1(n5759), .A2(n5789), .ZN(n7206) );
  OR2_X1 U6809 ( .A1(n5726), .A2(n7206), .ZN(n5760) );
  NOR2_X1 U6810 ( .A1(n8932), .A2(n7530), .ZN(n5763) );
  OAI22_X1 U6811 ( .A1(n7515), .A2(n5763), .B1(n7605), .B2(n7709), .ZN(n7603)
         );
  NAND2_X1 U6812 ( .A1(n5764), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U6813 ( .A1(n5713), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5768) );
  AND2_X1 U6814 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5765) );
  OR2_X1 U6815 ( .A1(n5765), .A2(n5782), .ZN(n7609) );
  NAND2_X1 U6816 ( .A1(n5734), .A2(n7609), .ZN(n5767) );
  NAND2_X1 U6817 ( .A1(n5735), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5766) );
  OR2_X1 U6818 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  NAND2_X1 U6819 ( .A1(n5773), .A2(n5772), .ZN(n7202) );
  OR2_X1 U6820 ( .A1(n5741), .A2(n7202), .ZN(n5779) );
  INV_X1 U6821 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7201) );
  OR2_X1 U6822 ( .A1(n5774), .A2(n7201), .ZN(n5777) );
  NAND2_X1 U6823 ( .A1(n5789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5776) );
  INV_X1 U6824 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5775) );
  NOR2_X1 U6825 ( .A1(n7717), .A2(n7669), .ZN(n5781) );
  NAND2_X1 U6826 ( .A1(n7717), .A2(n7669), .ZN(n5780) );
  NAND2_X1 U6827 ( .A1(n5764), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6828 ( .A1(n8596), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5787) );
  OR2_X1 U6829 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  NAND2_X1 U6830 ( .A1(n5800), .A2(n5784), .ZN(n7722) );
  NAND2_X1 U6831 ( .A1(n5734), .A2(n7722), .ZN(n5786) );
  NAND2_X1 U6832 ( .A1(n5735), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U6833 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  INV_X1 U6834 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5790) );
  XNOR2_X1 U6835 ( .A(n5791), .B(n5790), .ZN(n7207) );
  INV_X1 U6836 ( .A(n5792), .ZN(n5794) );
  XNOR2_X1 U6837 ( .A(n5794), .B(n5793), .ZN(n5795) );
  XNOR2_X1 U6838 ( .A(n5796), .B(n5795), .ZN(n7208) );
  OR2_X1 U6839 ( .A1(n7208), .A2(n5741), .ZN(n5798) );
  OR2_X1 U6840 ( .A1(n5774), .A2(n7209), .ZN(n5797) );
  OAI211_X1 U6841 ( .C1(n5726), .C2(n7207), .A(n5798), .B(n5797), .ZN(n7723)
         );
  INV_X1 U6842 ( .A(n7723), .ZN(n7906) );
  AND2_X1 U6843 ( .A1(n7915), .A2(n7906), .ZN(n5799) );
  OAI22_X1 U6844 ( .A1(n7715), .A2(n5799), .B1(n7906), .B2(n7915), .ZN(n7912)
         );
  NAND2_X1 U6845 ( .A1(n5764), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6846 ( .A1(n8596), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U6847 ( .A1(n5800), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6848 ( .A1(n5821), .A2(n5801), .ZN(n8901) );
  NAND2_X1 U6849 ( .A1(n5734), .A2(n8901), .ZN(n5803) );
  NAND2_X1 U6850 ( .A1(n5735), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5802) );
  NAND4_X1 U6851 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n7899)
         );
  XNOR2_X1 U6852 ( .A(n5807), .B(n5595), .ZN(n7210) );
  NAND2_X1 U6853 ( .A1(n7210), .A2(n8593), .ZN(n5811) );
  OR2_X1 U6854 ( .A1(n5818), .A2(n5685), .ZN(n5809) );
  AOI22_X1 U6855 ( .A1(n5994), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6862), .B2(
        n8944), .ZN(n5810) );
  INV_X1 U6856 ( .A(n8036), .ZN(n8902) );
  NAND2_X1 U6857 ( .A1(n7930), .A2(n8902), .ZN(n8495) );
  NAND2_X1 U6858 ( .A1(n8036), .A2(n7899), .ZN(n8496) );
  INV_X1 U6859 ( .A(n5812), .ZN(n5814) );
  NAND2_X1 U6860 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  AND2_X1 U6861 ( .A1(n5816), .A2(n5815), .ZN(n7215) );
  NAND2_X1 U6862 ( .A1(n7215), .A2(n8593), .ZN(n5820) );
  INV_X1 U6863 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U6864 ( .A1(n5818), .A2(n5817), .ZN(n5833) );
  NAND2_X1 U6865 ( .A1(n5833), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U6866 ( .A(n5860), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U6867 ( .A1(n5994), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6862), .B2(
        n10500), .ZN(n5819) );
  NAND2_X1 U6868 ( .A1(n5820), .A2(n5819), .ZN(n7934) );
  NAND2_X1 U6869 ( .A1(n8596), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U6870 ( .A1(n5764), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5825) );
  AND2_X1 U6871 ( .A1(n5821), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5822) );
  OR2_X1 U6872 ( .A1(n5822), .A2(n5865), .ZN(n7935) );
  NAND2_X1 U6873 ( .A1(n5734), .A2(n7935), .ZN(n5824) );
  NAND2_X1 U6874 ( .A1(n5735), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5823) );
  NAND4_X1 U6875 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n8929)
         );
  OR2_X1 U6876 ( .A1(n7934), .A2(n8929), .ZN(n7947) );
  NAND2_X1 U6877 ( .A1(n7934), .A2(n8929), .ZN(n5827) );
  NAND2_X1 U6878 ( .A1(n7947), .A2(n5827), .ZN(n8620) );
  OR2_X1 U6879 ( .A1(n8622), .A2(n8620), .ZN(n5828) );
  NAND2_X1 U6880 ( .A1(n7930), .A2(n8036), .ZN(n7926) );
  OR2_X1 U6881 ( .A1(n8620), .A2(n7926), .ZN(n7925) );
  AND2_X1 U6882 ( .A1(n7925), .A2(n7947), .ZN(n7944) );
  XNOR2_X1 U6883 ( .A(n5829), .B(n5830), .ZN(n7243) );
  NAND2_X1 U6884 ( .A1(n7243), .A2(n8593), .ZN(n5836) );
  INV_X1 U6885 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5859) );
  INV_X1 U6886 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U6887 ( .A1(n5859), .A2(n5831), .ZN(n5832) );
  OAI21_X1 U6888 ( .B1(n5833), .B2(n5832), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5834) );
  XNOR2_X1 U6889 ( .A(n5834), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U6890 ( .A1(n5994), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6862), .B2(
        n10530), .ZN(n5835) );
  NAND2_X1 U6891 ( .A1(n5836), .A2(n5835), .ZN(n8165) );
  NAND2_X1 U6892 ( .A1(n8596), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U6893 ( .A1(n5735), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5841) );
  OR2_X1 U6894 ( .A1(n5867), .A2(n5837), .ZN(n5838) );
  NAND2_X1 U6895 ( .A1(n5850), .A2(n5838), .ZN(n8135) );
  NAND2_X1 U6896 ( .A1(n5734), .A2(n8135), .ZN(n5840) );
  NAND2_X1 U6897 ( .A1(n5764), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6898 ( .A1(n8165), .A2(n8289), .ZN(n8502) );
  NAND2_X1 U6899 ( .A1(n8509), .A2(n8502), .ZN(n8625) );
  OR2_X1 U6900 ( .A1(n5847), .A2(n5685), .ZN(n5848) );
  XNOR2_X1 U6901 ( .A(n5848), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U6902 ( .A1(n5994), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6862), .B2(
        n10546), .ZN(n5849) );
  NAND2_X1 U6903 ( .A1(n8596), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6904 ( .A1(n5735), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6905 ( .A1(n5850), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6906 ( .A1(n5889), .A2(n5851), .ZN(n8285) );
  NAND2_X1 U6907 ( .A1(n5734), .A2(n8285), .ZN(n5853) );
  NAND2_X1 U6908 ( .A1(n5764), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5852) );
  OR2_X1 U6909 ( .A1(n5856), .A2(n8359), .ZN(n8511) );
  NAND2_X1 U6910 ( .A1(n5856), .A2(n8359), .ZN(n8512) );
  XNOR2_X1 U6911 ( .A(n5858), .B(n5857), .ZN(n7220) );
  NAND2_X1 U6912 ( .A1(n7220), .A2(n8593), .ZN(n5864) );
  NAND2_X1 U6913 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  NAND2_X1 U6914 ( .A1(n5861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U6915 ( .A(n5862), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U6916 ( .A1(n5994), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6862), .B2(
        n10514), .ZN(n5863) );
  NAND2_X1 U6917 ( .A1(n5864), .A2(n5863), .ZN(n8030) );
  NAND2_X1 U6918 ( .A1(n8596), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U6919 ( .A1(n5764), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5870) );
  NOR2_X1 U6920 ( .A1(n5865), .A2(n10187), .ZN(n5866) );
  OR2_X1 U6921 ( .A1(n5867), .A2(n5866), .ZN(n8003) );
  NAND2_X1 U6922 ( .A1(n5734), .A2(n8003), .ZN(n5869) );
  NAND2_X1 U6923 ( .A1(n5735), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5868) );
  OR2_X1 U6924 ( .A1(n8030), .A2(n8000), .ZN(n8128) );
  INV_X1 U6925 ( .A(n8128), .ZN(n5872) );
  NAND2_X1 U6926 ( .A1(n7924), .A2(n5873), .ZN(n5879) );
  INV_X1 U6927 ( .A(n5874), .ZN(n5877) );
  OR2_X1 U6928 ( .A1(n8030), .A2(n8133), .ZN(n8491) );
  NAND2_X1 U6929 ( .A1(n8030), .A2(n8133), .ZN(n8498) );
  INV_X1 U6930 ( .A(n8621), .ZN(n7945) );
  AND2_X1 U6931 ( .A1(n7945), .A2(n5875), .ZN(n5876) );
  INV_X1 U6932 ( .A(n8626), .ZN(n8115) );
  INV_X1 U6933 ( .A(n8289), .ZN(n8005) );
  OR2_X1 U6934 ( .A1(n8165), .A2(n8005), .ZN(n8114) );
  OR2_X1 U6935 ( .A1(n8115), .A2(n8114), .ZN(n8111) );
  INV_X1 U6936 ( .A(n8359), .ZN(n8928) );
  OR2_X1 U6937 ( .A1(n5856), .A2(n8928), .ZN(n5880) );
  AND2_X1 U6938 ( .A1(n8111), .A2(n5880), .ZN(n5881) );
  XNOR2_X1 U6939 ( .A(n5883), .B(n5882), .ZN(n7266) );
  NAND2_X1 U6940 ( .A1(n7266), .A2(n8593), .ZN(n5888) );
  NAND2_X1 U6941 ( .A1(n5884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5885) );
  MUX2_X1 U6942 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5885), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5886) );
  AND2_X1 U6943 ( .A1(n5886), .A2(n5019), .ZN(n10563) );
  AOI22_X1 U6944 ( .A1(n5994), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6862), .B2(
        n10563), .ZN(n5887) );
  NAND2_X1 U6945 ( .A1(n5888), .A2(n5887), .ZN(n8188) );
  NAND2_X1 U6946 ( .A1(n5764), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6947 ( .A1(n8596), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U6948 ( .A1(n5889), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U6949 ( .A1(n5905), .A2(n5890), .ZN(n8361) );
  NAND2_X1 U6950 ( .A1(n5734), .A2(n8361), .ZN(n5892) );
  NAND2_X1 U6951 ( .A1(n5735), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5891) );
  INV_X1 U6952 ( .A(n8400), .ZN(n8927) );
  NAND2_X1 U6953 ( .A1(n8188), .A2(n8927), .ZN(n5895) );
  OR2_X1 U6954 ( .A1(n8188), .A2(n8927), .ZN(n5896) );
  NAND2_X1 U6955 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  NAND2_X1 U6956 ( .A1(n5900), .A2(n5899), .ZN(n7276) );
  OR2_X1 U6957 ( .A1(n7276), .A2(n5741), .ZN(n5904) );
  NAND2_X1 U6958 ( .A1(n5019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5901) );
  MUX2_X1 U6959 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5901), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n5902) );
  AND2_X1 U6960 ( .A1(n5902), .A2(n5706), .ZN(n10579) );
  AOI22_X1 U6961 ( .A1(n5994), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6862), .B2(
        n10579), .ZN(n5903) );
  NAND2_X1 U6962 ( .A1(n8596), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U6963 ( .A1(n5735), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5909) );
  AND2_X1 U6964 ( .A1(n5905), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5906) );
  OR2_X1 U6965 ( .A1(n5906), .A2(n5919), .ZN(n8396) );
  NAND2_X1 U6966 ( .A1(n6112), .A2(n8396), .ZN(n5908) );
  NAND2_X1 U6967 ( .A1(n5764), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5907) );
  OR2_X1 U6968 ( .A1(n8402), .A2(n8926), .ZN(n8221) );
  INV_X1 U6969 ( .A(n8221), .ZN(n5911) );
  NAND2_X1 U6970 ( .A1(n8402), .A2(n8926), .ZN(n8220) );
  OR2_X1 U6971 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  NAND2_X1 U6972 ( .A1(n5915), .A2(n5914), .ZN(n7310) );
  OR2_X1 U6973 ( .A1(n7310), .A2(n5741), .ZN(n5917) );
  XNOR2_X1 U6974 ( .A(n5980), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U6975 ( .A1(n5994), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6862), .B2(
        n10597), .ZN(n5916) );
  NAND2_X1 U6976 ( .A1(n5917), .A2(n5916), .ZN(n8237) );
  NAND2_X1 U6977 ( .A1(n5764), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U6978 ( .A1(n8596), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5923) );
  OR2_X1 U6979 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  NAND2_X1 U6980 ( .A1(n5934), .A2(n5920), .ZN(n8870) );
  NAND2_X1 U6981 ( .A1(n6112), .A2(n8870), .ZN(n5922) );
  NAND2_X1 U6982 ( .A1(n5735), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U6983 ( .A(n8237), .B(n9169), .ZN(n8520) );
  NAND2_X1 U6984 ( .A1(n8235), .A2(n8520), .ZN(n5926) );
  NAND2_X1 U6985 ( .A1(n8237), .A2(n7079), .ZN(n5925) );
  OR2_X1 U6986 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U6987 ( .A1(n5930), .A2(n5929), .ZN(n7429) );
  OR2_X1 U6988 ( .A1(n7429), .A2(n5741), .ZN(n5933) );
  XNOR2_X1 U6989 ( .A(n5931), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U6990 ( .A1(n5994), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6862), .B2(
        n10613), .ZN(n5932) );
  NAND2_X1 U6991 ( .A1(n5764), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U6992 ( .A1(n8596), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U6993 ( .A1(n5934), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U6994 ( .A1(n5936), .A2(n5935), .ZN(n10828) );
  NAND2_X1 U6995 ( .A1(n6112), .A2(n10828), .ZN(n5938) );
  NAND2_X1 U6996 ( .A1(n5735), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5937) );
  NAND4_X1 U6997 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n8925)
         );
  AND2_X1 U6998 ( .A1(n10827), .A2(n8925), .ZN(n5942) );
  OR2_X1 U6999 ( .A1(n10827), .A2(n8925), .ZN(n5941) );
  OR2_X1 U7000 ( .A1(n8413), .A2(n9171), .ZN(n8530) );
  NAND2_X1 U7001 ( .A1(n8413), .A2(n9171), .ZN(n8531) );
  XNOR2_X1 U7002 ( .A(n5944), .B(n5943), .ZN(n7510) );
  NAND2_X1 U7003 ( .A1(n7510), .A2(n8593), .ZN(n5952) );
  INV_X1 U7004 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7005 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  NAND2_X1 U7006 ( .A1(n5947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  INV_X1 U7007 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7008 ( .A1(n5949), .A2(n5948), .ZN(n5961) );
  OR2_X1 U7009 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  AOI22_X1 U7010 ( .A1(n5994), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6862), .B2(
        n10645), .ZN(n5951) );
  NAND2_X1 U7011 ( .A1(n5764), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7012 ( .A1(n8596), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U7013 ( .A1(n5953), .A2(n10081), .ZN(n5954) );
  OR2_X1 U7014 ( .A1(n5966), .A2(n5954), .ZN(n9110) );
  NAND2_X1 U7015 ( .A1(n6112), .A2(n9110), .ZN(n5956) );
  NAND2_X1 U7016 ( .A1(n5735), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7017 ( .A1(n9243), .A2(n9095), .ZN(n8538) );
  INV_X1 U7018 ( .A(n9243), .ZN(n8846) );
  XNOR2_X1 U7019 ( .A(n5959), .B(n5960), .ZN(n7615) );
  NAND2_X1 U7020 ( .A1(n7615), .A2(n8593), .ZN(n5964) );
  NAND2_X1 U7021 ( .A1(n5961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7022 ( .A(n5962), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U7023 ( .A1(n5994), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6862), .B2(
        n10663), .ZN(n5963) );
  NAND2_X1 U7024 ( .A1(n8596), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7025 ( .A1(n5735), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5970) );
  NOR2_X1 U7026 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  OR2_X1 U7027 ( .A1(n5984), .A2(n5967), .ZN(n10857) );
  NAND2_X1 U7028 ( .A1(n6112), .A2(n10857), .ZN(n5969) );
  NAND2_X1 U7029 ( .A1(n5764), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7030 ( .A(n10852), .B(n9081), .ZN(n9092) );
  INV_X1 U7031 ( .A(n9092), .ZN(n9089) );
  INV_X1 U7032 ( .A(n5972), .ZN(n5974) );
  NAND2_X1 U7033 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U7034 ( .A1(n5976), .A2(n5975), .ZN(n7666) );
  INV_X1 U7035 ( .A(n5977), .ZN(n5978) );
  NAND2_X1 U7036 ( .A1(n5978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U7037 ( .A(n5993), .B(n5981), .ZN(n7027) );
  AOI22_X1 U7038 ( .A1(n5994), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6862), .B2(
        n7027), .ZN(n5982) );
  INV_X1 U7039 ( .A(n9232), .ZN(n8891) );
  NAND2_X1 U7040 ( .A1(n5764), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7041 ( .A1(n8596), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7042 ( .A1(n5984), .A2(n10096), .ZN(n5985) );
  NAND2_X1 U7043 ( .A1(n5985), .A2(n5997), .ZN(n9086) );
  NAND2_X1 U7044 ( .A1(n6112), .A2(n9086), .ZN(n5987) );
  NAND2_X1 U7045 ( .A1(n5735), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7046 ( .A1(n8891), .A2(n9094), .ZN(n5990) );
  XNOR2_X1 U7047 ( .A(n5992), .B(n5991), .ZN(n7780) );
  NAND2_X1 U7048 ( .A1(n7780), .A2(n8593), .ZN(n5996) );
  XNOR2_X1 U7049 ( .A(n6101), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6147) );
  AOI22_X1 U7050 ( .A1(n5994), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4941), .B2(
        n6862), .ZN(n5995) );
  NAND2_X1 U7051 ( .A1(n8596), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7052 ( .A1(n5764), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7053 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(n5997), .ZN(n5998) );
  NAND2_X1 U7054 ( .A1(n5998), .A2(n6007), .ZN(n9074) );
  NAND2_X1 U7055 ( .A1(n6112), .A2(n9074), .ZN(n6000) );
  NAND2_X1 U7056 ( .A1(n5735), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7057 ( .A1(n9226), .A2(n9063), .ZN(n9056) );
  INV_X1 U7058 ( .A(n9226), .ZN(n8829) );
  XNOR2_X1 U7059 ( .A(n6003), .B(n6004), .ZN(n7956) );
  NAND2_X1 U7060 ( .A1(n7956), .A2(n8593), .ZN(n6006) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7957) );
  OR2_X1 U7062 ( .A1(n5774), .A2(n7957), .ZN(n6005) );
  NAND2_X1 U7063 ( .A1(n5764), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7064 ( .A1(n8596), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7065 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6007), .ZN(n6008) );
  NAND2_X1 U7066 ( .A1(n6008), .A2(n5555), .ZN(n9067) );
  NAND2_X1 U7067 ( .A1(n6112), .A2(n9067), .ZN(n6010) );
  NAND2_X1 U7068 ( .A1(n5735), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7069 ( .A1(n9141), .A2(n9048), .ZN(n6134) );
  NAND2_X1 U7070 ( .A1(n9039), .A2(n6134), .ZN(n9058) );
  INV_X1 U7071 ( .A(n9058), .ZN(n9061) );
  INV_X1 U7072 ( .A(n9048), .ZN(n9072) );
  NOR2_X1 U7073 ( .A1(n9141), .A2(n9072), .ZN(n9043) );
  NAND2_X1 U7074 ( .A1(n6014), .A2(n6015), .ZN(n6016) );
  NAND2_X1 U7075 ( .A1(n6013), .A2(n6016), .ZN(n8026) );
  OR2_X1 U7076 ( .A1(n8026), .A2(n5741), .ZN(n6018) );
  INV_X1 U7077 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7982) );
  OR2_X1 U7078 ( .A1(n5774), .A2(n7982), .ZN(n6017) );
  NAND2_X1 U7079 ( .A1(n5764), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7080 ( .A1(n8596), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7081 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(n5555), .ZN(n6020) );
  INV_X1 U7082 ( .A(n6019), .ZN(n6030) );
  NAND2_X1 U7083 ( .A1(n6020), .A2(n6030), .ZN(n9052) );
  NAND2_X1 U7084 ( .A1(n6112), .A2(n9052), .ZN(n6022) );
  NAND2_X1 U7085 ( .A1(n5735), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6021) );
  NAND4_X1 U7086 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n9025)
         );
  NAND2_X1 U7087 ( .A1(n9053), .A2(n9025), .ZN(n6025) );
  NAND2_X1 U7088 ( .A1(n9024), .A2(n6025), .ZN(n8637) );
  INV_X1 U7089 ( .A(n8637), .ZN(n9044) );
  XNOR2_X1 U7090 ( .A(n6027), .B(n6026), .ZN(n8104) );
  NAND2_X1 U7091 ( .A1(n8104), .A2(n8593), .ZN(n6029) );
  INV_X1 U7092 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8106) );
  OR2_X1 U7093 ( .A1(n5774), .A2(n8106), .ZN(n6028) );
  NAND2_X1 U7094 ( .A1(n5764), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7095 ( .A1(n8596), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7096 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n6030), .ZN(n6031) );
  NAND2_X1 U7097 ( .A1(n6031), .A2(n6040), .ZN(n9032) );
  NAND2_X1 U7098 ( .A1(n6112), .A2(n9032), .ZN(n6033) );
  NAND2_X1 U7099 ( .A1(n5735), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6032) );
  NAND4_X1 U7100 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n8924)
         );
  XNOR2_X1 U7101 ( .A(n9033), .B(n8924), .ZN(n9019) );
  INV_X1 U7102 ( .A(n9019), .ZN(n9023) );
  NAND3_X1 U7103 ( .A1(n9022), .A2(n9023), .A3(n9024), .ZN(n9021) );
  NAND2_X1 U7104 ( .A1(n9033), .A2(n8924), .ZN(n8556) );
  NAND2_X1 U7105 ( .A1(n9021), .A2(n8556), .ZN(n9010) );
  XNOR2_X1 U7106 ( .A(n6036), .B(n6037), .ZN(n8216) );
  NAND2_X1 U7107 ( .A1(n8216), .A2(n8593), .ZN(n6039) );
  INV_X1 U7108 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8219) );
  OR2_X1 U7109 ( .A1(n5774), .A2(n8219), .ZN(n6038) );
  INV_X1 U7110 ( .A(n9016), .ZN(n9206) );
  NAND2_X1 U7111 ( .A1(n5764), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7112 ( .A1(n8596), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7113 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n6040), .ZN(n6041) );
  NAND2_X1 U7114 ( .A1(n6041), .A2(n6052), .ZN(n9015) );
  NAND2_X1 U7115 ( .A1(n6112), .A2(n9015), .ZN(n6043) );
  NAND2_X1 U7116 ( .A1(n5735), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6042) );
  NOR2_X1 U7117 ( .A1(n9206), .A2(n8878), .ZN(n6046) );
  XNOR2_X1 U7118 ( .A(n6047), .B(n6048), .ZN(n8271) );
  NAND2_X1 U7119 ( .A1(n8271), .A2(n8593), .ZN(n6050) );
  INV_X1 U7120 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8334) );
  OR2_X1 U7121 ( .A1(n5774), .A2(n8334), .ZN(n6049) );
  NAND2_X1 U7122 ( .A1(n5764), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7123 ( .A1(n8596), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6056) );
  INV_X1 U7124 ( .A(n6051), .ZN(n6064) );
  NAND2_X1 U7125 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n6052), .ZN(n6053) );
  NAND2_X1 U7126 ( .A1(n6064), .A2(n6053), .ZN(n9003) );
  NAND2_X1 U7127 ( .A1(n6112), .A2(n9003), .ZN(n6055) );
  NAND2_X1 U7128 ( .A1(n5735), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6054) );
  NAND4_X1 U7129 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n8987)
         );
  NAND2_X1 U7130 ( .A1(n9201), .A2(n8987), .ZN(n8640) );
  NOR2_X1 U7131 ( .A1(n9201), .A2(n8987), .ZN(n8639) );
  NAND2_X1 U7132 ( .A1(n6058), .A2(n6059), .ZN(n6060) );
  NAND2_X1 U7133 ( .A1(n6061), .A2(n6060), .ZN(n8447) );
  INV_X1 U7134 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8282) );
  OR2_X1 U7135 ( .A1(n5774), .A2(n8282), .ZN(n6062) );
  NAND2_X1 U7136 ( .A1(n5764), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7137 ( .A1(n8596), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7138 ( .A1(n6064), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7139 ( .A1(n6075), .A2(n6065), .ZN(n8992) );
  NAND2_X1 U7140 ( .A1(n6112), .A2(n8992), .ZN(n6067) );
  NAND2_X1 U7141 ( .A1(n5735), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6066) );
  INV_X1 U7142 ( .A(n9195), .ZN(n8985) );
  XNOR2_X1 U7143 ( .A(n6071), .B(n6070), .ZN(n8416) );
  NAND2_X1 U7144 ( .A1(n8416), .A2(n8593), .ZN(n6074) );
  INV_X1 U7145 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6072) );
  OR2_X1 U7146 ( .A1(n5774), .A2(n6072), .ZN(n6073) );
  NAND2_X1 U7147 ( .A1(n8596), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7148 ( .A1(n5764), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7149 ( .A1(n6075), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7150 ( .A1(n6077), .A2(n6076), .ZN(n8979) );
  NAND2_X1 U7151 ( .A1(n6112), .A2(n8979), .ZN(n6079) );
  NAND2_X1 U7152 ( .A1(n5735), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7153 ( .A1(n8973), .A2(n6082), .ZN(n6083) );
  NAND2_X1 U7154 ( .A1(n6085), .A2(n6084), .ZN(n6089) );
  INV_X1 U7155 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7156 ( .A1(n6087), .A2(n10122), .ZN(n6088) );
  NAND2_X1 U7157 ( .A1(n6089), .A2(n6088), .ZN(n6196) );
  MUX2_X1 U7158 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7195), .Z(n6197) );
  XNOR2_X1 U7159 ( .A(n6197), .B(n10017), .ZN(n6195) );
  NAND2_X1 U7160 ( .A1(n9996), .A2(n8593), .ZN(n6091) );
  INV_X1 U7161 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9270) );
  OR2_X1 U7162 ( .A1(n5774), .A2(n9270), .ZN(n6090) );
  NAND2_X1 U7163 ( .A1(n8596), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7164 ( .A1(n5764), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6098) );
  INV_X1 U7165 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6092) );
  AND2_X1 U7166 ( .A1(n6093), .A2(n6092), .ZN(n6111) );
  INV_X1 U7167 ( .A(n6111), .ZN(n8440) );
  NAND2_X1 U7168 ( .A1(n6094), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7169 ( .A1(n8440), .A2(n6095), .ZN(n8798) );
  NAND2_X1 U7170 ( .A1(n6112), .A2(n8798), .ZN(n6097) );
  NAND2_X1 U7171 ( .A1(n5735), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6096) );
  NAND4_X1 U7172 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n8966)
         );
  XNOR2_X1 U7173 ( .A(n7162), .B(n8795), .ZN(n6119) );
  NAND2_X1 U7174 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7175 ( .A1(n6106), .A2(n6103), .ZN(n6104) );
  NAND2_X1 U7176 ( .A1(n8649), .A2(n6149), .ZN(n8606) );
  INV_X1 U7177 ( .A(n6107), .ZN(n6108) );
  NAND2_X1 U7178 ( .A1(n6108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7179 ( .A1(n4941), .A2(n8659), .ZN(n7127) );
  OR2_X1 U7180 ( .A1(n7002), .A2(n8788), .ZN(n6110) );
  NAND2_X1 U7181 ( .A1(n5726), .A2(n6110), .ZN(n7148) );
  NAND2_X1 U7182 ( .A1(n8923), .A2(n9080), .ZN(n6117) );
  NAND2_X1 U7183 ( .A1(n6112), .A2(n6111), .ZN(n8600) );
  NAND2_X1 U7184 ( .A1(n8596), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7185 ( .A1(n5735), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7186 ( .A1(n5764), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6113) );
  INV_X1 U7187 ( .A(n8801), .ZN(n8922) );
  INV_X1 U7188 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7189 ( .A1(n7543), .A2(n6122), .ZN(n6123) );
  NAND2_X1 U7190 ( .A1(n6123), .A2(n8467), .ZN(n7526) );
  NAND2_X1 U7191 ( .A1(n8932), .A2(n7709), .ZN(n8483) );
  NAND2_X1 U7192 ( .A1(n7717), .A2(n7610), .ZN(n8484) );
  NAND2_X1 U7193 ( .A1(n8930), .A2(n7669), .ZN(n8487) );
  AND2_X1 U7194 ( .A1(n8484), .A2(n8487), .ZN(n8479) );
  NAND2_X1 U7195 ( .A1(n7915), .A2(n7723), .ZN(n8490) );
  INV_X1 U7196 ( .A(n7915), .ZN(n8895) );
  NAND2_X1 U7197 ( .A1(n8895), .A2(n7906), .ZN(n8488) );
  INV_X1 U7198 ( .A(n8620), .ZN(n7933) );
  INV_X1 U7199 ( .A(n8929), .ZN(n8899) );
  OR2_X1 U7200 ( .A1(n7934), .A2(n8899), .ZN(n7941) );
  NAND2_X1 U7201 ( .A1(n8491), .A2(n7941), .ZN(n8506) );
  INV_X1 U7202 ( .A(n8506), .ZN(n6125) );
  INV_X1 U7203 ( .A(n8511), .ZN(n6126) );
  OR2_X1 U7204 ( .A1(n8188), .A2(n8400), .ZN(n8515) );
  AND2_X1 U7205 ( .A1(n8188), .A2(n8400), .ZN(n8514) );
  NOR2_X1 U7206 ( .A1(n8402), .A2(n8868), .ZN(n8517) );
  INV_X1 U7207 ( .A(n8517), .ZN(n7076) );
  NAND2_X1 U7208 ( .A1(n8224), .A2(n7076), .ZN(n6128) );
  AND2_X1 U7209 ( .A1(n8402), .A2(n8868), .ZN(n8518) );
  INV_X1 U7210 ( .A(n8518), .ZN(n6127) );
  NAND2_X1 U7211 ( .A1(n6128), .A2(n6127), .ZN(n8234) );
  INV_X1 U7212 ( .A(n8520), .ZN(n8629) );
  NAND2_X1 U7213 ( .A1(n8237), .A2(n9169), .ZN(n8523) );
  INV_X1 U7214 ( .A(n8523), .ZN(n6129) );
  XNOR2_X1 U7215 ( .A(n10827), .B(n8925), .ZN(n9163) );
  NAND2_X1 U7216 ( .A1(n9164), .A2(n9163), .ZN(n9162) );
  INV_X1 U7217 ( .A(n8925), .ZN(n8915) );
  NOR2_X1 U7218 ( .A1(n10827), .A2(n8915), .ZN(n8525) );
  INV_X1 U7219 ( .A(n8525), .ZN(n8405) );
  AND2_X1 U7220 ( .A1(n8405), .A2(n8530), .ZN(n6131) );
  INV_X1 U7221 ( .A(n8531), .ZN(n6130) );
  NAND2_X1 U7222 ( .A1(n9114), .A2(n8633), .ZN(n6132) );
  NAND2_X1 U7223 ( .A1(n6132), .A2(n8534), .ZN(n9090) );
  OR2_X1 U7224 ( .A1(n10852), .A2(n9107), .ZN(n6133) );
  NAND2_X1 U7225 ( .A1(n9232), .A2(n9094), .ZN(n8537) );
  INV_X1 U7226 ( .A(n8547), .ZN(n9037) );
  INV_X1 U7227 ( .A(n9039), .ZN(n6135) );
  NAND2_X1 U7228 ( .A1(n6134), .A2(n9056), .ZN(n8548) );
  INV_X1 U7229 ( .A(n8548), .ZN(n9038) );
  OR2_X1 U7230 ( .A1(n6135), .A2(n9038), .ZN(n6136) );
  INV_X1 U7231 ( .A(n9025), .ZN(n9064) );
  OR2_X1 U7232 ( .A1(n9053), .A2(n9064), .ZN(n6139) );
  INV_X1 U7233 ( .A(n8924), .ZN(n9049) );
  NAND2_X1 U7234 ( .A1(n9033), .A2(n9049), .ZN(n6140) );
  NOR2_X1 U7235 ( .A1(n9016), .A2(n8878), .ZN(n8559) );
  INV_X1 U7236 ( .A(n8559), .ZN(n8459) );
  AND2_X1 U7237 ( .A1(n9016), .A2(n8878), .ZN(n8558) );
  INV_X1 U7238 ( .A(n8558), .ZN(n8458) );
  NAND2_X1 U7239 ( .A1(n6141), .A2(n8458), .ZN(n9004) );
  OR2_X1 U7240 ( .A1(n9201), .A2(n9012), .ZN(n6142) );
  NAND2_X1 U7241 ( .A1(n9004), .A2(n6142), .ZN(n6144) );
  NAND2_X1 U7242 ( .A1(n9201), .A2(n9012), .ZN(n6143) );
  OR2_X1 U7243 ( .A1(n9195), .A2(n8975), .ZN(n8613) );
  NAND2_X1 U7244 ( .A1(n9195), .A2(n8975), .ZN(n8612) );
  NOR2_X1 U7245 ( .A1(n8678), .A2(n8832), .ZN(n8568) );
  INV_X1 U7246 ( .A(n8568), .ZN(n8567) );
  AND2_X1 U7247 ( .A1(n8678), .A2(n8832), .ZN(n8569) );
  INV_X1 U7248 ( .A(n8569), .ZN(n8566) );
  NAND2_X1 U7249 ( .A1(n9185), .A2(n8976), .ZN(n8573) );
  NAND2_X1 U7250 ( .A1(n6145), .A2(n8573), .ZN(n6146) );
  OAI21_X1 U7251 ( .B1(n6146), .B2(n8795), .A(n7157), .ZN(n8784) );
  INV_X1 U7252 ( .A(n8784), .ZN(n6150) );
  NAND2_X1 U7253 ( .A1(n7958), .A2(n8655), .ZN(n6188) );
  NAND2_X1 U7254 ( .A1(n7179), .A2(n8344), .ZN(n7629) );
  INV_X1 U7255 ( .A(n8659), .ZN(n8105) );
  AND2_X1 U7256 ( .A1(n6149), .A2(n8105), .ZN(n6148) );
  OR2_X1 U7257 ( .A1(n7661), .A2(n8659), .ZN(n7172) );
  NAND2_X1 U7258 ( .A1(n8786), .A2(n5562), .ZN(n8686) );
  NAND2_X1 U7259 ( .A1(n6151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7260 ( .A1(n6181), .A2(n6182), .ZN(n6152) );
  INV_X1 U7261 ( .A(P2_B_REG_SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7262 ( .A(n8335), .B(n6156), .ZN(n6162) );
  NAND2_X1 U7263 ( .A1(n4969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6159) );
  MUX2_X1 U7264 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6159), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6161) );
  OAI21_X2 U7265 ( .B1(n6162), .B2(n8281), .A(n6166), .ZN(n6165) );
  NAND2_X1 U7266 ( .A1(n8437), .A2(n8335), .ZN(n6163) );
  INV_X1 U7267 ( .A(n6164), .ZN(n7037) );
  OR2_X1 U7268 ( .A1(n6165), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7269 ( .A1(n8281), .A2(n6166), .ZN(n6167) );
  AND2_X1 U7270 ( .A1(n7037), .A2(n9256), .ZN(n7126) );
  NOR2_X1 U7271 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6172) );
  NOR4_X1 U7272 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6171) );
  NOR4_X1 U7273 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6170) );
  NOR4_X1 U7274 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6169) );
  NAND4_X1 U7275 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n6178)
         );
  NOR4_X1 U7276 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6176) );
  NOR4_X1 U7277 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6175) );
  NOR4_X1 U7278 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6174) );
  NOR4_X1 U7279 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6173) );
  NAND4_X1 U7280 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n6177)
         );
  NOR2_X1 U7281 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  NOR2_X1 U7282 ( .A1(n8437), .A2(n8335), .ZN(n6180) );
  INV_X1 U7283 ( .A(n9255), .ZN(n7185) );
  NAND2_X1 U7284 ( .A1(n7129), .A2(n7185), .ZN(n6184) );
  INV_X1 U7285 ( .A(n9256), .ZN(n7130) );
  NOR2_X1 U7286 ( .A1(n4941), .A2(n8105), .ZN(n6185) );
  AND2_X1 U7287 ( .A1(n6149), .A2(n6185), .ZN(n6186) );
  INV_X1 U7288 ( .A(n7172), .ZN(n8156) );
  INV_X1 U7289 ( .A(n8649), .ZN(n8471) );
  NAND2_X1 U7290 ( .A1(n8156), .A2(n8471), .ZN(n6187) );
  NAND2_X1 U7291 ( .A1(n7037), .A2(n6187), .ZN(n6189) );
  NAND2_X1 U7292 ( .A1(n8590), .A2(n6188), .ZN(n7139) );
  NAND2_X1 U7293 ( .A1(n7520), .A2(n7139), .ZN(n7518) );
  AOI22_X1 U7294 ( .A1(n7130), .A2(n7520), .B1(n6189), .B2(n7518), .ZN(n6190)
         );
  NAND2_X1 U7295 ( .A1(n9175), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6191) );
  INV_X1 U7296 ( .A(n6192), .ZN(n6193) );
  NAND2_X1 U7297 ( .A1(n6196), .A2(n6195), .ZN(n6200) );
  INV_X1 U7298 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7299 ( .A1(n6198), .A2(n10017), .ZN(n6199) );
  MUX2_X1 U7300 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7195), .Z(n6255) );
  INV_X1 U7301 ( .A(SI_29_), .ZN(n6201) );
  NOR2_X1 U7302 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6204) );
  NOR2_X1 U7303 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6203) );
  NOR2_X2 U7304 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6247) );
  NOR2_X1 U7305 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6205) );
  NAND2_X1 U7306 ( .A1(n6227), .A2(n6212), .ZN(n6218) );
  NOR2_X1 U7307 ( .A1(n6214), .A2(n6213), .ZN(n6215) );
  NAND2_X2 U7308 ( .A1(n6215), .A2(n6216), .ZN(n9440) );
  NAND2_X1 U7309 ( .A1(n9262), .A2(n4938), .ZN(n6221) );
  AND2_X2 U7310 ( .A1(n6357), .A2(n5679), .ZN(n6372) );
  NAND2_X1 U7311 ( .A1(n6692), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6220) );
  AND2_X1 U7312 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  NAND2_X1 U7313 ( .A1(n6227), .A2(n6226), .ZN(n9987) );
  NAND2_X1 U7314 ( .A1(n6669), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7315 ( .A1(n6341), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7316 ( .A1(n6401), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6416) );
  NOR2_X1 U7317 ( .A1(n6416), .A2(n6415), .ZN(n6429) );
  NAND2_X1 U7318 ( .A1(n6429), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U7319 ( .A1(n6321), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6554) );
  INV_X1 U7320 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6553) );
  INV_X1 U7321 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7322 ( .A1(n6587), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6588) );
  INV_X1 U7323 ( .A(n6597), .ZN(n6230) );
  NAND2_X1 U7324 ( .A1(n6230), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6293) );
  INV_X1 U7325 ( .A(n6293), .ZN(n6231) );
  NAND2_X1 U7326 ( .A1(n6231), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6283) );
  INV_X1 U7327 ( .A(n6283), .ZN(n6232) );
  NAND2_X1 U7328 ( .A1(n6232), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6615) );
  INV_X1 U7329 ( .A(n6615), .ZN(n6233) );
  NAND2_X1 U7330 ( .A1(n6233), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6630) );
  INV_X1 U7331 ( .A(n6630), .ZN(n6234) );
  NAND2_X1 U7332 ( .A1(n6234), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6645) );
  INV_X1 U7333 ( .A(n6645), .ZN(n6235) );
  NAND2_X1 U7334 ( .A1(n6235), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6660) );
  INV_X1 U7335 ( .A(n6660), .ZN(n6236) );
  NAND2_X1 U7336 ( .A1(n6236), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6672) );
  INV_X1 U7337 ( .A(n6672), .ZN(n6237) );
  NAND2_X1 U7338 ( .A1(n6237), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9600) );
  OR2_X1 U7339 ( .A1(n6367), .A2(n9600), .ZN(n6242) );
  INV_X1 U7340 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6240) );
  OR2_X1 U7341 ( .A1(n6673), .A2(n6240), .ZN(n6241) );
  NAND4_X1 U7342 ( .A1(n6244), .A2(n6243), .A3(n6242), .A4(n6241), .ZN(n9634)
         );
  INV_X1 U7343 ( .A(n9634), .ZN(n6245) );
  NAND2_X1 U7344 ( .A1(n9560), .A2(n6245), .ZN(n6833) );
  INV_X1 U7345 ( .A(n6833), .ZN(n6252) );
  NOR2_X1 U7346 ( .A1(n9560), .A2(n6245), .ZN(n6764) );
  INV_X1 U7347 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7348 ( .A1(n4964), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6251) );
  MUX2_X1 U7349 ( .A(n6252), .B(n6764), .S(n7553), .Z(n6701) );
  NAND2_X1 U7350 ( .A1(n6253), .A2(SI_29_), .ZN(n6258) );
  INV_X1 U7351 ( .A(n6254), .ZN(n6256) );
  NAND2_X1 U7352 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  NAND2_X1 U7353 ( .A1(n6258), .A2(n6257), .ZN(n6685) );
  INV_X1 U7354 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8691) );
  INV_X1 U7355 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6259) );
  MUX2_X1 U7356 ( .A(n8691), .B(n6259), .S(n7195), .Z(n6260) );
  INV_X1 U7357 ( .A(SI_30_), .ZN(n10014) );
  NAND2_X1 U7358 ( .A1(n6260), .A2(n10014), .ZN(n6686) );
  INV_X1 U7359 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U7360 ( .A1(n6261), .A2(SI_30_), .ZN(n6262) );
  NAND2_X1 U7361 ( .A1(n6686), .A2(n6262), .ZN(n6687) );
  XNOR2_X1 U7362 ( .A(n6685), .B(n6687), .ZN(n8451) );
  NAND2_X1 U7363 ( .A1(n8451), .A2(n4939), .ZN(n6264) );
  NAND2_X1 U7364 ( .A1(n6692), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7365 ( .A1(n6669), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6267) );
  INV_X1 U7366 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9855) );
  OR2_X1 U7367 ( .A1(n6670), .A2(n9855), .ZN(n6266) );
  INV_X1 U7368 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9938) );
  OR2_X1 U7369 ( .A1(n6673), .A2(n9938), .ZN(n6265) );
  AND3_X1 U7370 ( .A1(n6267), .A2(n6266), .A3(n6265), .ZN(n9616) );
  OR2_X1 U7371 ( .A1(n9557), .A2(n9616), .ZN(n6729) );
  NAND2_X1 U7372 ( .A1(n6669), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6270) );
  INV_X1 U7373 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9851) );
  OR2_X1 U7374 ( .A1(n6670), .A2(n9851), .ZN(n6269) );
  INV_X1 U7375 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9936) );
  OR2_X1 U7376 ( .A1(n6673), .A2(n9936), .ZN(n6268) );
  AND3_X1 U7377 ( .A1(n6270), .A2(n6269), .A3(n6268), .ZN(n9567) );
  AND2_X1 U7378 ( .A1(n9557), .A2(n9616), .ZN(n6770) );
  INV_X1 U7379 ( .A(n6770), .ZN(n6684) );
  NAND2_X1 U7380 ( .A1(n9557), .A2(n9567), .ZN(n6766) );
  NAND2_X1 U7381 ( .A1(n8216), .A2(n4938), .ZN(n6272) );
  INV_X2 U7382 ( .A(n6393), .ZN(n6692) );
  NAND2_X1 U7383 ( .A1(n6692), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7384 ( .A1(n6669), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6278) );
  INV_X1 U7385 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9893) );
  OR2_X1 U7386 ( .A1(n6670), .A2(n9893), .ZN(n6277) );
  INV_X1 U7387 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7388 ( .A1(n6283), .A2(n6273), .ZN(n6274) );
  NAND2_X1 U7389 ( .A1(n6615), .A2(n6274), .ZN(n9711) );
  OR2_X1 U7390 ( .A1(n6599), .A2(n9711), .ZN(n6276) );
  INV_X1 U7391 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9956) );
  OR2_X1 U7392 ( .A1(n6673), .A2(n9956), .ZN(n6275) );
  NAND2_X1 U7393 ( .A1(n9889), .A2(n9729), .ZN(n9608) );
  NAND2_X1 U7394 ( .A1(n8104), .A2(n4939), .ZN(n6280) );
  NAND2_X1 U7395 ( .A1(n6692), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7396 ( .A1(n6669), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6287) );
  INV_X1 U7397 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9899) );
  OR2_X1 U7398 ( .A1(n6670), .A2(n9899), .ZN(n6286) );
  INV_X1 U7399 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7400 ( .A1(n6293), .A2(n6281), .ZN(n6282) );
  NAND2_X1 U7401 ( .A1(n6283), .A2(n6282), .ZN(n9734) );
  OR2_X1 U7402 ( .A1(n6599), .A2(n9734), .ZN(n6285) );
  INV_X1 U7403 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9959) );
  OR2_X1 U7404 ( .A1(n6673), .A2(n9959), .ZN(n6284) );
  NAND4_X1 U7405 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n9747)
         );
  INV_X1 U7406 ( .A(n9747), .ZN(n9717) );
  NAND2_X1 U7407 ( .A1(n9736), .A2(n9717), .ZN(n9606) );
  AND2_X1 U7408 ( .A1(n9608), .A2(n9606), .ZN(n6735) );
  INV_X1 U7409 ( .A(n6735), .ZN(n6288) );
  OR2_X1 U7410 ( .A1(n9889), .A2(n9729), .ZN(n6706) );
  OR2_X1 U7411 ( .A1(n9736), .A2(n9717), .ZN(n6298) );
  NAND2_X1 U7412 ( .A1(n6706), .A2(n6298), .ZN(n6751) );
  MUX2_X1 U7413 ( .A(n6288), .B(n6751), .S(n4933), .Z(n6624) );
  INV_X2 U7414 ( .A(n4938), .ZN(n6625) );
  NAND2_X1 U7415 ( .A1(n6692), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7416 ( .A1(n6669), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6297) );
  INV_X1 U7417 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9904) );
  OR2_X1 U7418 ( .A1(n6670), .A2(n9904), .ZN(n6296) );
  INV_X1 U7419 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7420 ( .A1(n6597), .A2(n6291), .ZN(n6292) );
  NAND2_X1 U7421 ( .A1(n6293), .A2(n6292), .ZN(n9755) );
  OR2_X1 U7422 ( .A1(n6599), .A2(n9755), .ZN(n6295) );
  INV_X1 U7423 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9963) );
  OR2_X1 U7424 ( .A1(n6673), .A2(n9963), .ZN(n6294) );
  NAND2_X1 U7425 ( .A1(n9754), .A2(n9771), .ZN(n6733) );
  OR2_X1 U7426 ( .A1(n9754), .A2(n9771), .ZN(n6822) );
  AND2_X1 U7427 ( .A1(n6298), .A2(n6822), .ZN(n6299) );
  MUX2_X1 U7428 ( .A(n6733), .B(n6299), .S(n7553), .Z(n6610) );
  OR2_X1 U7429 ( .A1(n7442), .A2(n6625), .ZN(n6309) );
  INV_X1 U7430 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6302) );
  AND4_X1 U7431 ( .A1(n6301), .A2(n6471), .A3(n6447), .A4(n6302), .ZN(n6303)
         );
  AND2_X1 U7432 ( .A1(n6300), .A2(n6303), .ZN(n6511) );
  INV_X1 U7433 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6304) );
  INV_X1 U7434 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7435 ( .A1(n6497), .A2(n6305), .ZN(n6500) );
  NAND2_X1 U7436 ( .A1(n6500), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6546) );
  INV_X1 U7437 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7438 ( .A1(n6546), .A2(n6315), .ZN(n6317) );
  NAND2_X1 U7439 ( .A1(n6317), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6307) );
  INV_X1 U7440 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6306) );
  XNOR2_X1 U7441 ( .A(n6307), .B(n6306), .ZN(n9543) );
  INV_X1 U7442 ( .A(n9543), .ZN(n10388) );
  AOI22_X1 U7443 ( .A1(n6692), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4934), .B2(
        n10388), .ZN(n6308) );
  NAND2_X1 U7444 ( .A1(n6590), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6314) );
  INV_X2 U7445 ( .A(n6669), .ZN(n6570) );
  INV_X1 U7446 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10384) );
  OR2_X1 U7447 ( .A1(n6570), .A2(n10384), .ZN(n6313) );
  INV_X1 U7448 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10381) );
  OR2_X1 U7449 ( .A1(n6670), .A2(n10381), .ZN(n6312) );
  OR2_X1 U7450 ( .A1(n6321), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7451 ( .A1(n6554), .A2(n6310), .ZN(n9408) );
  OR2_X1 U7452 ( .A1(n6599), .A2(n9408), .ZN(n6311) );
  NAND4_X1 U7453 ( .A1(n6314), .A2(n6313), .A3(n6312), .A4(n6311), .ZN(n9829)
         );
  INV_X1 U7454 ( .A(n9829), .ZN(n8427) );
  NAND2_X1 U7455 ( .A1(n9412), .A2(n8427), .ZN(n6748) );
  OR2_X1 U7456 ( .A1(n7429), .A2(n6625), .ZN(n6319) );
  OR2_X1 U7457 ( .A1(n6546), .A2(n6315), .ZN(n6316) );
  AOI22_X1 U7458 ( .A1(n6692), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4935), .B2(
        n10364), .ZN(n6318) );
  NAND2_X1 U7459 ( .A1(n6590), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6325) );
  INV_X1 U7460 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8210) );
  OR2_X1 U7461 ( .A1(n6570), .A2(n8210), .ZN(n6324) );
  INV_X1 U7462 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8300) );
  OR2_X1 U7463 ( .A1(n6670), .A2(n8300), .ZN(n6323) );
  OR2_X1 U7464 ( .A1(n5559), .A2(n6321), .ZN(n8431) );
  OR2_X1 U7465 ( .A1(n6599), .A2(n8431), .ZN(n6322) );
  NAND2_X1 U7466 ( .A1(n8433), .A2(n8371), .ZN(n6747) );
  NAND2_X1 U7467 ( .A1(n6748), .A2(n6747), .ZN(n6785) );
  OR2_X1 U7468 ( .A1(n9412), .A2(n8427), .ZN(n6710) );
  OR2_X1 U7469 ( .A1(n8433), .A2(n8371), .ZN(n6810) );
  NAND2_X1 U7470 ( .A1(n6710), .A2(n6810), .ZN(n6326) );
  MUX2_X1 U7471 ( .A(n6785), .B(n6326), .S(n7553), .Z(n6327) );
  INV_X1 U7472 ( .A(n6327), .ZN(n6545) );
  INV_X1 U7473 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6328) );
  OR2_X1 U7474 ( .A1(n6367), .A2(n6328), .ZN(n6333) );
  INV_X1 U7475 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6329) );
  OR2_X1 U7476 ( .A1(n6673), .A2(n6329), .ZN(n6332) );
  INV_X1 U7477 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6330) );
  OR2_X1 U7478 ( .A1(n6350), .A2(n6330), .ZN(n6331) );
  INV_X1 U7479 ( .A(n8450), .ZN(n6335) );
  NAND2_X1 U7480 ( .A1(n4939), .A2(n6335), .ZN(n6339) );
  NAND2_X1 U7481 ( .A1(n6372), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6338) );
  OR2_X1 U7482 ( .A1(n6336), .A2(n9985), .ZN(n6388) );
  XNOR2_X1 U7483 ( .A(n6388), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U7484 ( .A1(n4935), .A2(n9469), .ZN(n6337) );
  AND3_X2 U7485 ( .A1(n6339), .A2(n6338), .A3(n6337), .ZN(n10735) );
  NAND2_X1 U7486 ( .A1(n6340), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6345) );
  INV_X1 U7487 ( .A(n6350), .ZN(n6341) );
  INV_X1 U7488 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U7489 ( .A1(n6348), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7490 ( .A1(n7195), .A2(SI_0_), .ZN(n6346) );
  XNOR2_X1 U7491 ( .A(n6346), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U7492 ( .A1(n7351), .A2(n7774), .ZN(n6714) );
  NAND2_X1 U7493 ( .A1(n6340), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7494 ( .A1(n6348), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6353) );
  INV_X1 U7495 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7772) );
  INV_X1 U7496 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6349) );
  OR2_X1 U7497 ( .A1(n6350), .A2(n6349), .ZN(n6351) );
  NAND2_X1 U7498 ( .A1(n6666), .A2(n7196), .ZN(n6360) );
  NAND2_X1 U7499 ( .A1(n6372), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7500 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10302), .ZN(n6355) );
  XNOR2_X1 U7501 ( .A(n6355), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9452) );
  INV_X1 U7502 ( .A(n9452), .ZN(n6356) );
  AND3_X2 U7503 ( .A1(n6360), .A2(n6359), .A3(n6358), .ZN(n10725) );
  NAND2_X1 U7504 ( .A1(n10228), .A2(n10725), .ZN(n6788) );
  NAND2_X1 U7505 ( .A1(n6714), .A2(n6788), .ZN(n6362) );
  INV_X1 U7506 ( .A(n10228), .ZN(n10705) );
  NAND2_X1 U7507 ( .A1(n10705), .A2(n7777), .ZN(n6361) );
  NAND2_X1 U7508 ( .A1(n6362), .A2(n6361), .ZN(n10224) );
  INV_X1 U7509 ( .A(n10224), .ZN(n6365) );
  INV_X1 U7510 ( .A(n10735), .ZN(n9371) );
  NAND2_X1 U7511 ( .A1(n7767), .A2(n9371), .ZN(n6364) );
  NAND2_X1 U7512 ( .A1(n6669), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6371) );
  INV_X1 U7513 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6366) );
  OR2_X1 U7514 ( .A1(n6673), .A2(n6366), .ZN(n6370) );
  INV_X1 U7515 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9463) );
  OR2_X1 U7516 ( .A1(n6599), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6368) );
  AND4_X2 U7517 ( .A1(n6371), .A2(n6370), .A3(n6369), .A4(n6368), .ZN(n7560)
         );
  NAND2_X1 U7518 ( .A1(n6372), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6377) );
  INV_X1 U7519 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7520 ( .A1(n6388), .A2(n6373), .ZN(n6374) );
  NAND2_X1 U7521 ( .A1(n6374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6375) );
  XNOR2_X1 U7522 ( .A(n6375), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U7523 ( .A1(n4935), .A2(n9486), .ZN(n6376) );
  NAND2_X1 U7524 ( .A1(n7560), .A2(n7820), .ZN(n6716) );
  INV_X1 U7525 ( .A(n6716), .ZN(n6378) );
  OR2_X1 U7526 ( .A1(n7811), .A2(n6378), .ZN(n7837) );
  NAND2_X1 U7527 ( .A1(n6669), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6385) );
  INV_X1 U7528 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6379) );
  OR2_X1 U7529 ( .A1(n6673), .A2(n6379), .ZN(n6384) );
  INV_X1 U7530 ( .A(n6401), .ZN(n6382) );
  INV_X1 U7531 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7819) );
  INV_X1 U7532 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U7533 ( .A1(n7819), .A2(n6380), .ZN(n6381) );
  NAND2_X1 U7534 ( .A1(n6382), .A2(n6381), .ZN(n7831) );
  INV_X1 U7535 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6383) );
  NOR2_X1 U7536 ( .A1(n7202), .A2(n6625), .ZN(n6395) );
  INV_X1 U7537 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7203) );
  OR2_X1 U7538 ( .A1(n6386), .A2(n9985), .ZN(n6387) );
  AND2_X1 U7539 ( .A1(n6388), .A2(n6387), .ZN(n6390) );
  INV_X1 U7540 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7541 ( .A1(n6390), .A2(n6389), .ZN(n6407) );
  INV_X1 U7542 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U7543 ( .A1(n6391), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7544 ( .A1(n6407), .A2(n6392), .ZN(n9489) );
  AND2_X1 U7545 ( .A1(n6736), .A2(n6716), .ZN(n6396) );
  MUX2_X1 U7546 ( .A(n7837), .B(n6396), .S(n4933), .Z(n6400) );
  INV_X1 U7547 ( .A(n7834), .ZN(n10757) );
  NAND2_X1 U7548 ( .A1(n9426), .A2(n10757), .ZN(n6715) );
  INV_X1 U7549 ( .A(n6715), .ZN(n6399) );
  AND2_X1 U7550 ( .A1(n7836), .A2(n6715), .ZN(n6791) );
  NAND2_X1 U7551 ( .A1(n7811), .A2(n6791), .ZN(n6397) );
  MUX2_X1 U7552 ( .A(n6791), .B(n6397), .S(n4933), .Z(n6398) );
  NAND2_X1 U7553 ( .A1(n6341), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6406) );
  INV_X1 U7554 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7699) );
  OR2_X1 U7555 ( .A1(n6570), .A2(n7699), .ZN(n6405) );
  OAI21_X1 U7556 ( .B1(n6401), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6416), .ZN(
        n7703) );
  OR2_X1 U7557 ( .A1(n6599), .A2(n7703), .ZN(n6404) );
  INV_X1 U7558 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6402) );
  OR2_X1 U7559 ( .A1(n6673), .A2(n6402), .ZN(n6403) );
  OR2_X1 U7560 ( .A1(n7208), .A2(n6625), .ZN(n6410) );
  NAND2_X1 U7561 ( .A1(n6407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U7562 ( .A(n6408), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U7563 ( .A1(n6692), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4935), .B2(
        n9506), .ZN(n6409) );
  NAND2_X1 U7564 ( .A1(n7785), .A2(n7684), .ZN(n6738) );
  NAND2_X1 U7565 ( .A1(n7210), .A2(n4938), .ZN(n6414) );
  NAND2_X1 U7566 ( .A1(n6411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6412) );
  XNOR2_X1 U7567 ( .A(n6412), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U7568 ( .A1(n6692), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4935), .B2(
        n10313), .ZN(n6413) );
  NAND2_X1 U7569 ( .A1(n6414), .A2(n6413), .ZN(n7853) );
  NAND2_X1 U7570 ( .A1(n6341), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6422) );
  INV_X1 U7571 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7846) );
  OR2_X1 U7572 ( .A1(n6570), .A2(n7846), .ZN(n6421) );
  AND2_X1 U7573 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  OR2_X1 U7574 ( .A1(n6417), .A2(n6429), .ZN(n7742) );
  OR2_X1 U7575 ( .A1(n6599), .A2(n7742), .ZN(n6420) );
  INV_X1 U7576 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6418) );
  OR2_X1 U7577 ( .A1(n6673), .A2(n6418), .ZN(n6419) );
  OR2_X1 U7578 ( .A1(n7853), .A2(n7800), .ZN(n7794) );
  INV_X2 U7579 ( .A(n7684), .ZN(n7784) );
  INV_X1 U7580 ( .A(n6795), .ZN(n6460) );
  NAND2_X1 U7581 ( .A1(n7215), .A2(n4938), .ZN(n6428) );
  NAND2_X1 U7582 ( .A1(n6423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6424) );
  MUX2_X1 U7583 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6424), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n6426) );
  INV_X1 U7584 ( .A(n6300), .ZN(n6425) );
  AOI22_X1 U7585 ( .A1(n6692), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4934), .B2(
        n10325), .ZN(n6427) );
  NAND2_X1 U7586 ( .A1(n6590), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6435) );
  INV_X1 U7587 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9838) );
  OR2_X1 U7588 ( .A1(n6570), .A2(n9838), .ZN(n6434) );
  OR2_X1 U7589 ( .A1(n6429), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7590 ( .A1(n6440), .A2(n6430), .ZN(n9837) );
  OR2_X1 U7591 ( .A1(n6599), .A2(n9837), .ZN(n6433) );
  INV_X1 U7592 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6431) );
  OR2_X1 U7593 ( .A1(n6670), .A2(n6431), .ZN(n6432) );
  NAND2_X1 U7594 ( .A1(n9841), .A2(n7752), .ZN(n7858) );
  NAND2_X1 U7595 ( .A1(n7853), .A2(n7800), .ZN(n7789) );
  NAND2_X1 U7596 ( .A1(n7220), .A2(n4938), .ZN(n6437) );
  OR2_X1 U7597 ( .A1(n6300), .A2(n9985), .ZN(n6448) );
  XNOR2_X1 U7598 ( .A(n6448), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U7599 ( .A1(n6692), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4934), .B2(
        n10336), .ZN(n6436) );
  NAND2_X1 U7600 ( .A1(n6590), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6445) );
  INV_X1 U7601 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6438) );
  OR2_X1 U7602 ( .A1(n6670), .A2(n6438), .ZN(n6444) );
  INV_X1 U7603 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7989) );
  OR2_X1 U7604 ( .A1(n6570), .A2(n7989), .ZN(n6443) );
  NAND2_X1 U7605 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U7606 ( .A1(n6452), .A2(n6441), .ZN(n8058) );
  OR2_X1 U7607 ( .A1(n6599), .A2(n8058), .ZN(n6442) );
  OR2_X1 U7608 ( .A1(n8060), .A2(n8151), .ZN(n6465) );
  NAND2_X1 U7609 ( .A1(n8060), .A2(n8151), .ZN(n7860) );
  NAND2_X1 U7610 ( .A1(n6465), .A2(n7860), .ZN(n7984) );
  INV_X1 U7611 ( .A(n7984), .ZN(n7994) );
  OR2_X1 U7612 ( .A1(n9841), .A2(n7752), .ZN(n7791) );
  NAND3_X1 U7613 ( .A1(n6446), .A2(n7994), .A3(n7791), .ZN(n6459) );
  NAND2_X1 U7614 ( .A1(n7243), .A2(n4939), .ZN(n6451) );
  NAND2_X1 U7615 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND2_X1 U7616 ( .A1(n6449), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6469) );
  XNOR2_X1 U7617 ( .A(n6469), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9537) );
  AOI22_X1 U7618 ( .A1(n6692), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4934), .B2(
        n9537), .ZN(n6450) );
  NAND2_X1 U7619 ( .A1(n6590), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6458) );
  INV_X1 U7620 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7873) );
  OR2_X1 U7621 ( .A1(n6570), .A2(n7873), .ZN(n6457) );
  AND2_X1 U7622 ( .A1(n6452), .A2(n8149), .ZN(n6453) );
  OR2_X1 U7623 ( .A1(n6453), .A2(n6475), .ZN(n8148) );
  OR2_X1 U7624 ( .A1(n6599), .A2(n8148), .ZN(n6456) );
  INV_X1 U7625 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6454) );
  OR2_X1 U7626 ( .A1(n6670), .A2(n6454), .ZN(n6455) );
  NAND2_X1 U7627 ( .A1(n8142), .A2(n8138), .ZN(n7861) );
  NAND3_X1 U7628 ( .A1(n6459), .A2(n7861), .A3(n7860), .ZN(n6468) );
  OAI21_X1 U7629 ( .B1(n6460), .B2(n6736), .A(n7789), .ZN(n6462) );
  NAND2_X1 U7630 ( .A1(n7791), .A2(n7794), .ZN(n6712) );
  INV_X1 U7631 ( .A(n6712), .ZN(n6461) );
  OAI21_X1 U7632 ( .B1(n6463), .B2(n6462), .A(n6461), .ZN(n6464) );
  NAND3_X1 U7633 ( .A1(n6464), .A2(n7994), .A3(n7858), .ZN(n6466) );
  OR2_X1 U7634 ( .A1(n8142), .A2(n8138), .ZN(n7862) );
  NAND2_X1 U7635 ( .A1(n7862), .A2(n6465), .ZN(n6713) );
  INV_X1 U7636 ( .A(n6713), .ZN(n6741) );
  NAND2_X1 U7637 ( .A1(n6466), .A2(n6741), .ZN(n6467) );
  MUX2_X1 U7638 ( .A(n6468), .B(n6467), .S(n7553), .Z(n6526) );
  INV_X1 U7639 ( .A(n6526), .ZN(n6496) );
  NAND2_X1 U7640 ( .A1(n6469), .A2(n6301), .ZN(n6470) );
  NAND2_X1 U7641 ( .A1(n6470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U7642 ( .A1(n6472), .A2(n6471), .ZN(n6481) );
  OR2_X1 U7643 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  AOI22_X1 U7644 ( .A1(n6692), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4935), .B2(
        n10476), .ZN(n6474) );
  NAND2_X1 U7645 ( .A1(n6590), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6480) );
  INV_X1 U7646 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7888) );
  OR2_X1 U7647 ( .A1(n6570), .A2(n7888), .ZN(n6479) );
  NOR2_X1 U7648 ( .A1(n6475), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6476) );
  OR2_X1 U7649 ( .A1(n6485), .A2(n6476), .ZN(n8329) );
  OR2_X1 U7650 ( .A1(n6599), .A2(n8329), .ZN(n6478) );
  INV_X1 U7651 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9524) );
  OR2_X1 U7652 ( .A1(n6670), .A2(n9524), .ZN(n6477) );
  NAND2_X1 U7653 ( .A1(n8331), .A2(n8250), .ZN(n6744) );
  NAND2_X1 U7654 ( .A1(n7266), .A2(n4939), .ZN(n6484) );
  NAND2_X1 U7655 ( .A1(n6481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6482) );
  XNOR2_X1 U7656 ( .A(n6482), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U7657 ( .A1(n6692), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4934), .B2(
        n10360), .ZN(n6483) );
  NAND2_X1 U7658 ( .A1(n6341), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6491) );
  INV_X1 U7659 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8020) );
  OR2_X1 U7660 ( .A1(n6570), .A2(n8020), .ZN(n6490) );
  OR2_X1 U7661 ( .A1(n6485), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7662 ( .A1(n6516), .A2(n6486), .ZN(n8388) );
  OR2_X1 U7663 ( .A1(n6599), .A2(n8388), .ZN(n6489) );
  INV_X1 U7664 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6487) );
  OR2_X1 U7665 ( .A1(n6673), .A2(n6487), .ZN(n6488) );
  NAND4_X1 U7666 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n9421)
         );
  INV_X1 U7667 ( .A(n9421), .ZN(n8324) );
  NAND2_X1 U7668 ( .A1(n8390), .A2(n8324), .ZN(n7968) );
  NAND2_X1 U7669 ( .A1(n6744), .A2(n7861), .ZN(n6492) );
  NAND2_X1 U7670 ( .A1(n6492), .A2(n6801), .ZN(n6493) );
  NAND2_X1 U7671 ( .A1(n7968), .A2(n6493), .ZN(n6800) );
  INV_X1 U7672 ( .A(n6744), .ZN(n6494) );
  OR2_X1 U7673 ( .A1(n8390), .A2(n8324), .ZN(n6711) );
  OAI211_X1 U7674 ( .C1(n6494), .C2(n7862), .A(n6711), .B(n6801), .ZN(n6495)
         );
  MUX2_X1 U7675 ( .A(n6800), .B(n6495), .S(n4933), .Z(n6523) );
  AOI21_X1 U7676 ( .B1(n6496), .B2(n6744), .A(n6523), .ZN(n6543) );
  OR2_X1 U7677 ( .A1(n7310), .A2(n6625), .ZN(n6503) );
  NOR2_X1 U7678 ( .A1(n6497), .A2(n9985), .ZN(n6498) );
  MUX2_X1 U7679 ( .A(n9985), .B(n6498), .S(P1_IR_REG_13__SCAN_IN), .Z(n6499)
         );
  INV_X1 U7680 ( .A(n6499), .ZN(n6501) );
  AOI22_X1 U7681 ( .A1(n6692), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4934), .B2(
        n10433), .ZN(n6502) );
  AND2_X2 U7682 ( .A1(n6503), .A2(n6502), .ZN(n10815) );
  NAND2_X1 U7683 ( .A1(n6590), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6510) );
  INV_X1 U7684 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8079) );
  OR2_X1 U7685 ( .A1(n6570), .A2(n8079), .ZN(n6509) );
  NAND2_X1 U7686 ( .A1(n6518), .A2(n6504), .ZN(n6505) );
  NAND2_X1 U7687 ( .A1(n6506), .A2(n6505), .ZN(n8374) );
  OR2_X1 U7688 ( .A1(n6599), .A2(n8374), .ZN(n6508) );
  INV_X1 U7689 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9521) );
  OR2_X1 U7690 ( .A1(n6670), .A2(n9521), .ZN(n6507) );
  NAND4_X1 U7691 ( .A1(n6510), .A2(n6509), .A3(n6508), .A4(n6507), .ZN(n9419)
         );
  INV_X1 U7692 ( .A(n9419), .ZN(n8370) );
  NAND2_X1 U7693 ( .A1(n8376), .A2(n8370), .ZN(n6805) );
  OR2_X1 U7694 ( .A1(n7276), .A2(n6625), .ZN(n6514) );
  OR2_X1 U7695 ( .A1(n6511), .A2(n9985), .ZN(n6512) );
  XNOR2_X1 U7696 ( .A(n6512), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U7697 ( .A1(n6692), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4935), .B2(
        n10449), .ZN(n6513) );
  NAND2_X1 U7698 ( .A1(n6590), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6522) );
  INV_X1 U7699 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7976) );
  OR2_X1 U7700 ( .A1(n6570), .A2(n7976), .ZN(n6521) );
  NAND2_X1 U7701 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  NAND2_X1 U7702 ( .A1(n6518), .A2(n6517), .ZN(n8266) );
  OR2_X1 U7703 ( .A1(n6599), .A2(n8266), .ZN(n6520) );
  INV_X1 U7704 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9522) );
  OR2_X1 U7705 ( .A1(n6670), .A2(n9522), .ZN(n6519) );
  NAND4_X1 U7706 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n9420)
         );
  NAND2_X1 U7707 ( .A1(n8268), .A2(n8385), .ZN(n6804) );
  NAND4_X1 U7708 ( .A1(n6805), .A2(n4933), .A3(n7968), .A4(n6804), .ZN(n6542)
         );
  INV_X1 U7709 ( .A(n6801), .ZN(n6525) );
  INV_X1 U7710 ( .A(n6523), .ZN(n6524) );
  OAI21_X1 U7711 ( .B1(n6526), .B2(n6525), .A(n6524), .ZN(n6527) );
  OR2_X1 U7712 ( .A1(n8268), .A2(n8385), .ZN(n6745) );
  AND2_X1 U7713 ( .A1(n6745), .A2(n6711), .ZN(n6803) );
  NAND2_X1 U7714 ( .A1(n10815), .A2(n9419), .ZN(n6809) );
  NAND4_X1 U7715 ( .A1(n6527), .A2(n6803), .A3(n6809), .A4(n7553), .ZN(n6541)
         );
  NOR2_X1 U7716 ( .A1(n9420), .A2(n4933), .ZN(n6529) );
  NAND2_X1 U7717 ( .A1(n8370), .A2(n7553), .ZN(n6533) );
  INV_X1 U7718 ( .A(n6533), .ZN(n6528) );
  AOI21_X1 U7719 ( .B1(n8268), .B2(n6529), .A(n6528), .ZN(n6538) );
  NAND2_X1 U7720 ( .A1(n9420), .A2(n4933), .ZN(n6530) );
  NAND2_X1 U7721 ( .A1(n9419), .A2(n4933), .ZN(n6532) );
  OAI21_X1 U7722 ( .B1(n8268), .B2(n6530), .A(n6532), .ZN(n6531) );
  NAND2_X1 U7723 ( .A1(n10815), .A2(n6531), .ZN(n6537) );
  NOR2_X1 U7724 ( .A1(n6532), .A2(n8385), .ZN(n6535) );
  OAI21_X1 U7725 ( .B1(n9420), .B2(n6533), .A(n8268), .ZN(n6534) );
  OAI21_X1 U7726 ( .B1(n6535), .B2(n8268), .A(n6534), .ZN(n6536) );
  OAI211_X1 U7727 ( .C1(n10815), .C2(n6538), .A(n6537), .B(n6536), .ZN(n6539)
         );
  NOR2_X1 U7728 ( .A1(n8197), .A2(n6539), .ZN(n6540) );
  OAI211_X1 U7729 ( .C1(n6543), .C2(n6542), .A(n6541), .B(n6540), .ZN(n6544)
         );
  NAND2_X1 U7730 ( .A1(n6545), .A2(n6544), .ZN(n6562) );
  NAND2_X1 U7731 ( .A1(n7510), .A2(n4938), .ZN(n6551) );
  OAI21_X1 U7732 ( .B1(n6547), .B2(n9985), .A(n6546), .ZN(n6548) );
  OR2_X1 U7733 ( .A1(n6548), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7734 ( .A1(n6548), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6549) );
  AOI22_X1 U7735 ( .A1(n6692), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4934), .B2(
        n9546), .ZN(n6550) );
  NAND2_X1 U7736 ( .A1(n6590), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6559) );
  INV_X1 U7737 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6552) );
  OR2_X1 U7738 ( .A1(n6570), .A2(n6552), .ZN(n6558) );
  INV_X1 U7739 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9520) );
  OR2_X1 U7740 ( .A1(n6670), .A2(n9520), .ZN(n6557) );
  NAND2_X1 U7741 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NAND2_X1 U7742 ( .A1(n6568), .A2(n6555), .ZN(n9821) );
  OR2_X1 U7743 ( .A1(n6599), .A2(n9821), .ZN(n6556) );
  OR2_X1 U7744 ( .A1(n9930), .A2(n9403), .ZN(n6709) );
  AND2_X1 U7745 ( .A1(n6709), .A2(n6710), .ZN(n6811) );
  NAND2_X1 U7746 ( .A1(n9930), .A2(n9403), .ZN(n6749) );
  AND2_X1 U7747 ( .A1(n6749), .A2(n6748), .ZN(n6561) );
  INV_X1 U7748 ( .A(n6709), .ZN(n6560) );
  NAND2_X1 U7749 ( .A1(n7615), .A2(n4939), .ZN(n6566) );
  NAND2_X1 U7750 ( .A1(n6563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6564) );
  XNOR2_X1 U7751 ( .A(n6564), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U7752 ( .A1(n6692), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4935), .B2(
        n10399), .ZN(n6565) );
  AND2_X1 U7753 ( .A1(n6568), .A2(n6567), .ZN(n6569) );
  OR2_X1 U7754 ( .A1(n6569), .A2(n6581), .ZN(n9335) );
  INV_X1 U7755 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9926) );
  OR2_X1 U7756 ( .A1(n6670), .A2(n9926), .ZN(n6572) );
  INV_X1 U7757 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8313) );
  OR2_X1 U7758 ( .A1(n6570), .A2(n8313), .ZN(n6571) );
  AND2_X1 U7759 ( .A1(n6572), .A2(n6571), .ZN(n6574) );
  NAND2_X1 U7760 ( .A1(n6590), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6573) );
  OAI211_X1 U7761 ( .C1(n9335), .C2(n6599), .A(n6574), .B(n6573), .ZN(n9830)
         );
  INV_X1 U7762 ( .A(n9830), .ZN(n9324) );
  XNOR2_X1 U7763 ( .A(n9577), .B(n9324), .ZN(n9575) );
  INV_X1 U7764 ( .A(n9575), .ZN(n8308) );
  OR2_X1 U7765 ( .A1(n7666), .A2(n6625), .ZN(n6580) );
  INV_X1 U7766 ( .A(n6575), .ZN(n6576) );
  NAND2_X1 U7767 ( .A1(n6576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6577) );
  MUX2_X1 U7768 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6577), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n6578) );
  AND2_X1 U7769 ( .A1(n6578), .A2(n4964), .ZN(n10413) );
  AOI22_X1 U7770 ( .A1(n6692), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4935), .B2(
        n10413), .ZN(n6579) );
  NOR2_X1 U7771 ( .A1(n6581), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6582) );
  OR2_X1 U7772 ( .A1(n6587), .A2(n6582), .ZN(n9800) );
  AOI22_X1 U7773 ( .A1(n6341), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6669), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U7774 ( .A1(n6590), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6583) );
  OAI211_X1 U7775 ( .C1(n9800), .C2(n6599), .A(n6584), .B(n6583), .ZN(n9781)
         );
  INV_X1 U7776 ( .A(n9781), .ZN(n9332) );
  OR2_X1 U7777 ( .A1(n9919), .A2(n9332), .ZN(n6708) );
  OR2_X1 U7778 ( .A1(n9577), .A2(n9324), .ZN(n6815) );
  NAND2_X1 U7779 ( .A1(n7780), .A2(n4938), .ZN(n6586) );
  AOI22_X1 U7780 ( .A1(n6692), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10222), 
        .B2(n4935), .ZN(n6585) );
  OR2_X1 U7781 ( .A1(n6587), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6589) );
  AND2_X1 U7782 ( .A1(n6589), .A2(n6588), .ZN(n9792) );
  NAND2_X1 U7783 ( .A1(n9792), .A2(n5089), .ZN(n6593) );
  AOI22_X1 U7784 ( .A1(n6341), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6669), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U7785 ( .A1(n6590), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U7786 ( .A1(n9791), .A2(n9769), .ZN(n6821) );
  NAND2_X1 U7787 ( .A1(n9919), .A2(n9332), .ZN(n6750) );
  NAND3_X1 U7788 ( .A1(n6594), .A2(n6821), .A3(n6750), .ZN(n6604) );
  NAND2_X1 U7789 ( .A1(n7956), .A2(n4939), .ZN(n6596) );
  NAND2_X1 U7790 ( .A1(n6692), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U7791 ( .A1(n6669), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6603) );
  INV_X1 U7792 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9967) );
  OR2_X1 U7793 ( .A1(n6673), .A2(n9967), .ZN(n6602) );
  OAI21_X1 U7794 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n6598), .A(n6597), .ZN(
        n9763) );
  OR2_X1 U7795 ( .A1(n6599), .A2(n9763), .ZN(n6601) );
  INV_X1 U7796 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9910) );
  OR2_X1 U7797 ( .A1(n6670), .A2(n9910), .ZN(n6600) );
  OR2_X1 U7798 ( .A1(n9906), .A2(n9281), .ZN(n6823) );
  OR2_X1 U7799 ( .A1(n9791), .A2(n9769), .ZN(n6707) );
  NAND3_X1 U7800 ( .A1(n6604), .A2(n6823), .A3(n6707), .ZN(n6605) );
  NAND2_X1 U7801 ( .A1(n9906), .A2(n9281), .ZN(n9743) );
  AND2_X1 U7802 ( .A1(n6707), .A2(n6708), .ZN(n6817) );
  NAND2_X1 U7803 ( .A1(n9577), .A2(n9324), .ZN(n9806) );
  AND2_X1 U7804 ( .A1(n6750), .A2(n9806), .ZN(n6820) );
  NAND2_X1 U7805 ( .A1(n6606), .A2(n6820), .ZN(n6607) );
  NAND2_X1 U7806 ( .A1(n6817), .A2(n6607), .ZN(n6608) );
  NAND3_X1 U7807 ( .A1(n6608), .A2(n9743), .A3(n6821), .ZN(n6609) );
  NAND2_X1 U7808 ( .A1(n6822), .A2(n6733), .ZN(n9751) );
  NAND2_X1 U7809 ( .A1(n8271), .A2(n4938), .ZN(n6612) );
  NAND2_X1 U7810 ( .A1(n6692), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7811 ( .A1(n6669), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6621) );
  INV_X1 U7812 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6613) );
  OR2_X1 U7813 ( .A1(n6670), .A2(n6613), .ZN(n6620) );
  INV_X1 U7814 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U7815 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  NAND2_X1 U7816 ( .A1(n6630), .A2(n6616), .ZN(n9696) );
  OR2_X1 U7817 ( .A1(n6599), .A2(n9696), .ZN(n6619) );
  INV_X1 U7818 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6617) );
  OR2_X1 U7819 ( .A1(n6673), .A2(n6617), .ZN(n6618) );
  NAND4_X1 U7820 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n9679)
         );
  INV_X1 U7821 ( .A(n9679), .ZN(n9718) );
  OR2_X1 U7822 ( .A1(n9885), .A2(n9718), .ZN(n9609) );
  NAND2_X1 U7823 ( .A1(n9885), .A2(n9718), .ZN(n6753) );
  NAND2_X1 U7824 ( .A1(n9609), .A2(n6753), .ZN(n9700) );
  MUX2_X1 U7825 ( .A(n9608), .B(n6706), .S(n7553), .Z(n6622) );
  OAI211_X1 U7826 ( .C1(n6624), .C2(n6623), .A(n9694), .B(n6622), .ZN(n6637)
         );
  NAND2_X1 U7827 ( .A1(n6692), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U7828 ( .A1(n6669), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6636) );
  INV_X1 U7829 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6628) );
  OR2_X1 U7830 ( .A1(n6670), .A2(n6628), .ZN(n6635) );
  INV_X1 U7831 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U7832 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  NAND2_X1 U7833 ( .A1(n6645), .A2(n6631), .ZN(n9316) );
  OR2_X1 U7834 ( .A1(n6599), .A2(n9316), .ZN(n6634) );
  INV_X1 U7835 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6632) );
  OR2_X1 U7836 ( .A1(n6673), .A2(n6632), .ZN(n6633) );
  OR2_X1 U7837 ( .A1(n9879), .A2(n9702), .ZN(n6755) );
  NAND2_X1 U7838 ( .A1(n9879), .A2(n9702), .ZN(n9610) );
  AND3_X1 U7839 ( .A1(n6637), .A2(n9689), .A3(n9609), .ZN(n6641) );
  NAND2_X1 U7840 ( .A1(n6637), .A2(n6753), .ZN(n6639) );
  INV_X1 U7841 ( .A(n9610), .ZN(n6638) );
  AOI21_X1 U7842 ( .B1(n6639), .B2(n6755), .A(n6638), .ZN(n6640) );
  MUX2_X1 U7843 ( .A(n6641), .B(n6640), .S(n7553), .Z(n6654) );
  NAND2_X1 U7844 ( .A1(n8416), .A2(n4939), .ZN(n6643) );
  NAND2_X1 U7845 ( .A1(n6692), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U7846 ( .A1(n6669), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6650) );
  INV_X1 U7847 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9876) );
  OR2_X1 U7848 ( .A1(n6670), .A2(n9876), .ZN(n6649) );
  INV_X1 U7849 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U7850 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  NAND2_X1 U7851 ( .A1(n6660), .A2(n6646), .ZN(n9392) );
  INV_X1 U7852 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9950) );
  OR2_X1 U7853 ( .A1(n6673), .A2(n9950), .ZN(n6647) );
  NAND4_X1 U7854 ( .A1(n6650), .A2(n6649), .A3(n6648), .A4(n6647), .ZN(n9680)
         );
  INV_X1 U7855 ( .A(n9680), .ZN(n6651) );
  OR2_X1 U7856 ( .A1(n9672), .A2(n6651), .ZN(n6760) );
  INV_X1 U7857 ( .A(n6760), .ZN(n6653) );
  NAND2_X1 U7858 ( .A1(n9672), .A2(n6651), .ZN(n9611) );
  AND2_X1 U7859 ( .A1(n9611), .A2(n7553), .ZN(n6652) );
  OAI22_X1 U7860 ( .A1(n6654), .A2(n6653), .B1(n9665), .B2(n6652), .ZN(n6656)
         );
  NAND2_X1 U7861 ( .A1(n9611), .A2(n9610), .ZN(n6757) );
  NAND3_X1 U7862 ( .A1(n6757), .A2(n4933), .A3(n6760), .ZN(n6655) );
  NAND2_X1 U7863 ( .A1(n8438), .A2(n4938), .ZN(n6658) );
  NAND2_X1 U7864 ( .A1(n6692), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U7865 ( .A1(n6669), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6665) );
  INV_X1 U7866 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9946) );
  OR2_X1 U7867 ( .A1(n6673), .A2(n9946), .ZN(n6664) );
  INV_X1 U7868 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U7869 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  NAND2_X1 U7870 ( .A1(n6672), .A2(n6661), .ZN(n8776) );
  OR2_X1 U7871 ( .A1(n6367), .A2(n8776), .ZN(n6663) );
  INV_X1 U7872 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9870) );
  OR2_X1 U7873 ( .A1(n6670), .A2(n9870), .ZN(n6662) );
  OR2_X1 U7874 ( .A1(n9654), .A2(n9666), .ZN(n6761) );
  NAND2_X1 U7875 ( .A1(n9654), .A2(n9666), .ZN(n9612) );
  NAND2_X1 U7876 ( .A1(n9996), .A2(n4939), .ZN(n6668) );
  NAND2_X1 U7877 ( .A1(n6692), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U7878 ( .A1(n6669), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6677) );
  INV_X1 U7879 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9865) );
  OR2_X1 U7880 ( .A1(n6670), .A2(n9865), .ZN(n6676) );
  INV_X1 U7881 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6671) );
  XNOR2_X1 U7882 ( .A(n6672), .B(n6671), .ZN(n9627) );
  OR2_X1 U7883 ( .A1(n6367), .A2(n9627), .ZN(n6675) );
  INV_X1 U7884 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9943) );
  OR2_X1 U7885 ( .A1(n6673), .A2(n9943), .ZN(n6674) );
  OR2_X1 U7886 ( .A1(n9638), .A2(n9618), .ZN(n6758) );
  NAND2_X1 U7887 ( .A1(n9638), .A2(n9618), .ZN(n9613) );
  MUX2_X1 U7888 ( .A(n9612), .B(n6761), .S(n7553), .Z(n6678) );
  INV_X1 U7889 ( .A(n6764), .ZN(n6679) );
  MUX2_X1 U7890 ( .A(n9613), .B(n6758), .S(n4933), .Z(n6680) );
  NAND4_X1 U7891 ( .A1(n6768), .A2(n6684), .A3(n6766), .A4(n6683), .ZN(n6700)
         );
  OAI21_X1 U7892 ( .B1(n6685), .B2(n6687), .A(n6686), .ZN(n6691) );
  MUX2_X1 U7893 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7195), .Z(n6689) );
  INV_X1 U7894 ( .A(SI_31_), .ZN(n6688) );
  XNOR2_X1 U7895 ( .A(n6689), .B(n6688), .ZN(n6690) );
  NAND2_X1 U7896 ( .A1(n9257), .A2(n4938), .ZN(n6694) );
  NAND2_X1 U7897 ( .A1(n6692), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6693) );
  NOR2_X1 U7898 ( .A1(n9568), .A2(n9567), .ZN(n6771) );
  INV_X1 U7899 ( .A(n6771), .ZN(n6695) );
  AND2_X1 U7900 ( .A1(n9568), .A2(n9567), .ZN(n6772) );
  INV_X1 U7901 ( .A(n6772), .ZN(n6836) );
  NAND2_X1 U7902 ( .A1(n6695), .A2(n6836), .ZN(n6731) );
  INV_X1 U7903 ( .A(n6731), .ZN(n6699) );
  INV_X1 U7904 ( .A(n9567), .ZN(n7232) );
  INV_X1 U7905 ( .A(n9616), .ZN(n9416) );
  NAND2_X1 U7906 ( .A1(n7232), .A2(n9416), .ZN(n6696) );
  NAND2_X1 U7907 ( .A1(n9557), .A2(n6696), .ZN(n6697) );
  MUX2_X1 U7908 ( .A(n6697), .B(n6768), .S(n4933), .Z(n6698) );
  AOI21_X1 U7909 ( .B1(n6772), .B2(n7553), .A(n8028), .ZN(n6705) );
  INV_X1 U7910 ( .A(n9665), .ZN(n9661) );
  INV_X1 U7911 ( .A(n9787), .ZN(n6725) );
  NAND2_X1 U7912 ( .A1(n6709), .A2(n6749), .ZN(n9815) );
  INV_X1 U7913 ( .A(n9815), .ZN(n9828) );
  INV_X1 U7914 ( .A(n8076), .ZN(n8068) );
  INV_X1 U7915 ( .A(n8014), .ZN(n6722) );
  NAND2_X1 U7916 ( .A1(n6801), .A2(n6744), .ZN(n7886) );
  INV_X1 U7917 ( .A(n7886), .ZN(n7880) );
  INV_X1 U7918 ( .A(n7861), .ZN(n6719) );
  INV_X1 U7919 ( .A(n6714), .ZN(n7765) );
  NAND2_X1 U7920 ( .A1(n7351), .A2(n7774), .ZN(n6789) );
  NAND2_X1 U7921 ( .A1(n7765), .A2(n6789), .ZN(n10700) );
  NAND2_X1 U7922 ( .A1(n6736), .A2(n6715), .ZN(n7838) );
  NOR4_X1 U7923 ( .A1(n10700), .A2(n7838), .A3(n7809), .A4(n6848), .ZN(n6717)
         );
  AND2_X2 U7924 ( .A1(n6738), .A2(n6795), .ZN(n7788) );
  INV_X1 U7925 ( .A(n7557), .ZN(n10223) );
  XNOR2_X2 U7926 ( .A(n10228), .B(n10725), .ZN(n7766) );
  INV_X1 U7927 ( .A(n7766), .ZN(n7762) );
  NAND4_X1 U7928 ( .A1(n6717), .A2(n7788), .A3(n10223), .A4(n7762), .ZN(n6718)
         );
  INV_X1 U7929 ( .A(n7789), .ZN(n6794) );
  NAND2_X1 U7930 ( .A1(n7860), .A2(n7858), .ZN(n6740) );
  NOR4_X1 U7931 ( .A1(n6719), .A2(n6718), .A3(n6794), .A4(n6740), .ZN(n6720)
         );
  NAND4_X1 U7932 ( .A1(n7880), .A2(n6786), .A3(n7967), .A4(n6720), .ZN(n6721)
         );
  NOR4_X1 U7933 ( .A1(n8197), .A2(n8068), .A3(n6722), .A4(n6721), .ZN(n6723)
         );
  NAND4_X1 U7934 ( .A1(n9804), .A2(n9828), .A3(n8173), .A4(n6723), .ZN(n6724)
         );
  NOR4_X1 U7935 ( .A1(n9751), .A2(n6725), .A3(n9575), .A4(n6724), .ZN(n6726)
         );
  XNOR2_X1 U7936 ( .A(n9736), .B(n9747), .ZN(n9728) );
  NAND4_X1 U7937 ( .A1(n9715), .A2(n9766), .A3(n6726), .A4(n9728), .ZN(n6727)
         );
  NOR4_X1 U7938 ( .A1(n9661), .A2(n9700), .A3(n9590), .A4(n6727), .ZN(n6728)
         );
  NAND4_X1 U7939 ( .A1(n9614), .A2(n9630), .A3(n9648), .A4(n6728), .ZN(n6730)
         );
  INV_X1 U7940 ( .A(n6729), .ZN(n6832) );
  INV_X1 U7941 ( .A(n6774), .ZN(n6732) );
  NAND2_X1 U7942 ( .A1(n6733), .A2(n9743), .ZN(n6734) );
  NAND2_X1 U7943 ( .A1(n6734), .A2(n6822), .ZN(n9604) );
  AND3_X1 U7944 ( .A1(n6753), .A2(n6735), .A3(n9604), .ZN(n6828) );
  NAND2_X1 U7945 ( .A1(n6739), .A2(n7789), .ZN(n7795) );
  NAND2_X1 U7946 ( .A1(n7795), .A2(n6786), .ZN(n6743) );
  NAND2_X1 U7947 ( .A1(n6741), .A2(n6740), .ZN(n6797) );
  AND2_X1 U7948 ( .A1(n6797), .A2(n7861), .ZN(n6742) );
  NAND2_X1 U7949 ( .A1(n6743), .A2(n6742), .ZN(n7879) );
  NAND2_X1 U7950 ( .A1(n7879), .A2(n7880), .ZN(n7878) );
  NAND2_X1 U7951 ( .A1(n7878), .A2(n6744), .ZN(n8013) );
  NAND2_X1 U7952 ( .A1(n8013), .A2(n8014), .ZN(n8012) );
  NAND3_X1 U7953 ( .A1(n8012), .A2(n7967), .A3(n7968), .ZN(n7971) );
  NAND2_X1 U7954 ( .A1(n7971), .A2(n6745), .ZN(n8069) );
  AOI21_X2 U7955 ( .B1(n8069), .B2(n8076), .A(n6746), .ZN(n8202) );
  INV_X1 U7956 ( .A(n8197), .ZN(n8203) );
  NAND2_X1 U7957 ( .A1(n8202), .A2(n8203), .ZN(n8201) );
  NAND2_X1 U7958 ( .A1(n8201), .A2(n6747), .ZN(n8172) );
  NAND2_X1 U7959 ( .A1(n8172), .A2(n8173), .ZN(n8171) );
  NAND2_X1 U7960 ( .A1(n8171), .A2(n6748), .ZN(n9827) );
  NAND2_X1 U7961 ( .A1(n9827), .A2(n9828), .ZN(n9826) );
  NAND2_X1 U7962 ( .A1(n9807), .A2(n6750), .ZN(n9780) );
  NAND2_X1 U7963 ( .A1(n6751), .A2(n9608), .ZN(n6752) );
  NAND2_X1 U7964 ( .A1(n9609), .A2(n6752), .ZN(n6754) );
  NAND2_X1 U7965 ( .A1(n6754), .A2(n6753), .ZN(n6756) );
  NAND2_X1 U7966 ( .A1(n6756), .A2(n6755), .ZN(n6826) );
  AOI21_X1 U7967 ( .B1(n6828), .B2(n9605), .A(n6826), .ZN(n6765) );
  NAND2_X1 U7968 ( .A1(n9613), .A2(n9612), .ZN(n6759) );
  OR2_X1 U7969 ( .A1(n6759), .A2(n6757), .ZN(n6830) );
  INV_X1 U7970 ( .A(n6758), .ZN(n6763) );
  AOI21_X1 U7971 ( .B1(n6761), .B2(n6760), .A(n6759), .ZN(n6762) );
  NOR3_X1 U7972 ( .A1(n6764), .A2(n6763), .A3(n6762), .ZN(n6829) );
  OAI21_X1 U7973 ( .B1(n6765), .B2(n6830), .A(n6829), .ZN(n6767) );
  NAND3_X1 U7974 ( .A1(n6767), .A2(n6833), .A3(n6766), .ZN(n6769) );
  NAND2_X1 U7975 ( .A1(n6769), .A2(n6768), .ZN(n6773) );
  NOR2_X1 U7976 ( .A1(n6771), .A2(n6770), .ZN(n6835) );
  NAND2_X1 U7977 ( .A1(n6848), .A2(n7564), .ZN(n7568) );
  AOI211_X1 U7978 ( .C1(n6773), .C2(n6835), .A(n6772), .B(n7568), .ZN(n6775)
         );
  NOR2_X1 U7979 ( .A1(n6775), .A2(n6774), .ZN(n6776) );
  NAND2_X1 U7980 ( .A1(n7232), .A2(n10222), .ZN(n6777) );
  OAI21_X1 U7981 ( .B1(n9568), .B2(n6777), .A(n8109), .ZN(n6780) );
  NAND2_X1 U7982 ( .A1(n6784), .A2(n6783), .ZN(n6847) );
  INV_X1 U7983 ( .A(n6785), .ZN(n6814) );
  INV_X1 U7984 ( .A(n6786), .ZN(n6799) );
  INV_X1 U7985 ( .A(n6787), .ZN(n6793) );
  AOI21_X1 U7986 ( .B1(n6363), .B2(n10735), .A(n8028), .ZN(n6790) );
  NAND4_X1 U7987 ( .A1(n6791), .A2(n6790), .A3(n6789), .A4(n6788), .ZN(n6792)
         );
  NAND2_X1 U7988 ( .A1(n6793), .A2(n6792), .ZN(n6796) );
  AOI211_X1 U7989 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n5222), .ZN(n6798)
         );
  OAI21_X1 U7990 ( .B1(n6799), .B2(n6798), .A(n6797), .ZN(n6802) );
  AOI21_X1 U7991 ( .B1(n6802), .B2(n6801), .A(n6800), .ZN(n6807) );
  INV_X1 U7992 ( .A(n6803), .ZN(n6806) );
  OAI211_X1 U7993 ( .C1(n6807), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6808)
         );
  NAND3_X1 U7994 ( .A1(n6810), .A2(n6809), .A3(n6808), .ZN(n6813) );
  INV_X1 U7995 ( .A(n6811), .ZN(n6812) );
  AOI21_X1 U7996 ( .B1(n6814), .B2(n6813), .A(n6812), .ZN(n6816) );
  OAI21_X1 U7997 ( .B1(n6816), .B2(n5245), .A(n6815), .ZN(n6819) );
  INV_X1 U7998 ( .A(n6817), .ZN(n6818) );
  AOI21_X1 U7999 ( .B1(n6820), .B2(n6819), .A(n6818), .ZN(n6825) );
  INV_X1 U8000 ( .A(n6821), .ZN(n6824) );
  OAI211_X1 U8001 ( .C1(n6825), .C2(n6824), .A(n6823), .B(n6822), .ZN(n6827)
         );
  AOI21_X1 U8002 ( .B1(n6828), .B2(n6827), .A(n6826), .ZN(n6831) );
  OAI21_X1 U8003 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(n6834) );
  AOI21_X1 U8004 ( .B1(n6834), .B2(n6833), .A(n6832), .ZN(n6838) );
  INV_X1 U8005 ( .A(n6835), .ZN(n6837) );
  OAI21_X1 U8006 ( .B1(n6838), .B2(n6837), .A(n6836), .ZN(n6842) );
  NAND2_X1 U8007 ( .A1(n6839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6840) );
  MUX2_X1 U8008 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6840), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6841) );
  NAND2_X1 U8009 ( .A1(n6841), .A2(n4960), .ZN(n6856) );
  INV_X1 U8010 ( .A(n6856), .ZN(n7222) );
  NAND2_X1 U8011 ( .A1(n7222), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8195) );
  AOI21_X1 U8012 ( .B1(n6842), .B2(n7548), .A(n8195), .ZN(n6846) );
  NAND2_X1 U8013 ( .A1(n7961), .A2(n10222), .ZN(n10706) );
  INV_X1 U8014 ( .A(n10706), .ZN(n6843) );
  NAND2_X1 U8015 ( .A1(n6847), .A2(n5558), .ZN(n6860) );
  INV_X1 U8016 ( .A(n9440), .ZN(n9998) );
  INV_X1 U8017 ( .A(n9565), .ZN(n10298) );
  NAND2_X1 U8018 ( .A1(n9998), .A2(n10298), .ZN(n9431) );
  NAND2_X1 U8019 ( .A1(n7564), .A2(n9552), .ZN(n7550) );
  OR2_X1 U8020 ( .A1(n7346), .A2(n7550), .ZN(n10701) );
  NAND2_X1 U8021 ( .A1(n6851), .A2(n6850), .ZN(n6853) );
  NAND2_X1 U8022 ( .A1(n6853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6854) );
  NOR3_X1 U8023 ( .A1(n9431), .A2(n10701), .A3(n9983), .ZN(n6858) );
  OAI21_X1 U8024 ( .B1(n7564), .B2(n8195), .A(P1_B_REG_SCAN_IN), .ZN(n6857) );
  OR2_X1 U8025 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  NAND2_X1 U8026 ( .A1(n6860), .A2(n6859), .ZN(P1_U3242) );
  INV_X4 U8027 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U8028 ( .A1(n8590), .A2(n7239), .ZN(n6861) );
  INV_X1 U8029 ( .A(n7239), .ZN(n8217) );
  NAND2_X1 U8030 ( .A1(n6861), .A2(n7008), .ZN(n7005) );
  OR2_X1 U8031 ( .A1(n7005), .A2(n6862), .ZN(n6863) );
  NAND2_X1 U8032 ( .A1(n6863), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8033 ( .A(n10663), .ZN(n7635) );
  INV_X1 U8034 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10539) );
  INV_X1 U8035 ( .A(n8944), .ZN(n7212) );
  NAND2_X1 U8036 ( .A1(n6902), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6865) );
  INV_X1 U8037 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7331) );
  NOR2_X1 U8038 ( .A1(n7330), .A2(n7331), .ZN(n7329) );
  INV_X1 U8039 ( .A(n6865), .ZN(n6866) );
  INV_X1 U8040 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6867) );
  MUX2_X1 U8041 ( .A(n6867), .B(P2_REG2_REG_2__SCAN_IN), .S(n8449), .Z(n7315)
         );
  NOR2_X1 U8042 ( .A1(n7316), .A2(n7315), .ZN(n7314) );
  AOI21_X1 U8043 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n8449), .A(n7314), .ZN(
        n6868) );
  INV_X1 U8044 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7532) );
  INV_X1 U8045 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6869) );
  MUX2_X1 U8046 ( .A(n6869), .B(P2_REG2_REG_4__SCAN_IN), .S(n7406), .Z(n7409)
         );
  NAND2_X1 U8047 ( .A1(n10491), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10490) );
  INV_X1 U8048 ( .A(n8946), .ZN(n6871) );
  INV_X1 U8049 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6870) );
  MUX2_X1 U8050 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6870), .S(n8944), .Z(n8945)
         );
  AOI21_X1 U8051 ( .B1(n10490), .B2(n6871), .A(n8945), .ZN(n8950) );
  AOI21_X1 U8052 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7212), .A(n8950), .ZN(
        n6872) );
  XNOR2_X1 U8053 ( .A(n6872), .B(n10500), .ZN(n10507) );
  INV_X1 U8054 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10508) );
  INV_X1 U8055 ( .A(n10500), .ZN(n7218) );
  NAND2_X1 U8056 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7225), .ZN(n6874) );
  OAI21_X1 U8057 ( .B1(n7225), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6874), .ZN(
        n10524) );
  INV_X1 U8058 ( .A(n6874), .ZN(n6875) );
  NOR2_X1 U8059 ( .A1(n10539), .A2(n10540), .ZN(n10538) );
  NOR2_X1 U8060 ( .A1(n10530), .A2(n6876), .ZN(n6877) );
  NAND2_X1 U8061 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7247), .ZN(n6878) );
  OAI21_X1 U8062 ( .B1(n7247), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6878), .ZN(
        n10556) );
  NOR2_X1 U8063 ( .A1(n10557), .A2(n10556), .ZN(n10555) );
  INV_X1 U8064 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10572) );
  NOR2_X1 U8065 ( .A1(n10563), .A2(n6879), .ZN(n6880) );
  INV_X1 U8066 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6943) );
  XNOR2_X1 U8067 ( .A(n10579), .B(n6943), .ZN(n10591) );
  INV_X1 U8068 ( .A(n10579), .ZN(n7275) );
  NAND2_X1 U8069 ( .A1(n7275), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6881) );
  NAND2_X2 U8070 ( .A1(n10588), .A2(n6881), .ZN(n6882) );
  INV_X1 U8071 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10606) );
  INV_X1 U8072 ( .A(n6882), .ZN(n6883) );
  INV_X1 U8073 ( .A(n10613), .ZN(n7428) );
  NAND2_X1 U8074 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7428), .ZN(n6885) );
  OAI21_X1 U8075 ( .B1(n7428), .B2(P2_REG2_REG_14__SCAN_IN), .A(n6885), .ZN(
        n10623) );
  INV_X1 U8076 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10638) );
  NOR2_X1 U8077 ( .A1(n10629), .A2(n6888), .ZN(n6889) );
  MUX2_X1 U8078 ( .A(n6929), .B(P2_REG2_REG_16__SCAN_IN), .S(n10645), .Z(n6890) );
  INV_X1 U8079 ( .A(n6890), .ZN(n10654) );
  INV_X1 U8080 ( .A(n10645), .ZN(n7512) );
  INV_X1 U8081 ( .A(n6891), .ZN(n6892) );
  OR2_X2 U8082 ( .A1(n10663), .A2(n6891), .ZN(n7018) );
  INV_X1 U8083 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10674) );
  INV_X1 U8084 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9085) );
  OR2_X1 U8085 ( .A1(n7027), .A2(n9085), .ZN(n6894) );
  NAND2_X1 U8086 ( .A1(n7027), .A2(n9085), .ZN(n6893) );
  NAND2_X1 U8087 ( .A1(n6894), .A2(n6893), .ZN(n7020) );
  AOI21_X1 U8088 ( .B1(n7018), .B2(n9085), .A(n7027), .ZN(n6895) );
  INV_X1 U8089 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6896) );
  MUX2_X1 U8090 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n6896), .S(n4941), .Z(n6999)
         );
  XNOR2_X1 U8091 ( .A(n6897), .B(n6999), .ZN(n7017) );
  INV_X1 U8092 ( .A(n7005), .ZN(n6899) );
  OR2_X1 U8093 ( .A1(n7002), .A2(P2_U3151), .ZN(n9268) );
  INV_X1 U8094 ( .A(n9268), .ZN(n6898) );
  AND2_X1 U8095 ( .A1(n6899), .A2(n6898), .ZN(n7255) );
  INV_X1 U8096 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9154) );
  AOI22_X1 U8097 ( .A1(n10645), .A2(n9154), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n7512), .ZN(n10648) );
  NAND2_X1 U8098 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7428), .ZN(n6920) );
  INV_X1 U8099 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U8100 ( .A1(n10613), .A2(n6900), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7428), .ZN(n10616) );
  NAND2_X1 U8101 ( .A1(n7275), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6917) );
  INV_X1 U8102 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6901) );
  MUX2_X1 U8103 ( .A(n6901), .B(P2_REG1_REG_12__SCAN_IN), .S(n10579), .Z(
        n10581) );
  INV_X1 U8104 ( .A(n10563), .ZN(n7269) );
  NAND2_X1 U8105 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7247), .ZN(n6914) );
  INV_X1 U8106 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8160) );
  AOI22_X1 U8107 ( .A1(n10546), .A2(n8160), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7247), .ZN(n10549) );
  INV_X1 U8108 ( .A(n10530), .ZN(n7244) );
  NAND2_X1 U8109 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7225), .ZN(n6911) );
  INV_X1 U8110 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8034) );
  AOI22_X1 U8111 ( .A1(n10514), .A2(n8034), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7225), .ZN(n10517) );
  INV_X1 U8112 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6908) );
  INV_X1 U8113 ( .A(n8449), .ZN(n6968) );
  INV_X1 U8114 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6905) );
  INV_X1 U8115 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U8116 ( .A1(n5350), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6903) );
  AOI22_X1 U8117 ( .A1(n6864), .A2(n6903), .B1(n6902), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n7328) );
  NAND2_X1 U8118 ( .A1(n7328), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7327) );
  OAI21_X1 U8119 ( .B1(n7437), .B2(n6904), .A(n7327), .ZN(n7312) );
  MUX2_X1 U8120 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6905), .S(n8449), .Z(n7313)
         );
  NAND2_X1 U8121 ( .A1(n7312), .A2(n7313), .ZN(n7311) );
  OAI21_X1 U8122 ( .B1(n6968), .B2(n6905), .A(n7311), .ZN(n6906) );
  XNOR2_X1 U8123 ( .A(n6907), .B(n7207), .ZN(n10482) );
  NAND2_X1 U8124 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n10482), .ZN(n10481) );
  MUX2_X1 U8125 ( .A(n6908), .B(P2_REG1_REG_6__SCAN_IN), .S(n8944), .Z(n8937)
         );
  NAND2_X1 U8126 ( .A1(n6909), .A2(n7218), .ZN(n6910) );
  NAND2_X1 U8127 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n10499), .ZN(n10498) );
  NAND2_X1 U8128 ( .A1(n7244), .A2(n6912), .ZN(n6913) );
  NAND2_X1 U8129 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n10532), .ZN(n10531) );
  NAND2_X1 U8130 ( .A1(n7269), .A2(n6915), .ZN(n6916) );
  NAND2_X1 U8131 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10565), .ZN(n10564) );
  NAND2_X1 U8132 ( .A1(n7309), .A2(n6918), .ZN(n6919) );
  NAND2_X1 U8133 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10599), .ZN(n10598) );
  NAND2_X1 U8134 ( .A1(n6886), .A2(n6921), .ZN(n6922) );
  NAND2_X1 U8135 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10631), .ZN(n10630) );
  NAND2_X1 U8136 ( .A1(n7635), .A2(n6923), .ZN(n6924) );
  NAND2_X1 U8137 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10665), .ZN(n10664) );
  XNOR2_X1 U8138 ( .A(n7027), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n7023) );
  INV_X1 U8139 ( .A(n7027), .ZN(n7667) );
  AOI22_X1 U8140 ( .A1(n7022), .A2(n7023), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n7667), .ZN(n6925) );
  XNOR2_X1 U8141 ( .A(n4941), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6997) );
  XNOR2_X1 U8142 ( .A(n6925), .B(n6997), .ZN(n7014) );
  NAND2_X1 U8143 ( .A1(n7255), .A2(n8788), .ZN(n8939) );
  OR2_X1 U8144 ( .A1(n8788), .A2(n10674), .ZN(n6927) );
  NAND2_X1 U8145 ( .A1(n8788), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6926) );
  AND2_X1 U8146 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  NAND2_X1 U8147 ( .A1(n6928), .A2(n10663), .ZN(n6990) );
  XNOR2_X1 U8148 ( .A(n7635), .B(n6928), .ZN(n10668) );
  INV_X1 U8149 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6929) );
  OR2_X1 U8150 ( .A1(n8788), .A2(n6929), .ZN(n6931) );
  NAND2_X1 U8151 ( .A1(n8788), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8152 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  OR2_X1 U8153 ( .A1(n7512), .A2(n6932), .ZN(n6989) );
  XNOR2_X1 U8154 ( .A(n6932), .B(n10645), .ZN(n10651) );
  OR2_X1 U8155 ( .A1(n8788), .A2(n10638), .ZN(n6934) );
  NAND2_X1 U8156 ( .A1(n8788), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U8157 ( .A1(n6934), .A2(n6933), .ZN(n6935) );
  OR2_X1 U8158 ( .A1(n6886), .A2(n6935), .ZN(n6988) );
  XNOR2_X1 U8159 ( .A(n6935), .B(n10629), .ZN(n10634) );
  INV_X1 U8160 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6936) );
  OR2_X1 U8161 ( .A1(n8788), .A2(n6936), .ZN(n6938) );
  NAND2_X1 U8162 ( .A1(n8788), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8163 ( .A1(n6938), .A2(n6937), .ZN(n6939) );
  OR2_X1 U8164 ( .A1(n7428), .A2(n6939), .ZN(n6987) );
  XNOR2_X1 U8165 ( .A(n6939), .B(n10613), .ZN(n10619) );
  OR2_X1 U8166 ( .A1(n8788), .A2(n10606), .ZN(n6941) );
  NAND2_X1 U8167 ( .A1(n8788), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8168 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  OR2_X1 U8169 ( .A1(n7309), .A2(n6942), .ZN(n6986) );
  XNOR2_X1 U8170 ( .A(n6942), .B(n10597), .ZN(n10602) );
  OR2_X1 U8171 ( .A1(n8788), .A2(n6943), .ZN(n6945) );
  NAND2_X1 U8172 ( .A1(n8788), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8173 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  OR2_X1 U8174 ( .A1(n7275), .A2(n6946), .ZN(n6985) );
  XNOR2_X1 U8175 ( .A(n6946), .B(n10579), .ZN(n10585) );
  OR2_X1 U8176 ( .A1(n8788), .A2(n10572), .ZN(n6948) );
  NAND2_X1 U8177 ( .A1(n8788), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8178 ( .A1(n6948), .A2(n6947), .ZN(n6949) );
  OR2_X1 U8179 ( .A1(n7269), .A2(n6949), .ZN(n6984) );
  XNOR2_X1 U8180 ( .A(n6949), .B(n10563), .ZN(n10568) );
  INV_X1 U8181 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6950) );
  OR2_X1 U8182 ( .A1(n8788), .A2(n6950), .ZN(n6952) );
  NAND2_X1 U8183 ( .A1(n8788), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U8184 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  OR2_X1 U8185 ( .A1(n7247), .A2(n6953), .ZN(n6983) );
  XNOR2_X1 U8186 ( .A(n6953), .B(n10546), .ZN(n10552) );
  MUX2_X1 U8187 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8788), .Z(n6954) );
  OR2_X1 U8188 ( .A1(n6954), .A2(n7244), .ZN(n6982) );
  XNOR2_X1 U8189 ( .A(n6954), .B(n10530), .ZN(n10535) );
  MUX2_X1 U8190 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8788), .Z(n6955) );
  OR2_X1 U8191 ( .A1(n6955), .A2(n7225), .ZN(n6981) );
  XNOR2_X1 U8192 ( .A(n6955), .B(n10514), .ZN(n10520) );
  OR2_X1 U8193 ( .A1(n8788), .A2(n10508), .ZN(n6957) );
  NAND2_X1 U8194 ( .A1(n8788), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8195 ( .A1(n6957), .A2(n6956), .ZN(n6958) );
  OR2_X1 U8196 ( .A1(n7218), .A2(n6958), .ZN(n6980) );
  XNOR2_X1 U8197 ( .A(n6958), .B(n10500), .ZN(n10503) );
  MUX2_X1 U8198 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8788), .Z(n6979) );
  INV_X1 U8199 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6959) );
  OR2_X1 U8200 ( .A1(n8788), .A2(n6959), .ZN(n6961) );
  NAND2_X1 U8201 ( .A1(n8788), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U8202 ( .A1(n6961), .A2(n6960), .ZN(n6978) );
  MUX2_X1 U8203 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6967), .Z(n6965) );
  XNOR2_X1 U8204 ( .A(n6864), .B(n6965), .ZN(n7341) );
  OR2_X1 U8205 ( .A1(n6967), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U8206 ( .A1(n6967), .A2(n7437), .ZN(n6963) );
  NAND2_X1 U8207 ( .A1(n6964), .A2(n6963), .ZN(n7257) );
  NAND2_X1 U8208 ( .A1(n7257), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U8209 ( .A1(n7341), .A2(n7340), .ZN(n7339) );
  NAND2_X1 U8210 ( .A1(n6965), .A2(n7334), .ZN(n6966) );
  NAND2_X1 U8211 ( .A1(n7339), .A2(n6966), .ZN(n7323) );
  MUX2_X1 U8212 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6967), .Z(n6969) );
  XNOR2_X1 U8213 ( .A(n6969), .B(n6968), .ZN(n7322) );
  NAND2_X1 U8214 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U8215 ( .A1(n6969), .A2(n8449), .ZN(n6970) );
  NAND2_X1 U8216 ( .A1(n7321), .A2(n6970), .ZN(n7393) );
  OR2_X1 U8217 ( .A1(n8788), .A2(n7532), .ZN(n6972) );
  NAND2_X1 U8218 ( .A1(n8788), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8219 ( .A1(n6972), .A2(n6971), .ZN(n6973) );
  XNOR2_X1 U8220 ( .A(n6973), .B(n7206), .ZN(n7394) );
  OR2_X1 U8221 ( .A1(n7393), .A2(n7394), .ZN(n7391) );
  INV_X1 U8222 ( .A(n6973), .ZN(n6974) );
  NAND2_X1 U8223 ( .A1(n6974), .A2(n5359), .ZN(n6975) );
  NAND2_X1 U8224 ( .A1(n7391), .A2(n6975), .ZN(n7419) );
  MUX2_X1 U8225 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8788), .Z(n6976) );
  XNOR2_X1 U8226 ( .A(n6976), .B(n7406), .ZN(n7418) );
  OR2_X1 U8227 ( .A1(n7419), .A2(n7418), .ZN(n7421) );
  NAND2_X1 U8228 ( .A1(n6976), .A2(n7406), .ZN(n6977) );
  NAND2_X1 U8229 ( .A1(n7421), .A2(n6977), .ZN(n10486) );
  XNOR2_X1 U8230 ( .A(n6978), .B(n10483), .ZN(n10485) );
  AND2_X1 U8231 ( .A1(n10486), .A2(n10485), .ZN(n10487) );
  AOI21_X1 U8232 ( .B1(n7207), .B2(n6978), .A(n10487), .ZN(n8935) );
  XNOR2_X1 U8233 ( .A(n6979), .B(n8944), .ZN(n8934) );
  NAND2_X1 U8234 ( .A1(n8935), .A2(n8934), .ZN(n8933) );
  OAI21_X1 U8235 ( .B1(n6979), .B2(n7212), .A(n8933), .ZN(n10504) );
  NAND2_X1 U8236 ( .A1(n10503), .A2(n10504), .ZN(n10502) );
  NAND2_X1 U8237 ( .A1(n6980), .A2(n10502), .ZN(n10519) );
  NAND2_X1 U8238 ( .A1(n10520), .A2(n10519), .ZN(n10518) );
  NAND2_X1 U8239 ( .A1(n6981), .A2(n10518), .ZN(n10534) );
  NAND2_X1 U8240 ( .A1(n10535), .A2(n10534), .ZN(n10533) );
  NAND2_X1 U8241 ( .A1(n6982), .A2(n10533), .ZN(n10551) );
  NAND2_X1 U8242 ( .A1(n10552), .A2(n10551), .ZN(n10550) );
  NAND2_X1 U8243 ( .A1(n6983), .A2(n10550), .ZN(n10567) );
  NAND2_X1 U8244 ( .A1(n10568), .A2(n10567), .ZN(n10566) );
  NAND2_X1 U8245 ( .A1(n6984), .A2(n10566), .ZN(n10584) );
  NAND2_X1 U8246 ( .A1(n10585), .A2(n10584), .ZN(n10583) );
  NAND2_X1 U8247 ( .A1(n6985), .A2(n10583), .ZN(n10601) );
  NAND2_X1 U8248 ( .A1(n10602), .A2(n10601), .ZN(n10600) );
  NAND2_X1 U8249 ( .A1(n6986), .A2(n10600), .ZN(n10618) );
  NAND2_X1 U8250 ( .A1(n10619), .A2(n10618), .ZN(n10617) );
  NAND2_X1 U8251 ( .A1(n6987), .A2(n10617), .ZN(n10633) );
  NAND2_X1 U8252 ( .A1(n10634), .A2(n10633), .ZN(n10632) );
  NAND2_X1 U8253 ( .A1(n6988), .A2(n10632), .ZN(n10650) );
  NAND2_X1 U8254 ( .A1(n10651), .A2(n10650), .ZN(n10649) );
  NAND2_X1 U8255 ( .A1(n6989), .A2(n10649), .ZN(n10667) );
  NAND2_X1 U8256 ( .A1(n10668), .A2(n10667), .ZN(n10666) );
  NAND2_X1 U8257 ( .A1(n6990), .A2(n10666), .ZN(n6996) );
  INV_X1 U8258 ( .A(n6996), .ZN(n6994) );
  OR2_X1 U8259 ( .A1(n8788), .A2(n9085), .ZN(n6992) );
  NAND2_X1 U8260 ( .A1(n8788), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6991) );
  AND2_X1 U8261 ( .A1(n6992), .A2(n6991), .ZN(n6995) );
  INV_X1 U8262 ( .A(n6995), .ZN(n6993) );
  NAND2_X1 U8263 ( .A1(n6994), .A2(n6993), .ZN(n7025) );
  AND2_X1 U8264 ( .A1(n6996), .A2(n6995), .ZN(n7024) );
  AOI21_X1 U8265 ( .B1(n7027), .B2(n7025), .A(n7024), .ZN(n7001) );
  INV_X1 U8266 ( .A(n6997), .ZN(n6998) );
  MUX2_X1 U8267 ( .A(n6999), .B(n6998), .S(n8788), .Z(n7000) );
  XNOR2_X1 U8268 ( .A(n7001), .B(n7000), .ZN(n7012) );
  INV_X1 U8269 ( .A(n7002), .ZN(n8656) );
  NOR2_X2 U8270 ( .A1(n8931), .A2(n8656), .ZN(n10670) );
  NOR2_X1 U8271 ( .A1(n8788), .A2(P2_U3151), .ZN(n7003) );
  NAND2_X1 U8272 ( .A1(n7003), .A2(n7002), .ZN(n7004) );
  OR2_X1 U8273 ( .A1(n7005), .A2(n7004), .ZN(n7007) );
  OR2_X1 U8274 ( .A1(n7008), .A2(n9268), .ZN(n7006) );
  INV_X1 U8275 ( .A(n10662), .ZN(n7335) );
  INV_X1 U8276 ( .A(n7008), .ZN(n7009) );
  NOR2_X2 U8277 ( .A1(P2_U3150), .A2(n7009), .ZN(n10661) );
  NAND2_X1 U8278 ( .A1(n10661), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U8279 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8824) );
  OAI211_X1 U8280 ( .C1(n7335), .C2(n8655), .A(n7010), .B(n8824), .ZN(n7011)
         );
  INV_X1 U8281 ( .A(n7015), .ZN(n7016) );
  OAI21_X1 U8282 ( .B1(n7017), .B2(n10677), .A(n7016), .ZN(P2_U3201) );
  INV_X1 U8283 ( .A(n7018), .ZN(n7019) );
  OR2_X1 U8284 ( .A1(n7019), .A2(n10673), .ZN(n7021) );
  XNOR2_X1 U8285 ( .A(n7021), .B(n7020), .ZN(n7035) );
  INV_X1 U8286 ( .A(n7024), .ZN(n7026) );
  NAND2_X1 U8287 ( .A1(n7026), .A2(n7025), .ZN(n7032) );
  OAI21_X1 U8288 ( .B1(n7032), .B2(n8931), .A(n7335), .ZN(n7028) );
  NAND2_X1 U8289 ( .A1(n7028), .A2(n7027), .ZN(n7030) );
  NAND3_X1 U8290 ( .A1(n7032), .A2(n10670), .A3(n7667), .ZN(n7033) );
  NAND2_X1 U8291 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8886) );
  NOR2_X1 U8292 ( .A1(n7527), .A2(n8649), .ZN(n7036) );
  NAND2_X1 U8293 ( .A1(n7037), .A2(n7036), .ZN(n7039) );
  NAND2_X1 U8294 ( .A1(n8649), .A2(n7958), .ZN(n7038) );
  XNOR2_X1 U8295 ( .A(n4940), .B(n7723), .ZN(n7056) );
  NAND2_X1 U8296 ( .A1(n7042), .A2(n7041), .ZN(n7046) );
  NAND2_X1 U8297 ( .A1(n4991), .A2(n7046), .ZN(n7472) );
  NAND2_X1 U8298 ( .A1(n7474), .A2(n7432), .ZN(n7043) );
  AND2_X1 U8299 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  INV_X1 U8300 ( .A(n7046), .ZN(n7047) );
  XNOR2_X1 U8301 ( .A(n7050), .B(n7544), .ZN(n7048) );
  XNOR2_X1 U8302 ( .A(n7048), .B(n7538), .ZN(n7482) );
  INV_X1 U8303 ( .A(n7048), .ZN(n7049) );
  XNOR2_X1 U8304 ( .A(n4940), .B(n7709), .ZN(n7054) );
  XNOR2_X1 U8305 ( .A(n7054), .B(n7605), .ZN(n7504) );
  NAND2_X1 U8306 ( .A1(n7505), .A2(n7504), .ZN(n7503) );
  NAND2_X1 U8307 ( .A1(n7054), .A2(n8932), .ZN(n7595) );
  AND2_X1 U8308 ( .A1(n7594), .A2(n7595), .ZN(n7055) );
  XNOR2_X1 U8309 ( .A(n7056), .B(n7915), .ZN(n7618) );
  XNOR2_X1 U8310 ( .A(n8036), .B(n8794), .ZN(n7057) );
  XNOR2_X1 U8311 ( .A(n7057), .B(n7930), .ZN(n8893) );
  NAND2_X1 U8312 ( .A1(n8892), .A2(n7058), .ZN(n7895) );
  INV_X1 U8313 ( .A(n7895), .ZN(n7060) );
  XNOR2_X1 U8314 ( .A(n7934), .B(n8794), .ZN(n7061) );
  XNOR2_X1 U8315 ( .A(n7061), .B(n8899), .ZN(n7894) );
  NAND2_X1 U8316 ( .A1(n7060), .A2(n7059), .ZN(n7897) );
  NAND2_X1 U8317 ( .A1(n7061), .A2(n8899), .ZN(n7062) );
  XOR2_X1 U8318 ( .A(n8794), .B(n8030), .Z(n8001) );
  NOR2_X1 U8319 ( .A1(n8001), .A2(n8000), .ZN(n7064) );
  NAND2_X1 U8320 ( .A1(n8001), .A2(n8000), .ZN(n7063) );
  XNOR2_X1 U8321 ( .A(n8165), .B(n8794), .ZN(n7065) );
  XOR2_X1 U8322 ( .A(n8289), .B(n7065), .Z(n8096) );
  INV_X1 U8323 ( .A(n7065), .ZN(n7066) );
  XNOR2_X1 U8324 ( .A(n5856), .B(n8794), .ZN(n7067) );
  NAND2_X1 U8325 ( .A1(n7068), .A2(n7067), .ZN(n8351) );
  XNOR2_X1 U8326 ( .A(n8188), .B(n7474), .ZN(n7074) );
  XNOR2_X1 U8327 ( .A(n7074), .B(n8400), .ZN(n8352) );
  INV_X1 U8328 ( .A(n8352), .ZN(n7071) );
  OR2_X1 U8329 ( .A1(n8928), .A2(n7071), .ZN(n7070) );
  NOR2_X1 U8330 ( .A1(n7071), .A2(n8351), .ZN(n7072) );
  MUX2_X1 U8331 ( .A(n8220), .B(n7076), .S(n8794), .Z(n8394) );
  XOR2_X1 U8332 ( .A(n8794), .B(n8402), .Z(n7077) );
  XNOR2_X1 U8333 ( .A(n8237), .B(n8794), .ZN(n7078) );
  XNOR2_X1 U8334 ( .A(n7078), .B(n7079), .ZN(n8864) );
  INV_X1 U8335 ( .A(n7078), .ZN(n7080) );
  NAND2_X1 U8336 ( .A1(n8863), .A2(n7081), .ZN(n8806) );
  INV_X1 U8337 ( .A(n8806), .ZN(n7083) );
  XNOR2_X1 U8338 ( .A(n10827), .B(n8794), .ZN(n7084) );
  XNOR2_X1 U8339 ( .A(n7084), .B(n8915), .ZN(n8809) );
  INV_X1 U8340 ( .A(n8809), .ZN(n7082) );
  XNOR2_X1 U8341 ( .A(n8413), .B(n8794), .ZN(n7087) );
  XNOR2_X1 U8342 ( .A(n7087), .B(n9171), .ZN(n8908) );
  NAND2_X1 U8343 ( .A1(n8910), .A2(n7088), .ZN(n8840) );
  XNOR2_X1 U8344 ( .A(n9243), .B(n8794), .ZN(n7089) );
  XOR2_X1 U8345 ( .A(n9095), .B(n7089), .Z(n8839) );
  NAND2_X1 U8346 ( .A1(n8840), .A2(n8839), .ZN(n8838) );
  INV_X1 U8347 ( .A(n7089), .ZN(n7090) );
  INV_X1 U8348 ( .A(n9095), .ZN(n10844) );
  NAND2_X1 U8349 ( .A1(n7090), .A2(n10844), .ZN(n7091) );
  NAND2_X1 U8350 ( .A1(n8838), .A2(n7091), .ZN(n10849) );
  INV_X1 U8351 ( .A(n10849), .ZN(n7093) );
  XNOR2_X1 U8352 ( .A(n8536), .B(n8794), .ZN(n7094) );
  XNOR2_X1 U8353 ( .A(n7094), .B(n9081), .ZN(n10848) );
  INV_X1 U8354 ( .A(n10848), .ZN(n7092) );
  INV_X1 U8355 ( .A(n7094), .ZN(n7095) );
  XNOR2_X1 U8356 ( .A(n9232), .B(n8794), .ZN(n7098) );
  XNOR2_X1 U8357 ( .A(n7098), .B(n9094), .ZN(n8882) );
  INV_X1 U8358 ( .A(n7098), .ZN(n7099) );
  NAND2_X1 U8359 ( .A1(n7099), .A2(n10846), .ZN(n7100) );
  NAND2_X1 U8360 ( .A1(n8884), .A2(n7100), .ZN(n8823) );
  XNOR2_X1 U8361 ( .A(n9071), .B(n8794), .ZN(n8822) );
  NAND2_X1 U8362 ( .A1(n8823), .A2(n8822), .ZN(n8821) );
  INV_X1 U8363 ( .A(n8822), .ZN(n7101) );
  INV_X1 U8364 ( .A(n9063), .ZN(n9083) );
  NAND2_X1 U8365 ( .A1(n7101), .A2(n9083), .ZN(n7102) );
  XNOR2_X1 U8366 ( .A(n9141), .B(n8794), .ZN(n7104) );
  XNOR2_X1 U8367 ( .A(n7104), .B(n9048), .ZN(n8857) );
  NAND2_X1 U8368 ( .A1(n7104), .A2(n9048), .ZN(n7105) );
  XNOR2_X1 U8369 ( .A(n9053), .B(n8794), .ZN(n7106) );
  XNOR2_X1 U8370 ( .A(n7106), .B(n9025), .ZN(n8663) );
  XNOR2_X1 U8371 ( .A(n9033), .B(n8794), .ZN(n7108) );
  XNOR2_X1 U8372 ( .A(n7108), .B(n8924), .ZN(n8876) );
  NAND2_X1 U8373 ( .A1(n8874), .A2(n8876), .ZN(n8875) );
  INV_X1 U8374 ( .A(n7108), .ZN(n7109) );
  NAND2_X1 U8375 ( .A1(n7109), .A2(n8924), .ZN(n7110) );
  XNOR2_X1 U8376 ( .A(n9016), .B(n8794), .ZN(n7112) );
  NAND2_X1 U8377 ( .A1(n8815), .A2(n8878), .ZN(n7115) );
  INV_X1 U8378 ( .A(n7111), .ZN(n7113) );
  NAND2_X1 U8379 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U8380 ( .A1(n7115), .A2(n7114), .ZN(n8847) );
  XNOR2_X1 U8381 ( .A(n9201), .B(n8794), .ZN(n7116) );
  XNOR2_X1 U8382 ( .A(n7116), .B(n8987), .ZN(n8848) );
  NAND2_X1 U8383 ( .A1(n8847), .A2(n8848), .ZN(n8670) );
  NAND2_X1 U8384 ( .A1(n7116), .A2(n9012), .ZN(n8669) );
  XNOR2_X1 U8385 ( .A(n8678), .B(n7474), .ZN(n7117) );
  NAND2_X1 U8386 ( .A1(n7117), .A2(n8988), .ZN(n8672) );
  INV_X1 U8387 ( .A(n8672), .ZN(n7120) );
  XNOR2_X1 U8388 ( .A(n9195), .B(n8794), .ZN(n7122) );
  NAND2_X1 U8389 ( .A1(n7122), .A2(n8975), .ZN(n8671) );
  INV_X1 U8390 ( .A(n7117), .ZN(n7118) );
  NAND2_X1 U8391 ( .A1(n7118), .A2(n8832), .ZN(n8673) );
  AND2_X1 U8392 ( .A1(n8671), .A2(n8673), .ZN(n7119) );
  AND2_X1 U8393 ( .A1(n8669), .A2(n7121), .ZN(n7125) );
  INV_X1 U8394 ( .A(n7121), .ZN(n7124) );
  XNOR2_X1 U8395 ( .A(n7122), .B(n8999), .ZN(n8831) );
  AND2_X1 U8396 ( .A1(n8831), .A2(n8672), .ZN(n7123) );
  XNOR2_X1 U8397 ( .A(n9185), .B(n8794), .ZN(n8790) );
  XNOR2_X1 U8398 ( .A(n8790), .B(n8976), .ZN(n8792) );
  XNOR2_X1 U8399 ( .A(n8793), .B(n8792), .ZN(n7155) );
  NAND2_X1 U8400 ( .A1(n7126), .A2(n7129), .ZN(n7184) );
  INV_X1 U8401 ( .A(n8344), .ZN(n9173) );
  OR2_X1 U8402 ( .A1(n9173), .A2(n8590), .ZN(n7128) );
  OAI21_X1 U8403 ( .B1(n7184), .B2(n7128), .A(n7178), .ZN(n7133) );
  NAND3_X1 U8404 ( .A1(n6164), .A2(n7130), .A3(n7129), .ZN(n7181) );
  INV_X1 U8405 ( .A(n7178), .ZN(n7131) );
  NAND2_X1 U8406 ( .A1(n7181), .A2(n7131), .ZN(n7140) );
  AND2_X1 U8407 ( .A1(n7140), .A2(n7185), .ZN(n7132) );
  INV_X1 U8408 ( .A(n7184), .ZN(n7134) );
  NAND2_X1 U8409 ( .A1(n7134), .A2(n7187), .ZN(n7136) );
  INV_X1 U8410 ( .A(n7187), .ZN(n7135) );
  NAND3_X1 U8411 ( .A1(n8576), .A2(n7178), .A3(n8344), .ZN(n7137) );
  NAND2_X1 U8412 ( .A1(n7137), .A2(n10831), .ZN(n7180) );
  NAND2_X1 U8413 ( .A1(n7184), .A2(n7180), .ZN(n7142) );
  AND2_X1 U8414 ( .A1(n7138), .A2(n7239), .ZN(n7141) );
  NAND4_X1 U8415 ( .A1(n7142), .A2(n7141), .A3(n7140), .A4(n7139), .ZN(n7143)
         );
  NAND2_X1 U8416 ( .A1(n7143), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7145) );
  NOR2_X1 U8417 ( .A1(n7179), .A2(n9255), .ZN(n8657) );
  NAND2_X1 U8418 ( .A1(n7181), .A2(n8657), .ZN(n7144) );
  INV_X1 U8419 ( .A(n8657), .ZN(n7146) );
  OR2_X1 U8420 ( .A1(n7181), .A2(n7146), .ZN(n7149) );
  INV_X1 U8421 ( .A(n7148), .ZN(n7147) );
  INV_X1 U8423 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10007) );
  OAI22_X1 U8424 ( .A1(n8898), .A2(n4936), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10007), .ZN(n7151) );
  NOR2_X2 U8425 ( .A1(n7149), .A2(n7148), .ZN(n10845) );
  NOR2_X1 U8426 ( .A1(n8914), .A2(n8832), .ZN(n7150) );
  AOI211_X1 U8427 ( .C1(n8969), .C2(n10856), .A(n7151), .B(n7150), .ZN(n7152)
         );
  OAI21_X1 U8428 ( .B1(n7155), .B2(n8907), .A(n7154), .ZN(P2_U3154) );
  NAND2_X1 U8429 ( .A1(n8803), .A2(n4936), .ZN(n7156) );
  NAND2_X1 U8430 ( .A1(n9262), .A2(n8593), .ZN(n7159) );
  INV_X1 U8431 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9264) );
  OR2_X1 U8432 ( .A1(n5774), .A2(n9264), .ZN(n7158) );
  XNOR2_X1 U8433 ( .A(n8608), .B(n4931), .ZN(n7171) );
  INV_X1 U8434 ( .A(n7529), .ZN(n8120) );
  NAND2_X1 U8435 ( .A1(n7171), .A2(n8120), .ZN(n7170) );
  NAND2_X1 U8436 ( .A1(n8782), .A2(n4936), .ZN(n7161) );
  NAND2_X1 U8437 ( .A1(n7163), .A2(n9103), .ZN(n7169) );
  NAND2_X1 U8438 ( .A1(n5764), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7166) );
  NAND2_X1 U8439 ( .A1(n8596), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7165) );
  NAND2_X1 U8440 ( .A1(n5735), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7164) );
  INV_X1 U8441 ( .A(n8587), .ZN(n8921) );
  AND2_X1 U8442 ( .A1(n5726), .A2(P2_B_REG_SCAN_IN), .ZN(n7167) );
  NOR2_X1 U8443 ( .A1(n9106), .A2(n7167), .ZN(n8955) );
  AOI22_X1 U8444 ( .A1(n8921), .A2(n8955), .B1(n9080), .B2(n4937), .ZN(n7168)
         );
  NAND2_X1 U8445 ( .A1(n8454), .A2(n7174), .ZN(n7176) );
  NAND2_X1 U8446 ( .A1(n9175), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8447 ( .A1(n7177), .A2(n5554), .ZN(P2_U3488) );
  AND2_X1 U8448 ( .A1(n7179), .A2(n7178), .ZN(n7183) );
  INV_X1 U8449 ( .A(n7180), .ZN(n7182) );
  NAND2_X1 U8450 ( .A1(n7186), .A2(n10843), .ZN(n7193) );
  NAND2_X1 U8451 ( .A1(n7188), .A2(n7187), .ZN(n9249) );
  INV_X1 U8452 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7189) );
  NOR2_X1 U8453 ( .A1(n10843), .A2(n7189), .ZN(n7190) );
  NAND2_X1 U8454 ( .A1(n7193), .A2(n7192), .ZN(P2_U3456) );
  INV_X1 U8455 ( .A(n7572), .ZN(n7194) );
  INV_X2 U8456 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U8457 ( .A(n9469), .ZN(n9446) );
  NAND2_X1 U8458 ( .A1(n7195), .A2(P1_U3086), .ZN(n8027) );
  NOR2_X2 U8459 ( .A1(n7195), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9997) );
  INV_X1 U8460 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7265) );
  OAI222_X1 U8461 ( .A1(n9446), .A2(P1_U3086), .B1(n8027), .B2(n8450), .C1(
        n8445), .C2(n7265), .ZN(P1_U3353) );
  INV_X2 U8462 ( .A(n9267), .ZN(n9266) );
  INV_X1 U8463 ( .A(n7196), .ZN(n7199) );
  INV_X1 U8464 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7197) );
  AND2_X1 U8465 ( .A1(n7195), .A2(P2_U3151), .ZN(n9260) );
  INV_X2 U8466 ( .A(n9260), .ZN(n9263) );
  OAI222_X1 U8467 ( .A1(n9266), .A2(n7199), .B1(n7334), .B2(P2_U3151), .C1(
        n7197), .C2(n9263), .ZN(P2_U3294) );
  AOI22_X1 U8468 ( .A1(n9997), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9452), .ZN(n7198) );
  OAI21_X1 U8469 ( .B1(n7199), .B2(n8027), .A(n7198), .ZN(P1_U3354) );
  AOI22_X1 U8470 ( .A1(n9486), .A2(P1_STATE_REG_SCAN_IN), .B1(n9997), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n7200) );
  OAI21_X1 U8471 ( .B1(n7205), .B2(n8027), .A(n7200), .ZN(P1_U3352) );
  OAI222_X1 U8472 ( .A1(n9266), .A2(n7202), .B1(n7406), .B2(P2_U3151), .C1(
        n7201), .C2(n9263), .ZN(P2_U3291) );
  OAI222_X1 U8473 ( .A1(n8445), .A2(n7203), .B1(n8027), .B2(n7202), .C1(
        P1_U3086), .C2(n9489), .ZN(P1_U3351) );
  INV_X1 U8474 ( .A(n9506), .ZN(n7204) );
  OAI222_X1 U8475 ( .A1(n7204), .A2(P1_U3086), .B1(n8027), .B2(n7208), .C1(
        n8445), .C2(n5592), .ZN(P1_U3350) );
  OAI222_X1 U8476 ( .A1(n9263), .A2(n5580), .B1(n7206), .B2(P2_U3151), .C1(
        n9266), .C2(n7205), .ZN(P2_U3292) );
  OAI222_X1 U8477 ( .A1(n9263), .A2(n7209), .B1(n9266), .B2(n7208), .C1(
        P2_U3151), .C2(n7207), .ZN(P2_U3290) );
  INV_X1 U8478 ( .A(n7210), .ZN(n7213) );
  INV_X1 U8479 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7211) );
  OAI222_X1 U8480 ( .A1(n9266), .A2(n7213), .B1(n7212), .B2(P2_U3151), .C1(
        n7211), .C2(n9263), .ZN(P2_U3289) );
  INV_X1 U8481 ( .A(n10313), .ZN(n7214) );
  INV_X1 U8482 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7263) );
  OAI222_X1 U8483 ( .A1(n7214), .A2(P1_U3086), .B1(n8445), .B2(n7263), .C1(
        n7213), .C2(n10000), .ZN(P1_U3349) );
  INV_X1 U8484 ( .A(n7215), .ZN(n7219) );
  AOI22_X1 U8485 ( .A1(n10325), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9997), .ZN(n7216) );
  OAI21_X1 U8486 ( .B1(n7219), .B2(n8027), .A(n7216), .ZN(P1_U3348) );
  INV_X1 U8487 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7217) );
  OAI222_X1 U8488 ( .A1(n9266), .A2(n7219), .B1(n7218), .B2(P2_U3151), .C1(
        n7217), .C2(n9263), .ZN(P2_U3288) );
  INV_X1 U8489 ( .A(n7220), .ZN(n7224) );
  AOI22_X1 U8490 ( .A1(n10336), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9997), .ZN(n7221) );
  OAI21_X1 U8491 ( .B1(n7224), .B2(n8027), .A(n7221), .ZN(P1_U3347) );
  INV_X1 U8492 ( .A(n9430), .ZN(n7223) );
  NAND2_X1 U8493 ( .A1(n9983), .A2(n8195), .ZN(n9429) );
  NOR2_X1 U8494 ( .A1(n10683), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8495 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7237) );
  OAI222_X1 U8496 ( .A1(n7225), .A2(P2_U3151), .B1(n9266), .B2(n7224), .C1(
        n9263), .C2(n7237), .ZN(P2_U3287) );
  INV_X1 U8497 ( .A(n6165), .ZN(n7226) );
  INV_X1 U8498 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n7227) );
  NOR2_X1 U8499 ( .A1(n7279), .A2(n7227), .ZN(P2_U3261) );
  INV_X1 U8500 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n7228) );
  NOR2_X1 U8501 ( .A1(n7279), .A2(n7228), .ZN(P2_U3258) );
  INV_X1 U8502 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n7229) );
  NOR2_X1 U8503 ( .A1(n7279), .A2(n7229), .ZN(P2_U3260) );
  INV_X1 U8504 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n7230) );
  NOR2_X1 U8505 ( .A1(n7279), .A2(n7230), .ZN(P2_U3249) );
  INV_X1 U8506 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n7231) );
  NOR2_X1 U8507 ( .A1(n7279), .A2(n7231), .ZN(P2_U3259) );
  INV_X1 U8508 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U8509 ( .A1(n7232), .A2(P1_U3973), .ZN(n7233) );
  OAI21_X1 U8510 ( .B1(P1_U3973), .B2(n7234), .A(n7233), .ZN(P1_U3585) );
  INV_X1 U8511 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7245) );
  NAND2_X1 U8512 ( .A1(n8327), .A2(P1_U3973), .ZN(n7235) );
  OAI21_X1 U8513 ( .B1(n7245), .B2(P1_U3973), .A(n7235), .ZN(P1_U3563) );
  INV_X1 U8514 ( .A(n8151), .ZN(n8044) );
  NAND2_X1 U8515 ( .A1(n8044), .A2(P1_U3973), .ZN(n7236) );
  OAI21_X1 U8516 ( .B1(n7237), .B2(P1_U3973), .A(n7236), .ZN(P1_U3562) );
  INV_X1 U8517 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U8518 ( .A1(n9830), .A2(P1_U3973), .ZN(n7238) );
  OAI21_X1 U8519 ( .B1(n7636), .B2(P1_U3973), .A(n7238), .ZN(P1_U3571) );
  NAND4_X1 U8520 ( .A1(n8437), .A2(n8335), .A3(P2_STATE_REG_SCAN_IN), .A4(
        n7239), .ZN(n7240) );
  OAI21_X1 U8521 ( .B1(n7279), .B2(P2_D_REG_0__SCAN_IN), .A(n7240), .ZN(n7241)
         );
  INV_X1 U8522 ( .A(n7241), .ZN(P2_U3376) );
  AOI22_X1 U8523 ( .A1(n10476), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9997), .ZN(n7242) );
  OAI21_X1 U8524 ( .B1(n7248), .B2(n8027), .A(n7242), .ZN(P1_U3345) );
  INV_X1 U8525 ( .A(n7243), .ZN(n7249) );
  OAI222_X1 U8526 ( .A1(n9266), .A2(n7249), .B1(n9263), .B2(n7245), .C1(
        P2_U3151), .C2(n7244), .ZN(P2_U3286) );
  INV_X1 U8527 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7246) );
  OAI222_X1 U8528 ( .A1(n9266), .A2(n7248), .B1(n7247), .B2(P2_U3151), .C1(
        n7246), .C2(n9263), .ZN(P2_U3285) );
  INV_X1 U8529 ( .A(n9537), .ZN(n7250) );
  INV_X1 U8530 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7278) );
  OAI222_X1 U8531 ( .A1(n7250), .A2(P1_U3086), .B1(n8445), .B2(n7278), .C1(
        n7249), .C2(n10000), .ZN(P1_U3346) );
  INV_X1 U8532 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U8533 ( .A1(n9809), .A2(P1_U3973), .ZN(n7251) );
  OAI21_X1 U8534 ( .B1(n7782), .B2(P1_U3973), .A(n7251), .ZN(P1_U3573) );
  INV_X1 U8535 ( .A(n7252), .ZN(n7537) );
  NAND2_X1 U8536 ( .A1(n7537), .A2(P2_U3893), .ZN(n7253) );
  OAI21_X1 U8537 ( .B1(P2_U3893), .B2(n5566), .A(n7253), .ZN(P2_U3491) );
  NAND2_X1 U8538 ( .A1(n8931), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7254) );
  OAI21_X1 U8539 ( .B1(n9171), .B2(n8931), .A(n7254), .ZN(P2_U3506) );
  INV_X1 U8540 ( .A(n10670), .ZN(n7404) );
  INV_X1 U8541 ( .A(n7255), .ZN(n7256) );
  NAND2_X1 U8542 ( .A1(n7404), .A2(n7256), .ZN(n7259) );
  OAI21_X1 U8543 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7257), .A(n7340), .ZN(n7258) );
  AOI22_X1 U8544 ( .A1(n7259), .A2(n7258), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n7261) );
  NAND2_X1 U8545 ( .A1(n10661), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n7260) );
  OAI211_X1 U8546 ( .C1(n7335), .C2(n5350), .A(n7261), .B(n7260), .ZN(P2_U3182) );
  NAND2_X1 U8547 ( .A1(n7899), .A2(P2_U3893), .ZN(n7262) );
  OAI21_X1 U8548 ( .B1(P2_U3893), .B2(n7263), .A(n7262), .ZN(P2_U3497) );
  NAND2_X1 U8549 ( .A1(n7538), .A2(P2_U3893), .ZN(n7264) );
  OAI21_X1 U8550 ( .B1(P2_U3893), .B2(n7265), .A(n7264), .ZN(P2_U3493) );
  INV_X1 U8551 ( .A(n7266), .ZN(n7270) );
  AOI22_X1 U8552 ( .A1(n10360), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9997), .ZN(n7267) );
  OAI21_X1 U8553 ( .B1(n7270), .B2(n8027), .A(n7267), .ZN(P1_U3344) );
  AOI22_X1 U8554 ( .A1(n10449), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9997), .ZN(n7268) );
  OAI21_X1 U8555 ( .B1(n7276), .B2(n8027), .A(n7268), .ZN(P1_U3343) );
  INV_X1 U8556 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7271) );
  OAI222_X1 U8557 ( .A1(n9263), .A2(n7271), .B1(n9266), .B2(n7270), .C1(
        P2_U3151), .C2(n7269), .ZN(P2_U3284) );
  INV_X1 U8558 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7273) );
  NAND2_X1 U8559 ( .A1(n8000), .A2(P2_U3893), .ZN(n7272) );
  OAI21_X1 U8560 ( .B1(P2_U3893), .B2(n7273), .A(n7272), .ZN(P2_U3499) );
  INV_X1 U8561 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7274) );
  OAI222_X1 U8562 ( .A1(n9266), .A2(n7276), .B1(n7275), .B2(P2_U3151), .C1(
        n7274), .C2(n9263), .ZN(P2_U3283) );
  NAND2_X1 U8563 ( .A1(n8005), .A2(P2_U3893), .ZN(n7277) );
  OAI21_X1 U8564 ( .B1(P2_U3893), .B2(n7278), .A(n7277), .ZN(P2_U3500) );
  CLKBUF_X2 U8565 ( .A(n7279), .Z(n7305) );
  INV_X1 U8566 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n7280) );
  NOR2_X1 U8567 ( .A1(n7305), .A2(n7280), .ZN(P2_U3262) );
  INV_X1 U8568 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n7281) );
  NOR2_X1 U8569 ( .A1(n7305), .A2(n7281), .ZN(P2_U3234) );
  INV_X1 U8570 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n7282) );
  NOR2_X1 U8571 ( .A1(n7305), .A2(n7282), .ZN(P2_U3256) );
  INV_X1 U8572 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n7283) );
  NOR2_X1 U8573 ( .A1(n7305), .A2(n7283), .ZN(P2_U3257) );
  INV_X1 U8574 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n7284) );
  NOR2_X1 U8575 ( .A1(n7305), .A2(n7284), .ZN(P2_U3254) );
  INV_X1 U8576 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n7285) );
  NOR2_X1 U8577 ( .A1(n7305), .A2(n7285), .ZN(P2_U3253) );
  INV_X1 U8578 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n7286) );
  NOR2_X1 U8579 ( .A1(n7305), .A2(n7286), .ZN(P2_U3252) );
  INV_X1 U8580 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7287) );
  NOR2_X1 U8581 ( .A1(n7305), .A2(n7287), .ZN(P2_U3251) );
  INV_X1 U8582 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n7288) );
  NOR2_X1 U8583 ( .A1(n7305), .A2(n7288), .ZN(P2_U3250) );
  INV_X1 U8584 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n7289) );
  NOR2_X1 U8585 ( .A1(n7305), .A2(n7289), .ZN(P2_U3255) );
  INV_X1 U8586 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n7290) );
  NOR2_X1 U8587 ( .A1(n7305), .A2(n7290), .ZN(P2_U3248) );
  INV_X1 U8588 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n7291) );
  NOR2_X1 U8589 ( .A1(n7305), .A2(n7291), .ZN(P2_U3247) );
  INV_X1 U8590 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n7292) );
  NOR2_X1 U8591 ( .A1(n7305), .A2(n7292), .ZN(P2_U3246) );
  INV_X1 U8592 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n7293) );
  NOR2_X1 U8593 ( .A1(n7305), .A2(n7293), .ZN(P2_U3245) );
  INV_X1 U8594 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n7294) );
  NOR2_X1 U8595 ( .A1(n7305), .A2(n7294), .ZN(P2_U3243) );
  INV_X1 U8596 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7295) );
  NOR2_X1 U8597 ( .A1(n7305), .A2(n7295), .ZN(P2_U3242) );
  INV_X1 U8598 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n7296) );
  NOR2_X1 U8599 ( .A1(n7305), .A2(n7296), .ZN(P2_U3241) );
  INV_X1 U8600 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n7297) );
  NOR2_X1 U8601 ( .A1(n7305), .A2(n7297), .ZN(P2_U3240) );
  INV_X1 U8602 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n7298) );
  NOR2_X1 U8603 ( .A1(n7305), .A2(n7298), .ZN(P2_U3239) );
  INV_X1 U8604 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n7299) );
  NOR2_X1 U8605 ( .A1(n7305), .A2(n7299), .ZN(P2_U3238) );
  INV_X1 U8606 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n7300) );
  NOR2_X1 U8607 ( .A1(n7305), .A2(n7300), .ZN(P2_U3237) );
  INV_X1 U8608 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n7301) );
  NOR2_X1 U8609 ( .A1(n7305), .A2(n7301), .ZN(P2_U3236) );
  INV_X1 U8610 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n7302) );
  NOR2_X1 U8611 ( .A1(n7305), .A2(n7302), .ZN(P2_U3235) );
  INV_X1 U8612 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n7303) );
  NOR2_X1 U8613 ( .A1(n7305), .A2(n7303), .ZN(P2_U3263) );
  INV_X1 U8614 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n7304) );
  NOR2_X1 U8615 ( .A1(n7305), .A2(n7304), .ZN(P2_U3244) );
  NAND2_X1 U8616 ( .A1(n8895), .A2(P2_U3893), .ZN(n7306) );
  OAI21_X1 U8617 ( .B1(P2_U3893), .B2(n5592), .A(n7306), .ZN(P2_U3496) );
  AOI22_X1 U8618 ( .A1(n10433), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9997), .ZN(n7307) );
  OAI21_X1 U8619 ( .B1(n7310), .B2(n8027), .A(n7307), .ZN(P1_U3342) );
  INV_X1 U8620 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7308) );
  OAI222_X1 U8621 ( .A1(n9266), .A2(n7310), .B1(n7309), .B2(P2_U3151), .C1(
        n7308), .C2(n9263), .ZN(P2_U3282) );
  INV_X1 U8622 ( .A(n10661), .ZN(n7424) );
  INV_X1 U8623 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7326) );
  OAI21_X1 U8624 ( .B1(n7313), .B2(n7312), .A(n7311), .ZN(n7320) );
  AOI21_X1 U8625 ( .B1(n7316), .B2(n7315), .A(n7314), .ZN(n7317) );
  NOR2_X1 U8626 ( .A1(n10677), .A2(n7317), .ZN(n7319) );
  INV_X1 U8627 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10211) );
  OAI22_X1 U8628 ( .A1(n7335), .A2(n8449), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10211), .ZN(n7318) );
  AOI211_X1 U8629 ( .C1(n10671), .C2(n7320), .A(n7319), .B(n7318), .ZN(n7325)
         );
  OAI211_X1 U8630 ( .C1(n7323), .C2(n7322), .A(n7321), .B(n10670), .ZN(n7324)
         );
  OAI211_X1 U8631 ( .C1(n7424), .C2(n7326), .A(n7325), .B(n7324), .ZN(P2_U3184) );
  INV_X1 U8632 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7344) );
  OAI21_X1 U8633 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n7328), .A(n7327), .ZN(
        n7338) );
  AOI21_X1 U8634 ( .B1(n7331), .B2(n7330), .A(n7329), .ZN(n7332) );
  NOR2_X1 U8635 ( .A1(n10677), .A2(n7332), .ZN(n7337) );
  INV_X1 U8636 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7333) );
  OAI22_X1 U8637 ( .A1(n7335), .A2(n7334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7333), .ZN(n7336) );
  AOI211_X1 U8638 ( .C1(n10671), .C2(n7338), .A(n7337), .B(n7336), .ZN(n7343)
         );
  OAI211_X1 U8639 ( .C1(n7341), .C2(n7340), .A(n10670), .B(n7339), .ZN(n7342)
         );
  OAI211_X1 U8640 ( .C1(n7424), .C2(n7344), .A(n7343), .B(n7342), .ZN(P2_U3183) );
  INV_X1 U8641 ( .A(n7346), .ZN(n7345) );
  OAI22_X1 U8643 ( .A1(n10705), .A2(n7349), .B1(n10725), .B2(n7350), .ZN(n7356) );
  INV_X1 U8644 ( .A(n7351), .ZN(n7768) );
  NAND3_X1 U8645 ( .A1(n7346), .A2(n7550), .A3(n7383), .ZN(n7451) );
  OAI22_X1 U8646 ( .A1(n7768), .A2(n7350), .B1(n7448), .B2(n7774), .ZN(n7348)
         );
  NOR2_X1 U8647 ( .A1(n7348), .A2(n7451), .ZN(n7352) );
  NOR2_X1 U8648 ( .A1(n7348), .A2(n7347), .ZN(n8682) );
  AOI222_X1 U8649 ( .A1(n7351), .A2(n7453), .B1(n7554), .B2(n8722), .C1(n5118), 
        .C2(n10302), .ZN(n8681) );
  NOR2_X1 U8650 ( .A1(n8682), .A2(n8681), .ZN(n8680) );
  INV_X2 U8651 ( .A(n7448), .ZN(n7491) );
  AOI22_X1 U8652 ( .A1(n8722), .A2(n10228), .B1(n7777), .B2(n7491), .ZN(n7353)
         );
  XNOR2_X1 U8653 ( .A(n7353), .B(n7451), .ZN(n7354) );
  AOI21_X1 U8654 ( .B1(n7356), .B2(n7355), .A(n7461), .ZN(n7390) );
  NAND2_X1 U8655 ( .A1(n8448), .A2(P1_B_REG_SCAN_IN), .ZN(n7358) );
  MUX2_X1 U8656 ( .A(n7358), .B(P1_B_REG_SCAN_IN), .S(n7357), .Z(n7359) );
  INV_X1 U8657 ( .A(n8417), .ZN(n7361) );
  NAND2_X1 U8658 ( .A1(n7361), .A2(n8448), .ZN(n9982) );
  OAI21_X1 U8659 ( .B1(n9980), .B2(P1_D_REG_1__SCAN_IN), .A(n9982), .ZN(n7576)
         );
  INV_X1 U8660 ( .A(n7576), .ZN(n7695) );
  INV_X1 U8661 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U8662 ( .A1(n7372), .A2(n7360), .ZN(n7363) );
  NAND2_X1 U8663 ( .A1(n7361), .A2(n8273), .ZN(n7362) );
  NOR2_X1 U8664 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n7367) );
  NOR4_X1 U8665 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n7366) );
  NOR4_X1 U8666 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n7365) );
  NOR4_X1 U8667 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n7364) );
  NAND4_X1 U8668 ( .A1(n7367), .A2(n7366), .A3(n7365), .A4(n7364), .ZN(n7374)
         );
  NOR4_X1 U8669 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n7371) );
  NOR4_X1 U8670 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n7370) );
  NOR4_X1 U8671 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n7369) );
  NOR4_X1 U8672 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n7368) );
  NAND4_X1 U8673 ( .A1(n7371), .A2(n7370), .A3(n7369), .A4(n7368), .ZN(n7373)
         );
  OAI21_X1 U8674 ( .B1(n7374), .B2(n7373), .A(n7372), .ZN(n7574) );
  NAND2_X1 U8675 ( .A1(n10814), .A2(n7568), .ZN(n7379) );
  NOR2_X1 U8676 ( .A1(n7379), .A2(n9983), .ZN(n7375) );
  INV_X1 U8677 ( .A(n7377), .ZN(n7382) );
  OR2_X1 U8678 ( .A1(n10701), .A2(n9983), .ZN(n7380) );
  NOR2_X1 U8679 ( .A1(n7382), .A2(n7380), .ZN(n7387) );
  NAND2_X1 U8680 ( .A1(n7387), .A2(n9440), .ZN(n9404) );
  OR2_X1 U8681 ( .A1(n10702), .A2(n7961), .ZN(n7701) );
  NOR2_X1 U8682 ( .A1(n7701), .A2(n9983), .ZN(n7376) );
  NAND2_X1 U8683 ( .A1(n7377), .A2(n7376), .ZN(n7378) );
  AOI22_X1 U8684 ( .A1(n9372), .A2(n6363), .B1(n9411), .B2(n7777), .ZN(n7389)
         );
  NAND3_X1 U8685 ( .A1(n7380), .A2(n7379), .A3(n7701), .ZN(n7381) );
  NAND2_X1 U8686 ( .A1(n7382), .A2(n7381), .ZN(n7385) );
  OR2_X1 U8687 ( .A1(n7568), .A2(n7548), .ZN(n7384) );
  AND2_X1 U8688 ( .A1(n7384), .A2(n7383), .ZN(n7573) );
  NAND2_X1 U8689 ( .A1(n7385), .A2(n7573), .ZN(n7443) );
  INV_X1 U8690 ( .A(n7443), .ZN(n7386) );
  NAND2_X1 U8691 ( .A1(n7386), .A2(n7572), .ZN(n9373) );
  AND2_X2 U8692 ( .A1(n7387), .A2(n9998), .ZN(n9406) );
  AOI22_X1 U8693 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n9373), .B1(n9406), .B2(
        n7351), .ZN(n7388) );
  OAI211_X1 U8694 ( .C1(n7390), .C2(n9414), .A(n7389), .B(n7388), .ZN(P1_U3222) );
  INV_X1 U8695 ( .A(n7391), .ZN(n7392) );
  AOI21_X1 U8696 ( .B1(n7394), .B2(n7393), .A(n7392), .ZN(n7405) );
  NOR2_X1 U8697 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10178), .ZN(n7507) );
  XOR2_X1 U8698 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7395), .Z(n7400) );
  INV_X1 U8699 ( .A(n7396), .ZN(n7397) );
  AOI21_X1 U8700 ( .B1(n7532), .B2(n7398), .A(n7397), .ZN(n7399) );
  OAI22_X1 U8701 ( .A1(n7400), .A2(n8939), .B1(n10677), .B2(n7399), .ZN(n7401)
         );
  AOI211_X1 U8702 ( .C1(n5359), .C2(n10662), .A(n7507), .B(n7401), .ZN(n7403)
         );
  NAND2_X1 U8703 ( .A1(n10661), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n7402) );
  OAI211_X1 U8704 ( .C1(n7405), .C2(n7404), .A(n7403), .B(n7402), .ZN(P2_U3185) );
  INV_X1 U8705 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7425) );
  INV_X1 U8706 ( .A(n7406), .ZN(n7417) );
  INV_X1 U8707 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7407) );
  NOR2_X1 U8708 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7407), .ZN(n7599) );
  AOI21_X1 U8709 ( .B1(n7410), .B2(n7409), .A(n7408), .ZN(n7415) );
  AOI21_X1 U8710 ( .B1(n7413), .B2(n7412), .A(n7411), .ZN(n7414) );
  OAI22_X1 U8711 ( .A1(n7415), .A2(n10677), .B1(n8939), .B2(n7414), .ZN(n7416)
         );
  AOI211_X1 U8712 ( .C1(n7417), .C2(n10662), .A(n7599), .B(n7416), .ZN(n7423)
         );
  NAND2_X1 U8713 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  NAND3_X1 U8714 ( .A1(n7421), .A2(n10670), .A3(n7420), .ZN(n7422) );
  OAI211_X1 U8715 ( .C1(n7425), .C2(n7424), .A(n7423), .B(n7422), .ZN(P2_U3186) );
  AOI22_X1 U8716 ( .A1(n10364), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9997), .ZN(n7426) );
  OAI21_X1 U8717 ( .B1(n7429), .B2(n8027), .A(n7426), .ZN(P1_U3341) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7427) );
  OAI222_X1 U8719 ( .A1(n9266), .A2(n7429), .B1(n7428), .B2(P2_U3151), .C1(
        n7427), .C2(n9263), .ZN(P2_U3281) );
  INV_X1 U8720 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U8721 ( .A1(n7537), .A2(n7432), .ZN(n8472) );
  AND2_X1 U8722 ( .A1(n7044), .A2(n8472), .ZN(n8463) );
  INV_X1 U8723 ( .A(n8463), .ZN(n7430) );
  OAI21_X1 U8724 ( .B1(n9103), .B2(n9182), .A(n7430), .ZN(n7431) );
  OR2_X1 U8725 ( .A1(n7041), .A2(n9106), .ZN(n7634) );
  OAI211_X1 U8726 ( .C1(n8344), .C2(n7432), .A(n7431), .B(n7634), .ZN(n7435)
         );
  NAND2_X1 U8727 ( .A1(n7435), .A2(n10843), .ZN(n7433) );
  OAI21_X1 U8728 ( .B1(n10843), .B2(n7434), .A(n7433), .ZN(P2_U3390) );
  NAND2_X1 U8729 ( .A1(n7435), .A2(n8349), .ZN(n7436) );
  OAI21_X1 U8730 ( .B1(n8349), .B2(n7437), .A(n7436), .ZN(P2_U3459) );
  NAND2_X1 U8731 ( .A1(n7626), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7485) );
  NAND2_X1 U8732 ( .A1(n7485), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7439) );
  AOI22_X1 U8733 ( .A1(n7631), .A2(n10853), .B1(n10847), .B2(n7040), .ZN(n7438) );
  OAI211_X1 U8734 ( .C1(n8463), .C2(n8907), .A(n7439), .B(n7438), .ZN(P2_U3172) );
  INV_X1 U8735 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7440) );
  OAI222_X1 U8736 ( .A1(n9266), .A2(n7442), .B1(n6886), .B2(P2_U3151), .C1(
        n7440), .C2(n9263), .ZN(P2_U3280) );
  INV_X1 U8737 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7441) );
  OAI222_X1 U8738 ( .A1(P1_U3086), .A2(n9543), .B1(n10000), .B2(n7442), .C1(
        n7441), .C2(n8445), .ZN(P1_U3340) );
  NAND2_X1 U8739 ( .A1(n7443), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7444) );
  AOI22_X1 U8740 ( .A1(n10226), .A2(n8722), .B1(n7820), .B2(n7491), .ZN(n7445)
         );
  XNOR2_X1 U8741 ( .A(n7445), .B(n8767), .ZN(n7490) );
  OR2_X1 U8742 ( .A1(n7560), .A2(n7349), .ZN(n7447) );
  NAND2_X1 U8743 ( .A1(n7820), .A2(n8722), .ZN(n7446) );
  NAND2_X1 U8744 ( .A1(n7447), .A2(n7446), .ZN(n7488) );
  XNOR2_X1 U8745 ( .A(n7490), .B(n7488), .ZN(n7464) );
  NAND2_X1 U8746 ( .A1(n6363), .A2(n8722), .ZN(n7450) );
  OR2_X1 U8747 ( .A1(n10735), .A2(n7448), .ZN(n7449) );
  NAND2_X1 U8748 ( .A1(n7450), .A2(n7449), .ZN(n7452) );
  INV_X1 U8749 ( .A(n7451), .ZN(n9288) );
  XNOR2_X1 U8750 ( .A(n7452), .B(n9288), .ZN(n7456) );
  NAND2_X1 U8751 ( .A1(n6363), .A2(n7453), .ZN(n7455) );
  OR2_X1 U8752 ( .A1(n10735), .A2(n7350), .ZN(n7454) );
  AND2_X1 U8753 ( .A1(n7455), .A2(n7454), .ZN(n7457) );
  NAND2_X1 U8754 ( .A1(n7456), .A2(n7457), .ZN(n7462) );
  INV_X1 U8755 ( .A(n7456), .ZN(n7459) );
  INV_X1 U8756 ( .A(n7457), .ZN(n7458) );
  NAND2_X1 U8757 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  AND2_X1 U8758 ( .A1(n7462), .A2(n7460), .ZN(n9368) );
  NAND2_X1 U8759 ( .A1(n9367), .A2(n7462), .ZN(n7463) );
  NAND2_X1 U8760 ( .A1(n7463), .A2(n7464), .ZN(n7497) );
  OAI21_X1 U8761 ( .B1(n7464), .B2(n7463), .A(n7497), .ZN(n7465) );
  NAND2_X1 U8762 ( .A1(n7465), .A2(n9390), .ZN(n7470) );
  NAND2_X1 U8763 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9460) );
  INV_X1 U8764 ( .A(n9460), .ZN(n7468) );
  INV_X1 U8765 ( .A(n9406), .ZN(n9318) );
  OAI22_X1 U8766 ( .A1(n9318), .A2(n7767), .B1(n7466), .B2(n9404), .ZN(n7467)
         );
  AOI211_X1 U8767 ( .C1(n7820), .C2(n9411), .A(n7468), .B(n7467), .ZN(n7469)
         );
  OAI211_X1 U8768 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9409), .A(n7470), .B(
        n7469), .ZN(P1_U3218) );
  NAND2_X1 U8769 ( .A1(n9680), .A2(P1_U3973), .ZN(n7471) );
  OAI21_X1 U8770 ( .B1(n6072), .B2(P1_U3973), .A(n7471), .ZN(P1_U3580) );
  INV_X1 U8771 ( .A(n7536), .ZN(n7473) );
  OAI21_X1 U8772 ( .B1(n7631), .B2(n7474), .A(n7473), .ZN(n7476) );
  AOI21_X1 U8773 ( .B1(n7472), .B2(n7476), .A(n7475), .ZN(n7480) );
  INV_X1 U8774 ( .A(n10853), .ZN(n8920) );
  AOI22_X1 U8775 ( .A1(n10847), .A2(n7538), .B1(n10845), .B2(n7537), .ZN(n7477) );
  OAI21_X1 U8776 ( .B1(n8920), .B2(n7590), .A(n7477), .ZN(n7478) );
  AOI21_X1 U8777 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7485), .A(n7478), .ZN(
        n7479) );
  OAI21_X1 U8778 ( .B1(n7480), .B2(n8907), .A(n7479), .ZN(P2_U3162) );
  AOI21_X1 U8779 ( .B1(n7482), .B2(n7481), .A(n5028), .ZN(n7487) );
  AOI22_X1 U8780 ( .A1(n10847), .A2(n8932), .B1(n10845), .B2(n7040), .ZN(n7483) );
  OAI21_X1 U8781 ( .B1(n7544), .B2(n8920), .A(n7483), .ZN(n7484) );
  AOI21_X1 U8782 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7485), .A(n7484), .ZN(
        n7486) );
  OAI21_X1 U8783 ( .B1(n7487), .B2(n8907), .A(n7486), .ZN(P2_U3177) );
  INV_X1 U8784 ( .A(n7488), .ZN(n7489) );
  NAND2_X1 U8785 ( .A1(n7490), .A2(n7489), .ZN(n7495) );
  AND2_X1 U8786 ( .A1(n7497), .A2(n7495), .ZN(n7499) );
  NAND2_X1 U8787 ( .A1(n9426), .A2(n8722), .ZN(n7493) );
  NAND2_X1 U8788 ( .A1(n7834), .A2(n7491), .ZN(n7492) );
  NAND2_X1 U8789 ( .A1(n7493), .A2(n7492), .ZN(n7494) );
  XNOR2_X1 U8790 ( .A(n7494), .B(n8767), .ZN(n7674) );
  AOI22_X1 U8791 ( .A1(n9426), .A2(n7453), .B1(n8722), .B2(n7834), .ZN(n7677)
         );
  XNOR2_X1 U8792 ( .A(n7674), .B(n7677), .ZN(n7498) );
  NAND2_X1 U8793 ( .A1(n7497), .A2(n7496), .ZN(n7675) );
  OAI211_X1 U8794 ( .C1(n7499), .C2(n7498), .A(n9390), .B(n7675), .ZN(n7502)
         );
  AND2_X1 U8795 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10682) );
  OAI22_X1 U8796 ( .A1(n9318), .A2(n7560), .B1(n7785), .B2(n9404), .ZN(n7500)
         );
  AOI211_X1 U8797 ( .C1(n7834), .C2(n9411), .A(n10682), .B(n7500), .ZN(n7501)
         );
  OAI211_X1 U8798 ( .C1(n9409), .C2(n7831), .A(n7502), .B(n7501), .ZN(P1_U3230) );
  OAI211_X1 U8799 ( .C1(n7505), .C2(n7504), .A(n7503), .B(n10854), .ZN(n7509)
         );
  OAI22_X1 U8800 ( .A1(n8920), .A2(n7709), .B1(n7717), .B2(n8898), .ZN(n7506)
         );
  AOI211_X1 U8801 ( .C1(n10845), .C2(n7538), .A(n7507), .B(n7506), .ZN(n7508)
         );
  OAI211_X1 U8802 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7626), .A(n7509), .B(
        n7508), .ZN(P2_U3158) );
  INV_X1 U8803 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7511) );
  INV_X1 U8804 ( .A(n7510), .ZN(n7513) );
  INV_X1 U8805 ( .A(n9546), .ZN(n10423) );
  OAI222_X1 U8806 ( .A1(n8445), .A2(n7511), .B1(n8027), .B2(n7513), .C1(n10423), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8807 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7514) );
  OAI222_X1 U8808 ( .A1(n9263), .A2(n7514), .B1(n9266), .B2(n7513), .C1(
        P2_U3151), .C2(n7512), .ZN(P2_U3279) );
  XNOR2_X1 U8809 ( .A(n7515), .B(n8618), .ZN(n7516) );
  OAI222_X1 U8810 ( .A1(n9106), .A2(n7717), .B1(n9170), .B2(n7517), .C1(n9168), 
        .C2(n7516), .ZN(n7710) );
  INV_X1 U8811 ( .A(n7710), .ZN(n7535) );
  INV_X1 U8812 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U8813 ( .A1(n7037), .A2(n7519), .ZN(n7523) );
  INV_X1 U8814 ( .A(n7520), .ZN(n7521) );
  NAND2_X1 U8815 ( .A1(n9256), .A2(n7521), .ZN(n7522) );
  NAND2_X1 U8816 ( .A1(n7523), .A2(n7522), .ZN(n7524) );
  NAND2_X1 U8817 ( .A1(n7525), .A2(n7524), .ZN(n7628) );
  INV_X2 U8818 ( .A(n10837), .ZN(n10839) );
  OAI21_X1 U8819 ( .B1(n7526), .B2(n8618), .A(n7606), .ZN(n7712) );
  AND2_X1 U8820 ( .A1(n7527), .A2(n8649), .ZN(n7721) );
  INV_X1 U8821 ( .A(n7721), .ZN(n7528) );
  NAND2_X1 U8822 ( .A1(n7529), .A2(n7528), .ZN(n10835) );
  AOI22_X1 U8823 ( .A1(n9112), .A2(n7530), .B1(n9111), .B2(n10178), .ZN(n7531)
         );
  OAI21_X1 U8824 ( .B1(n7532), .B2(n10837), .A(n7531), .ZN(n7533) );
  AOI21_X1 U8825 ( .B1(n7712), .B2(n9115), .A(n7533), .ZN(n7534) );
  OAI21_X1 U8826 ( .B1(n7535), .B2(n10839), .A(n7534), .ZN(P2_U3230) );
  XNOR2_X1 U8827 ( .A(n8462), .B(n7044), .ZN(n7588) );
  XNOR2_X1 U8828 ( .A(n8462), .B(n7536), .ZN(n7539) );
  AOI222_X1 U8829 ( .A1(n9103), .A2(n7539), .B1(n7538), .B2(n9082), .C1(n7537), 
        .C2(n9080), .ZN(n7584) );
  OAI21_X1 U8830 ( .B1(n9165), .B2(n7588), .A(n7584), .ZN(n7592) );
  INV_X1 U8831 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7540) );
  OAI22_X1 U8832 ( .A1(n9249), .A2(n7590), .B1(n10843), .B2(n7540), .ZN(n7541)
         );
  AOI21_X1 U8833 ( .B1(n7592), .B2(n10843), .A(n7541), .ZN(n7542) );
  INV_X1 U8834 ( .A(n7542), .ZN(P2_U3393) );
  XNOR2_X1 U8835 ( .A(n7543), .B(n6122), .ZN(n7663) );
  NOR2_X1 U8836 ( .A1(n7544), .A2(n8344), .ZN(n7662) );
  XNOR2_X1 U8837 ( .A(n7545), .B(n6122), .ZN(n7546) );
  OAI222_X1 U8838 ( .A1(n9106), .A2(n7605), .B1(n9170), .B2(n7041), .C1(n9168), 
        .C2(n7546), .ZN(n7659) );
  AOI211_X1 U8839 ( .C1(n7663), .C2(n9182), .A(n7662), .B(n7659), .ZN(n10742)
         );
  NAND2_X1 U8840 ( .A1(n9175), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7547) );
  OAI21_X1 U8841 ( .B1(n10742), .B2(n9175), .A(n7547), .ZN(P2_U3461) );
  INV_X1 U8842 ( .A(n7548), .ZN(n7549) );
  NAND2_X1 U8843 ( .A1(n7550), .A2(n7549), .ZN(n7551) );
  AND2_X1 U8844 ( .A1(n7551), .A2(n10702), .ZN(n7552) );
  NAND2_X1 U8845 ( .A1(n7552), .A2(n10701), .ZN(n8207) );
  OR2_X1 U8846 ( .A1(n7553), .A2(n7563), .ZN(n10731) );
  NAND2_X1 U8847 ( .A1(n7351), .A2(n7554), .ZN(n7761) );
  NAND2_X1 U8848 ( .A1(n7766), .A2(n7761), .ZN(n7556) );
  NAND2_X1 U8849 ( .A1(n10705), .A2(n10725), .ZN(n7555) );
  NAND2_X1 U8850 ( .A1(n7556), .A2(n7555), .ZN(n10219) );
  NAND2_X1 U8851 ( .A1(n10219), .A2(n7557), .ZN(n7559) );
  NAND2_X1 U8852 ( .A1(n7767), .A2(n10735), .ZN(n7558) );
  NAND2_X1 U8853 ( .A1(n7559), .A2(n7558), .ZN(n7808) );
  NAND2_X1 U8854 ( .A1(n7560), .A2(n10744), .ZN(n7561) );
  NAND2_X1 U8855 ( .A1(n9426), .A2(n7834), .ZN(n7562) );
  XOR2_X1 U8856 ( .A(n7787), .B(n7788), .Z(n7708) );
  NAND2_X1 U8857 ( .A1(n6848), .A2(n7563), .ZN(n7566) );
  NAND2_X1 U8858 ( .A1(n7564), .A2(n10222), .ZN(n7565) );
  OAI21_X1 U8859 ( .B1(n7788), .B2(n6787), .A(n7567), .ZN(n7570) );
  INV_X1 U8860 ( .A(n7800), .ZN(n9424) );
  INV_X1 U8861 ( .A(n7568), .ZN(n7569) );
  AOI222_X1 U8862 ( .A1(n10230), .A2(n7570), .B1(n9424), .B2(n10225), .C1(
        n9426), .C2(n10227), .ZN(n7698) );
  OAI21_X1 U8863 ( .B1(n7830), .B2(n7784), .A(n9562), .ZN(n7571) );
  AND2_X1 U8864 ( .A1(n7830), .A2(n7784), .ZN(n7851) );
  OR2_X1 U8865 ( .A1(n7571), .A2(n7851), .ZN(n7700) );
  OAI211_X1 U8866 ( .C1(n10810), .C2(n7708), .A(n7698), .B(n7700), .ZN(n7582)
         );
  NAND3_X1 U8867 ( .A1(n7574), .A2(n7573), .A3(n7572), .ZN(n7693) );
  NAND2_X1 U8868 ( .A1(n7576), .A2(n7575), .ZN(n7577) );
  INV_X1 U8869 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9480) );
  OAI22_X1 U8870 ( .A1(n9928), .A2(n7784), .B1(n10819), .B2(n9480), .ZN(n7578)
         );
  AOI21_X1 U8871 ( .B1(n7582), .B2(n10819), .A(n7578), .ZN(n7579) );
  INV_X1 U8872 ( .A(n7579), .ZN(P1_U3527) );
  NAND2_X1 U8873 ( .A1(n10823), .A2(n9931), .ZN(n9977) );
  OAI22_X1 U8874 ( .A1(n9977), .A2(n7784), .B1(n10823), .B2(n6402), .ZN(n7581)
         );
  AOI21_X1 U8875 ( .B1(n7582), .B2(n10823), .A(n7581), .ZN(n7583) );
  INV_X1 U8876 ( .A(n7583), .ZN(P1_U3468) );
  INV_X1 U8877 ( .A(n9115), .ZN(n9101) );
  MUX2_X1 U8878 ( .A(n7331), .B(n7584), .S(n10837), .Z(n7587) );
  AOI22_X1 U8879 ( .A1(n9112), .A2(n7585), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9111), .ZN(n7586) );
  OAI211_X1 U8880 ( .C1(n7588), .C2(n9101), .A(n7587), .B(n7586), .ZN(P2_U3232) );
  INV_X1 U8881 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7589) );
  OAI22_X1 U8882 ( .A1(n7590), .A2(n9158), .B1(n8349), .B2(n7589), .ZN(n7591)
         );
  AOI21_X1 U8883 ( .B1(n7592), .B2(n8349), .A(n7591), .ZN(n7593) );
  INV_X1 U8884 ( .A(n7593), .ZN(P2_U3460) );
  INV_X1 U8885 ( .A(n7609), .ZN(n7602) );
  INV_X1 U8886 ( .A(n7619), .ZN(n7597) );
  AOI21_X1 U8887 ( .B1(n7503), .B2(n7595), .A(n7594), .ZN(n7596) );
  OAI21_X1 U8888 ( .B1(n7597), .B2(n7596), .A(n10854), .ZN(n7601) );
  OAI22_X1 U8889 ( .A1(n8920), .A2(n7669), .B1(n7915), .B2(n8898), .ZN(n7598)
         );
  AOI211_X1 U8890 ( .C1(n10845), .C2(n8932), .A(n7599), .B(n7598), .ZN(n7600)
         );
  OAI211_X1 U8891 ( .C1(n7602), .C2(n7626), .A(n7601), .B(n7600), .ZN(P2_U3170) );
  XNOR2_X1 U8892 ( .A(n7603), .B(n5252), .ZN(n7604) );
  OAI222_X1 U8893 ( .A1(n9106), .A2(n7915), .B1(n9170), .B2(n7605), .C1(n7604), 
        .C2(n9168), .ZN(n7670) );
  INV_X1 U8894 ( .A(n7670), .ZN(n7614) );
  NAND3_X1 U8895 ( .A1(n7606), .A2(n8486), .A3(n5252), .ZN(n7607) );
  NAND2_X1 U8896 ( .A1(n7608), .A2(n7607), .ZN(n7672) );
  AOI22_X1 U8897 ( .A1(n9112), .A2(n7610), .B1(n9111), .B2(n7609), .ZN(n7611)
         );
  OAI21_X1 U8898 ( .B1(n6869), .B2(n10837), .A(n7611), .ZN(n7612) );
  AOI21_X1 U8899 ( .B1(n7672), .B2(n9115), .A(n7612), .ZN(n7613) );
  OAI21_X1 U8900 ( .B1(n7614), .B2(n10839), .A(n7613), .ZN(P2_U3229) );
  INV_X1 U8901 ( .A(n7615), .ZN(n7637) );
  AOI22_X1 U8902 ( .A1(n10399), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9997), .ZN(n7616) );
  OAI21_X1 U8903 ( .B1(n7637), .B2(n8027), .A(n7616), .ZN(P1_U3338) );
  AOI22_X1 U8904 ( .A1(n10413), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9997), .ZN(n7617) );
  OAI21_X1 U8905 ( .B1(n7666), .B2(n8027), .A(n7617), .ZN(P1_U3337) );
  INV_X1 U8906 ( .A(n7722), .ZN(n7627) );
  AND3_X1 U8907 ( .A1(n7619), .A2(n7618), .A3(n7053), .ZN(n7620) );
  OAI21_X1 U8908 ( .B1(n7621), .B2(n7620), .A(n10854), .ZN(n7625) );
  NAND2_X1 U8909 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10495) );
  INV_X1 U8910 ( .A(n10495), .ZN(n7623) );
  OAI22_X1 U8911 ( .A1(n8920), .A2(n7906), .B1(n8914), .B2(n7717), .ZN(n7622)
         );
  AOI211_X1 U8912 ( .C1(n10847), .C2(n7899), .A(n7623), .B(n7622), .ZN(n7624)
         );
  OAI211_X1 U8913 ( .C1(n7627), .C2(n7626), .A(n7625), .B(n7624), .ZN(P2_U3167) );
  NOR3_X1 U8914 ( .A1(n8463), .A2(n7629), .A3(n7628), .ZN(n7630) );
  AOI21_X1 U8915 ( .B1(n9111), .B2(P2_REG3_REG_0__SCAN_IN), .A(n7630), .ZN(
        n7633) );
  AOI22_X1 U8916 ( .A1(n10839), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9112), .B2(
        n7631), .ZN(n7632) );
  OAI211_X1 U8917 ( .C1(n10839), .C2(n7634), .A(n7633), .B(n7632), .ZN(
        P2_U3233) );
  OAI222_X1 U8918 ( .A1(n9266), .A2(n7637), .B1(n9263), .B2(n7636), .C1(
        P2_U3151), .C2(n7635), .ZN(P2_U3278) );
  NOR2_X1 U8919 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7638) );
  AOI21_X1 U8920 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7638), .ZN(n10297) );
  NOR2_X1 U8921 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7639) );
  AOI21_X1 U8922 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7639), .ZN(n10294) );
  NOR2_X1 U8923 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7640) );
  AOI21_X1 U8924 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7640), .ZN(n10291) );
  NOR2_X1 U8925 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7641) );
  AOI21_X1 U8926 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7641), .ZN(n10288) );
  NOR2_X1 U8927 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7642) );
  AOI21_X1 U8928 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7642), .ZN(n10285) );
  NOR2_X1 U8929 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7643) );
  AOI21_X1 U8930 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7643), .ZN(n10282) );
  NOR2_X1 U8931 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7644) );
  AOI21_X1 U8932 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7644), .ZN(n10279) );
  NOR2_X1 U8933 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7645) );
  AOI21_X1 U8934 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7645), .ZN(n10276) );
  NOR2_X1 U8935 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7646) );
  AOI21_X1 U8936 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7646), .ZN(n10273) );
  NOR2_X1 U8937 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7647) );
  AOI21_X1 U8938 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7647), .ZN(n10270) );
  NOR2_X1 U8939 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7648) );
  AOI21_X1 U8940 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7648), .ZN(n10267) );
  NOR2_X1 U8941 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7649) );
  AOI21_X1 U8942 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7649), .ZN(n10264) );
  NOR2_X1 U8943 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7650) );
  AOI21_X1 U8944 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7650), .ZN(n10261) );
  NOR2_X1 U8945 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7651) );
  AOI21_X1 U8946 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7651), .ZN(n10258) );
  NAND2_X1 U8947 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10244) );
  INV_X1 U8948 ( .A(n10244), .ZN(n7652) );
  INV_X1 U8949 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U8950 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  AOI22_X1 U8951 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7652), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10243), .ZN(n10249) );
  NAND2_X1 U8952 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7653) );
  OAI21_X1 U8953 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7653), .ZN(n10248) );
  NOR2_X1 U8954 ( .A1(n10249), .A2(n10248), .ZN(n10247) );
  AOI21_X1 U8955 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10247), .ZN(n10252) );
  NAND2_X1 U8956 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7654) );
  OAI21_X1 U8957 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7654), .ZN(n10251) );
  NOR2_X1 U8958 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  AOI21_X1 U8959 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10250), .ZN(n10255) );
  NOR2_X1 U8960 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7655) );
  AOI21_X1 U8961 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7655), .ZN(n10254) );
  NAND2_X1 U8962 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  OAI21_X1 U8963 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10253), .ZN(n10257) );
  NAND2_X1 U8964 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U8965 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10256), .ZN(n10260) );
  NAND2_X1 U8966 ( .A1(n10261), .A2(n10260), .ZN(n10259) );
  OAI21_X1 U8967 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10259), .ZN(n10263) );
  NAND2_X1 U8968 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  OAI21_X1 U8969 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10262), .ZN(n10266) );
  NAND2_X1 U8970 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  OAI21_X1 U8971 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10265), .ZN(n10269) );
  NAND2_X1 U8972 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  OAI21_X1 U8973 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10268), .ZN(n10272) );
  NAND2_X1 U8974 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  OAI21_X1 U8975 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10271), .ZN(n10275) );
  NAND2_X1 U8976 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  OAI21_X1 U8977 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10274), .ZN(n10278) );
  NAND2_X1 U8978 ( .A1(n10279), .A2(n10278), .ZN(n10277) );
  OAI21_X1 U8979 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10277), .ZN(n10281) );
  NAND2_X1 U8980 ( .A1(n10282), .A2(n10281), .ZN(n10280) );
  OAI21_X1 U8981 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10280), .ZN(n10284) );
  NAND2_X1 U8982 ( .A1(n10285), .A2(n10284), .ZN(n10283) );
  OAI21_X1 U8983 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10283), .ZN(n10287) );
  NAND2_X1 U8984 ( .A1(n10288), .A2(n10287), .ZN(n10286) );
  OAI21_X1 U8985 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10286), .ZN(n10290) );
  NAND2_X1 U8986 ( .A1(n10291), .A2(n10290), .ZN(n10289) );
  OAI21_X1 U8987 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10289), .ZN(n10293) );
  NAND2_X1 U8988 ( .A1(n10294), .A2(n10293), .ZN(n10292) );
  OAI21_X1 U8989 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10292), .ZN(n10296) );
  NAND2_X1 U8990 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  OAI21_X1 U8991 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10295), .ZN(n7658) );
  XNOR2_X1 U8992 ( .A(n7656), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7657) );
  XNOR2_X1 U8993 ( .A(n7658), .B(n7657), .ZN(ADD_1068_U4) );
  NOR2_X1 U8994 ( .A1(n10829), .A2(n10211), .ZN(n7660) );
  AOI211_X1 U8995 ( .C1(n7662), .C2(n7661), .A(n7660), .B(n7659), .ZN(n7665)
         );
  AOI22_X1 U8996 ( .A1(n7663), .A2(n9115), .B1(n10839), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n7664) );
  OAI21_X1 U8997 ( .B1(n7665), .B2(n10839), .A(n7664), .ZN(P2_U3231) );
  INV_X1 U8998 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7668) );
  OAI222_X1 U8999 ( .A1(n9263), .A2(n7668), .B1(P2_U3151), .B2(n7667), .C1(
        n7666), .C2(n9266), .ZN(P2_U3277) );
  NOR2_X1 U9000 ( .A1(n7669), .A2(n8344), .ZN(n7671) );
  AOI211_X1 U9001 ( .C1(n9182), .C2(n7672), .A(n7671), .B(n7670), .ZN(n10754)
         );
  NAND2_X1 U9002 ( .A1(n9175), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7673) );
  OAI21_X1 U9003 ( .B1(n10754), .B2(n9175), .A(n7673), .ZN(P2_U3463) );
  INV_X1 U9004 ( .A(n7674), .ZN(n7676) );
  OAI21_X1 U9005 ( .B1(n7677), .B2(n7676), .A(n7675), .ZN(n7680) );
  AOI22_X1 U9006 ( .A1(n9425), .A2(n8722), .B1(n7684), .B2(n7491), .ZN(n7678)
         );
  XOR2_X1 U9007 ( .A(n8767), .B(n7678), .Z(n7679) );
  INV_X1 U9008 ( .A(n7729), .ZN(n7681) );
  NOR2_X1 U9009 ( .A1(n7728), .A2(n7681), .ZN(n7682) );
  AOI22_X1 U9010 ( .A1(n9425), .A2(n7453), .B1(n8722), .B2(n7684), .ZN(n7730)
         );
  XNOR2_X1 U9011 ( .A(n7682), .B(n7730), .ZN(n7691) );
  NAND2_X1 U9012 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9477) );
  INV_X1 U9013 ( .A(n9477), .ZN(n7683) );
  AOI21_X1 U9014 ( .B1(n9406), .B2(n9426), .A(n7683), .ZN(n7689) );
  NAND2_X1 U9015 ( .A1(n9411), .A2(n7684), .ZN(n7688) );
  INV_X1 U9016 ( .A(n7703), .ZN(n7685) );
  NAND2_X1 U9017 ( .A1(n9395), .A2(n7685), .ZN(n7687) );
  OR2_X1 U9018 ( .A1(n9404), .A2(n7800), .ZN(n7686) );
  NAND4_X1 U9019 ( .A1(n7689), .A2(n7688), .A3(n7687), .A4(n7686), .ZN(n7690)
         );
  AOI21_X1 U9020 ( .B1(n7691), .B2(n9390), .A(n7690), .ZN(n7692) );
  INV_X1 U9021 ( .A(n7692), .ZN(P1_U3227) );
  INV_X1 U9022 ( .A(n7693), .ZN(n7696) );
  NAND3_X1 U9023 ( .A1(n7696), .A2(n7695), .A3(n7694), .ZN(n7697) );
  NAND2_X1 U9024 ( .A1(n8207), .A2(n7763), .ZN(n10233) );
  MUX2_X1 U9025 ( .A(n7699), .B(n7698), .S(n10712), .Z(n7707) );
  INV_X1 U9026 ( .A(n7700), .ZN(n7705) );
  INV_X1 U9027 ( .A(n7701), .ZN(n7702) );
  OAI22_X1 U9028 ( .A1(n10237), .A2(n7784), .B1(n10709), .B2(n7703), .ZN(n7704) );
  AOI21_X1 U9029 ( .B1(n7705), .B2(n9844), .A(n7704), .ZN(n7706) );
  OAI211_X1 U9030 ( .C1(n7708), .C2(n9835), .A(n7707), .B(n7706), .ZN(P1_U3288) );
  INV_X1 U9031 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7714) );
  NOR2_X1 U9032 ( .A1(n7709), .A2(n8344), .ZN(n7711) );
  AOI211_X1 U9033 ( .C1(n9182), .C2(n7712), .A(n7711), .B(n7710), .ZN(n10752)
         );
  OR2_X1 U9034 ( .A1(n10752), .A2(n9175), .ZN(n7713) );
  OAI21_X1 U9035 ( .B1(n8349), .B2(n7714), .A(n7713), .ZN(P2_U3462) );
  XNOR2_X1 U9036 ( .A(n7715), .B(n8617), .ZN(n7720) );
  OAI21_X1 U9037 ( .B1(n7716), .B2(n8617), .A(n7916), .ZN(n7909) );
  OAI22_X1 U9038 ( .A1(n7930), .A2(n9106), .B1(n7717), .B2(n9170), .ZN(n7718)
         );
  AOI21_X1 U9039 ( .B1(n7909), .B2(n8120), .A(n7718), .ZN(n7719) );
  OAI21_X1 U9040 ( .B1(n7720), .B2(n9168), .A(n7719), .ZN(n7907) );
  INV_X1 U9041 ( .A(n7907), .ZN(n7727) );
  AND2_X1 U9042 ( .A1(n10837), .A2(n7721), .ZN(n8443) );
  AOI22_X1 U9043 ( .A1(n9112), .A2(n7723), .B1(n9111), .B2(n7722), .ZN(n7724)
         );
  OAI21_X1 U9044 ( .B1(n6959), .B2(n10837), .A(n7724), .ZN(n7725) );
  AOI21_X1 U9045 ( .B1(n7909), .B2(n8443), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9046 ( .B1(n7727), .B2(n10839), .A(n7726), .ZN(P2_U3228) );
  NAND2_X1 U9047 ( .A1(n7853), .A2(n7491), .ZN(n7732) );
  OR2_X1 U9048 ( .A1(n7800), .A2(n7350), .ZN(n7731) );
  NAND2_X1 U9049 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  XNOR2_X1 U9050 ( .A(n7733), .B(n7451), .ZN(n7736) );
  NAND2_X1 U9051 ( .A1(n7853), .A2(n8722), .ZN(n7735) );
  OR2_X1 U9052 ( .A1(n7800), .A2(n7349), .ZN(n7734) );
  NAND2_X1 U9053 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  INV_X1 U9054 ( .A(n7736), .ZN(n7739) );
  INV_X1 U9055 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U9056 ( .A1(n7739), .A2(n7738), .ZN(n7750) );
  NAND2_X1 U9057 ( .A1(n5029), .A2(n7750), .ZN(n7740) );
  XNOR2_X1 U9058 ( .A(n7751), .B(n7740), .ZN(n7748) );
  NAND2_X1 U9059 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10317) );
  INV_X1 U9060 ( .A(n10317), .ZN(n7741) );
  AOI21_X1 U9061 ( .B1(n9406), .B2(n9425), .A(n7741), .ZN(n7746) );
  NAND2_X1 U9062 ( .A1(n9411), .A2(n7853), .ZN(n7745) );
  INV_X1 U9063 ( .A(n7742), .ZN(n7852) );
  NAND2_X1 U9064 ( .A1(n9395), .A2(n7852), .ZN(n7744) );
  OR2_X1 U9065 ( .A1(n9404), .A2(n7752), .ZN(n7743) );
  NAND4_X1 U9066 ( .A1(n7746), .A2(n7745), .A3(n7744), .A4(n7743), .ZN(n7747)
         );
  AOI21_X1 U9067 ( .B1(n7748), .B2(n9390), .A(n7747), .ZN(n7749) );
  INV_X1 U9068 ( .A(n7749), .ZN(P1_U3239) );
  AOI22_X1 U9069 ( .A1(n9841), .A2(n7491), .B1(n8722), .B2(n9423), .ZN(n7753)
         );
  XOR2_X1 U9070 ( .A(n8767), .B(n7753), .Z(n8043) );
  AOI22_X1 U9071 ( .A1(n9841), .A2(n8722), .B1(n7453), .B2(n9423), .ZN(n8041)
         );
  XNOR2_X1 U9072 ( .A(n8043), .B(n5402), .ZN(n7754) );
  XNOR2_X1 U9073 ( .A(n8042), .B(n7754), .ZN(n7760) );
  NAND2_X1 U9074 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10333) );
  INV_X1 U9075 ( .A(n10333), .ZN(n7756) );
  NOR2_X1 U9076 ( .A1(n9404), .A2(n8151), .ZN(n7755) );
  AOI211_X1 U9077 ( .C1(n9406), .C2(n9424), .A(n7756), .B(n7755), .ZN(n7757)
         );
  OAI21_X1 U9078 ( .B1(n9409), .B2(n9837), .A(n7757), .ZN(n7758) );
  AOI21_X1 U9079 ( .B1(n9841), .B2(n9411), .A(n7758), .ZN(n7759) );
  OAI21_X1 U9080 ( .B1(n7760), .B2(n9414), .A(n7759), .ZN(P1_U3213) );
  XNOR2_X1 U9081 ( .A(n7762), .B(n7761), .ZN(n10723) );
  INV_X1 U9082 ( .A(n7763), .ZN(n7764) );
  NAND2_X1 U9083 ( .A1(n10235), .A2(n7764), .ZN(n8215) );
  XNOR2_X1 U9084 ( .A(n7766), .B(n7765), .ZN(n7770) );
  OAI22_X1 U9085 ( .A1(n7768), .A2(n9770), .B1(n7767), .B2(n10704), .ZN(n7769)
         );
  AOI21_X1 U9086 ( .B1(n7770), .B2(n10230), .A(n7769), .ZN(n7771) );
  OAI21_X1 U9087 ( .B1(n10723), .B2(n8207), .A(n7771), .ZN(n10726) );
  NAND2_X1 U9088 ( .A1(n10726), .A2(n10712), .ZN(n7779) );
  INV_X1 U9089 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9428) );
  OAI22_X1 U9090 ( .A1(n10235), .A2(n9428), .B1(n7772), .B2(n10709), .ZN(n7776) );
  INV_X1 U9091 ( .A(n10221), .ZN(n7773) );
  OAI211_X1 U9092 ( .C1(n10725), .C2(n7774), .A(n7773), .B(n9562), .ZN(n10724)
         );
  NOR2_X1 U9093 ( .A1(n9739), .A2(n10724), .ZN(n7775) );
  AOI211_X1 U9094 ( .C1(n9840), .C2(n7777), .A(n7776), .B(n7775), .ZN(n7778)
         );
  OAI211_X1 U9095 ( .C1(n10723), .C2(n8215), .A(n7779), .B(n7778), .ZN(
        P1_U3292) );
  INV_X1 U9096 ( .A(n7780), .ZN(n7783) );
  INV_X1 U9097 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7781) );
  OAI222_X1 U9098 ( .A1(n9552), .A2(P1_U3086), .B1(n10000), .B2(n7783), .C1(
        n7781), .C2(n8445), .ZN(P1_U3336) );
  OAI222_X1 U9099 ( .A1(n8655), .A2(P2_U3151), .B1(n9266), .B2(n7783), .C1(
        n9263), .C2(n7782), .ZN(P2_U3276) );
  NAND2_X1 U9100 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U9101 ( .A1(n7794), .A2(n7789), .ZN(n7848) );
  OR2_X1 U9102 ( .A1(n7853), .A2(n9424), .ZN(n7790) );
  NAND2_X1 U9103 ( .A1(n7847), .A2(n7790), .ZN(n7792) );
  NAND2_X1 U9104 ( .A1(n7791), .A2(n7858), .ZN(n7798) );
  NAND2_X1 U9105 ( .A1(n7792), .A2(n7798), .ZN(n7868) );
  OAI21_X1 U9106 ( .B1(n7792), .B2(n7798), .A(n7868), .ZN(n9843) );
  INV_X1 U9107 ( .A(n7853), .ZN(n10767) );
  NAND2_X1 U9108 ( .A1(n7851), .A2(n10767), .ZN(n7850) );
  AOI21_X1 U9109 ( .B1(n7850), .B2(n9841), .A(n9819), .ZN(n7793) );
  AND2_X1 U9110 ( .A1(n7793), .A2(n7986), .ZN(n9845) );
  NAND2_X1 U9111 ( .A1(n7795), .A2(n7794), .ZN(n7797) );
  OR2_X1 U9112 ( .A1(n7797), .A2(n7798), .ZN(n7859) );
  INV_X1 U9113 ( .A(n7859), .ZN(n7796) );
  AOI21_X1 U9114 ( .B1(n7798), .B2(n7797), .A(n7796), .ZN(n7799) );
  OAI222_X1 U9115 ( .A1(n10704), .A2(n8151), .B1(n9770), .B2(n7800), .C1(
        n10716), .C2(n7799), .ZN(n9836) );
  AOI211_X1 U9116 ( .C1(n10806), .C2(n9843), .A(n9845), .B(n9836), .ZN(n7807)
         );
  INV_X1 U9117 ( .A(n9928), .ZN(n8093) );
  NOR2_X1 U9118 ( .A1(n10819), .A2(n6431), .ZN(n7801) );
  AOI21_X1 U9119 ( .B1(n9841), .B2(n8093), .A(n7801), .ZN(n7802) );
  OAI21_X1 U9120 ( .B1(n7807), .B2(n10818), .A(n7802), .ZN(P1_U3529) );
  INV_X1 U9121 ( .A(n9977), .ZN(n7805) );
  INV_X1 U9122 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7803) );
  NOR2_X1 U9123 ( .A1(n10823), .A2(n7803), .ZN(n7804) );
  AOI21_X1 U9124 ( .B1(n9841), .B2(n7805), .A(n7804), .ZN(n7806) );
  OAI21_X1 U9125 ( .B1(n7807), .B2(n10820), .A(n7806), .ZN(P1_U3474) );
  XNOR2_X1 U9126 ( .A(n7809), .B(n7808), .ZN(n10747) );
  INV_X1 U9127 ( .A(n8207), .ZN(n10738) );
  NAND2_X1 U9128 ( .A1(n10747), .A2(n10738), .ZN(n7817) );
  INV_X1 U9129 ( .A(n7809), .ZN(n7810) );
  XNOR2_X1 U9130 ( .A(n7811), .B(n7810), .ZN(n7815) );
  NAND2_X1 U9131 ( .A1(n6363), .A2(n10227), .ZN(n7813) );
  NAND2_X1 U9132 ( .A1(n9426), .A2(n10225), .ZN(n7812) );
  NAND2_X1 U9133 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  AOI21_X1 U9134 ( .B1(n7815), .B2(n10230), .A(n7814), .ZN(n7816) );
  AND2_X1 U9135 ( .A1(n7817), .A2(n7816), .ZN(n10749) );
  INV_X1 U9136 ( .A(n8215), .ZN(n7824) );
  AOI21_X1 U9137 ( .B1(n10220), .B2(n7820), .A(n9819), .ZN(n7818) );
  NAND2_X1 U9138 ( .A1(n7818), .A2(n7827), .ZN(n10743) );
  INV_X1 U9139 ( .A(n10709), .ZN(n9822) );
  AOI22_X1 U9140 ( .A1(n4932), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9822), .B2(
        n7819), .ZN(n7822) );
  NAND2_X1 U9141 ( .A1(n9840), .A2(n7820), .ZN(n7821) );
  OAI211_X1 U9142 ( .C1(n10743), .C2(n9739), .A(n7822), .B(n7821), .ZN(n7823)
         );
  AOI21_X1 U9143 ( .B1(n10747), .B2(n7824), .A(n7823), .ZN(n7825) );
  OAI21_X1 U9144 ( .B1(n10749), .B2(n4932), .A(n7825), .ZN(P1_U3290) );
  XNOR2_X1 U9145 ( .A(n7826), .B(n7838), .ZN(n10759) );
  NAND2_X1 U9146 ( .A1(n7827), .A2(n7834), .ZN(n7828) );
  NAND2_X1 U9147 ( .A1(n7828), .A2(n9562), .ZN(n7829) );
  OR2_X1 U9148 ( .A1(n7830), .A2(n7829), .ZN(n10755) );
  INV_X1 U9149 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7832) );
  OAI22_X1 U9150 ( .A1(n10235), .A2(n7832), .B1(n7831), .B2(n10709), .ZN(n7833) );
  AOI21_X1 U9151 ( .B1(n9840), .B2(n7834), .A(n7833), .ZN(n7835) );
  OAI21_X1 U9152 ( .B1(n10755), .B2(n9739), .A(n7835), .ZN(n7842) );
  NAND2_X1 U9153 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  XNOR2_X1 U9154 ( .A(n7839), .B(n7838), .ZN(n7840) );
  AOI222_X1 U9155 ( .A1(n10230), .A2(n7840), .B1(n9425), .B2(n10225), .C1(
        n10226), .C2(n10227), .ZN(n10756) );
  NOR2_X1 U9156 ( .A1(n10756), .A2(n4932), .ZN(n7841) );
  AOI211_X1 U9157 ( .C1(n9842), .C2(n10759), .A(n7842), .B(n7841), .ZN(n7843)
         );
  INV_X1 U9158 ( .A(n7843), .ZN(P1_U3289) );
  XOR2_X1 U9159 ( .A(n7844), .B(n7848), .Z(n7845) );
  AOI222_X1 U9160 ( .A1(n10230), .A2(n7845), .B1(n9423), .B2(n10225), .C1(
        n9425), .C2(n10227), .ZN(n10766) );
  MUX2_X1 U9161 ( .A(n7846), .B(n10766), .S(n10712), .Z(n7857) );
  OAI21_X1 U9162 ( .B1(n7849), .B2(n7848), .A(n7847), .ZN(n10769) );
  OAI211_X1 U9163 ( .C1(n7851), .C2(n10767), .A(n9562), .B(n7850), .ZN(n10765)
         );
  AOI22_X1 U9164 ( .A1(n9840), .A2(n7853), .B1(n7852), .B2(n9822), .ZN(n7854)
         );
  OAI21_X1 U9165 ( .B1(n10765), .B2(n9739), .A(n7854), .ZN(n7855) );
  AOI21_X1 U9166 ( .B1(n10769), .B2(n9842), .A(n7855), .ZN(n7856) );
  NAND2_X1 U9167 ( .A1(n7857), .A2(n7856), .ZN(P1_U3287) );
  NAND2_X1 U9168 ( .A1(n7859), .A2(n7858), .ZN(n7993) );
  NAND2_X1 U9169 ( .A1(n7993), .A2(n7994), .ZN(n7992) );
  NAND2_X1 U9170 ( .A1(n7992), .A2(n7860), .ZN(n7864) );
  NAND2_X1 U9171 ( .A1(n7862), .A2(n7861), .ZN(n7870) );
  INV_X1 U9172 ( .A(n7870), .ZN(n7863) );
  XNOR2_X1 U9173 ( .A(n7864), .B(n7863), .ZN(n7866) );
  NOR2_X1 U9174 ( .A1(n8151), .A2(n9770), .ZN(n7865) );
  AOI21_X1 U9175 ( .B1(n7866), .B2(n10230), .A(n7865), .ZN(n10783) );
  OR2_X1 U9176 ( .A1(n9841), .A2(n9423), .ZN(n7867) );
  NAND2_X1 U9177 ( .A1(n7868), .A2(n7867), .ZN(n7985) );
  OR2_X1 U9178 ( .A1(n8060), .A2(n8044), .ZN(n7869) );
  NAND2_X1 U9179 ( .A1(n7983), .A2(n7869), .ZN(n7871) );
  NAND2_X1 U9180 ( .A1(n7871), .A2(n7870), .ZN(n7885) );
  OAI21_X1 U9181 ( .B1(n7871), .B2(n7870), .A(n7885), .ZN(n10786) );
  INV_X1 U9182 ( .A(n8142), .ZN(n10784) );
  XNOR2_X1 U9183 ( .A(n7987), .B(n10784), .ZN(n7872) );
  INV_X1 U9184 ( .A(n8250), .ZN(n9422) );
  AOI22_X1 U9185 ( .A1(n7872), .A2(n9562), .B1(n10225), .B2(n9422), .ZN(n10782) );
  OAI22_X1 U9186 ( .A1(n10712), .A2(n7873), .B1(n8148), .B2(n10709), .ZN(n7874) );
  AOI21_X1 U9187 ( .B1(n8142), .B2(n9840), .A(n7874), .ZN(n7875) );
  OAI21_X1 U9188 ( .B1(n10782), .B2(n9739), .A(n7875), .ZN(n7876) );
  AOI21_X1 U9189 ( .B1(n10786), .B2(n9842), .A(n7876), .ZN(n7877) );
  OAI21_X1 U9190 ( .B1(n10783), .B2(n4932), .A(n7877), .ZN(P1_U3284) );
  OAI21_X1 U9191 ( .B1(n7880), .B2(n7879), .A(n7878), .ZN(n7883) );
  NAND2_X1 U9192 ( .A1(n9421), .A2(n10225), .ZN(n7881) );
  OAI21_X1 U9193 ( .B1(n8138), .B2(n9770), .A(n7881), .ZN(n7882) );
  AOI21_X1 U9194 ( .B1(n7883), .B2(n10230), .A(n7882), .ZN(n10792) );
  OR2_X1 U9195 ( .A1(n8142), .A2(n8327), .ZN(n7884) );
  NAND2_X1 U9196 ( .A1(n7885), .A2(n7884), .ZN(n7887) );
  OAI21_X1 U9197 ( .B1(n7887), .B2(n7886), .A(n7963), .ZN(n10795) );
  NAND2_X1 U9198 ( .A1(n10795), .A2(n9842), .ZN(n7893) );
  OAI22_X1 U9199 ( .A1(n10712), .A2(n7888), .B1(n8329), .B2(n10709), .ZN(n7891) );
  INV_X1 U9200 ( .A(n8331), .ZN(n10793) );
  INV_X1 U9201 ( .A(n7975), .ZN(n8019) );
  OAI211_X1 U9202 ( .C1(n10793), .C2(n7889), .A(n8019), .B(n9562), .ZN(n10791)
         );
  NOR2_X1 U9203 ( .A1(n10791), .A2(n9739), .ZN(n7890) );
  AOI211_X1 U9204 ( .C1(n9840), .C2(n8331), .A(n7891), .B(n7890), .ZN(n7892)
         );
  OAI211_X1 U9205 ( .C1(n4932), .C2(n10792), .A(n7893), .B(n7892), .ZN(
        P1_U3283) );
  NAND2_X1 U9206 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  AOI21_X1 U9207 ( .B1(n7897), .B2(n7896), .A(n8907), .ZN(n7905) );
  NAND2_X1 U9208 ( .A1(n10856), .A2(n7935), .ZN(n7903) );
  NAND2_X1 U9209 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10511) );
  INV_X1 U9210 ( .A(n10511), .ZN(n7898) );
  AOI21_X1 U9211 ( .B1(n10847), .B2(n8000), .A(n7898), .ZN(n7902) );
  NAND2_X1 U9212 ( .A1(n10853), .A2(n7934), .ZN(n7901) );
  NAND2_X1 U9213 ( .A1(n10845), .A2(n7899), .ZN(n7900) );
  NAND4_X1 U9214 ( .A1(n7903), .A2(n7902), .A3(n7901), .A4(n7900), .ZN(n7904)
         );
  OR2_X1 U9215 ( .A1(n7905), .A2(n7904), .ZN(P2_U3153) );
  INV_X1 U9216 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7911) );
  NOR2_X1 U9217 ( .A1(n7906), .A2(n8344), .ZN(n7908) );
  AOI211_X1 U9218 ( .C1(n8156), .C2(n7909), .A(n7908), .B(n7907), .ZN(n10762)
         );
  OR2_X1 U9219 ( .A1(n10762), .A2(n9175), .ZN(n7910) );
  OAI21_X1 U9220 ( .B1(n8349), .B2(n7911), .A(n7910), .ZN(P2_U3464) );
  OR2_X1 U9221 ( .A1(n7912), .A2(n8622), .ZN(n7927) );
  INV_X1 U9222 ( .A(n7927), .ZN(n7913) );
  AOI21_X1 U9223 ( .B1(n8622), .B2(n7912), .A(n7913), .ZN(n7914) );
  OAI222_X1 U9224 ( .A1(n9106), .A2(n8899), .B1(n9170), .B2(n7915), .C1(n9168), 
        .C2(n7914), .ZN(n8037) );
  INV_X1 U9225 ( .A(n8037), .ZN(n7923) );
  NAND3_X1 U9226 ( .A1(n7916), .A2(n8490), .A3(n5254), .ZN(n7917) );
  NAND2_X1 U9227 ( .A1(n7918), .A2(n7917), .ZN(n8039) );
  NOR2_X1 U9228 ( .A1(n8981), .A2(n8036), .ZN(n7921) );
  INV_X1 U9229 ( .A(n8901), .ZN(n7919) );
  OAI22_X1 U9230 ( .A1(n10837), .A2(n6870), .B1(n7919), .B2(n10829), .ZN(n7920) );
  AOI211_X1 U9231 ( .C1(n8039), .C2(n9115), .A(n7921), .B(n7920), .ZN(n7922)
         );
  OAI21_X1 U9232 ( .B1(n7923), .B2(n10839), .A(n7922), .ZN(P2_U3227) );
  AND2_X1 U9233 ( .A1(n7924), .A2(n7925), .ZN(n7948) );
  NAND3_X1 U9234 ( .A1(n7927), .A2(n8620), .A3(n7926), .ZN(n7928) );
  AND2_X1 U9235 ( .A1(n7948), .A2(n7928), .ZN(n7929) );
  OAI222_X1 U9236 ( .A1(n9106), .A2(n8133), .B1(n9170), .B2(n7930), .C1(n9168), 
        .C2(n7929), .ZN(n8063) );
  INV_X1 U9237 ( .A(n8063), .ZN(n7940) );
  INV_X1 U9238 ( .A(n7942), .ZN(n7931) );
  AOI21_X1 U9239 ( .B1(n7933), .B2(n7932), .A(n7931), .ZN(n8065) );
  INV_X1 U9240 ( .A(n7934), .ZN(n8499) );
  NOR2_X1 U9241 ( .A1(n8981), .A2(n8499), .ZN(n7938) );
  INV_X1 U9242 ( .A(n7935), .ZN(n7936) );
  OAI22_X1 U9243 ( .A1(n10837), .A2(n10508), .B1(n7936), .B2(n10829), .ZN(
        n7937) );
  AOI211_X1 U9244 ( .C1(n8065), .C2(n9115), .A(n7938), .B(n7937), .ZN(n7939)
         );
  OAI21_X1 U9245 ( .B1(n7940), .B2(n10839), .A(n7939), .ZN(P2_U3226) );
  NAND2_X1 U9246 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  XNOR2_X1 U9247 ( .A(n7943), .B(n8621), .ZN(n8029) );
  INV_X1 U9248 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U9249 ( .A1(n7924), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U9250 ( .A1(n7946), .A2(n7945), .ZN(n8129) );
  NAND3_X1 U9251 ( .A1(n7948), .A2(n8621), .A3(n7947), .ZN(n7949) );
  NAND2_X1 U9252 ( .A1(n8129), .A2(n7949), .ZN(n7952) );
  NAND2_X1 U9253 ( .A1(n8929), .A2(n9080), .ZN(n7950) );
  OAI21_X1 U9254 ( .B1(n8289), .B2(n9106), .A(n7950), .ZN(n7951) );
  AOI21_X1 U9255 ( .B1(n7952), .B2(n9103), .A(n7951), .ZN(n8033) );
  MUX2_X1 U9256 ( .A(n7953), .B(n8033), .S(n10837), .Z(n7955) );
  AOI22_X1 U9257 ( .A1(n9112), .A2(n8030), .B1(n9111), .B2(n8003), .ZN(n7954)
         );
  OAI211_X1 U9258 ( .C1(n8029), .C2(n9101), .A(n7955), .B(n7954), .ZN(P2_U3225) );
  INV_X1 U9259 ( .A(n7956), .ZN(n7960) );
  OAI222_X1 U9260 ( .A1(n9266), .A2(n7960), .B1(n7958), .B2(P2_U3151), .C1(
        n7957), .C2(n9263), .ZN(P2_U3275) );
  INV_X1 U9261 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7959) );
  OAI222_X1 U9262 ( .A1(P1_U3086), .A2(n7961), .B1(n10000), .B2(n7960), .C1(
        n7959), .C2(n8445), .ZN(P1_U3335) );
  OR2_X1 U9263 ( .A1(n8331), .A2(n9422), .ZN(n7962) );
  NAND2_X1 U9264 ( .A1(n7963), .A2(n7962), .ZN(n8011) );
  NAND2_X1 U9265 ( .A1(n8390), .A2(n9421), .ZN(n7964) );
  NAND2_X1 U9266 ( .A1(n8011), .A2(n7964), .ZN(n7966) );
  OR2_X1 U9267 ( .A1(n8390), .A2(n9421), .ZN(n7965) );
  NAND2_X1 U9268 ( .A1(n7966), .A2(n7965), .ZN(n8072) );
  XOR2_X1 U9269 ( .A(n8072), .B(n7967), .Z(n10807) );
  INV_X1 U9270 ( .A(n10807), .ZN(n7981) );
  INV_X1 U9271 ( .A(n7967), .ZN(n7970) );
  NAND2_X1 U9272 ( .A1(n8012), .A2(n7968), .ZN(n7969) );
  NAND2_X1 U9273 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  NAND3_X1 U9274 ( .A1(n7972), .A2(n7971), .A3(n10230), .ZN(n7974) );
  AOI22_X1 U9275 ( .A1(n10227), .A2(n9421), .B1(n9419), .B2(n10225), .ZN(n7973) );
  NAND2_X1 U9276 ( .A1(n7974), .A2(n7973), .ZN(n10805) );
  INV_X1 U9277 ( .A(n8390), .ZN(n8090) );
  OAI211_X1 U9278 ( .C1(n10803), .C2(n8018), .A(n9562), .B(n8080), .ZN(n10802)
         );
  OAI22_X1 U9279 ( .A1(n10712), .A2(n7976), .B1(n8266), .B2(n10709), .ZN(n7977) );
  AOI21_X1 U9280 ( .B1(n8268), .B2(n9840), .A(n7977), .ZN(n7978) );
  OAI21_X1 U9281 ( .B1(n10802), .B2(n9739), .A(n7978), .ZN(n7979) );
  AOI21_X1 U9282 ( .B1(n10805), .B2(n10235), .A(n7979), .ZN(n7980) );
  OAI21_X1 U9283 ( .B1(n7981), .B2(n9835), .A(n7980), .ZN(P1_U3281) );
  OAI222_X1 U9284 ( .A1(n9266), .A2(n8026), .B1(n8471), .B2(P2_U3151), .C1(
        n7982), .C2(n9263), .ZN(P2_U3274) );
  OAI21_X1 U9285 ( .B1(n7985), .B2(n7984), .A(n7983), .ZN(n10777) );
  AOI21_X1 U9286 ( .B1(n7986), .B2(n8060), .A(n9819), .ZN(n7988) );
  NAND2_X1 U9287 ( .A1(n7988), .A2(n7987), .ZN(n10774) );
  OAI22_X1 U9288 ( .A1(n10712), .A2(n7989), .B1(n8058), .B2(n10709), .ZN(n7990) );
  AOI21_X1 U9289 ( .B1(n8060), .B2(n9840), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9290 ( .B1(n10774), .B2(n9739), .A(n7991), .ZN(n7997) );
  OAI21_X1 U9291 ( .B1(n7994), .B2(n7993), .A(n7992), .ZN(n7995) );
  AOI222_X1 U9292 ( .A1(n10230), .A2(n7995), .B1(n8327), .B2(n10225), .C1(
        n9423), .C2(n10227), .ZN(n10775) );
  NOR2_X1 U9293 ( .A1(n10775), .A2(n4932), .ZN(n7996) );
  AOI211_X1 U9294 ( .C1(n9842), .C2(n10777), .A(n7997), .B(n7996), .ZN(n7998)
         );
  INV_X1 U9295 ( .A(n7998), .ZN(P1_U3285) );
  XNOR2_X1 U9296 ( .A(n8001), .B(n8000), .ZN(n8002) );
  XNOR2_X1 U9297 ( .A(n7999), .B(n8002), .ZN(n8010) );
  NAND2_X1 U9298 ( .A1(n10856), .A2(n8003), .ZN(n8007) );
  NAND2_X1 U9299 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10527) );
  INV_X1 U9300 ( .A(n10527), .ZN(n8004) );
  AOI21_X1 U9301 ( .B1(n10847), .B2(n8005), .A(n8004), .ZN(n8006) );
  OAI211_X1 U9302 ( .C1(n8899), .C2(n8914), .A(n8007), .B(n8006), .ZN(n8008)
         );
  AOI21_X1 U9303 ( .B1(n8030), .B2(n10853), .A(n8008), .ZN(n8009) );
  OAI21_X1 U9304 ( .B1(n8010), .B2(n8907), .A(n8009), .ZN(P2_U3161) );
  XNOR2_X1 U9305 ( .A(n8011), .B(n8014), .ZN(n8086) );
  OAI21_X1 U9306 ( .B1(n8014), .B2(n8013), .A(n8012), .ZN(n8016) );
  OAI22_X1 U9307 ( .A1(n8385), .A2(n10704), .B1(n8250), .B2(n9770), .ZN(n8015)
         );
  AOI21_X1 U9308 ( .B1(n8016), .B2(n10230), .A(n8015), .ZN(n8017) );
  OAI21_X1 U9309 ( .B1(n8086), .B2(n8207), .A(n8017), .ZN(n8087) );
  NAND2_X1 U9310 ( .A1(n8087), .A2(n10712), .ZN(n8024) );
  AOI211_X1 U9311 ( .C1(n8390), .C2(n8019), .A(n9819), .B(n8018), .ZN(n8088)
         );
  NOR2_X1 U9312 ( .A1(n8090), .A2(n10237), .ZN(n8022) );
  OAI22_X1 U9313 ( .A1(n10712), .A2(n8020), .B1(n8388), .B2(n10709), .ZN(n8021) );
  AOI211_X1 U9314 ( .C1(n8088), .C2(n9844), .A(n8022), .B(n8021), .ZN(n8023)
         );
  OAI211_X1 U9315 ( .C1(n8086), .C2(n8215), .A(n8024), .B(n8023), .ZN(P1_U3282) );
  INV_X1 U9316 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8025) );
  OAI222_X1 U9317 ( .A1(P1_U3086), .A2(n8028), .B1(n8027), .B2(n8026), .C1(
        n8025), .C2(n8445), .ZN(P1_U3334) );
  OR2_X1 U9318 ( .A1(n8029), .A2(n9165), .ZN(n8032) );
  NAND2_X1 U9319 ( .A1(n8030), .A2(n9173), .ZN(n8031) );
  OR2_X1 U9320 ( .A1(n8349), .A2(n8034), .ZN(n8035) );
  OAI21_X1 U9321 ( .B1(n10781), .B2(n9175), .A(n8035), .ZN(P2_U3467) );
  NOR2_X1 U9322 ( .A1(n8036), .A2(n8344), .ZN(n8038) );
  AOI211_X1 U9323 ( .C1(n9182), .C2(n8039), .A(n8038), .B(n8037), .ZN(n10764)
         );
  NAND2_X1 U9324 ( .A1(n9175), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8040) );
  OAI21_X1 U9325 ( .B1(n10764), .B2(n9175), .A(n8040), .ZN(P2_U3465) );
  OAI22_X1 U9326 ( .A1(n5342), .A2(n7350), .B1(n8151), .B2(n7349), .ZN(n8054)
         );
  AOI22_X1 U9327 ( .A1(n8060), .A2(n7491), .B1(n8722), .B2(n8044), .ZN(n8045)
         );
  XNOR2_X1 U9328 ( .A(n8045), .B(n7451), .ZN(n8048) );
  INV_X1 U9329 ( .A(n8048), .ZN(n8046) );
  NAND2_X1 U9330 ( .A1(n8049), .A2(n8048), .ZN(n8143) );
  INV_X1 U9331 ( .A(n8054), .ZN(n8051) );
  INV_X1 U9332 ( .A(n8144), .ZN(n8052) );
  AOI21_X1 U9333 ( .B1(n8054), .B2(n8053), .A(n8052), .ZN(n8062) );
  NAND2_X1 U9334 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10349) );
  INV_X1 U9335 ( .A(n10349), .ZN(n8056) );
  NOR2_X1 U9336 ( .A1(n9404), .A2(n8138), .ZN(n8055) );
  AOI211_X1 U9337 ( .C1(n9406), .C2(n9423), .A(n8056), .B(n8055), .ZN(n8057)
         );
  OAI21_X1 U9338 ( .B1(n9409), .B2(n8058), .A(n8057), .ZN(n8059) );
  AOI21_X1 U9339 ( .B1(n8060), .B2(n9411), .A(n8059), .ZN(n8061) );
  OAI21_X1 U9340 ( .B1(n8062), .B2(n9414), .A(n8061), .ZN(P1_U3221) );
  INV_X1 U9341 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8067) );
  NOR2_X1 U9342 ( .A1(n8499), .A2(n8344), .ZN(n8064) );
  AOI211_X1 U9343 ( .C1(n8065), .C2(n9182), .A(n8064), .B(n8063), .ZN(n10773)
         );
  OR2_X1 U9344 ( .A1(n10773), .A2(n9175), .ZN(n8066) );
  OAI21_X1 U9345 ( .B1(n8349), .B2(n8067), .A(n8066), .ZN(P2_U3466) );
  XNOR2_X1 U9346 ( .A(n8069), .B(n8068), .ZN(n8070) );
  AOI222_X1 U9347 ( .A1(n10230), .A2(n8070), .B1(n9418), .B2(n10225), .C1(
        n9420), .C2(n10227), .ZN(n10813) );
  NAND2_X1 U9348 ( .A1(n8268), .A2(n9420), .ZN(n8071) );
  OR2_X1 U9349 ( .A1(n8268), .A2(n9420), .ZN(n8073) );
  AND2_X1 U9350 ( .A1(n8075), .A2(n8076), .ZN(n10811) );
  INV_X1 U9351 ( .A(n10811), .ZN(n8078) );
  NAND3_X1 U9352 ( .A1(n8078), .A2(n9842), .A3(n8077), .ZN(n8085) );
  OAI22_X1 U9353 ( .A1(n10712), .A2(n8079), .B1(n8374), .B2(n10709), .ZN(n8083) );
  INV_X1 U9354 ( .A(n8080), .ZN(n8081) );
  OAI211_X1 U9355 ( .C1(n10815), .C2(n8081), .A(n5022), .B(n9562), .ZN(n10812)
         );
  NOR2_X1 U9356 ( .A1(n10812), .A2(n9739), .ZN(n8082) );
  AOI211_X1 U9357 ( .C1(n9840), .C2(n8376), .A(n8083), .B(n8082), .ZN(n8084)
         );
  OAI211_X1 U9358 ( .C1(n4932), .C2(n10813), .A(n8085), .B(n8084), .ZN(
        P1_U3280) );
  INV_X1 U9359 ( .A(n10731), .ZN(n10746) );
  INV_X1 U9360 ( .A(n8086), .ZN(n8089) );
  AOI211_X1 U9361 ( .C1(n10746), .C2(n8089), .A(n8088), .B(n8087), .ZN(n8095)
         );
  OAI22_X1 U9362 ( .A1(n8090), .A2(n9977), .B1(n10823), .B2(n6487), .ZN(n8091)
         );
  INV_X1 U9363 ( .A(n8091), .ZN(n8092) );
  OAI21_X1 U9364 ( .B1(n8095), .B2(n10820), .A(n8092), .ZN(P1_U3486) );
  INV_X1 U9365 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9525) );
  AOI22_X1 U9366 ( .A1(n8390), .A2(n8093), .B1(n10818), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n8094) );
  OAI21_X1 U9367 ( .B1(n8095), .B2(n10818), .A(n8094), .ZN(P1_U3533) );
  XNOR2_X1 U9368 ( .A(n8097), .B(n8096), .ZN(n8103) );
  NAND2_X1 U9369 ( .A1(n10856), .A2(n8135), .ZN(n8100) );
  NAND2_X1 U9370 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10543) );
  INV_X1 U9371 ( .A(n10543), .ZN(n8098) );
  AOI21_X1 U9372 ( .B1(n10847), .B2(n8928), .A(n8098), .ZN(n8099) );
  OAI211_X1 U9373 ( .C1(n8133), .C2(n8914), .A(n8100), .B(n8099), .ZN(n8101)
         );
  AOI21_X1 U9374 ( .B1(n8165), .B2(n10853), .A(n8101), .ZN(n8102) );
  OAI21_X1 U9375 ( .B1(n8103), .B2(n8907), .A(n8102), .ZN(P2_U3171) );
  INV_X1 U9376 ( .A(n8104), .ZN(n8108) );
  OAI222_X1 U9377 ( .A1(n9263), .A2(n8106), .B1(n9266), .B2(n8108), .C1(
        P2_U3151), .C2(n8105), .ZN(P2_U3273) );
  INV_X1 U9378 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8107) );
  OAI222_X1 U9379 ( .A1(n8109), .A2(P1_U3086), .B1(n10000), .B2(n8108), .C1(
        n8107), .C2(n8445), .ZN(P1_U3333) );
  XNOR2_X1 U9380 ( .A(n8110), .B(n8626), .ZN(n8157) );
  OAI22_X1 U9381 ( .A1(n8289), .A2(n9170), .B1(n8400), .B2(n9106), .ZN(n8119)
         );
  AND2_X1 U9382 ( .A1(n8112), .A2(n8111), .ZN(n8117) );
  NAND2_X1 U9383 ( .A1(n8129), .A2(n8128), .ZN(n8113) );
  NAND2_X1 U9384 ( .A1(n8113), .A2(n8625), .ZN(n8131) );
  NAND3_X1 U9385 ( .A1(n8131), .A2(n8115), .A3(n8114), .ZN(n8116) );
  AOI21_X1 U9386 ( .B1(n8117), .B2(n8116), .A(n9168), .ZN(n8118) );
  AOI211_X1 U9387 ( .C1(n8120), .C2(n8157), .A(n8119), .B(n8118), .ZN(n8159)
         );
  INV_X1 U9388 ( .A(n5856), .ZN(n8122) );
  AOI22_X1 U9389 ( .A1(n10839), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n9111), .B2(
        n8285), .ZN(n8121) );
  OAI21_X1 U9390 ( .B1(n8122), .B2(n8981), .A(n8121), .ZN(n8123) );
  AOI21_X1 U9391 ( .B1(n8157), .B2(n8443), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9392 ( .B1(n8159), .B2(n10839), .A(n8124), .ZN(P2_U3223) );
  OR2_X1 U9393 ( .A1(n8125), .A2(n8625), .ZN(n8127) );
  NAND2_X1 U9394 ( .A1(n8125), .A2(n8625), .ZN(n8126) );
  NAND2_X1 U9395 ( .A1(n8127), .A2(n8126), .ZN(n8162) );
  NAND3_X1 U9396 ( .A1(n8129), .A2(n5281), .A3(n8128), .ZN(n8130) );
  AND2_X1 U9397 ( .A1(n8131), .A2(n8130), .ZN(n8132) );
  OAI222_X1 U9398 ( .A1(n9106), .A2(n8359), .B1(n9170), .B2(n8133), .C1(n9168), 
        .C2(n8132), .ZN(n8163) );
  INV_X1 U9399 ( .A(n8163), .ZN(n8134) );
  MUX2_X1 U9400 ( .A(n10539), .B(n8134), .S(n10837), .Z(n8137) );
  AOI22_X1 U9401 ( .A1(n8165), .A2(n9112), .B1(n9111), .B2(n8135), .ZN(n8136)
         );
  OAI211_X1 U9402 ( .C1(n9101), .C2(n8162), .A(n8137), .B(n8136), .ZN(P2_U3224) );
  NAND2_X1 U9403 ( .A1(n8142), .A2(n7491), .ZN(n8140) );
  OR2_X1 U9404 ( .A1(n8138), .A2(n7350), .ZN(n8139) );
  NAND2_X1 U9405 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  XNOR2_X1 U9406 ( .A(n8141), .B(n8767), .ZN(n8244) );
  AOI22_X1 U9407 ( .A1(n8142), .A2(n8722), .B1(n7453), .B2(n8327), .ZN(n8242)
         );
  XNOR2_X1 U9408 ( .A(n8244), .B(n8242), .ZN(n8146) );
  NAND2_X1 U9409 ( .A1(n8145), .A2(n8146), .ZN(n8246) );
  OAI21_X1 U9410 ( .B1(n8146), .B2(n8145), .A(n8246), .ZN(n8147) );
  NAND2_X1 U9411 ( .A1(n8147), .A2(n9390), .ZN(n8155) );
  INV_X1 U9412 ( .A(n8148), .ZN(n8153) );
  NOR2_X1 U9413 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8149), .ZN(n9504) );
  AOI21_X1 U9414 ( .B1(n9372), .B2(n9422), .A(n9504), .ZN(n8150) );
  OAI21_X1 U9415 ( .B1(n8151), .B2(n9318), .A(n8150), .ZN(n8152) );
  AOI21_X1 U9416 ( .B1(n8153), .B2(n9395), .A(n8152), .ZN(n8154) );
  OAI211_X1 U9417 ( .C1(n10784), .C2(n9398), .A(n8155), .B(n8154), .ZN(
        P1_U3231) );
  AOI22_X1 U9418 ( .A1(n8157), .A2(n8156), .B1(n9173), .B2(n5856), .ZN(n8158)
         );
  AND2_X1 U9419 ( .A1(n8159), .A2(n8158), .ZN(n10799) );
  OR2_X1 U9420 ( .A1(n8349), .A2(n8160), .ZN(n8161) );
  OAI21_X1 U9421 ( .B1(n10799), .B2(n9175), .A(n8161), .ZN(P2_U3469) );
  INV_X1 U9422 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8167) );
  NOR2_X1 U9423 ( .A1(n8162), .A2(n9165), .ZN(n8164) );
  AOI211_X1 U9424 ( .C1(n9173), .C2(n8165), .A(n8164), .B(n8163), .ZN(n10790)
         );
  OR2_X1 U9425 ( .A1(n10790), .A2(n9175), .ZN(n8166) );
  OAI21_X1 U9426 ( .B1(n8349), .B2(n8167), .A(n8166), .ZN(P2_U3468) );
  NAND2_X1 U9427 ( .A1(n8376), .A2(n9419), .ZN(n8168) );
  NAND2_X1 U9428 ( .A1(n8198), .A2(n8197), .ZN(n8200) );
  NAND2_X1 U9429 ( .A1(n8433), .A2(n9418), .ZN(n8170) );
  NAND2_X1 U9430 ( .A1(n8200), .A2(n8170), .ZN(n8304) );
  XNOR2_X1 U9431 ( .A(n8304), .B(n8173), .ZN(n8276) );
  INV_X1 U9432 ( .A(n8276), .ZN(n8183) );
  OAI21_X1 U9433 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8174) );
  NAND2_X1 U9434 ( .A1(n8174), .A2(n10230), .ZN(n8177) );
  OAI22_X1 U9435 ( .A1(n8371), .A2(n9770), .B1(n9403), .B2(n10704), .ZN(n8175)
         );
  INV_X1 U9436 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U9437 ( .A1(n8177), .A2(n8176), .ZN(n8274) );
  AOI211_X1 U9438 ( .C1(n9412), .C2(n8208), .A(n9819), .B(n9816), .ZN(n8275)
         );
  NAND2_X1 U9439 ( .A1(n8275), .A2(n9844), .ZN(n8180) );
  INV_X1 U9440 ( .A(n9408), .ZN(n8178) );
  AOI22_X1 U9441 ( .A1(n4932), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8178), .B2(
        n9822), .ZN(n8179) );
  OAI211_X1 U9442 ( .C1(n5338), .C2(n10237), .A(n8180), .B(n8179), .ZN(n8181)
         );
  AOI21_X1 U9443 ( .B1(n10712), .B2(n8274), .A(n8181), .ZN(n8182) );
  OAI21_X1 U9444 ( .B1(n8183), .B2(n9835), .A(n8182), .ZN(P1_U3278) );
  XNOR2_X1 U9445 ( .A(n8184), .B(n8628), .ZN(n8185) );
  OAI222_X1 U9446 ( .A1(n9106), .A2(n8868), .B1(n9170), .B2(n8359), .C1(n9168), 
        .C2(n8185), .ZN(n8229) );
  INV_X1 U9447 ( .A(n8229), .ZN(n8193) );
  OAI21_X1 U9448 ( .B1(n8187), .B2(n8628), .A(n8186), .ZN(n8231) );
  INV_X1 U9449 ( .A(n8188), .ZN(n8364) );
  NOR2_X1 U9450 ( .A1(n8364), .A2(n8981), .ZN(n8191) );
  INV_X1 U9451 ( .A(n8361), .ZN(n8189) );
  OAI22_X1 U9452 ( .A1(n10837), .A2(n10572), .B1(n8189), .B2(n10829), .ZN(
        n8190) );
  AOI211_X1 U9453 ( .C1(n8231), .C2(n9115), .A(n8191), .B(n8190), .ZN(n8192)
         );
  OAI21_X1 U9454 ( .B1(n8193), .B2(n10839), .A(n8192), .ZN(P2_U3222) );
  INV_X1 U9455 ( .A(n8216), .ZN(n8196) );
  NAND2_X1 U9456 ( .A1(n9997), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8194) );
  OAI211_X1 U9457 ( .C1(n8196), .C2(n10000), .A(n8195), .B(n8194), .ZN(
        P1_U3332) );
  OR2_X1 U9458 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  NAND2_X1 U9459 ( .A1(n8200), .A2(n8199), .ZN(n8293) );
  OAI21_X1 U9460 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8205) );
  OAI22_X1 U9461 ( .A1(n8370), .A2(n9770), .B1(n8427), .B2(n10704), .ZN(n8204)
         );
  AOI21_X1 U9462 ( .B1(n8205), .B2(n10230), .A(n8204), .ZN(n8206) );
  OAI21_X1 U9463 ( .B1(n8293), .B2(n8207), .A(n8206), .ZN(n8294) );
  NAND2_X1 U9464 ( .A1(n8294), .A2(n10235), .ZN(n8214) );
  INV_X1 U9465 ( .A(n8208), .ZN(n8209) );
  AOI211_X1 U9466 ( .C1(n8433), .C2(n5022), .A(n9819), .B(n8209), .ZN(n8295)
         );
  NOR2_X1 U9467 ( .A1(n8302), .A2(n10237), .ZN(n8212) );
  OAI22_X1 U9468 ( .A1(n10712), .A2(n8210), .B1(n8431), .B2(n10709), .ZN(n8211) );
  AOI211_X1 U9469 ( .C1(n8295), .C2(n9844), .A(n8212), .B(n8211), .ZN(n8213)
         );
  OAI211_X1 U9470 ( .C1(n8293), .C2(n8215), .A(n8214), .B(n8213), .ZN(P1_U3279) );
  NAND2_X1 U9471 ( .A1(n8216), .A2(n9267), .ZN(n8218) );
  NAND2_X1 U9472 ( .A1(n8217), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8661) );
  OAI211_X1 U9473 ( .C1(n8219), .C2(n9263), .A(n8218), .B(n8661), .ZN(P2_U3272) );
  XNOR2_X1 U9474 ( .A(n8222), .B(n5009), .ZN(n8223) );
  OAI222_X1 U9475 ( .A1(n9170), .A2(n8400), .B1(n9106), .B2(n9169), .C1(n8223), 
        .C2(n9168), .ZN(n8337) );
  INV_X1 U9476 ( .A(n8337), .ZN(n8228) );
  XNOR2_X1 U9477 ( .A(n8224), .B(n5009), .ZN(n8338) );
  INV_X1 U9478 ( .A(n8402), .ZN(n8343) );
  AOI22_X1 U9479 ( .A1(n10839), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9111), .B2(
        n8396), .ZN(n8225) );
  OAI21_X1 U9480 ( .B1(n8343), .B2(n8981), .A(n8225), .ZN(n8226) );
  AOI21_X1 U9481 ( .B1(n8338), .B2(n9115), .A(n8226), .ZN(n8227) );
  OAI21_X1 U9482 ( .B1(n8228), .B2(n10839), .A(n8227), .ZN(P2_U3221) );
  INV_X1 U9483 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8233) );
  NOR2_X1 U9484 ( .A1(n8364), .A2(n8344), .ZN(n8230) );
  AOI211_X1 U9485 ( .C1(n9182), .C2(n8231), .A(n8230), .B(n8229), .ZN(n10801)
         );
  OR2_X1 U9486 ( .A1(n10801), .A2(n9175), .ZN(n8232) );
  OAI21_X1 U9487 ( .B1(n8349), .B2(n8233), .A(n8232), .ZN(P2_U3470) );
  XNOR2_X1 U9488 ( .A(n8234), .B(n8520), .ZN(n8345) );
  XNOR2_X1 U9489 ( .A(n8235), .B(n8520), .ZN(n8236) );
  OAI222_X1 U9490 ( .A1(n9106), .A2(n8915), .B1(n9170), .B2(n8868), .C1(n9168), 
        .C2(n8236), .ZN(n8347) );
  INV_X1 U9491 ( .A(n8237), .ZN(n8873) );
  INV_X1 U9492 ( .A(n8870), .ZN(n8238) );
  OAI22_X1 U9493 ( .A1(n8873), .A2(n10831), .B1(n8238), .B2(n10829), .ZN(n8239) );
  OAI21_X1 U9494 ( .B1(n8347), .B2(n8239), .A(n10837), .ZN(n8241) );
  NAND2_X1 U9495 ( .A1(n10839), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8240) );
  OAI211_X1 U9496 ( .C1(n8345), .C2(n9101), .A(n8241), .B(n8240), .ZN(P2_U3220) );
  INV_X1 U9497 ( .A(n8242), .ZN(n8243) );
  OR2_X1 U9498 ( .A1(n8244), .A2(n8243), .ZN(n8245) );
  NAND2_X1 U9499 ( .A1(n8331), .A2(n7491), .ZN(n8248) );
  OR2_X1 U9500 ( .A1(n8250), .A2(n7350), .ZN(n8247) );
  NAND2_X1 U9501 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  XNOR2_X1 U9502 ( .A(n8249), .B(n8767), .ZN(n8319) );
  NAND2_X1 U9503 ( .A1(n8331), .A2(n8722), .ZN(n8252) );
  OR2_X1 U9504 ( .A1(n8250), .A2(n7349), .ZN(n8251) );
  NAND2_X1 U9505 ( .A1(n8252), .A2(n8251), .ZN(n8323) );
  NOR2_X1 U9506 ( .A1(n8319), .A2(n8323), .ZN(n8258) );
  NAND2_X1 U9507 ( .A1(n8390), .A2(n7491), .ZN(n8254) );
  NAND2_X1 U9508 ( .A1(n9421), .A2(n8722), .ZN(n8253) );
  NAND2_X1 U9509 ( .A1(n8254), .A2(n8253), .ZN(n8255) );
  XNOR2_X1 U9510 ( .A(n8255), .B(n9288), .ZN(n8260) );
  AND2_X1 U9511 ( .A1(n9421), .A2(n7453), .ZN(n8256) );
  AOI21_X1 U9512 ( .B1(n8390), .B2(n8722), .A(n8256), .ZN(n8259) );
  NOR2_X1 U9513 ( .A1(n8260), .A2(n8259), .ZN(n8382) );
  AOI21_X1 U9514 ( .B1(n8319), .B2(n8323), .A(n8382), .ZN(n8257) );
  OAI22_X1 U9515 ( .A1(n10803), .A2(n7350), .B1(n8385), .B2(n7349), .ZN(n8367)
         );
  NAND2_X1 U9516 ( .A1(n8268), .A2(n7491), .ZN(n8262) );
  NAND2_X1 U9517 ( .A1(n9420), .A2(n8722), .ZN(n8261) );
  NAND2_X1 U9518 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  XNOR2_X1 U9519 ( .A(n8263), .B(n7451), .ZN(n8368) );
  XOR2_X1 U9520 ( .A(n8367), .B(n8368), .Z(n8365) );
  XOR2_X1 U9521 ( .A(n8366), .B(n8365), .Z(n8270) );
  NAND2_X1 U9522 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n10463) );
  OAI21_X1 U9523 ( .B1(n9404), .B2(n8370), .A(n10463), .ZN(n8264) );
  AOI21_X1 U9524 ( .B1(n9406), .B2(n9421), .A(n8264), .ZN(n8265) );
  OAI21_X1 U9525 ( .B1(n9409), .B2(n8266), .A(n8265), .ZN(n8267) );
  AOI21_X1 U9526 ( .B1(n8268), .B2(n9411), .A(n8267), .ZN(n8269) );
  OAI21_X1 U9527 ( .B1(n8270), .B2(n9414), .A(n8269), .ZN(P1_U3224) );
  INV_X1 U9528 ( .A(n8271), .ZN(n8336) );
  INV_X1 U9529 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8272) );
  OAI222_X1 U9530 ( .A1(n8273), .A2(P1_U3086), .B1(n10000), .B2(n8336), .C1(
        n8272), .C2(n8445), .ZN(P1_U3331) );
  INV_X1 U9531 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8277) );
  AOI211_X1 U9532 ( .C1(n8276), .C2(n10806), .A(n8275), .B(n8274), .ZN(n8279)
         );
  MUX2_X1 U9533 ( .A(n8277), .B(n8279), .S(n10823), .Z(n8278) );
  OAI21_X1 U9534 ( .B1(n5338), .B2(n9977), .A(n8278), .ZN(P1_U3498) );
  MUX2_X1 U9535 ( .A(n10381), .B(n8279), .S(n10819), .Z(n8280) );
  OAI21_X1 U9536 ( .B1(n5338), .B2(n9928), .A(n8280), .ZN(P1_U3537) );
  INV_X1 U9537 ( .A(n8281), .ZN(n8283) );
  OAI222_X1 U9538 ( .A1(n9266), .A2(n8447), .B1(P2_U3151), .B2(n8283), .C1(
        n8282), .C2(n9263), .ZN(P2_U3270) );
  AOI21_X1 U9539 ( .B1(n8928), .B2(n8284), .A(n4930), .ZN(n8292) );
  NAND2_X1 U9540 ( .A1(n10856), .A2(n8285), .ZN(n8288) );
  NAND2_X1 U9541 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10560) );
  INV_X1 U9542 ( .A(n10560), .ZN(n8286) );
  AOI21_X1 U9543 ( .B1(n10847), .B2(n8927), .A(n8286), .ZN(n8287) );
  OAI211_X1 U9544 ( .C1(n8289), .C2(n8914), .A(n8288), .B(n8287), .ZN(n8290)
         );
  AOI21_X1 U9545 ( .B1(n5856), .B2(n10853), .A(n8290), .ZN(n8291) );
  OAI21_X1 U9546 ( .B1(n8292), .B2(n8907), .A(n8291), .ZN(P2_U3157) );
  INV_X1 U9547 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8297) );
  INV_X1 U9548 ( .A(n8293), .ZN(n8296) );
  AOI211_X1 U9549 ( .C1(n8296), .C2(n10746), .A(n8295), .B(n8294), .ZN(n8299)
         );
  MUX2_X1 U9550 ( .A(n8297), .B(n8299), .S(n10823), .Z(n8298) );
  OAI21_X1 U9551 ( .B1(n8302), .B2(n9977), .A(n8298), .ZN(P1_U3495) );
  MUX2_X1 U9552 ( .A(n8300), .B(n8299), .S(n10819), .Z(n8301) );
  OAI21_X1 U9553 ( .B1(n8302), .B2(n9928), .A(n8301), .ZN(P1_U3536) );
  OR2_X1 U9554 ( .A1(n9412), .A2(n9829), .ZN(n8303) );
  NAND2_X1 U9555 ( .A1(n8304), .A2(n8303), .ZN(n8306) );
  NAND2_X1 U9556 ( .A1(n9412), .A2(n9829), .ZN(n8305) );
  INV_X1 U9557 ( .A(n9403), .ZN(n9417) );
  NAND2_X1 U9558 ( .A1(n9930), .A2(n9417), .ZN(n8307) );
  XNOR2_X1 U9559 ( .A(n9576), .B(n8308), .ZN(n9925) );
  INV_X1 U9560 ( .A(n9925), .ZN(n8318) );
  INV_X1 U9561 ( .A(n8309), .ZN(n8311) );
  INV_X1 U9562 ( .A(n9805), .ZN(n8310) );
  AOI21_X1 U9563 ( .B1(n8311), .B2(n9575), .A(n8310), .ZN(n8312) );
  OAI222_X1 U9564 ( .A1(n10704), .A2(n9332), .B1(n9770), .B2(n9403), .C1(
        n10716), .C2(n8312), .ZN(n9923) );
  NAND2_X1 U9565 ( .A1(n9923), .A2(n10235), .ZN(n8317) );
  INV_X1 U9566 ( .A(n9930), .ZN(n9825) );
  NAND2_X1 U9567 ( .A1(n9825), .A2(n9816), .ZN(n9817) );
  AOI211_X1 U9568 ( .C1(n9577), .C2(n9817), .A(n9819), .B(n5344), .ZN(n9924)
         );
  INV_X1 U9569 ( .A(n9577), .ZN(n9978) );
  NOR2_X1 U9570 ( .A1(n9978), .A2(n10237), .ZN(n8315) );
  OAI22_X1 U9571 ( .A1(n10712), .A2(n8313), .B1(n9335), .B2(n10709), .ZN(n8314) );
  AOI211_X1 U9572 ( .C1(n9924), .C2(n9844), .A(n8315), .B(n8314), .ZN(n8316)
         );
  OAI211_X1 U9573 ( .C1(n8318), .C2(n9835), .A(n8317), .B(n8316), .ZN(P1_U3276) );
  INV_X1 U9574 ( .A(n8319), .ZN(n8320) );
  NAND2_X1 U9575 ( .A1(n8321), .A2(n8320), .ZN(n8379) );
  OAI21_X1 U9576 ( .B1(n8321), .B2(n8320), .A(n8379), .ZN(n8322) );
  NOR2_X1 U9577 ( .A1(n8322), .A2(n8323), .ZN(n8381) );
  AOI21_X1 U9578 ( .B1(n8323), .B2(n8322), .A(n8381), .ZN(n8333) );
  NAND2_X1 U9579 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10477) );
  INV_X1 U9580 ( .A(n10477), .ZN(n8326) );
  NOR2_X1 U9581 ( .A1(n9404), .A2(n8324), .ZN(n8325) );
  AOI211_X1 U9582 ( .C1(n9406), .C2(n8327), .A(n8326), .B(n8325), .ZN(n8328)
         );
  OAI21_X1 U9583 ( .B1(n9409), .B2(n8329), .A(n8328), .ZN(n8330) );
  AOI21_X1 U9584 ( .B1(n8331), .B2(n9411), .A(n8330), .ZN(n8332) );
  OAI21_X1 U9585 ( .B1(n8333), .B2(n9414), .A(n8332), .ZN(P1_U3217) );
  OAI222_X1 U9586 ( .A1(n9266), .A2(n8336), .B1(P2_U3151), .B2(n8335), .C1(
        n8334), .C2(n9263), .ZN(P2_U3271) );
  AOI21_X1 U9587 ( .B1(n9182), .B2(n8338), .A(n8337), .ZN(n8340) );
  MUX2_X1 U9588 ( .A(n6901), .B(n8340), .S(n8349), .Z(n8339) );
  OAI21_X1 U9589 ( .B1(n8343), .B2(n9158), .A(n8339), .ZN(P2_U3471) );
  INV_X1 U9590 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8341) );
  MUX2_X1 U9591 ( .A(n8341), .B(n8340), .S(n10843), .Z(n8342) );
  OAI21_X1 U9592 ( .B1(n8343), .B2(n9249), .A(n8342), .ZN(P2_U3426) );
  OAI22_X1 U9593 ( .A1(n8345), .A2(n9165), .B1(n8873), .B2(n8344), .ZN(n8346)
         );
  NOR2_X1 U9594 ( .A1(n8347), .A2(n8346), .ZN(n10825) );
  INV_X1 U9595 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8348) );
  OR2_X1 U9596 ( .A1(n8349), .A2(n8348), .ZN(n8350) );
  OAI21_X1 U9597 ( .B1(n10825), .B2(n9175), .A(n8350), .ZN(P2_U3472) );
  INV_X1 U9598 ( .A(n8351), .ZN(n8353) );
  NOR3_X1 U9599 ( .A1(n4930), .A2(n8353), .A3(n8352), .ZN(n8356) );
  INV_X1 U9600 ( .A(n8354), .ZN(n8355) );
  OAI21_X1 U9601 ( .B1(n8356), .B2(n8355), .A(n10854), .ZN(n8363) );
  NAND2_X1 U9602 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10576) );
  INV_X1 U9603 ( .A(n10576), .ZN(n8357) );
  AOI21_X1 U9604 ( .B1(n10847), .B2(n8926), .A(n8357), .ZN(n8358) );
  OAI21_X1 U9605 ( .B1(n8359), .B2(n8914), .A(n8358), .ZN(n8360) );
  AOI21_X1 U9606 ( .B1(n8361), .B2(n10856), .A(n8360), .ZN(n8362) );
  OAI211_X1 U9607 ( .C1(n8364), .C2(n8920), .A(n8363), .B(n8362), .ZN(P2_U3176) );
  AOI22_X1 U9608 ( .A1(n8376), .A2(n7491), .B1(n8722), .B2(n9419), .ZN(n8369)
         );
  XNOR2_X1 U9609 ( .A(n8369), .B(n7451), .ZN(n8421) );
  OAI22_X1 U9610 ( .A1(n10815), .A2(n7350), .B1(n8370), .B2(n7349), .ZN(n8422)
         );
  XNOR2_X1 U9611 ( .A(n8421), .B(n8422), .ZN(n8419) );
  XOR2_X1 U9612 ( .A(n8420), .B(n8419), .Z(n8378) );
  NAND2_X1 U9613 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n10446) );
  OAI21_X1 U9614 ( .B1(n9404), .B2(n8371), .A(n10446), .ZN(n8372) );
  AOI21_X1 U9615 ( .B1(n9406), .B2(n9420), .A(n8372), .ZN(n8373) );
  OAI21_X1 U9616 ( .B1(n9409), .B2(n8374), .A(n8373), .ZN(n8375) );
  AOI21_X1 U9617 ( .B1(n8376), .B2(n9411), .A(n8375), .ZN(n8377) );
  OAI21_X1 U9618 ( .B1(n8378), .B2(n9414), .A(n8377), .ZN(P1_U3234) );
  INV_X1 U9619 ( .A(n8379), .ZN(n8380) );
  NOR2_X1 U9620 ( .A1(n8381), .A2(n8380), .ZN(n8384) );
  NOR2_X1 U9621 ( .A1(n8382), .A2(n5024), .ZN(n8383) );
  XNOR2_X1 U9622 ( .A(n8384), .B(n8383), .ZN(n8392) );
  NAND2_X1 U9623 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10361) );
  OAI21_X1 U9624 ( .B1(n9404), .B2(n8385), .A(n10361), .ZN(n8386) );
  AOI21_X1 U9625 ( .B1(n9406), .B2(n9422), .A(n8386), .ZN(n8387) );
  OAI21_X1 U9626 ( .B1(n9409), .B2(n8388), .A(n8387), .ZN(n8389) );
  AOI21_X1 U9627 ( .B1(n8390), .B2(n9411), .A(n8389), .ZN(n8391) );
  OAI21_X1 U9628 ( .B1(n8392), .B2(n9414), .A(n8391), .ZN(P1_U3236) );
  NAND2_X1 U9629 ( .A1(n5023), .A2(n8394), .ZN(n8395) );
  XNOR2_X1 U9630 ( .A(n8393), .B(n8395), .ZN(n8404) );
  NAND2_X1 U9631 ( .A1(n10856), .A2(n8396), .ZN(n8399) );
  NAND2_X1 U9632 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10594) );
  INV_X1 U9633 ( .A(n10594), .ZN(n8397) );
  AOI21_X1 U9634 ( .B1(n10847), .B2(n7079), .A(n8397), .ZN(n8398) );
  OAI211_X1 U9635 ( .C1(n8400), .C2(n8914), .A(n8399), .B(n8398), .ZN(n8401)
         );
  AOI21_X1 U9636 ( .B1(n8402), .B2(n10853), .A(n8401), .ZN(n8403) );
  OAI21_X1 U9637 ( .B1(n8404), .B2(n8907), .A(n8403), .ZN(P2_U3164) );
  NAND2_X1 U9638 ( .A1(n9162), .A2(n8405), .ZN(n8406) );
  XNOR2_X1 U9639 ( .A(n8406), .B(n8615), .ZN(n9252) );
  NAND2_X1 U9640 ( .A1(n8407), .A2(n8615), .ZN(n8408) );
  NAND3_X1 U9641 ( .A1(n8409), .A2(n9103), .A3(n8408), .ZN(n8411) );
  AOI22_X1 U9642 ( .A1(n10844), .A2(n9082), .B1(n9080), .B2(n8925), .ZN(n8410)
         );
  NAND2_X1 U9643 ( .A1(n8411), .A2(n8410), .ZN(n9248) );
  MUX2_X1 U9644 ( .A(n9248), .B(P2_REG2_REG_15__SCAN_IN), .S(n10839), .Z(n8412) );
  INV_X1 U9645 ( .A(n8412), .ZN(n8415) );
  AOI22_X1 U9646 ( .A1(n8413), .A2(n9112), .B1(n9111), .B2(n8917), .ZN(n8414)
         );
  OAI211_X1 U9647 ( .C1(n9252), .C2(n9101), .A(n8415), .B(n8414), .ZN(P2_U3218) );
  INV_X1 U9648 ( .A(n8416), .ZN(n8436) );
  AOI22_X1 U9649 ( .A1(n8417), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9997), .ZN(n8418) );
  OAI21_X1 U9650 ( .B1(n8436), .B2(n10000), .A(n8418), .ZN(P1_U3329) );
  INV_X1 U9651 ( .A(n8422), .ZN(n8423) );
  AOI22_X1 U9652 ( .A1(n8433), .A2(n7491), .B1(n8722), .B2(n9418), .ZN(n8425)
         );
  XNOR2_X1 U9653 ( .A(n8425), .B(n8767), .ZN(n8693) );
  AOI22_X1 U9654 ( .A1(n8433), .A2(n8722), .B1(n7453), .B2(n9418), .ZN(n8692)
         );
  XNOR2_X1 U9655 ( .A(n8693), .B(n8692), .ZN(n8426) );
  XNOR2_X1 U9656 ( .A(n8694), .B(n8426), .ZN(n8435) );
  NAND2_X1 U9657 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10377) );
  INV_X1 U9658 ( .A(n10377), .ZN(n8429) );
  NOR2_X1 U9659 ( .A1(n9404), .A2(n8427), .ZN(n8428) );
  AOI211_X1 U9660 ( .C1(n9406), .C2(n9419), .A(n8429), .B(n8428), .ZN(n8430)
         );
  OAI21_X1 U9661 ( .B1(n9409), .B2(n8431), .A(n8430), .ZN(n8432) );
  AOI21_X1 U9662 ( .B1(n8433), .B2(n9411), .A(n8432), .ZN(n8434) );
  OAI21_X1 U9663 ( .B1(n8435), .B2(n9414), .A(n8434), .ZN(P1_U3215) );
  OAI222_X1 U9664 ( .A1(P2_U3151), .A2(n8437), .B1(n9266), .B2(n8436), .C1(
        n9263), .C2(n6072), .ZN(P2_U3269) );
  INV_X1 U9665 ( .A(n8438), .ZN(n8789) );
  AOI22_X1 U9666 ( .A1(n10298), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9997), .ZN(n8439) );
  OAI21_X1 U9667 ( .B1(n8789), .B2(n10000), .A(n8439), .ZN(P1_U3328) );
  NOR2_X1 U9668 ( .A1(n10829), .A2(n8440), .ZN(n8958) );
  AOI21_X1 U9669 ( .B1(n10839), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8958), .ZN(
        n8441) );
  OAI21_X1 U9670 ( .B1(n8588), .B2(n8981), .A(n8441), .ZN(n8442) );
  AOI21_X1 U9671 ( .B1(n7171), .B2(n8443), .A(n8442), .ZN(n8444) );
  OAI21_X1 U9672 ( .B1(n5547), .B2(n10839), .A(n8444), .ZN(P2_U3204) );
  INV_X1 U9673 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8446) );
  OAI222_X1 U9674 ( .A1(n8448), .A2(P1_U3086), .B1(n10000), .B2(n8447), .C1(
        n8446), .C2(n8445), .ZN(P1_U3330) );
  OAI222_X1 U9675 ( .A1(n9263), .A2(n5572), .B1(n9266), .B2(n8450), .C1(
        P2_U3151), .C2(n8449), .ZN(P2_U3293) );
  NAND2_X1 U9676 ( .A1(n8451), .A2(n8593), .ZN(n8453) );
  OR2_X1 U9677 ( .A1(n5774), .A2(n8691), .ZN(n8452) );
  NAND2_X1 U9678 ( .A1(n8586), .A2(n8587), .ZN(n8589) );
  NAND2_X1 U9679 ( .A1(n8454), .A2(n8801), .ZN(n8455) );
  NOR2_X1 U9680 ( .A1(n8605), .A2(n8590), .ZN(n8601) );
  NAND2_X1 U9681 ( .A1(n8601), .A2(n4937), .ZN(n8457) );
  NAND2_X1 U9682 ( .A1(n8457), .A2(n8456), .ZN(n8579) );
  MUX2_X1 U9683 ( .A(n9201), .B(n8987), .S(n8576), .Z(n8562) );
  OR2_X1 U9684 ( .A1(n9039), .A2(n8590), .ZN(n8460) );
  AND2_X1 U9685 ( .A1(n8637), .A2(n8460), .ZN(n8552) );
  NAND3_X1 U9686 ( .A1(n9039), .A2(n8590), .A3(n8547), .ZN(n8461) );
  OAI21_X1 U9687 ( .B1(n8548), .B2(n8590), .A(n8461), .ZN(n8546) );
  INV_X1 U9688 ( .A(n9078), .ZN(n8635) );
  MUX2_X1 U9689 ( .A(n9107), .B(n8536), .S(n8576), .Z(n8542) );
  AND2_X1 U9690 ( .A1(n8463), .A2(n8462), .ZN(n8619) );
  NAND2_X1 U9691 ( .A1(n8483), .A2(n8464), .ZN(n8466) );
  NOR2_X1 U9692 ( .A1(n8466), .A2(n8576), .ZN(n8465) );
  OAI21_X1 U9693 ( .B1(n8619), .B2(n7543), .A(n8465), .ZN(n8482) );
  INV_X1 U9694 ( .A(n8466), .ZN(n8469) );
  NAND2_X1 U9695 ( .A1(n8470), .A2(n8576), .ZN(n8468) );
  OAI211_X1 U9696 ( .C1(n8469), .C2(n8576), .A(n8468), .B(n6121), .ZN(n8480)
         );
  INV_X1 U9697 ( .A(n8470), .ZN(n8477) );
  NAND2_X1 U9698 ( .A1(n7044), .A2(n8471), .ZN(n8474) );
  NAND3_X1 U9699 ( .A1(n8474), .A2(n8473), .A3(n8472), .ZN(n8476) );
  NAND4_X1 U9700 ( .A1(n8477), .A2(n8476), .A3(n8576), .A4(n8475), .ZN(n8478)
         );
  AND3_X1 U9701 ( .A1(n8480), .A2(n8479), .A3(n8478), .ZN(n8481) );
  NAND2_X1 U9702 ( .A1(n8482), .A2(n8481), .ZN(n8489) );
  INV_X1 U9703 ( .A(n8483), .ZN(n8485) );
  NAND2_X1 U9704 ( .A1(n8509), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U9705 ( .A1(n8502), .A2(n8498), .ZN(n8492) );
  MUX2_X1 U9706 ( .A(n8493), .B(n8492), .S(n8576), .Z(n8494) );
  INV_X1 U9707 ( .A(n8494), .ZN(n8507) );
  MUX2_X1 U9708 ( .A(n8496), .B(n8495), .S(n8576), .Z(n8497) );
  OAI21_X1 U9709 ( .B1(n8499), .B2(n8929), .A(n8498), .ZN(n8500) );
  NAND2_X1 U9710 ( .A1(n8507), .A2(n8500), .ZN(n8501) );
  NAND4_X1 U9711 ( .A1(n8510), .A2(n8512), .A3(n8502), .A4(n8501), .ZN(n8503)
         );
  NAND3_X1 U9712 ( .A1(n8503), .A2(n8511), .A3(n8515), .ZN(n8505) );
  NAND2_X1 U9713 ( .A1(n8507), .A2(n8506), .ZN(n8508) );
  NAND4_X1 U9714 ( .A1(n8511), .A2(n8510), .A3(n8509), .A4(n8508), .ZN(n8513)
         );
  NAND2_X1 U9715 ( .A1(n8513), .A2(n8512), .ZN(n8516) );
  MUX2_X1 U9716 ( .A(n8518), .B(n8517), .S(n8590), .Z(n8519) );
  NOR2_X1 U9717 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U9718 ( .A1(n8873), .A2(n7079), .ZN(n8522) );
  MUX2_X1 U9719 ( .A(n8523), .B(n8522), .S(n8576), .Z(n8524) );
  AND2_X1 U9720 ( .A1(n10827), .A2(n8915), .ZN(n8526) );
  MUX2_X1 U9721 ( .A(n8526), .B(n8525), .S(n8590), .Z(n8527) );
  INV_X1 U9722 ( .A(n8527), .ZN(n8528) );
  NAND3_X1 U9723 ( .A1(n8529), .A2(n8615), .A3(n8528), .ZN(n8533) );
  MUX2_X1 U9724 ( .A(n8531), .B(n8530), .S(n8576), .Z(n8532) );
  NAND3_X1 U9725 ( .A1(n8633), .A2(n8533), .A3(n8532), .ZN(n8543) );
  MUX2_X1 U9726 ( .A(n8538), .B(n8534), .S(n8590), .Z(n8535) );
  INV_X1 U9727 ( .A(n8538), .ZN(n8539) );
  AND2_X1 U9728 ( .A1(n10852), .A2(n8539), .ZN(n8540) );
  OR3_X1 U9729 ( .A1(n8543), .A2(n8542), .A3(n8635), .ZN(n8544) );
  NAND3_X1 U9730 ( .A1(n8546), .A2(n8545), .A3(n8544), .ZN(n8551) );
  OR3_X1 U9731 ( .A1(n8548), .A2(n8590), .A3(n8547), .ZN(n8550) );
  NAND3_X1 U9732 ( .A1(n8548), .A2(n8590), .A3(n9039), .ZN(n8549) );
  NAND4_X1 U9733 ( .A1(n8552), .A2(n8551), .A3(n8550), .A4(n8549), .ZN(n8555)
         );
  INV_X1 U9734 ( .A(n9053), .ZN(n9215) );
  MUX2_X1 U9735 ( .A(n9064), .B(n9215), .S(n8590), .Z(n8553) );
  NAND2_X1 U9736 ( .A1(n8553), .A2(n9024), .ZN(n8554) );
  MUX2_X1 U9737 ( .A(n9033), .B(n8924), .S(n8576), .Z(n8557) );
  MUX2_X1 U9738 ( .A(n8559), .B(n8558), .S(n8576), .Z(n8560) );
  AOI21_X1 U9739 ( .B1(n8640), .B2(n8562), .A(n8561), .ZN(n8565) );
  XOR2_X1 U9740 ( .A(n8999), .B(n9195), .Z(n8564) );
  MUX2_X1 U9741 ( .A(n8612), .B(n8613), .S(n8576), .Z(n8563) );
  OAI21_X1 U9742 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8571) );
  MUX2_X1 U9743 ( .A(n8569), .B(n8568), .S(n8576), .Z(n8570) );
  AOI21_X1 U9744 ( .B1(n8571), .B2(n8978), .A(n8570), .ZN(n8575) );
  NAND2_X1 U9745 ( .A1(n8572), .A2(n8573), .ZN(n8962) );
  MUX2_X1 U9746 ( .A(n8573), .B(n8572), .S(n8576), .Z(n8574) );
  OAI21_X1 U9747 ( .B1(n8575), .B2(n8962), .A(n8574), .ZN(n8580) );
  NAND2_X1 U9748 ( .A1(n8579), .A2(n8580), .ZN(n8578) );
  MUX2_X1 U9749 ( .A(n4937), .B(n8803), .S(n8576), .Z(n8577) );
  NAND2_X1 U9750 ( .A1(n8578), .A2(n8577), .ZN(n8584) );
  INV_X1 U9751 ( .A(n8579), .ZN(n8582) );
  INV_X1 U9752 ( .A(n8580), .ZN(n8581) );
  NAND2_X1 U9753 ( .A1(n8582), .A2(n8581), .ZN(n8583) );
  NAND2_X1 U9754 ( .A1(n8584), .A2(n8583), .ZN(n8585) );
  NAND2_X1 U9755 ( .A1(n8585), .A2(n4931), .ZN(n8602) );
  INV_X1 U9756 ( .A(n8602), .ZN(n8591) );
  NAND2_X1 U9757 ( .A1(n8588), .A2(n8922), .ZN(n8607) );
  NAND2_X1 U9758 ( .A1(n8592), .A2(n8607), .ZN(n8645) );
  OAI211_X1 U9759 ( .C1(n8591), .C2(n8645), .A(n8590), .B(n8589), .ZN(n8604)
         );
  INV_X1 U9760 ( .A(n8592), .ZN(n8652) );
  NAND2_X1 U9761 ( .A1(n9257), .A2(n8593), .ZN(n8595) );
  OR2_X1 U9762 ( .A1(n5774), .A2(n7234), .ZN(n8594) );
  NAND2_X1 U9763 ( .A1(n5764), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U9764 ( .A1(n8596), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U9765 ( .A1(n5735), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8597) );
  NAND4_X1 U9766 ( .A1(n8600), .A2(n8599), .A3(n8598), .A4(n8597), .ZN(n8956)
         );
  NOR2_X1 U9767 ( .A1(n9178), .A2(n8956), .ZN(n8647) );
  AOI211_X1 U9768 ( .C1(n8602), .C2(n8601), .A(n8652), .B(n8647), .ZN(n8603)
         );
  AOI21_X1 U9769 ( .B1(n8604), .B2(n8603), .A(n6149), .ZN(n8611) );
  INV_X1 U9770 ( .A(n9178), .ZN(n8651) );
  INV_X1 U9771 ( .A(n8956), .ZN(n8609) );
  NOR2_X1 U9772 ( .A1(n8651), .A2(n8609), .ZN(n8646) );
  INV_X1 U9773 ( .A(n8646), .ZN(n8610) );
  INV_X1 U9774 ( .A(n8962), .ZN(n8964) );
  INV_X1 U9775 ( .A(n8978), .ZN(n8972) );
  INV_X1 U9776 ( .A(n8615), .ZN(n8631) );
  NOR2_X1 U9777 ( .A1(n6121), .A2(n5252), .ZN(n8616) );
  AND4_X1 U9778 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n8623)
         );
  NAND4_X1 U9779 ( .A1(n8623), .A2(n8622), .A3(n8621), .A4(n8620), .ZN(n8624)
         );
  NOR3_X1 U9780 ( .A1(n8626), .A2(n8625), .A3(n8624), .ZN(n8627) );
  NAND4_X1 U9781 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n5009), .ZN(n8630)
         );
  NOR3_X1 U9782 ( .A1(n8631), .A2(n5168), .A3(n8630), .ZN(n8632) );
  NAND2_X1 U9783 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  NOR2_X1 U9784 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  NAND4_X1 U9785 ( .A1(n8637), .A2(n9071), .A3(n8636), .A4(n9092), .ZN(n8638)
         );
  INV_X1 U9786 ( .A(n8639), .ZN(n8641) );
  NAND2_X1 U9787 ( .A1(n8641), .A2(n8640), .ZN(n9005) );
  NAND4_X1 U9788 ( .A1(n8994), .A2(n5563), .A3(n9005), .A4(n9019), .ZN(n8642)
         );
  NOR2_X1 U9789 ( .A1(n8972), .A2(n8642), .ZN(n8643) );
  NAND3_X1 U9790 ( .A1(n8795), .A2(n8964), .A3(n8643), .ZN(n8644) );
  INV_X1 U9791 ( .A(n8647), .ZN(n8648) );
  OAI21_X1 U9792 ( .B1(n8650), .B2(n8649), .A(n8648), .ZN(n8653) );
  AOI22_X1 U9793 ( .A1(n8653), .A2(n6149), .B1(n8652), .B2(n8651), .ZN(n8654)
         );
  NAND3_X1 U9794 ( .A1(n8657), .A2(n8656), .A3(n8788), .ZN(n8658) );
  OAI211_X1 U9795 ( .C1(n8659), .C2(n8661), .A(n8658), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8660) );
  XOR2_X1 U9796 ( .A(n8663), .B(n8662), .Z(n8668) );
  NAND2_X1 U9797 ( .A1(n10856), .A2(n9052), .ZN(n8665) );
  AOI22_X1 U9798 ( .A1(n10847), .A2(n8924), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8664) );
  OAI211_X1 U9799 ( .C1(n9048), .C2(n8914), .A(n8665), .B(n8664), .ZN(n8666)
         );
  AOI21_X1 U9800 ( .B1(n9053), .B2(n10853), .A(n8666), .ZN(n8667) );
  OAI21_X1 U9801 ( .B1(n8668), .B2(n8907), .A(n8667), .ZN(P2_U3163) );
  NAND2_X1 U9802 ( .A1(n8670), .A2(n8669), .ZN(n8830) );
  NAND2_X1 U9803 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U9804 ( .A1(n10856), .A2(n8979), .ZN(n8676) );
  AOI22_X1 U9805 ( .A1(n10845), .A2(n8999), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8675) );
  OAI211_X1 U9806 ( .C1(n8976), .C2(n8898), .A(n8676), .B(n8675), .ZN(n8677)
         );
  AOI21_X1 U9807 ( .B1(n8678), .B2(n10853), .A(n8677), .ZN(n8679) );
  INV_X1 U9808 ( .A(n9373), .ZN(n8685) );
  AND2_X1 U9809 ( .A1(n8682), .A2(n8681), .ZN(n9441) );
  OR3_X1 U9810 ( .A1(n8680), .A2(n9441), .A3(n9414), .ZN(n8684) );
  AOI22_X1 U9811 ( .A1(n9372), .A2(n10228), .B1(n9411), .B2(n7554), .ZN(n8683)
         );
  OAI211_X1 U9812 ( .C1(n8685), .C2(n10708), .A(n8684), .B(n8683), .ZN(
        P1_U3232) );
  NAND2_X1 U9813 ( .A1(n8686), .A2(n10843), .ZN(n8689) );
  INV_X1 U9814 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8687) );
  OR2_X1 U9815 ( .A1(n10843), .A2(n8687), .ZN(n8688) );
  OAI21_X1 U9816 ( .B1(n8782), .B2(n9249), .A(n5548), .ZN(P2_U3455) );
  INV_X1 U9817 ( .A(n8451), .ZN(n9993) );
  OAI222_X1 U9818 ( .A1(n9263), .A2(n8691), .B1(n9266), .B2(n9993), .C1(
        P2_U3151), .C2(n8690), .ZN(P2_U3265) );
  AOI22_X1 U9819 ( .A1(n9412), .A2(n7491), .B1(n8722), .B2(n9829), .ZN(n8695)
         );
  XNOR2_X1 U9820 ( .A(n8695), .B(n8767), .ZN(n9400) );
  AOI22_X1 U9821 ( .A1(n9412), .A2(n8722), .B1(n7453), .B2(n9829), .ZN(n9399)
         );
  OAI22_X1 U9822 ( .A1(n9825), .A2(n7350), .B1(n9403), .B2(n7349), .ZN(n8699)
         );
  NAND2_X1 U9823 ( .A1(n9930), .A2(n7491), .ZN(n8697) );
  NAND2_X1 U9824 ( .A1(n9417), .A2(n8722), .ZN(n8696) );
  NAND2_X1 U9825 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  XNOR2_X1 U9826 ( .A(n8698), .B(n7451), .ZN(n8700) );
  XOR2_X1 U9827 ( .A(n8699), .B(n8700), .Z(n9323) );
  NAND2_X1 U9828 ( .A1(n9322), .A2(n9323), .ZN(n8702) );
  NAND2_X1 U9829 ( .A1(n9577), .A2(n7491), .ZN(n8704) );
  NAND2_X1 U9830 ( .A1(n9830), .A2(n8722), .ZN(n8703) );
  NAND2_X1 U9831 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  XNOR2_X1 U9832 ( .A(n8705), .B(n8767), .ZN(n8706) );
  AOI22_X1 U9833 ( .A1(n9577), .A2(n8722), .B1(n7453), .B2(n9830), .ZN(n8707)
         );
  XNOR2_X1 U9834 ( .A(n8706), .B(n8707), .ZN(n9331) );
  INV_X1 U9835 ( .A(n8706), .ZN(n8708) );
  NAND2_X1 U9836 ( .A1(n8708), .A2(n8707), .ZN(n8712) );
  AOI22_X1 U9837 ( .A1(n9919), .A2(n7491), .B1(n8722), .B2(n9781), .ZN(n8710)
         );
  XNOR2_X1 U9838 ( .A(n8710), .B(n8767), .ZN(n8711) );
  INV_X1 U9839 ( .A(n8711), .ZN(n8713) );
  AND2_X1 U9840 ( .A1(n9331), .A2(n8711), .ZN(n8714) );
  INV_X1 U9841 ( .A(n9919), .ZN(n9803) );
  OAI22_X1 U9842 ( .A1(n9803), .A2(n7350), .B1(n9332), .B2(n7349), .ZN(n9380)
         );
  AOI22_X1 U9843 ( .A1(n9791), .A2(n7491), .B1(n8722), .B2(n9809), .ZN(n8716)
         );
  XNOR2_X1 U9844 ( .A(n8716), .B(n8767), .ZN(n8718) );
  AOI22_X1 U9845 ( .A1(n9791), .A2(n8722), .B1(n7453), .B2(n9809), .ZN(n8717)
         );
  XNOR2_X1 U9846 ( .A(n8718), .B(n8717), .ZN(n9279) );
  NAND2_X1 U9847 ( .A1(n9906), .A2(n7491), .ZN(n8720) );
  OR2_X1 U9848 ( .A1(n9281), .A2(n7350), .ZN(n8719) );
  NAND2_X1 U9849 ( .A1(n8720), .A2(n8719), .ZN(n8721) );
  XNOR2_X1 U9850 ( .A(n8721), .B(n8767), .ZN(n8723) );
  AOI22_X1 U9851 ( .A1(n9906), .A2(n8722), .B1(n7453), .B2(n9782), .ZN(n8724)
         );
  XNOR2_X1 U9852 ( .A(n8723), .B(n8724), .ZN(n9352) );
  INV_X1 U9853 ( .A(n8723), .ZN(n8725) );
  NAND2_X1 U9854 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  NOR2_X1 U9855 ( .A1(n9771), .A2(n7350), .ZN(n8727) );
  AOI21_X1 U9856 ( .B1(n9754), .B2(n7491), .A(n8727), .ZN(n8728) );
  XNOR2_X1 U9857 ( .A(n8728), .B(n7451), .ZN(n8731) );
  OAI22_X1 U9858 ( .A1(n9965), .A2(n7350), .B1(n9771), .B2(n7349), .ZN(n8729)
         );
  XNOR2_X1 U9859 ( .A(n8731), .B(n8729), .ZN(n9306) );
  NAND2_X1 U9860 ( .A1(n9305), .A2(n9306), .ZN(n8733) );
  INV_X1 U9861 ( .A(n8729), .ZN(n8730) );
  NAND2_X1 U9862 ( .A1(n8731), .A2(n8730), .ZN(n8732) );
  AOI22_X1 U9863 ( .A1(n9736), .A2(n7491), .B1(n8722), .B2(n9747), .ZN(n8734)
         );
  XNOR2_X1 U9864 ( .A(n8734), .B(n8767), .ZN(n8735) );
  AOI22_X1 U9865 ( .A1(n9889), .A2(n7491), .B1(n8722), .B2(n9587), .ZN(n8737)
         );
  XNOR2_X1 U9866 ( .A(n8737), .B(n8767), .ZN(n8744) );
  AOI22_X1 U9867 ( .A1(n9889), .A2(n8722), .B1(n7453), .B2(n9587), .ZN(n8743)
         );
  XNOR2_X1 U9868 ( .A(n8744), .B(n8743), .ZN(n9339) );
  NAND2_X1 U9869 ( .A1(n9885), .A2(n7491), .ZN(n8739) );
  NAND2_X1 U9870 ( .A1(n9679), .A2(n8722), .ZN(n8738) );
  NAND2_X1 U9871 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  XNOR2_X1 U9872 ( .A(n8740), .B(n7451), .ZN(n8746) );
  NAND2_X1 U9873 ( .A1(n9885), .A2(n8722), .ZN(n8742) );
  NAND2_X1 U9874 ( .A1(n9679), .A2(n7453), .ZN(n8741) );
  NAND2_X1 U9875 ( .A1(n8742), .A2(n8741), .ZN(n8747) );
  NAND2_X1 U9876 ( .A1(n8746), .A2(n8747), .ZN(n9342) );
  INV_X1 U9877 ( .A(n9342), .ZN(n8745) );
  OR2_X1 U9878 ( .A1(n9339), .A2(n8745), .ZN(n8752) );
  NAND2_X1 U9879 ( .A1(n8744), .A2(n8743), .ZN(n9340) );
  OR2_X1 U9880 ( .A1(n8745), .A2(n9340), .ZN(n8750) );
  INV_X1 U9881 ( .A(n8746), .ZN(n8749) );
  INV_X1 U9882 ( .A(n8747), .ZN(n8748) );
  NAND2_X1 U9883 ( .A1(n8749), .A2(n8748), .ZN(n9343) );
  OAI22_X1 U9884 ( .A1(n9685), .A2(n7350), .B1(n9702), .B2(n7349), .ZN(n8760)
         );
  NAND2_X1 U9885 ( .A1(n9879), .A2(n7491), .ZN(n8754) );
  OR2_X1 U9886 ( .A1(n9702), .A2(n7350), .ZN(n8753) );
  NAND2_X1 U9887 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  XNOR2_X1 U9888 ( .A(n8755), .B(n8767), .ZN(n8761) );
  XOR2_X1 U9889 ( .A(n8760), .B(n8761), .Z(n9314) );
  AND2_X1 U9890 ( .A1(n9680), .A2(n7453), .ZN(n8756) );
  AOI21_X1 U9891 ( .B1(n9672), .B2(n8722), .A(n8756), .ZN(n8763) );
  NAND2_X1 U9892 ( .A1(n9672), .A2(n7491), .ZN(n8758) );
  NAND2_X1 U9893 ( .A1(n9680), .A2(n8722), .ZN(n8757) );
  NAND2_X1 U9894 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  XNOR2_X1 U9895 ( .A(n8759), .B(n8767), .ZN(n8765) );
  XOR2_X1 U9896 ( .A(n8763), .B(n8765), .Z(n9386) );
  NOR2_X1 U9897 ( .A1(n8761), .A2(n8760), .ZN(n9387) );
  NOR2_X1 U9898 ( .A1(n9386), .A2(n9387), .ZN(n8762) );
  INV_X1 U9899 ( .A(n8763), .ZN(n8764) );
  NAND2_X1 U9900 ( .A1(n8765), .A2(n8764), .ZN(n8771) );
  AOI22_X1 U9901 ( .A1(n9654), .A2(n7491), .B1(n8722), .B2(n9633), .ZN(n8766)
         );
  XOR2_X1 U9902 ( .A(n8767), .B(n8766), .Z(n8769) );
  OAI22_X1 U9903 ( .A1(n9948), .A2(n7350), .B1(n9666), .B2(n7349), .ZN(n8768)
         );
  NOR2_X1 U9904 ( .A1(n8769), .A2(n8768), .ZN(n9300) );
  AOI21_X1 U9905 ( .B1(n8769), .B2(n8768), .A(n9300), .ZN(n8770) );
  AOI21_X1 U9906 ( .B1(n9389), .B2(n8771), .A(n8770), .ZN(n8775) );
  INV_X1 U9907 ( .A(n8770), .ZN(n8773) );
  INV_X1 U9908 ( .A(n8771), .ZN(n8772) );
  NOR2_X1 U9909 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  OAI21_X1 U9910 ( .B1(n8775), .B2(n9295), .A(n9390), .ZN(n8780) );
  INV_X1 U9911 ( .A(n8776), .ZN(n9655) );
  AOI22_X1 U9912 ( .A1(n9406), .A2(n9680), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8777) );
  OAI21_X1 U9913 ( .B1(n9618), .B2(n9404), .A(n8777), .ZN(n8778) );
  AOI21_X1 U9914 ( .B1(n9655), .B2(n9395), .A(n8778), .ZN(n8779) );
  OAI211_X1 U9915 ( .C1(n9948), .C2(n9398), .A(n8780), .B(n8779), .ZN(P1_U3214) );
  AOI22_X1 U9916 ( .A1(n10839), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9111), .B2(
        n8798), .ZN(n8781) );
  OAI21_X1 U9917 ( .B1(n8782), .B2(n8981), .A(n8781), .ZN(n8783) );
  AOI21_X1 U9918 ( .B1(n8784), .B2(n9115), .A(n8783), .ZN(n8785) );
  OAI21_X1 U9919 ( .B1(n8786), .B2(n10839), .A(n8785), .ZN(P2_U3205) );
  OAI222_X1 U9920 ( .A1(n9266), .A2(n8789), .B1(n8788), .B2(P2_U3151), .C1(
        n8787), .C2(n9263), .ZN(P2_U3268) );
  OAI21_X1 U9921 ( .B1(n8793), .B2(n8792), .A(n8791), .ZN(n8797) );
  XNOR2_X1 U9922 ( .A(n8795), .B(n8794), .ZN(n8796) );
  XNOR2_X1 U9923 ( .A(n8797), .B(n8796), .ZN(n8805) );
  NAND2_X1 U9924 ( .A1(n10856), .A2(n8798), .ZN(n8800) );
  AOI22_X1 U9925 ( .A1(n10845), .A2(n8923), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8799) );
  OAI211_X1 U9926 ( .C1(n8801), .C2(n8898), .A(n8800), .B(n8799), .ZN(n8802)
         );
  AOI21_X1 U9927 ( .B1(n8803), .B2(n10853), .A(n8802), .ZN(n8804) );
  OAI21_X1 U9928 ( .B1(n8805), .B2(n8907), .A(n8804), .ZN(P2_U3160) );
  INV_X1 U9929 ( .A(n8807), .ZN(n8808) );
  AOI21_X1 U9930 ( .B1(n8809), .B2(n8806), .A(n8808), .ZN(n8814) );
  INV_X1 U9931 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10110) );
  OAI22_X1 U9932 ( .A1(n8898), .A2(n9171), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10110), .ZN(n8811) );
  NOR2_X1 U9933 ( .A1(n8914), .A2(n9169), .ZN(n8810) );
  AOI211_X1 U9934 ( .C1(n10828), .C2(n10856), .A(n8811), .B(n8810), .ZN(n8813)
         );
  NAND2_X1 U9935 ( .A1(n10827), .A2(n10853), .ZN(n8812) );
  OAI211_X1 U9936 ( .C1(n8814), .C2(n8907), .A(n8813), .B(n8812), .ZN(P2_U3155) );
  XNOR2_X1 U9937 ( .A(n8815), .B(n9026), .ZN(n8820) );
  INV_X1 U9938 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10066) );
  OAI22_X1 U9939 ( .A1(n8898), .A2(n9012), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10066), .ZN(n8817) );
  NOR2_X1 U9940 ( .A1(n8914), .A2(n9049), .ZN(n8816) );
  AOI211_X1 U9941 ( .C1(n9015), .C2(n10856), .A(n8817), .B(n8816), .ZN(n8819)
         );
  NAND2_X1 U9942 ( .A1(n9016), .A2(n10853), .ZN(n8818) );
  OAI211_X1 U9943 ( .C1(n8820), .C2(n8907), .A(n8819), .B(n8818), .ZN(P2_U3156) );
  OAI211_X1 U9944 ( .C1(n8823), .C2(n8822), .A(n8821), .B(n10854), .ZN(n8828)
         );
  NAND2_X1 U9945 ( .A1(n10845), .A2(n10846), .ZN(n8825) );
  OAI211_X1 U9946 ( .C1(n9048), .C2(n8898), .A(n8825), .B(n8824), .ZN(n8826)
         );
  AOI21_X1 U9947 ( .B1(n9074), .B2(n10856), .A(n8826), .ZN(n8827) );
  OAI211_X1 U9948 ( .C1(n8829), .C2(n8920), .A(n8828), .B(n8827), .ZN(P2_U3159) );
  XOR2_X1 U9949 ( .A(n8831), .B(n8830), .Z(n8837) );
  OAI22_X1 U9950 ( .A1(n8898), .A2(n8832), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10192), .ZN(n8834) );
  NOR2_X1 U9951 ( .A1(n8914), .A2(n9012), .ZN(n8833) );
  AOI211_X1 U9952 ( .C1(n8992), .C2(n10856), .A(n8834), .B(n8833), .ZN(n8836)
         );
  NAND2_X1 U9953 ( .A1(n9195), .A2(n10853), .ZN(n8835) );
  OAI211_X1 U9954 ( .C1(n8837), .C2(n8907), .A(n8836), .B(n8835), .ZN(P2_U3165) );
  OAI211_X1 U9955 ( .C1(n8840), .C2(n8839), .A(n8838), .B(n10854), .ZN(n8845)
         );
  NAND2_X1 U9956 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10658) );
  INV_X1 U9957 ( .A(n10658), .ZN(n8841) );
  AOI21_X1 U9958 ( .B1(n10847), .B2(n9081), .A(n8841), .ZN(n8842) );
  OAI21_X1 U9959 ( .B1(n9171), .B2(n8914), .A(n8842), .ZN(n8843) );
  AOI21_X1 U9960 ( .B1(n9110), .B2(n10856), .A(n8843), .ZN(n8844) );
  OAI211_X1 U9961 ( .C1(n8846), .C2(n8920), .A(n8845), .B(n8844), .ZN(P2_U3166) );
  XOR2_X1 U9962 ( .A(n8848), .B(n8847), .Z(n8853) );
  INV_X1 U9963 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10085) );
  OAI22_X1 U9964 ( .A1(n8898), .A2(n8975), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10085), .ZN(n8850) );
  NOR2_X1 U9965 ( .A1(n8914), .A2(n8878), .ZN(n8849) );
  AOI211_X1 U9966 ( .C1(n9003), .C2(n10856), .A(n8850), .B(n8849), .ZN(n8852)
         );
  NAND2_X1 U9967 ( .A1(n9201), .A2(n10853), .ZN(n8851) );
  OAI211_X1 U9968 ( .C1(n8853), .C2(n8907), .A(n8852), .B(n8851), .ZN(P2_U3169) );
  INV_X1 U9969 ( .A(n8854), .ZN(n8855) );
  AOI21_X1 U9970 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8862) );
  NAND2_X1 U9971 ( .A1(n10856), .A2(n9067), .ZN(n8859) );
  AOI22_X1 U9972 ( .A1(n10847), .A2(n9025), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8858) );
  OAI211_X1 U9973 ( .C1(n9063), .C2(n8914), .A(n8859), .B(n8858), .ZN(n8860)
         );
  AOI21_X1 U9974 ( .B1(n9141), .B2(n10853), .A(n8860), .ZN(n8861) );
  OAI21_X1 U9975 ( .B1(n8862), .B2(n8907), .A(n8861), .ZN(P2_U3173) );
  OAI211_X1 U9976 ( .C1(n8865), .C2(n8864), .A(n8863), .B(n10854), .ZN(n8872)
         );
  NAND2_X1 U9977 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10610) );
  INV_X1 U9978 ( .A(n10610), .ZN(n8866) );
  AOI21_X1 U9979 ( .B1(n10847), .B2(n8925), .A(n8866), .ZN(n8867) );
  OAI21_X1 U9980 ( .B1(n8868), .B2(n8914), .A(n8867), .ZN(n8869) );
  AOI21_X1 U9981 ( .B1(n8870), .B2(n10856), .A(n8869), .ZN(n8871) );
  OAI211_X1 U9982 ( .C1(n8873), .C2(n8920), .A(n8872), .B(n8871), .ZN(P2_U3174) );
  OAI211_X1 U9983 ( .C1(n8874), .C2(n8876), .A(n8875), .B(n10854), .ZN(n8881)
         );
  AOI22_X1 U9984 ( .A1(n10845), .A2(n9025), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8877) );
  OAI21_X1 U9985 ( .B1(n8878), .B2(n8898), .A(n8877), .ZN(n8879) );
  AOI21_X1 U9986 ( .B1(n9032), .B2(n10856), .A(n8879), .ZN(n8880) );
  OAI211_X1 U9987 ( .C1(n5205), .C2(n8920), .A(n8881), .B(n8880), .ZN(P2_U3175) );
  AOI21_X1 U9988 ( .B1(n8883), .B2(n8882), .A(n8907), .ZN(n8885) );
  NAND2_X1 U9989 ( .A1(n8885), .A2(n8884), .ZN(n8890) );
  NAND2_X1 U9990 ( .A1(n10845), .A2(n9081), .ZN(n8887) );
  OAI211_X1 U9991 ( .C1(n9063), .C2(n8898), .A(n8887), .B(n8886), .ZN(n8888)
         );
  AOI21_X1 U9992 ( .B1(n9086), .B2(n10856), .A(n8888), .ZN(n8889) );
  OAI211_X1 U9993 ( .C1(n8891), .C2(n8920), .A(n8890), .B(n8889), .ZN(P2_U3178) );
  OAI211_X1 U9994 ( .C1(n8894), .C2(n8893), .A(n8892), .B(n10854), .ZN(n8906)
         );
  NAND2_X1 U9995 ( .A1(n10845), .A2(n8895), .ZN(n8897) );
  INV_X1 U9996 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U9997 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10210), .ZN(n8943) );
  INV_X1 U9998 ( .A(n8943), .ZN(n8896) );
  OAI211_X1 U9999 ( .C1(n8899), .C2(n8898), .A(n8897), .B(n8896), .ZN(n8900)
         );
  INV_X1 U10000 ( .A(n8900), .ZN(n8905) );
  NAND2_X1 U10001 ( .A1(n10856), .A2(n8901), .ZN(n8904) );
  NAND2_X1 U10002 ( .A1(n10853), .A2(n8902), .ZN(n8903) );
  NAND4_X1 U10003 ( .A1(n8906), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(
        P2_U3179) );
  AOI21_X1 U10004 ( .B1(n8909), .B2(n8908), .A(n8907), .ZN(n8911) );
  NAND2_X1 U10005 ( .A1(n8911), .A2(n8910), .ZN(n8919) );
  NAND2_X1 U10006 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10642)
         );
  INV_X1 U10007 ( .A(n10642), .ZN(n8912) );
  AOI21_X1 U10008 ( .B1(n10847), .B2(n10844), .A(n8912), .ZN(n8913) );
  OAI21_X1 U10009 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8916) );
  AOI21_X1 U10010 ( .B1(n8917), .B2(n10856), .A(n8916), .ZN(n8918) );
  OAI211_X1 U10011 ( .C1(n9250), .C2(n8920), .A(n8919), .B(n8918), .ZN(
        P2_U3181) );
  MUX2_X1 U10012 ( .A(n8956), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8931), .Z(
        P2_U3522) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8921), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8922), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10015 ( .A(n4937), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8931), .Z(
        P2_U3519) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8923), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8988), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10018 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8999), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10019 ( .A(n8987), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8931), .Z(
        P2_U3515) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9026), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10021 ( .A(n8924), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8931), .Z(
        P2_U3513) );
  MUX2_X1 U10022 ( .A(n9025), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8931), .Z(
        P2_U3512) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9072), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9083), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n10846), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9081), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n10844), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10028 ( .A(n8925), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8931), .Z(
        P2_U3505) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n7079), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8926), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8927), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8928), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10033 ( .A(n8929), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8931), .Z(
        P2_U3498) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8930), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10035 ( .A(n8932), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8931), .Z(
        P2_U3494) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7040), .S(P2_U3893), .Z(
        P2_U3492) );
  OAI21_X1 U10037 ( .B1(n8935), .B2(n8934), .A(n8933), .ZN(n8936) );
  NAND2_X1 U10038 ( .A1(n8936), .A2(n10670), .ZN(n8954) );
  INV_X1 U10039 ( .A(n8937), .ZN(n8938) );
  NAND3_X1 U10040 ( .A1(n5026), .A2(n10481), .A3(n8938), .ZN(n8940) );
  AOI21_X1 U10041 ( .B1(n8941), .B2(n8940), .A(n8939), .ZN(n8942) );
  AOI211_X1 U10042 ( .C1(n8944), .C2(n10662), .A(n8943), .B(n8942), .ZN(n8953)
         );
  NAND2_X1 U10043 ( .A1(n10661), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8952) );
  INV_X1 U10044 ( .A(n10490), .ZN(n8948) );
  INV_X1 U10045 ( .A(n8945), .ZN(n8947) );
  NOR3_X1 U10046 ( .A1(n8948), .A2(n8947), .A3(n8946), .ZN(n8949) );
  INV_X1 U10047 ( .A(n10677), .ZN(n10492) );
  OAI21_X1 U10048 ( .B1(n8950), .B2(n8949), .A(n10492), .ZN(n8951) );
  NAND4_X1 U10049 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(
        P2_U3188) );
  NAND2_X1 U10050 ( .A1(n8956), .A2(n8955), .ZN(n9176) );
  INV_X1 U10051 ( .A(n9176), .ZN(n8957) );
  NOR3_X1 U10052 ( .A1(n10839), .A2(n8958), .A3(n8957), .ZN(n8961) );
  NOR2_X1 U10053 ( .A1(n10837), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8959) );
  OAI22_X1 U10054 ( .A1(n9178), .A2(n8981), .B1(n8961), .B2(n8959), .ZN(
        P2_U3202) );
  NOR2_X1 U10055 ( .A1(n10837), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8960) );
  OAI22_X1 U10056 ( .A1(n9181), .A2(n8981), .B1(n8961), .B2(n8960), .ZN(
        P2_U3203) );
  XNOR2_X1 U10057 ( .A(n8963), .B(n8962), .ZN(n9188) );
  INV_X1 U10058 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8968) );
  XNOR2_X1 U10059 ( .A(n8965), .B(n8964), .ZN(n8967) );
  AOI222_X1 U10060 ( .A1(n9103), .A2(n8967), .B1(n4937), .B2(n9082), .C1(n8988), .C2(n9080), .ZN(n9183) );
  MUX2_X1 U10061 ( .A(n8968), .B(n9183), .S(n10837), .Z(n8971) );
  AOI22_X1 U10062 ( .A1(n9185), .A2(n9112), .B1(n9111), .B2(n8969), .ZN(n8970)
         );
  OAI211_X1 U10063 ( .C1(n9188), .C2(n9101), .A(n8971), .B(n8970), .ZN(
        P2_U3206) );
  XNOR2_X1 U10064 ( .A(n8973), .B(n8972), .ZN(n8974) );
  OAI222_X1 U10065 ( .A1(n9106), .A2(n8976), .B1(n9170), .B2(n8975), .C1(n9168), .C2(n8974), .ZN(n9125) );
  INV_X1 U10066 ( .A(n9125), .ZN(n8984) );
  XNOR2_X1 U10067 ( .A(n8977), .B(n8978), .ZN(n9126) );
  AOI22_X1 U10068 ( .A1(n10839), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9111), 
        .B2(n8979), .ZN(n8980) );
  OAI21_X1 U10069 ( .B1(n9192), .B2(n8981), .A(n8980), .ZN(n8982) );
  AOI21_X1 U10070 ( .B1(n9126), .B2(n9115), .A(n8982), .ZN(n8983) );
  OAI21_X1 U10071 ( .B1(n8984), .B2(n10839), .A(n8983), .ZN(P2_U3207) );
  NOR2_X1 U10072 ( .A1(n8985), .A2(n10831), .ZN(n8991) );
  XNOR2_X1 U10073 ( .A(n8986), .B(n8994), .ZN(n8989) );
  AOI222_X1 U10074 ( .A1(n9103), .A2(n8989), .B1(n8988), .B2(n9082), .C1(n8987), .C2(n9080), .ZN(n9193) );
  INV_X1 U10075 ( .A(n9193), .ZN(n8990) );
  AOI211_X1 U10076 ( .C1(n9111), .C2(n8992), .A(n8991), .B(n8990), .ZN(n8996)
         );
  XNOR2_X1 U10077 ( .A(n8993), .B(n8994), .ZN(n9196) );
  AOI22_X1 U10078 ( .A1(n9196), .A2(n9115), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10839), .ZN(n8995) );
  OAI21_X1 U10079 ( .B1(n8996), .B2(n10839), .A(n8995), .ZN(P2_U3208) );
  INV_X1 U10080 ( .A(n9201), .ZN(n8997) );
  NOR2_X1 U10081 ( .A1(n8997), .A2(n10831), .ZN(n9002) );
  XOR2_X1 U10082 ( .A(n9005), .B(n8998), .Z(n9000) );
  AOI222_X1 U10083 ( .A1(n9103), .A2(n9000), .B1(n8999), .B2(n9082), .C1(n9026), .C2(n9080), .ZN(n9199) );
  INV_X1 U10084 ( .A(n9199), .ZN(n9001) );
  AOI211_X1 U10085 ( .C1(n9111), .C2(n9003), .A(n9002), .B(n9001), .ZN(n9007)
         );
  XNOR2_X1 U10086 ( .A(n9004), .B(n9005), .ZN(n9202) );
  AOI22_X1 U10087 ( .A1(n9202), .A2(n9115), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10839), .ZN(n9006) );
  OAI21_X1 U10088 ( .B1(n9007), .B2(n10839), .A(n9006), .ZN(P2_U3209) );
  XNOR2_X1 U10089 ( .A(n9008), .B(n9009), .ZN(n9207) );
  INV_X1 U10090 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9014) );
  XNOR2_X1 U10091 ( .A(n9010), .B(n9009), .ZN(n9011) );
  OAI222_X1 U10092 ( .A1(n9170), .A2(n9049), .B1(n9106), .B2(n9012), .C1(n9011), .C2(n9168), .ZN(n9205) );
  INV_X1 U10093 ( .A(n9205), .ZN(n9013) );
  MUX2_X1 U10094 ( .A(n9014), .B(n9013), .S(n10837), .Z(n9018) );
  AOI22_X1 U10095 ( .A1(n9016), .A2(n9112), .B1(n9111), .B2(n9015), .ZN(n9017)
         );
  OAI211_X1 U10096 ( .C1(n9207), .C2(n9101), .A(n9018), .B(n9017), .ZN(
        P2_U3210) );
  XNOR2_X1 U10097 ( .A(n9020), .B(n9019), .ZN(n9211) );
  INV_X1 U10098 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U10099 ( .A1(n9021), .A2(n9103), .ZN(n9029) );
  AOI21_X1 U10100 ( .B1(n9022), .B2(n9024), .A(n9023), .ZN(n9028) );
  AOI22_X1 U10101 ( .A1(n9026), .A2(n9082), .B1(n9080), .B2(n9025), .ZN(n9027)
         );
  OAI21_X1 U10102 ( .B1(n9029), .B2(n9028), .A(n9027), .ZN(n9210) );
  INV_X1 U10103 ( .A(n9210), .ZN(n9030) );
  MUX2_X1 U10104 ( .A(n9031), .B(n9030), .S(n10837), .Z(n9035) );
  AOI22_X1 U10105 ( .A1(n9033), .A2(n9112), .B1(n9111), .B2(n9032), .ZN(n9034)
         );
  OAI211_X1 U10106 ( .C1(n9211), .C2(n9101), .A(n9035), .B(n9034), .ZN(
        P2_U3211) );
  OR2_X1 U10107 ( .A1(n9036), .A2(n9037), .ZN(n9057) );
  NAND2_X1 U10108 ( .A1(n9057), .A2(n9038), .ZN(n9040) );
  NAND3_X1 U10109 ( .A1(n9040), .A2(n9044), .A3(n9039), .ZN(n9041) );
  NAND2_X1 U10110 ( .A1(n9042), .A2(n9041), .ZN(n9216) );
  INV_X1 U10111 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9051) );
  INV_X1 U10112 ( .A(n9022), .ZN(n9046) );
  NOR3_X1 U10113 ( .A1(n4967), .A2(n9044), .A3(n9043), .ZN(n9045) );
  NOR2_X1 U10114 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  OAI222_X1 U10115 ( .A1(n9106), .A2(n9049), .B1(n9170), .B2(n9048), .C1(n9168), .C2(n9047), .ZN(n9214) );
  INV_X1 U10116 ( .A(n9214), .ZN(n9050) );
  MUX2_X1 U10117 ( .A(n9051), .B(n9050), .S(n10837), .Z(n9055) );
  AOI22_X1 U10118 ( .A1(n9053), .A2(n9112), .B1(n9111), .B2(n9052), .ZN(n9054)
         );
  OAI211_X1 U10119 ( .C1(n9216), .C2(n9101), .A(n9055), .B(n9054), .ZN(
        P2_U3212) );
  NAND2_X1 U10120 ( .A1(n9057), .A2(n9056), .ZN(n9059) );
  XNOR2_X1 U10121 ( .A(n9059), .B(n9058), .ZN(n9221) );
  INV_X1 U10122 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9066) );
  AOI21_X1 U10123 ( .B1(n9061), .B2(n9060), .A(n4967), .ZN(n9062) );
  OAI222_X1 U10124 ( .A1(n9106), .A2(n9064), .B1(n9170), .B2(n9063), .C1(n9168), .C2(n9062), .ZN(n9219) );
  INV_X1 U10125 ( .A(n9219), .ZN(n9065) );
  MUX2_X1 U10126 ( .A(n9066), .B(n9065), .S(n10837), .Z(n9069) );
  AOI22_X1 U10127 ( .A1(n9141), .A2(n9112), .B1(n9111), .B2(n9067), .ZN(n9068)
         );
  OAI211_X1 U10128 ( .C1(n9221), .C2(n9101), .A(n9069), .B(n9068), .ZN(
        P2_U3213) );
  XNOR2_X1 U10129 ( .A(n9036), .B(n9071), .ZN(n9229) );
  XOR2_X1 U10130 ( .A(n9071), .B(n9070), .Z(n9073) );
  AOI222_X1 U10131 ( .A1(n9103), .A2(n9073), .B1(n9072), .B2(n9082), .C1(
        n10846), .C2(n9080), .ZN(n9224) );
  MUX2_X1 U10132 ( .A(n6896), .B(n9224), .S(n10837), .Z(n9076) );
  AOI22_X1 U10133 ( .A1(n9226), .A2(n9112), .B1(n9111), .B2(n9074), .ZN(n9075)
         );
  OAI211_X1 U10134 ( .C1(n9229), .C2(n9101), .A(n9076), .B(n9075), .ZN(
        P2_U3214) );
  XNOR2_X1 U10135 ( .A(n9077), .B(n9078), .ZN(n9235) );
  XNOR2_X1 U10136 ( .A(n9079), .B(n9078), .ZN(n9084) );
  AOI222_X1 U10137 ( .A1(n9103), .A2(n9084), .B1(n9083), .B2(n9082), .C1(n9081), .C2(n9080), .ZN(n9230) );
  MUX2_X1 U10138 ( .A(n9085), .B(n9230), .S(n10837), .Z(n9088) );
  AOI22_X1 U10139 ( .A1(n9232), .A2(n9112), .B1(n9111), .B2(n9086), .ZN(n9087)
         );
  OAI211_X1 U10140 ( .C1(n9235), .C2(n9101), .A(n9088), .B(n9087), .ZN(
        P2_U3215) );
  XNOR2_X1 U10141 ( .A(n9090), .B(n9089), .ZN(n9238) );
  INV_X1 U10142 ( .A(n9238), .ZN(n9102) );
  INV_X1 U10143 ( .A(n9091), .ZN(n9093) );
  AOI21_X1 U10144 ( .B1(n9093), .B2(n9092), .A(n9168), .ZN(n9098) );
  OAI22_X1 U10145 ( .A1(n9095), .A2(n9170), .B1(n9094), .B2(n9106), .ZN(n9096)
         );
  AOI21_X1 U10146 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9236) );
  MUX2_X1 U10147 ( .A(n10674), .B(n9236), .S(n10837), .Z(n9100) );
  AOI22_X1 U10148 ( .A1(n10852), .A2(n9112), .B1(n9111), .B2(n10857), .ZN(
        n9099) );
  OAI211_X1 U10149 ( .C1(n9102), .C2(n9101), .A(n9100), .B(n9099), .ZN(
        P2_U3216) );
  OAI211_X1 U10150 ( .C1(n9105), .C2(n9113), .A(n9104), .B(n9103), .ZN(n9109)
         );
  OR2_X1 U10151 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  OAI211_X1 U10152 ( .C1(n9171), .C2(n9170), .A(n9109), .B(n9108), .ZN(n9153)
         );
  AOI21_X1 U10153 ( .B1(n9111), .B2(n9110), .A(n9153), .ZN(n9118) );
  AOI22_X1 U10154 ( .A1(n9243), .A2(n9112), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n10839), .ZN(n9117) );
  XNOR2_X1 U10155 ( .A(n9114), .B(n9113), .ZN(n9245) );
  NAND2_X1 U10156 ( .A1(n9245), .A2(n9115), .ZN(n9116) );
  OAI211_X1 U10157 ( .C1(n9118), .C2(n10839), .A(n9117), .B(n9116), .ZN(
        P2_U3217) );
  NOR2_X1 U10158 ( .A1(n9175), .A2(n9176), .ZN(n9120) );
  AOI21_X1 U10159 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9175), .A(n9120), .ZN(
        n9119) );
  OAI21_X1 U10160 ( .B1(n9178), .B2(n9158), .A(n9119), .ZN(P2_U3490) );
  AOI21_X1 U10161 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9175), .A(n9120), .ZN(
        n9121) );
  OAI21_X1 U10162 ( .B1(n9181), .B2(n9158), .A(n9121), .ZN(P2_U3489) );
  INV_X1 U10163 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9122) );
  MUX2_X1 U10164 ( .A(n9183), .B(n9122), .S(n9175), .Z(n9124) );
  NAND2_X1 U10165 ( .A1(n9185), .A2(n7174), .ZN(n9123) );
  OAI211_X1 U10166 ( .C1(n9188), .C2(n9159), .A(n9124), .B(n9123), .ZN(
        P2_U3486) );
  AOI21_X1 U10167 ( .B1(n9126), .B2(n9182), .A(n9125), .ZN(n9189) );
  INV_X1 U10168 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9127) );
  MUX2_X1 U10169 ( .A(n9189), .B(n9127), .S(n9175), .Z(n9128) );
  OAI21_X1 U10170 ( .B1(n9192), .B2(n9158), .A(n9128), .ZN(P2_U3485) );
  INV_X1 U10171 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U10172 ( .A(n9193), .B(n9129), .S(n9175), .Z(n9131) );
  INV_X1 U10173 ( .A(n9159), .ZN(n9155) );
  AOI22_X1 U10174 ( .A1(n9196), .A2(n9155), .B1(n7174), .B2(n9195), .ZN(n9130)
         );
  NAND2_X1 U10175 ( .A1(n9131), .A2(n9130), .ZN(P2_U3484) );
  INV_X1 U10176 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9132) );
  MUX2_X1 U10177 ( .A(n9199), .B(n9132), .S(n9175), .Z(n9134) );
  AOI22_X1 U10178 ( .A1(n9202), .A2(n9155), .B1(n7174), .B2(n9201), .ZN(n9133)
         );
  NAND2_X1 U10179 ( .A1(n9134), .A2(n9133), .ZN(P2_U3483) );
  MUX2_X1 U10180 ( .A(n9205), .B(P2_REG1_REG_23__SCAN_IN), .S(n9175), .Z(n9136) );
  OAI22_X1 U10181 ( .A1(n9207), .A2(n9159), .B1(n9206), .B2(n9158), .ZN(n9135)
         );
  OR2_X1 U10182 ( .A1(n9136), .A2(n9135), .ZN(P2_U3482) );
  MUX2_X1 U10183 ( .A(n9210), .B(P2_REG1_REG_22__SCAN_IN), .S(n9175), .Z(n9138) );
  OAI22_X1 U10184 ( .A1(n9211), .A2(n9159), .B1(n5205), .B2(n9158), .ZN(n9137)
         );
  OR2_X1 U10185 ( .A1(n9138), .A2(n9137), .ZN(P2_U3481) );
  MUX2_X1 U10186 ( .A(n9214), .B(P2_REG1_REG_21__SCAN_IN), .S(n9175), .Z(n9140) );
  OAI22_X1 U10187 ( .A1(n9216), .A2(n9159), .B1(n9215), .B2(n9158), .ZN(n9139)
         );
  OR2_X1 U10188 ( .A1(n9140), .A2(n9139), .ZN(P2_U3480) );
  MUX2_X1 U10189 ( .A(n9219), .B(P2_REG1_REG_20__SCAN_IN), .S(n9175), .Z(n9143) );
  INV_X1 U10190 ( .A(n9141), .ZN(n9220) );
  OAI22_X1 U10191 ( .A1(n9221), .A2(n9159), .B1(n9220), .B2(n9158), .ZN(n9142)
         );
  OR2_X1 U10192 ( .A1(n9143), .A2(n9142), .ZN(P2_U3479) );
  INV_X1 U10193 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9144) );
  MUX2_X1 U10194 ( .A(n9224), .B(n9144), .S(n9175), .Z(n9146) );
  NAND2_X1 U10195 ( .A1(n9226), .A2(n7174), .ZN(n9145) );
  OAI211_X1 U10196 ( .C1(n9229), .C2(n9159), .A(n9146), .B(n9145), .ZN(
        P2_U3478) );
  INV_X1 U10197 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9147) );
  MUX2_X1 U10198 ( .A(n9230), .B(n9147), .S(n9175), .Z(n9149) );
  NAND2_X1 U10199 ( .A1(n9232), .A2(n7174), .ZN(n9148) );
  OAI211_X1 U10200 ( .C1(n9235), .C2(n9159), .A(n9149), .B(n9148), .ZN(
        P2_U3477) );
  INV_X1 U10201 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9150) );
  MUX2_X1 U10202 ( .A(n9236), .B(n9150), .S(n9175), .Z(n9152) );
  AOI22_X1 U10203 ( .A1(n9238), .A2(n9155), .B1(n7174), .B2(n10852), .ZN(n9151) );
  NAND2_X1 U10204 ( .A1(n9152), .A2(n9151), .ZN(P2_U3476) );
  INV_X1 U10205 ( .A(n9153), .ZN(n9242) );
  MUX2_X1 U10206 ( .A(n9242), .B(n9154), .S(n9175), .Z(n9157) );
  AOI22_X1 U10207 ( .A1(n9245), .A2(n9155), .B1(n7174), .B2(n9243), .ZN(n9156)
         );
  NAND2_X1 U10208 ( .A1(n9157), .A2(n9156), .ZN(P2_U3475) );
  MUX2_X1 U10209 ( .A(n9248), .B(P2_REG1_REG_15__SCAN_IN), .S(n9175), .Z(n9161) );
  OAI22_X1 U10210 ( .A1(n9252), .A2(n9159), .B1(n9250), .B2(n9158), .ZN(n9160)
         );
  OR2_X1 U10211 ( .A1(n9161), .A2(n9160), .ZN(P2_U3474) );
  OAI21_X1 U10212 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n10826) );
  NOR2_X1 U10213 ( .A1(n10826), .A2(n9165), .ZN(n9172) );
  XNOR2_X1 U10214 ( .A(n9166), .B(n5168), .ZN(n9167) );
  OAI222_X1 U10215 ( .A1(n9106), .A2(n9171), .B1(n9170), .B2(n9169), .C1(n9168), .C2(n9167), .ZN(n10833) );
  AOI211_X1 U10216 ( .C1(n9173), .C2(n10827), .A(n9172), .B(n10833), .ZN(
        n10842) );
  NAND2_X1 U10217 ( .A1(n9175), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9174) );
  OAI21_X1 U10218 ( .B1(n10842), .B2(n9175), .A(n9174), .ZN(P2_U3473) );
  NOR2_X1 U10219 ( .A1(n10840), .A2(n9176), .ZN(n9179) );
  AOI21_X1 U10220 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n10840), .A(n9179), .ZN(
        n9177) );
  OAI21_X1 U10221 ( .B1(n9178), .B2(n9249), .A(n9177), .ZN(P2_U3458) );
  AOI21_X1 U10222 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n10840), .A(n9179), .ZN(
        n9180) );
  OAI21_X1 U10223 ( .B1(n9181), .B2(n9249), .A(n9180), .ZN(P2_U3457) );
  NAND2_X1 U10224 ( .A1(n10843), .A2(n9182), .ZN(n9251) );
  INV_X1 U10225 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9184) );
  MUX2_X1 U10226 ( .A(n9184), .B(n9183), .S(n10843), .Z(n9187) );
  NAND2_X1 U10227 ( .A1(n9185), .A2(n7191), .ZN(n9186) );
  OAI211_X1 U10228 ( .C1(n9188), .C2(n9251), .A(n9187), .B(n9186), .ZN(
        P2_U3454) );
  INV_X1 U10229 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U10230 ( .A(n9190), .B(n9189), .S(n10843), .Z(n9191) );
  OAI21_X1 U10231 ( .B1(n9192), .B2(n9249), .A(n9191), .ZN(P2_U3453) );
  INV_X1 U10232 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9194) );
  MUX2_X1 U10233 ( .A(n9194), .B(n9193), .S(n10843), .Z(n9198) );
  INV_X1 U10234 ( .A(n9251), .ZN(n9244) );
  AOI22_X1 U10235 ( .A1(n9196), .A2(n9244), .B1(n7191), .B2(n9195), .ZN(n9197)
         );
  NAND2_X1 U10236 ( .A1(n9198), .A2(n9197), .ZN(P2_U3452) );
  INV_X1 U10237 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9200) );
  MUX2_X1 U10238 ( .A(n9200), .B(n9199), .S(n10843), .Z(n9204) );
  AOI22_X1 U10239 ( .A1(n9202), .A2(n9244), .B1(n7191), .B2(n9201), .ZN(n9203)
         );
  NAND2_X1 U10240 ( .A1(n9204), .A2(n9203), .ZN(P2_U3451) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9205), .S(n10843), .Z(
        n9209) );
  OAI22_X1 U10242 ( .A1(n9207), .A2(n9251), .B1(n9206), .B2(n9249), .ZN(n9208)
         );
  OR2_X1 U10243 ( .A1(n9209), .A2(n9208), .ZN(P2_U3450) );
  MUX2_X1 U10244 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9210), .S(n10843), .Z(
        n9213) );
  OAI22_X1 U10245 ( .A1(n9211), .A2(n9251), .B1(n5205), .B2(n9249), .ZN(n9212)
         );
  OR2_X1 U10246 ( .A1(n9213), .A2(n9212), .ZN(P2_U3449) );
  MUX2_X1 U10247 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9214), .S(n10843), .Z(
        n9218) );
  OAI22_X1 U10248 ( .A1(n9216), .A2(n9251), .B1(n9215), .B2(n9249), .ZN(n9217)
         );
  OR2_X1 U10249 ( .A1(n9218), .A2(n9217), .ZN(P2_U3448) );
  MUX2_X1 U10250 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9219), .S(n10843), .Z(
        n9223) );
  OAI22_X1 U10251 ( .A1(n9221), .A2(n9251), .B1(n9220), .B2(n9249), .ZN(n9222)
         );
  OR2_X1 U10252 ( .A1(n9223), .A2(n9222), .ZN(P2_U3447) );
  INV_X1 U10253 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9225) );
  MUX2_X1 U10254 ( .A(n9225), .B(n9224), .S(n10843), .Z(n9228) );
  NAND2_X1 U10255 ( .A1(n9226), .A2(n7191), .ZN(n9227) );
  OAI211_X1 U10256 ( .C1(n9229), .C2(n9251), .A(n9228), .B(n9227), .ZN(
        P2_U3446) );
  INV_X1 U10257 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U10258 ( .A(n9231), .B(n9230), .S(n10843), .Z(n9234) );
  NAND2_X1 U10259 ( .A1(n9232), .A2(n7191), .ZN(n9233) );
  OAI211_X1 U10260 ( .C1(n9235), .C2(n9251), .A(n9234), .B(n9233), .ZN(
        P2_U3444) );
  INV_X1 U10261 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9237) );
  MUX2_X1 U10262 ( .A(n9237), .B(n9236), .S(n10843), .Z(n9240) );
  AOI22_X1 U10263 ( .A1(n9238), .A2(n9244), .B1(n7191), .B2(n10852), .ZN(n9239) );
  NAND2_X1 U10264 ( .A1(n9240), .A2(n9239), .ZN(P2_U3441) );
  INV_X1 U10265 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9241) );
  MUX2_X1 U10266 ( .A(n9242), .B(n9241), .S(n10840), .Z(n9247) );
  AOI22_X1 U10267 ( .A1(n9245), .A2(n9244), .B1(n7191), .B2(n9243), .ZN(n9246)
         );
  NAND2_X1 U10268 ( .A1(n9247), .A2(n9246), .ZN(P2_U3438) );
  MUX2_X1 U10269 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9248), .S(n10843), .Z(
        n9254) );
  OAI22_X1 U10270 ( .A1(n9252), .A2(n9251), .B1(n9250), .B2(n9249), .ZN(n9253)
         );
  OR2_X1 U10271 ( .A1(n9254), .A2(n9253), .ZN(P2_U3435) );
  MUX2_X1 U10272 ( .A(n9256), .B(P2_D_REG_1__SCAN_IN), .S(n9255), .Z(P2_U3377)
         );
  INV_X1 U10273 ( .A(n9257), .ZN(n9990) );
  NOR4_X1 U10274 ( .A1(n9258), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5685), .ZN(n9259) );
  AOI21_X1 U10275 ( .B1(n9260), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9259), .ZN(
        n9261) );
  OAI21_X1 U10276 ( .B1(n9990), .B2(n9266), .A(n9261), .ZN(P2_U3264) );
  INV_X1 U10277 ( .A(n9262), .ZN(n9995) );
  OAI222_X1 U10278 ( .A1(n9266), .A2(n9995), .B1(n9265), .B2(P2_U3151), .C1(
        n9264), .C2(n9263), .ZN(P2_U3266) );
  NAND2_X1 U10279 ( .A1(n9996), .A2(n9267), .ZN(n9269) );
  OAI211_X1 U10280 ( .C1(n9263), .C2(n9270), .A(n9269), .B(n9268), .ZN(
        P2_U3267) );
  MUX2_X1 U10281 ( .A(n9271), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XOR2_X1 U10282 ( .A(n9339), .B(n9272), .Z(n9277) );
  AOI22_X1 U10283 ( .A1(n9372), .A2(n9679), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9274) );
  NAND2_X1 U10284 ( .A1(n9406), .A2(n9747), .ZN(n9273) );
  OAI211_X1 U10285 ( .C1(n9409), .C2(n9711), .A(n9274), .B(n9273), .ZN(n9275)
         );
  AOI21_X1 U10286 ( .B1(n9889), .B2(n9411), .A(n9275), .ZN(n9276) );
  OAI21_X1 U10287 ( .B1(n9277), .B2(n9414), .A(n9276), .ZN(P1_U3216) );
  XOR2_X1 U10288 ( .A(n9279), .B(n9278), .Z(n9285) );
  NAND2_X1 U10289 ( .A1(n9781), .A2(n9406), .ZN(n9280) );
  NAND2_X1 U10290 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9550) );
  OAI211_X1 U10291 ( .C1(n9281), .C2(n9404), .A(n9280), .B(n9550), .ZN(n9282)
         );
  AOI21_X1 U10292 ( .B1(n9792), .B2(n9395), .A(n9282), .ZN(n9284) );
  NAND2_X1 U10293 ( .A1(n9791), .A2(n9411), .ZN(n9283) );
  OAI211_X1 U10294 ( .C1(n9285), .C2(n9414), .A(n9284), .B(n9283), .ZN(
        P1_U3219) );
  NAND2_X1 U10295 ( .A1(n9638), .A2(n7491), .ZN(n9287) );
  OR2_X1 U10296 ( .A1(n9618), .A2(n7350), .ZN(n9286) );
  NAND2_X1 U10297 ( .A1(n9287), .A2(n9286), .ZN(n9289) );
  XNOR2_X1 U10298 ( .A(n9289), .B(n9288), .ZN(n9292) );
  NAND2_X1 U10299 ( .A1(n9638), .A2(n8722), .ZN(n9290) );
  OAI21_X1 U10300 ( .B1(n9618), .B2(n7349), .A(n9290), .ZN(n9291) );
  XNOR2_X1 U10301 ( .A(n9292), .B(n9291), .ZN(n9299) );
  INV_X1 U10302 ( .A(n9300), .ZN(n9293) );
  NAND2_X1 U10303 ( .A1(n9293), .A2(n9390), .ZN(n9294) );
  NAND3_X1 U10304 ( .A1(n9295), .A2(n9390), .A3(n9299), .ZN(n9303) );
  AOI22_X1 U10305 ( .A1(n9372), .A2(n9634), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9297) );
  NAND2_X1 U10306 ( .A1(n9406), .A2(n9633), .ZN(n9296) );
  OAI211_X1 U10307 ( .C1(n9409), .C2(n9627), .A(n9297), .B(n9296), .ZN(n9298)
         );
  AOI21_X1 U10308 ( .B1(n9638), .B2(n9411), .A(n9298), .ZN(n9302) );
  NAND3_X1 U10309 ( .A1(n9300), .A2(n9299), .A3(n9390), .ZN(n9301) );
  NAND4_X1 U10310 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(
        P1_U3220) );
  XOR2_X1 U10311 ( .A(n9306), .B(n9305), .Z(n9311) );
  AOI22_X1 U10312 ( .A1(n9372), .A2(n9747), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9308) );
  NAND2_X1 U10313 ( .A1(n9406), .A2(n9782), .ZN(n9307) );
  OAI211_X1 U10314 ( .C1(n9409), .C2(n9755), .A(n9308), .B(n9307), .ZN(n9309)
         );
  AOI21_X1 U10315 ( .B1(n9754), .B2(n9411), .A(n9309), .ZN(n9310) );
  OAI21_X1 U10316 ( .B1(n9311), .B2(n9414), .A(n9310), .ZN(P1_U3223) );
  OAI21_X1 U10317 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9315) );
  NAND2_X1 U10318 ( .A1(n9315), .A2(n9390), .ZN(n9321) );
  INV_X1 U10319 ( .A(n9316), .ZN(n9683) );
  AOI22_X1 U10320 ( .A1(n9372), .A2(n9680), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9317) );
  OAI21_X1 U10321 ( .B1(n9718), .B2(n9318), .A(n9317), .ZN(n9319) );
  AOI21_X1 U10322 ( .B1(n9683), .B2(n9395), .A(n9319), .ZN(n9320) );
  OAI211_X1 U10323 ( .C1(n9685), .C2(n9398), .A(n9321), .B(n9320), .ZN(
        P1_U3225) );
  XOR2_X1 U10324 ( .A(n9322), .B(n9323), .Z(n9329) );
  NAND2_X1 U10325 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10430)
         );
  OAI21_X1 U10326 ( .B1(n9404), .B2(n9324), .A(n10430), .ZN(n9325) );
  AOI21_X1 U10327 ( .B1(n9406), .B2(n9829), .A(n9325), .ZN(n9326) );
  OAI21_X1 U10328 ( .B1(n9409), .B2(n9821), .A(n9326), .ZN(n9327) );
  AOI21_X1 U10329 ( .B1(n9930), .B2(n9411), .A(n9327), .ZN(n9328) );
  OAI21_X1 U10330 ( .B1(n9329), .B2(n9414), .A(n9328), .ZN(P1_U3226) );
  XOR2_X1 U10331 ( .A(n9330), .B(n9331), .Z(n9338) );
  NAND2_X1 U10332 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10401)
         );
  OAI21_X1 U10333 ( .B1(n9332), .B2(n9404), .A(n10401), .ZN(n9333) );
  AOI21_X1 U10334 ( .B1(n9406), .B2(n9417), .A(n9333), .ZN(n9334) );
  OAI21_X1 U10335 ( .B1(n9409), .B2(n9335), .A(n9334), .ZN(n9336) );
  AOI21_X1 U10336 ( .B1(n9577), .B2(n9411), .A(n9336), .ZN(n9337) );
  OAI21_X1 U10337 ( .B1(n9338), .B2(n9414), .A(n9337), .ZN(P1_U3228) );
  OR2_X1 U10338 ( .A1(n9272), .A2(n9339), .ZN(n9341) );
  NAND2_X1 U10339 ( .A1(n9341), .A2(n9340), .ZN(n9345) );
  NAND2_X1 U10340 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  XNOR2_X1 U10341 ( .A(n9345), .B(n9344), .ZN(n9350) );
  INV_X1 U10342 ( .A(n9702), .ZN(n9592) );
  AOI22_X1 U10343 ( .A1(n9372), .A2(n9592), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9347) );
  NAND2_X1 U10344 ( .A1(n9406), .A2(n9587), .ZN(n9346) );
  OAI211_X1 U10345 ( .C1(n9409), .C2(n9696), .A(n9347), .B(n9346), .ZN(n9348)
         );
  AOI21_X1 U10346 ( .B1(n9885), .B2(n9411), .A(n9348), .ZN(n9349) );
  OAI21_X1 U10347 ( .B1(n9350), .B2(n9414), .A(n9349), .ZN(P1_U3229) );
  XOR2_X1 U10348 ( .A(n9352), .B(n9351), .Z(n9357) );
  NAND2_X1 U10349 ( .A1(n9809), .A2(n9406), .ZN(n9354) );
  INV_X1 U10350 ( .A(n9771), .ZN(n9583) );
  AOI22_X1 U10351 ( .A1(n9372), .A2(n9583), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9353) );
  OAI211_X1 U10352 ( .C1(n9409), .C2(n9763), .A(n9354), .B(n9353), .ZN(n9355)
         );
  AOI21_X1 U10353 ( .B1(n9906), .B2(n9411), .A(n9355), .ZN(n9356) );
  OAI21_X1 U10354 ( .B1(n9357), .B2(n9414), .A(n9356), .ZN(P1_U3233) );
  NAND2_X1 U10355 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  XOR2_X1 U10356 ( .A(n9361), .B(n9360), .Z(n9366) );
  AOI22_X1 U10357 ( .A1(n9372), .A2(n9587), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9363) );
  NAND2_X1 U10358 ( .A1(n9406), .A2(n9583), .ZN(n9362) );
  OAI211_X1 U10359 ( .C1(n9409), .C2(n9734), .A(n9363), .B(n9362), .ZN(n9364)
         );
  AOI21_X1 U10360 ( .B1(n9736), .B2(n9411), .A(n9364), .ZN(n9365) );
  OAI21_X1 U10361 ( .B1(n9366), .B2(n9414), .A(n9365), .ZN(P1_U3235) );
  INV_X1 U10362 ( .A(n9367), .ZN(n9370) );
  NOR3_X1 U10363 ( .A1(n7461), .A2(n4945), .A3(n9368), .ZN(n9369) );
  OAI21_X1 U10364 ( .B1(n9370), .B2(n9369), .A(n9390), .ZN(n9376) );
  AOI22_X1 U10365 ( .A1(n9372), .A2(n10226), .B1(n9411), .B2(n9371), .ZN(n9375) );
  AOI22_X1 U10366 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n9373), .B1(n9406), .B2(
        n10228), .ZN(n9374) );
  NAND3_X1 U10367 ( .A1(n9376), .A2(n9375), .A3(n9374), .ZN(P1_U3237) );
  NAND2_X1 U10368 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  XOR2_X1 U10369 ( .A(n9380), .B(n9379), .Z(n9385) );
  NAND2_X1 U10370 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10417)
         );
  OAI21_X1 U10371 ( .B1(n9769), .B2(n9404), .A(n10417), .ZN(n9381) );
  AOI21_X1 U10372 ( .B1(n9406), .B2(n9830), .A(n9381), .ZN(n9382) );
  OAI21_X1 U10373 ( .B1(n9409), .B2(n9800), .A(n9382), .ZN(n9383) );
  AOI21_X1 U10374 ( .B1(n9919), .B2(n9411), .A(n9383), .ZN(n9384) );
  OAI21_X1 U10375 ( .B1(n9385), .B2(n9414), .A(n9384), .ZN(P1_U3238) );
  INV_X1 U10376 ( .A(n9312), .ZN(n9388) );
  OAI21_X1 U10377 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9391) );
  NAND3_X1 U10378 ( .A1(n9391), .A2(n9390), .A3(n9389), .ZN(n9397) );
  INV_X1 U10379 ( .A(n9392), .ZN(n9671) );
  AOI22_X1 U10380 ( .A1(n9406), .A2(n9592), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9393) );
  OAI21_X1 U10381 ( .B1(n9666), .B2(n9404), .A(n9393), .ZN(n9394) );
  AOI21_X1 U10382 ( .B1(n9671), .B2(n9395), .A(n9394), .ZN(n9396) );
  OAI211_X1 U10383 ( .C1(n9952), .C2(n9398), .A(n9397), .B(n9396), .ZN(
        P1_U3240) );
  XNOR2_X1 U10384 ( .A(n9400), .B(n9399), .ZN(n9401) );
  XNOR2_X1 U10385 ( .A(n9402), .B(n9401), .ZN(n9415) );
  NAND2_X1 U10386 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10389)
         );
  OAI21_X1 U10387 ( .B1(n9404), .B2(n9403), .A(n10389), .ZN(n9405) );
  AOI21_X1 U10388 ( .B1(n9406), .B2(n9418), .A(n9405), .ZN(n9407) );
  OAI21_X1 U10389 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n9410) );
  AOI21_X1 U10390 ( .B1(n9412), .B2(n9411), .A(n9410), .ZN(n9413) );
  OAI21_X1 U10391 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(P1_U3241) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9416), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10393 ( .A(n9634), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9427), .Z(
        P1_U3583) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9595), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9633), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9592), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10397 ( .A(n9679), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9427), .Z(
        P1_U3578) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9587), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10399 ( .A(n9747), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9427), .Z(
        P1_U3576) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9583), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9782), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10402 ( .A(n9781), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9427), .Z(
        P1_U3572) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9417), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10404 ( .A(n9829), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9427), .Z(
        P1_U3569) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9418), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10406 ( .A(n9419), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9427), .Z(
        P1_U3567) );
  MUX2_X1 U10407 ( .A(n9420), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9427), .Z(
        P1_U3566) );
  MUX2_X1 U10408 ( .A(n9421), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9427), .Z(
        P1_U3565) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9422), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9423), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9424), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9425), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10413 ( .A(n9426), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9427), .Z(
        P1_U3558) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10226), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10415 ( .A(n6363), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9427), .Z(
        P1_U3556) );
  MUX2_X1 U10416 ( .A(n10228), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9427), .Z(
        P1_U3555) );
  MUX2_X1 U10417 ( .A(n7351), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9427), .Z(
        P1_U3554) );
  MUX2_X1 U10418 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9428), .S(n9452), .Z(n9433)
         );
  AND2_X1 U10419 ( .A1(n10302), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U10420 ( .A1(n9430), .A2(n9429), .ZN(n10304) );
  OR2_X1 U10421 ( .A1(n10304), .A2(n9431), .ZN(n10470) );
  NAND2_X1 U10422 ( .A1(n9433), .A2(n9432), .ZN(n9449) );
  OAI211_X1 U10423 ( .C1(n9433), .C2(n9432), .A(n10685), .B(n9449), .ZN(n9439)
         );
  MUX2_X1 U10424 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6349), .S(n9452), .Z(n9435)
         );
  AND2_X1 U10425 ( .A1(n10302), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9434) );
  OR2_X1 U10426 ( .A1(n10304), .A2(n10298), .ZN(n10466) );
  NAND2_X1 U10427 ( .A1(n9435), .A2(n9434), .ZN(n9454) );
  OAI211_X1 U10428 ( .C1(n9435), .C2(n9434), .A(n10689), .B(n9454), .ZN(n9438)
         );
  AOI22_X1 U10429 ( .A1(n10683), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9437) );
  INV_X1 U10430 ( .A(n10461), .ZN(n10693) );
  NAND2_X1 U10431 ( .A1(n10693), .A2(n9452), .ZN(n9436) );
  NAND4_X1 U10432 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(
        P1_U3244) );
  NOR2_X1 U10433 ( .A1(n9440), .A2(n10298), .ZN(n10300) );
  INV_X1 U10434 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10714) );
  NOR2_X1 U10435 ( .A1(n9440), .A2(n10714), .ZN(n10299) );
  XOR2_X1 U10436 ( .A(n10302), .B(n10299), .Z(n9443) );
  OAI21_X1 U10437 ( .B1(n8680), .B2(n9441), .A(n10300), .ZN(n9442) );
  OAI211_X1 U10438 ( .C1(n10300), .C2(n9443), .A(n9442), .B(P1_U3973), .ZN(
        n10697) );
  NAND2_X1 U10439 ( .A1(n10683), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U10440 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9444) );
  OAI211_X1 U10441 ( .C1(n10461), .C2(n9446), .A(n9445), .B(n9444), .ZN(n9447)
         );
  INV_X1 U10442 ( .A(n9447), .ZN(n9459) );
  INV_X1 U10443 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10236) );
  MUX2_X1 U10444 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10236), .S(n9469), .Z(n9451) );
  NAND2_X1 U10445 ( .A1(n9452), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U10446 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  NAND2_X1 U10447 ( .A1(n9451), .A2(n9450), .ZN(n9471) );
  OAI211_X1 U10448 ( .C1(n9451), .C2(n9450), .A(n10685), .B(n9471), .ZN(n9458)
         );
  MUX2_X1 U10449 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6330), .S(n9469), .Z(n9456)
         );
  NAND2_X1 U10450 ( .A1(n9452), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U10451 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  NAND2_X1 U10452 ( .A1(n9456), .A2(n9455), .ZN(n9465) );
  OAI211_X1 U10453 ( .C1(n9456), .C2(n9455), .A(n10689), .B(n9465), .ZN(n9457)
         );
  NAND4_X1 U10454 ( .A1(n10697), .A2(n9459), .A3(n9458), .A4(n9457), .ZN(
        P1_U3245) );
  INV_X1 U10455 ( .A(n10683), .ZN(n10480) );
  INV_X1 U10456 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9461) );
  OAI21_X1 U10457 ( .B1(n10480), .B2(n9461), .A(n9460), .ZN(n9462) );
  AOI21_X1 U10458 ( .B1(n9486), .B2(n10693), .A(n9462), .ZN(n9476) );
  XNOR2_X1 U10459 ( .A(n9486), .B(n9463), .ZN(n9467) );
  NAND2_X1 U10460 ( .A1(n9469), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U10461 ( .A1(n9465), .A2(n9464), .ZN(n9466) );
  NAND2_X1 U10462 ( .A1(n9466), .A2(n9467), .ZN(n9482) );
  OAI211_X1 U10463 ( .C1(n9467), .C2(n9466), .A(n10689), .B(n9482), .ZN(n9475)
         );
  INV_X1 U10464 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9468) );
  XNOR2_X1 U10465 ( .A(n9486), .B(n9468), .ZN(n9473) );
  NAND2_X1 U10466 ( .A1(n9469), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U10467 ( .A1(n9471), .A2(n9470), .ZN(n9472) );
  NAND2_X1 U10468 ( .A1(n9472), .A2(n9473), .ZN(n9488) );
  OAI211_X1 U10469 ( .C1(n9473), .C2(n9472), .A(n10685), .B(n9488), .ZN(n9474)
         );
  NAND3_X1 U10470 ( .A1(n9476), .A2(n9475), .A3(n9474), .ZN(P1_U3246) );
  INV_X1 U10471 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9478) );
  OAI21_X1 U10472 ( .B1(n10480), .B2(n9478), .A(n9477), .ZN(n9479) );
  AOI21_X1 U10473 ( .B1(n9506), .B2(n10693), .A(n9479), .ZN(n9495) );
  MUX2_X1 U10474 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9480), .S(n9506), .Z(n9485)
         );
  NAND2_X1 U10475 ( .A1(n9486), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U10476 ( .A1(n9482), .A2(n9481), .ZN(n10690) );
  XNOR2_X1 U10477 ( .A(n9489), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U10478 ( .A1(n10690), .A2(n10691), .ZN(n10688) );
  INV_X1 U10479 ( .A(n9489), .ZN(n10692) );
  NAND2_X1 U10480 ( .A1(n10692), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U10481 ( .A1(n10688), .A2(n9483), .ZN(n9484) );
  NAND2_X1 U10482 ( .A1(n9484), .A2(n9485), .ZN(n9508) );
  OAI211_X1 U10483 ( .C1(n9485), .C2(n9484), .A(n10689), .B(n9508), .ZN(n9494)
         );
  MUX2_X1 U10484 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7699), .S(n9506), .Z(n9492)
         );
  NAND2_X1 U10485 ( .A1(n9486), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U10486 ( .A1(n9488), .A2(n9487), .ZN(n10686) );
  XNOR2_X1 U10487 ( .A(n9489), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10687) );
  NAND2_X1 U10488 ( .A1(n10686), .A2(n10687), .ZN(n10684) );
  NAND2_X1 U10489 ( .A1(n10692), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U10490 ( .A1(n10684), .A2(n9490), .ZN(n9491) );
  NAND2_X1 U10491 ( .A1(n9491), .A2(n9492), .ZN(n9498) );
  OAI211_X1 U10492 ( .C1(n9492), .C2(n9491), .A(n10685), .B(n9498), .ZN(n9493)
         );
  NAND3_X1 U10493 ( .A1(n9495), .A2(n9494), .A3(n9493), .ZN(P1_U3248) );
  NOR2_X1 U10494 ( .A1(n9537), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9496) );
  AOI21_X1 U10495 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9537), .A(n9496), .ZN(
        n9502) );
  NAND2_X1 U10496 ( .A1(n9506), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U10497 ( .A1(n9498), .A2(n9497), .ZN(n10308) );
  MUX2_X1 U10498 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7846), .S(n10313), .Z(
        n10309) );
  AND2_X1 U10499 ( .A1(n10308), .A2(n10309), .ZN(n10306) );
  AOI21_X1 U10500 ( .B1(n10313), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10306), .ZN(
        n10327) );
  NAND2_X1 U10501 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n10325), .ZN(n9499) );
  OAI21_X1 U10502 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n10325), .A(n9499), .ZN(
        n10328) );
  NOR2_X1 U10503 ( .A1(n10327), .A2(n10328), .ZN(n10326) );
  AOI21_X1 U10504 ( .B1(n10325), .B2(P1_REG2_REG_7__SCAN_IN), .A(n10326), .ZN(
        n10338) );
  NAND2_X1 U10505 ( .A1(n10336), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9500) );
  OAI21_X1 U10506 ( .B1(n10336), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9500), .ZN(
        n10339) );
  NOR2_X1 U10507 ( .A1(n10338), .A2(n10339), .ZN(n10337) );
  AOI21_X1 U10508 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10336), .A(n10337), .ZN(
        n9501) );
  NAND2_X1 U10509 ( .A1(n9502), .A2(n9501), .ZN(n9536) );
  OAI21_X1 U10510 ( .B1(n9502), .B2(n9501), .A(n9536), .ZN(n9503) );
  NAND2_X1 U10511 ( .A1(n9503), .A2(n10685), .ZN(n9519) );
  AOI21_X1 U10512 ( .B1(n10683), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9504), .ZN(
        n9518) );
  NOR2_X1 U10513 ( .A1(n9537), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9505) );
  AOI21_X1 U10514 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9537), .A(n9505), .ZN(
        n9514) );
  NAND2_X1 U10515 ( .A1(n9506), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U10516 ( .A1(n9508), .A2(n9507), .ZN(n10311) );
  INV_X1 U10517 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10770) );
  MUX2_X1 U10518 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10770), .S(n10313), .Z(
        n10312) );
  NAND2_X1 U10519 ( .A1(n10311), .A2(n10312), .ZN(n10310) );
  NAND2_X1 U10520 ( .A1(n10313), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9509) );
  AND2_X1 U10521 ( .A1(n10310), .A2(n9509), .ZN(n10321) );
  NAND2_X1 U10522 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n10325), .ZN(n9510) );
  OAI21_X1 U10523 ( .B1(n10325), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9510), .ZN(
        n10320) );
  NOR2_X1 U10524 ( .A1(n10321), .A2(n10320), .ZN(n10322) );
  AOI21_X1 U10525 ( .B1(n10325), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10322), .ZN(
        n10342) );
  OR2_X1 U10526 ( .A1(n10336), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U10527 ( .A1(n10336), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U10528 ( .A1(n9512), .A2(n9511), .ZN(n10343) );
  NOR2_X1 U10529 ( .A1(n10342), .A2(n10343), .ZN(n10341) );
  AOI21_X1 U10530 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10336), .A(n10341), .ZN(
        n9513) );
  NAND2_X1 U10531 ( .A1(n9514), .A2(n9513), .ZN(n9523) );
  OAI21_X1 U10532 ( .B1(n9514), .B2(n9513), .A(n9523), .ZN(n9515) );
  NAND2_X1 U10533 ( .A1(n9515), .A2(n10689), .ZN(n9517) );
  NAND2_X1 U10534 ( .A1(n10693), .A2(n9537), .ZN(n9516) );
  NAND4_X1 U10535 ( .A1(n9519), .A2(n9518), .A3(n9517), .A4(n9516), .ZN(
        P1_U3252) );
  OR2_X1 U10536 ( .A1(n10399), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9529) );
  XNOR2_X1 U10537 ( .A(n10399), .B(n9926), .ZN(n10397) );
  XNOR2_X1 U10538 ( .A(n9546), .B(n9520), .ZN(n10421) );
  MUX2_X1 U10539 ( .A(n9521), .B(P1_REG1_REG_13__SCAN_IN), .S(n10433), .Z(
        n10440) );
  OR2_X1 U10540 ( .A1(n10449), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9526) );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9522), .S(n10449), .Z(
        n10451) );
  OAI21_X1 U10542 ( .B1(n9537), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9523), .ZN(
        n10469) );
  MUX2_X1 U10543 ( .A(n9524), .B(P1_REG1_REG_10__SCAN_IN), .S(n10476), .Z(
        n10468) );
  NOR2_X1 U10544 ( .A1(n10469), .A2(n10468), .ZN(n10467) );
  AOI21_X1 U10545 ( .B1(n10476), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10467), 
        .ZN(n10357) );
  MUX2_X1 U10546 ( .A(n9525), .B(P1_REG1_REG_11__SCAN_IN), .S(n10360), .Z(
        n10356) );
  NOR2_X1 U10547 ( .A1(n10357), .A2(n10356), .ZN(n10355) );
  AOI21_X1 U10548 ( .B1(n10360), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10355), 
        .ZN(n10452) );
  NAND2_X1 U10549 ( .A1(n10451), .A2(n10452), .ZN(n10450) );
  NAND2_X1 U10550 ( .A1(n9526), .A2(n10450), .ZN(n10439) );
  NOR2_X1 U10551 ( .A1(n10440), .A2(n10439), .ZN(n10438) );
  AOI21_X1 U10552 ( .B1(n10433), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10438), 
        .ZN(n10367) );
  XNOR2_X1 U10553 ( .A(n10364), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10366) );
  NOR2_X1 U10554 ( .A1(n10367), .A2(n10366), .ZN(n10365) );
  AOI21_X1 U10555 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10364), .A(n10365), 
        .ZN(n9527) );
  NOR2_X1 U10556 ( .A1(n9527), .A2(n9543), .ZN(n9528) );
  XNOR2_X1 U10557 ( .A(n9543), .B(n9527), .ZN(n10382) );
  NOR2_X1 U10558 ( .A1(n10381), .A2(n10382), .ZN(n10380) );
  NOR2_X1 U10559 ( .A1(n9528), .A2(n10380), .ZN(n10422) );
  NAND2_X1 U10560 ( .A1(n10421), .A2(n10422), .ZN(n10420) );
  OAI21_X1 U10561 ( .B1(n9546), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10420), .ZN(
        n10396) );
  NAND2_X1 U10562 ( .A1(n10397), .A2(n10396), .ZN(n10395) );
  AND2_X1 U10563 ( .A1(n9529), .A2(n10395), .ZN(n10404) );
  NAND2_X1 U10564 ( .A1(n10413), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9531) );
  OAI21_X1 U10565 ( .B1(n10413), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9531), .ZN(
        n10405) );
  INV_X1 U10566 ( .A(n10405), .ZN(n9530) );
  NAND2_X1 U10567 ( .A1(n10404), .A2(n9530), .ZN(n10408) );
  NAND2_X1 U10568 ( .A1(n10408), .A2(n9531), .ZN(n9533) );
  XNOR2_X1 U10569 ( .A(n9552), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9532) );
  XNOR2_X1 U10570 ( .A(n9533), .B(n9532), .ZN(n9556) );
  NAND2_X1 U10571 ( .A1(n10413), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9547) );
  OAI21_X1 U10572 ( .B1(n10413), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9547), .ZN(
        n10410) );
  NOR2_X1 U10573 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10399), .ZN(n9534) );
  AOI21_X1 U10574 ( .B1(n10399), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9534), .ZN(
        n10394) );
  NOR2_X1 U10575 ( .A1(n10449), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9535) );
  AOI21_X1 U10576 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10449), .A(n9535), .ZN(
        n10456) );
  OAI21_X1 U10577 ( .B1(n9537), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9536), .ZN(
        n10473) );
  NAND2_X1 U10578 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10476), .ZN(n9538) );
  OAI21_X1 U10579 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10476), .A(n9538), .ZN(
        n10472) );
  NOR2_X1 U10580 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  AOI21_X1 U10581 ( .B1(n10476), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10471), 
        .ZN(n10354) );
  NAND2_X1 U10582 ( .A1(n10360), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9539) );
  OAI21_X1 U10583 ( .B1(n10360), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9539), .ZN(
        n10353) );
  NOR2_X1 U10584 ( .A1(n10354), .A2(n10353), .ZN(n10352) );
  AOI21_X1 U10585 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10360), .A(n10352), 
        .ZN(n10455) );
  NAND2_X1 U10586 ( .A1(n10456), .A2(n10455), .ZN(n10454) );
  OAI21_X1 U10587 ( .B1(n10449), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10454), 
        .ZN(n10435) );
  NAND2_X1 U10588 ( .A1(n10433), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9540) );
  OAI21_X1 U10589 ( .B1(n10433), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9540), .ZN(
        n10436) );
  NOR2_X1 U10590 ( .A1(n10435), .A2(n10436), .ZN(n10434) );
  AOI21_X1 U10591 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10433), .A(n10434), 
        .ZN(n10370) );
  NAND2_X1 U10592 ( .A1(n10364), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9541) );
  OAI21_X1 U10593 ( .B1(n10364), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9541), .ZN(
        n10371) );
  NOR2_X1 U10594 ( .A1(n10370), .A2(n10371), .ZN(n10369) );
  AOI21_X1 U10595 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10364), .A(n10369), 
        .ZN(n9542) );
  NOR2_X1 U10596 ( .A1(n9542), .A2(n9543), .ZN(n9544) );
  XNOR2_X1 U10597 ( .A(n9543), .B(n9542), .ZN(n10385) );
  NOR2_X1 U10598 ( .A1(n10384), .A2(n10385), .ZN(n10383) );
  NOR2_X1 U10599 ( .A1(n9544), .A2(n10383), .ZN(n10426) );
  NAND2_X1 U10600 ( .A1(n9546), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9545) );
  OAI21_X1 U10601 ( .B1(n9546), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9545), .ZN(
        n10425) );
  NOR2_X1 U10602 ( .A1(n10426), .A2(n10425), .ZN(n10424) );
  AOI21_X1 U10603 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9546), .A(n10424), .ZN(
        n10393) );
  NAND2_X1 U10604 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  OAI21_X1 U10605 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10399), .A(n10392), 
        .ZN(n10409) );
  OR2_X1 U10606 ( .A1(n10410), .A2(n10409), .ZN(n10412) );
  NAND2_X1 U10607 ( .A1(n10412), .A2(n9547), .ZN(n9549) );
  XNOR2_X1 U10608 ( .A(n10222), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9548) );
  XNOR2_X1 U10609 ( .A(n9549), .B(n9548), .ZN(n9554) );
  NAND2_X1 U10610 ( .A1(n10683), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9551) );
  OAI211_X1 U10611 ( .C1(n10461), .C2(n9552), .A(n9551), .B(n9550), .ZN(n9553)
         );
  AOI21_X1 U10612 ( .B1(n10685), .B2(n9554), .A(n9553), .ZN(n9555) );
  OAI21_X1 U10613 ( .B1(n9556), .B2(n10466), .A(n9555), .ZN(P1_U3262) );
  NAND2_X1 U10614 ( .A1(n9774), .A2(n9965), .ZN(n9732) );
  NOR2_X2 U10615 ( .A1(n9640), .A2(n9560), .ZN(n9599) );
  NAND2_X1 U10616 ( .A1(n9940), .A2(n9599), .ZN(n9571) );
  INV_X1 U10617 ( .A(P1_B_REG_SCAN_IN), .ZN(n9564) );
  OR2_X1 U10618 ( .A1(n9565), .A2(n9564), .ZN(n9566) );
  NAND2_X1 U10619 ( .A1(n10225), .A2(n9566), .ZN(n9617) );
  NOR2_X1 U10620 ( .A1(n9853), .A2(n4932), .ZN(n9573) );
  NOR2_X1 U10621 ( .A1(n9561), .A2(n10237), .ZN(n9569) );
  AOI211_X1 U10622 ( .C1(n4932), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9573), .B(
        n9569), .ZN(n9570) );
  OAI21_X1 U10623 ( .B1(n9850), .B2(n9739), .A(n9570), .ZN(P1_U3263) );
  OAI211_X1 U10624 ( .C1(n9940), .C2(n9599), .A(n9562), .B(n9571), .ZN(n9854)
         );
  NOR2_X1 U10625 ( .A1(n9940), .A2(n10237), .ZN(n9572) );
  AOI211_X1 U10626 ( .C1(n4932), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9573), .B(
        n9572), .ZN(n9574) );
  OAI21_X1 U10627 ( .B1(n9854), .B2(n9739), .A(n9574), .ZN(P1_U3264) );
  INV_X1 U10628 ( .A(n9797), .ZN(n9578) );
  OR2_X1 U10629 ( .A1(n9919), .A2(n9781), .ZN(n9579) );
  NAND2_X1 U10630 ( .A1(n9791), .A2(n9809), .ZN(n9580) );
  OR2_X1 U10631 ( .A1(n9906), .A2(n9782), .ZN(n9582) );
  NAND2_X1 U10632 ( .A1(n9762), .A2(n9582), .ZN(n9750) );
  NAND2_X1 U10633 ( .A1(n9750), .A2(n9751), .ZN(n9585) );
  OR2_X1 U10634 ( .A1(n9754), .A2(n9583), .ZN(n9584) );
  NAND2_X1 U10635 ( .A1(n9736), .A2(n9747), .ZN(n9586) );
  OR2_X1 U10636 ( .A1(n9885), .A2(n9679), .ZN(n9588) );
  NAND2_X1 U10637 ( .A1(n9589), .A2(n9588), .ZN(n9690) );
  NAND2_X1 U10638 ( .A1(n9879), .A2(n9592), .ZN(n9593) );
  OR2_X1 U10639 ( .A1(n9672), .A2(n9680), .ZN(n9594) );
  AOI211_X1 U10640 ( .C1(n9560), .C2(n9640), .A(n9819), .B(n9599), .ZN(n9857)
         );
  NOR2_X1 U10641 ( .A1(n9860), .A2(n10237), .ZN(n9603) );
  INV_X1 U10642 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9601) );
  OAI22_X1 U10643 ( .A1(n10712), .A2(n9601), .B1(n9600), .B2(n10709), .ZN(
        n9602) );
  AOI211_X1 U10644 ( .C1(n9857), .C2(n9844), .A(n9603), .B(n9602), .ZN(n9623)
         );
  NAND2_X1 U10645 ( .A1(n9727), .A2(n9728), .ZN(n9607) );
  NAND2_X1 U10646 ( .A1(n9678), .A2(n9610), .ZN(n9664) );
  NAND2_X1 U10647 ( .A1(n9664), .A2(n9665), .ZN(n9663) );
  NAND2_X1 U10648 ( .A1(n9615), .A2(n10230), .ZN(n9621) );
  INV_X1 U10649 ( .A(n9619), .ZN(n9620) );
  NAND2_X1 U10650 ( .A1(n9621), .A2(n9620), .ZN(n9858) );
  NAND2_X1 U10651 ( .A1(n9858), .A2(n10235), .ZN(n9622) );
  OAI211_X1 U10652 ( .C1(n9835), .C2(n9861), .A(n9623), .B(n9622), .ZN(
        P1_U3356) );
  NAND2_X1 U10653 ( .A1(n9624), .A2(n9630), .ZN(n9625) );
  NAND2_X1 U10654 ( .A1(n9864), .A2(n9842), .ZN(n9644) );
  INV_X1 U10655 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9628) );
  OAI22_X1 U10656 ( .A1(n10712), .A2(n9628), .B1(n9627), .B2(n10709), .ZN(
        n9629) );
  AOI21_X1 U10657 ( .B1(n9638), .B2(n9840), .A(n9629), .ZN(n9643) );
  XNOR2_X1 U10658 ( .A(n9631), .B(n9630), .ZN(n9632) );
  NAND2_X1 U10659 ( .A1(n9632), .A2(n10230), .ZN(n9636) );
  AOI22_X1 U10660 ( .A1(n10225), .A2(n9634), .B1(n9633), .B2(n10227), .ZN(
        n9635) );
  NAND2_X1 U10661 ( .A1(n9636), .A2(n9635), .ZN(n9862) );
  NAND2_X1 U10662 ( .A1(n9862), .A2(n10235), .ZN(n9642) );
  AOI21_X1 U10663 ( .B1(n9638), .B2(n9637), .A(n9819), .ZN(n9639) );
  AND2_X1 U10664 ( .A1(n9640), .A2(n9639), .ZN(n9863) );
  NAND2_X1 U10665 ( .A1(n9863), .A2(n9844), .ZN(n9641) );
  NAND4_X1 U10666 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(
        P1_U3265) );
  XNOR2_X1 U10667 ( .A(n9645), .B(n9648), .ZN(n9869) );
  INV_X1 U10668 ( .A(n9869), .ZN(n9660) );
  OAI21_X1 U10669 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9649) );
  NAND2_X1 U10670 ( .A1(n9649), .A2(n10230), .ZN(n9651) );
  AOI22_X1 U10671 ( .A1(n9595), .A2(n10225), .B1(n10227), .B2(n9680), .ZN(
        n9650) );
  NAND2_X1 U10672 ( .A1(n9651), .A2(n9650), .ZN(n9867) );
  AOI211_X1 U10673 ( .C1(n9654), .C2(n9669), .A(n9819), .B(n9653), .ZN(n9868)
         );
  NAND2_X1 U10674 ( .A1(n9868), .A2(n9844), .ZN(n9657) );
  AOI22_X1 U10675 ( .A1(n4932), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9655), .B2(
        n9822), .ZN(n9656) );
  OAI211_X1 U10676 ( .C1(n9948), .C2(n10237), .A(n9657), .B(n9656), .ZN(n9658)
         );
  AOI21_X1 U10677 ( .B1(n9867), .B2(n10235), .A(n9658), .ZN(n9659) );
  OAI21_X1 U10678 ( .B1(n9660), .B2(n9835), .A(n9659), .ZN(P1_U3266) );
  XNOR2_X1 U10679 ( .A(n9662), .B(n9661), .ZN(n9874) );
  OAI21_X1 U10680 ( .B1(n9665), .B2(n9664), .A(n9663), .ZN(n9668) );
  OAI22_X1 U10681 ( .A1(n9702), .A2(n9770), .B1(n9666), .B2(n10704), .ZN(n9667) );
  AOI21_X1 U10682 ( .B1(n9668), .B2(n10230), .A(n9667), .ZN(n9873) );
  INV_X1 U10683 ( .A(n9873), .ZN(n9676) );
  INV_X1 U10684 ( .A(n9682), .ZN(n9670) );
  OAI211_X1 U10685 ( .C1(n9952), .C2(n9670), .A(n9562), .B(n9669), .ZN(n9872)
         );
  AOI22_X1 U10686 ( .A1(n4932), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9671), .B2(
        n9822), .ZN(n9674) );
  NAND2_X1 U10687 ( .A1(n9672), .A2(n9840), .ZN(n9673) );
  OAI211_X1 U10688 ( .C1(n9872), .C2(n9739), .A(n9674), .B(n9673), .ZN(n9675)
         );
  AOI21_X1 U10689 ( .B1(n9676), .B2(n10235), .A(n9675), .ZN(n9677) );
  OAI21_X1 U10690 ( .B1(n9874), .B2(n9835), .A(n9677), .ZN(P1_U3267) );
  OAI21_X1 U10691 ( .B1(n5560), .B2(n9689), .A(n9678), .ZN(n9681) );
  AOI222_X1 U10692 ( .A1(n10230), .A2(n9681), .B1(n9680), .B2(n10225), .C1(
        n9679), .C2(n10227), .ZN(n9882) );
  OAI211_X1 U10693 ( .C1(n9685), .C2(n9695), .A(n9562), .B(n9682), .ZN(n9881)
         );
  INV_X1 U10694 ( .A(n9881), .ZN(n9687) );
  AOI22_X1 U10695 ( .A1(n4932), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9683), .B2(
        n9822), .ZN(n9684) );
  OAI21_X1 U10696 ( .B1(n9685), .B2(n10237), .A(n9684), .ZN(n9686) );
  AOI21_X1 U10697 ( .B1(n9687), .B2(n9844), .A(n9686), .ZN(n9692) );
  NAND2_X1 U10698 ( .A1(n9690), .A2(n9689), .ZN(n9878) );
  NAND3_X1 U10699 ( .A1(n9688), .A2(n9878), .A3(n9842), .ZN(n9691) );
  OAI211_X1 U10700 ( .C1(n9882), .C2(n4932), .A(n9692), .B(n9691), .ZN(
        P1_U3268) );
  XNOR2_X1 U10701 ( .A(n9693), .B(n9694), .ZN(n9888) );
  AOI211_X1 U10702 ( .C1(n9885), .C2(n9720), .A(n9819), .B(n9695), .ZN(n9884)
         );
  INV_X1 U10703 ( .A(n9885), .ZN(n9699) );
  INV_X1 U10704 ( .A(n9696), .ZN(n9697) );
  AOI22_X1 U10705 ( .A1(n4932), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9697), .B2(
        n9822), .ZN(n9698) );
  OAI21_X1 U10706 ( .B1(n9699), .B2(n10237), .A(n9698), .ZN(n9707) );
  AOI21_X1 U10707 ( .B1(n9701), .B2(n9700), .A(n10716), .ZN(n9705) );
  OAI22_X1 U10708 ( .A1(n9729), .A2(n9770), .B1(n9702), .B2(n10704), .ZN(n9703) );
  AOI21_X1 U10709 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9887) );
  NOR2_X1 U10710 ( .A1(n9887), .A2(n4932), .ZN(n9706) );
  AOI211_X1 U10711 ( .C1(n9884), .C2(n9844), .A(n9707), .B(n9706), .ZN(n9708)
         );
  OAI21_X1 U10712 ( .B1(n9888), .B2(n9835), .A(n9708), .ZN(P1_U3269) );
  INV_X1 U10713 ( .A(n9715), .ZN(n9710) );
  OAI21_X1 U10714 ( .B1(n4977), .B2(n9710), .A(n9709), .ZN(n9892) );
  NAND2_X1 U10715 ( .A1(n9892), .A2(n9842), .ZN(n9725) );
  INV_X1 U10716 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9712) );
  OAI22_X1 U10717 ( .A1(n10712), .A2(n9712), .B1(n9711), .B2(n10709), .ZN(
        n9713) );
  AOI21_X1 U10718 ( .B1(n9889), .B2(n9840), .A(n9713), .ZN(n9724) );
  XOR2_X1 U10719 ( .A(n9714), .B(n9715), .Z(n9716) );
  OAI222_X1 U10720 ( .A1(n10704), .A2(n9718), .B1(n9770), .B2(n9717), .C1(
        n9716), .C2(n10716), .ZN(n9890) );
  NAND2_X1 U10721 ( .A1(n9890), .A2(n10235), .ZN(n9723) );
  AOI21_X1 U10722 ( .B1(n9889), .B2(n9733), .A(n9819), .ZN(n9721) );
  NAND2_X1 U10723 ( .A1(n9891), .A2(n9844), .ZN(n9722) );
  NAND4_X1 U10724 ( .A1(n9725), .A2(n9724), .A3(n9723), .A4(n9722), .ZN(
        P1_U3270) );
  XNOR2_X1 U10725 ( .A(n5031), .B(n9728), .ZN(n9897) );
  XNOR2_X1 U10726 ( .A(n9728), .B(n9727), .ZN(n9731) );
  OAI22_X1 U10727 ( .A1(n9771), .A2(n9770), .B1(n9729), .B2(n10704), .ZN(n9730) );
  AOI21_X1 U10728 ( .B1(n9731), .B2(n10230), .A(n9730), .ZN(n9896) );
  INV_X1 U10729 ( .A(n9896), .ZN(n9741) );
  INV_X1 U10730 ( .A(n9732), .ZN(n9752) );
  OAI211_X1 U10731 ( .C1(n9961), .C2(n9752), .A(n9562), .B(n9733), .ZN(n9895)
         );
  INV_X1 U10732 ( .A(n9734), .ZN(n9735) );
  AOI22_X1 U10733 ( .A1(n4932), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9735), .B2(
        n9822), .ZN(n9738) );
  NAND2_X1 U10734 ( .A1(n9736), .A2(n9840), .ZN(n9737) );
  OAI211_X1 U10735 ( .C1(n9895), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9740)
         );
  AOI21_X1 U10736 ( .B1(n9741), .B2(n10235), .A(n9740), .ZN(n9742) );
  OAI21_X1 U10737 ( .B1(n9897), .B2(n9835), .A(n9742), .ZN(P1_U3271) );
  NAND2_X1 U10738 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  XNOR2_X1 U10739 ( .A(n9745), .B(n9751), .ZN(n9746) );
  OR2_X1 U10740 ( .A1(n9746), .A2(n10716), .ZN(n9749) );
  AOI22_X1 U10741 ( .A1(n9782), .A2(n10227), .B1(n10225), .B2(n9747), .ZN(
        n9748) );
  NAND2_X1 U10742 ( .A1(n9749), .A2(n9748), .ZN(n9901) );
  INV_X1 U10743 ( .A(n9901), .ZN(n9761) );
  XNOR2_X1 U10744 ( .A(n9750), .B(n9751), .ZN(n9903) );
  NAND2_X1 U10745 ( .A1(n9903), .A2(n9842), .ZN(n9760) );
  INV_X1 U10746 ( .A(n9774), .ZN(n9753) );
  AOI211_X1 U10747 ( .C1(n9754), .C2(n9753), .A(n9819), .B(n9752), .ZN(n9902)
         );
  INV_X1 U10748 ( .A(n9755), .ZN(n9756) );
  AOI22_X1 U10749 ( .A1(n4932), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9756), .B2(
        n9822), .ZN(n9757) );
  OAI21_X1 U10750 ( .B1(n9965), .B2(n10237), .A(n9757), .ZN(n9758) );
  AOI21_X1 U10751 ( .B1(n9902), .B2(n9844), .A(n9758), .ZN(n9759) );
  OAI211_X1 U10752 ( .C1(n4932), .C2(n9761), .A(n9760), .B(n9759), .ZN(
        P1_U3272) );
  OAI21_X1 U10753 ( .B1(n5545), .B2(n9581), .A(n9762), .ZN(n9909) );
  NAND2_X1 U10754 ( .A1(n9909), .A2(n9842), .ZN(n9778) );
  INV_X1 U10755 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9764) );
  OAI22_X1 U10756 ( .A1(n10712), .A2(n9764), .B1(n9763), .B2(n10709), .ZN(
        n9765) );
  AOI21_X1 U10757 ( .B1(n9906), .B2(n9840), .A(n9765), .ZN(n9777) );
  XOR2_X1 U10758 ( .A(n9767), .B(n9766), .Z(n9768) );
  OAI222_X1 U10759 ( .A1(n10704), .A2(n9771), .B1(n9770), .B2(n9769), .C1(
        n9768), .C2(n10716), .ZN(n9907) );
  NAND2_X1 U10760 ( .A1(n9907), .A2(n10235), .ZN(n9776) );
  NAND2_X1 U10761 ( .A1(n9906), .A2(n9789), .ZN(n9772) );
  NAND2_X1 U10762 ( .A1(n9772), .A2(n9562), .ZN(n9773) );
  NOR2_X1 U10763 ( .A1(n9774), .A2(n9773), .ZN(n9908) );
  NAND2_X1 U10764 ( .A1(n9908), .A2(n9844), .ZN(n9775) );
  NAND4_X1 U10765 ( .A1(n9778), .A2(n9777), .A3(n9776), .A4(n9775), .ZN(
        P1_U3273) );
  OAI21_X1 U10766 ( .B1(n9787), .B2(n9780), .A(n9779), .ZN(n9783) );
  AOI222_X1 U10767 ( .A1(n10230), .A2(n9783), .B1(n9782), .B2(n10225), .C1(
        n9781), .C2(n10227), .ZN(n9912) );
  INV_X1 U10768 ( .A(n9784), .ZN(n9785) );
  AOI21_X1 U10769 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9915) );
  NAND2_X1 U10770 ( .A1(n9915), .A2(n9842), .ZN(n9796) );
  INV_X1 U10771 ( .A(n9788), .ZN(n9798) );
  INV_X1 U10772 ( .A(n9789), .ZN(n9790) );
  AOI211_X1 U10773 ( .C1(n9791), .C2(n9798), .A(n9819), .B(n9790), .ZN(n9914)
         );
  AOI22_X1 U10774 ( .A1(n4932), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9792), .B2(
        n9822), .ZN(n9793) );
  OAI21_X1 U10775 ( .B1(n9558), .B2(n10237), .A(n9793), .ZN(n9794) );
  AOI21_X1 U10776 ( .B1(n9914), .B2(n9844), .A(n9794), .ZN(n9795) );
  OAI211_X1 U10777 ( .C1(n4932), .C2(n9912), .A(n9796), .B(n9795), .ZN(
        P1_U3274) );
  XOR2_X1 U10778 ( .A(n9797), .B(n9804), .Z(n9922) );
  AOI211_X1 U10779 ( .C1(n9919), .C2(n9799), .A(n9819), .B(n9788), .ZN(n9918)
         );
  INV_X1 U10780 ( .A(n9800), .ZN(n9801) );
  AOI22_X1 U10781 ( .A1(n4932), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9801), .B2(
        n9822), .ZN(n9802) );
  OAI21_X1 U10782 ( .B1(n9803), .B2(n10237), .A(n9802), .ZN(n9812) );
  NAND3_X1 U10783 ( .A1(n5242), .A2(n9806), .A3(n9805), .ZN(n9808) );
  NAND2_X1 U10784 ( .A1(n9808), .A2(n9807), .ZN(n9810) );
  AOI222_X1 U10785 ( .A1(n10230), .A2(n9810), .B1(n9809), .B2(n10225), .C1(
        n9830), .C2(n10227), .ZN(n9921) );
  NOR2_X1 U10786 ( .A1(n9921), .A2(n4932), .ZN(n9811) );
  AOI211_X1 U10787 ( .C1(n9918), .C2(n9844), .A(n9812), .B(n9811), .ZN(n9813)
         );
  OAI21_X1 U10788 ( .B1(n9835), .B2(n9922), .A(n9813), .ZN(P1_U3275) );
  XNOR2_X1 U10789 ( .A(n9814), .B(n9815), .ZN(n9934) );
  INV_X1 U10790 ( .A(n9816), .ZN(n9820) );
  INV_X1 U10791 ( .A(n9817), .ZN(n9818) );
  AOI211_X1 U10792 ( .C1(n9930), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9929)
         );
  INV_X1 U10793 ( .A(n9821), .ZN(n9823) );
  AOI22_X1 U10794 ( .A1(n4932), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9823), .B2(
        n9822), .ZN(n9824) );
  OAI21_X1 U10795 ( .B1(n9825), .B2(n10237), .A(n9824), .ZN(n9833) );
  OAI21_X1 U10796 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9831) );
  AOI222_X1 U10797 ( .A1(n10230), .A2(n9831), .B1(n9830), .B2(n10225), .C1(
        n9829), .C2(n10227), .ZN(n9933) );
  NOR2_X1 U10798 ( .A1(n9933), .A2(n4932), .ZN(n9832) );
  AOI211_X1 U10799 ( .C1(n9929), .C2(n9844), .A(n9833), .B(n9832), .ZN(n9834)
         );
  OAI21_X1 U10800 ( .B1(n9835), .B2(n9934), .A(n9834), .ZN(P1_U3277) );
  NAND2_X1 U10801 ( .A1(n9836), .A2(n10235), .ZN(n9849) );
  OAI22_X1 U10802 ( .A1(n10712), .A2(n9838), .B1(n9837), .B2(n10709), .ZN(
        n9839) );
  AOI21_X1 U10803 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9848) );
  NAND2_X1 U10804 ( .A1(n9843), .A2(n9842), .ZN(n9847) );
  NAND2_X1 U10805 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  NAND4_X1 U10806 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(
        P1_U3286) );
  MUX2_X1 U10807 ( .A(n9851), .B(n9935), .S(n10819), .Z(n9852) );
  OAI21_X1 U10808 ( .B1(n9561), .B2(n9928), .A(n9852), .ZN(P1_U3553) );
  AND2_X1 U10809 ( .A1(n9854), .A2(n9853), .ZN(n9937) );
  MUX2_X1 U10810 ( .A(n9855), .B(n9937), .S(n10819), .Z(n9856) );
  OAI21_X1 U10811 ( .B1(n9940), .B2(n9928), .A(n9856), .ZN(P1_U3552) );
  INV_X1 U10812 ( .A(n9560), .ZN(n9860) );
  INV_X1 U10813 ( .A(n9857), .ZN(n9859) );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9941), .S(n10819), .Z(
        P1_U3551) );
  MUX2_X1 U10815 ( .A(n9865), .B(n9942), .S(n10819), .Z(n9866) );
  OAI21_X1 U10816 ( .B1(n9944), .B2(n9928), .A(n9866), .ZN(P1_U3550) );
  AOI211_X1 U10817 ( .C1(n9869), .C2(n10806), .A(n9868), .B(n9867), .ZN(n9945)
         );
  MUX2_X1 U10818 ( .A(n9870), .B(n9945), .S(n10819), .Z(n9871) );
  OAI21_X1 U10819 ( .B1(n9948), .B2(n9928), .A(n9871), .ZN(P1_U3549) );
  OAI211_X1 U10820 ( .C1(n9874), .C2(n10810), .A(n9873), .B(n9872), .ZN(n9875)
         );
  INV_X1 U10821 ( .A(n9875), .ZN(n9949) );
  MUX2_X1 U10822 ( .A(n9949), .B(n9876), .S(n10818), .Z(n9877) );
  OAI21_X1 U10823 ( .B1(n9952), .B2(n9928), .A(n9877), .ZN(P1_U3548) );
  NAND3_X1 U10824 ( .A1(n9688), .A2(n10806), .A3(n9878), .ZN(n9883) );
  NAND2_X1 U10825 ( .A1(n9879), .A2(n9931), .ZN(n9880) );
  NAND4_X1 U10826 ( .A1(n9883), .A2(n9882), .A3(n9881), .A4(n9880), .ZN(n9953)
         );
  MUX2_X1 U10827 ( .A(n9953), .B(P1_REG1_REG_25__SCAN_IN), .S(n10818), .Z(
        P1_U3547) );
  AOI21_X1 U10828 ( .B1(n9931), .B2(n9885), .A(n9884), .ZN(n9886) );
  OAI211_X1 U10829 ( .C1(n9888), .C2(n10810), .A(n9887), .B(n9886), .ZN(n9954)
         );
  MUX2_X1 U10830 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9954), .S(n10819), .Z(
        P1_U3546) );
  AOI211_X1 U10831 ( .C1(n9892), .C2(n10806), .A(n9891), .B(n9890), .ZN(n9955)
         );
  MUX2_X1 U10832 ( .A(n9893), .B(n9955), .S(n10819), .Z(n9894) );
  OAI21_X1 U10833 ( .B1(n9559), .B2(n9928), .A(n9894), .ZN(P1_U3545) );
  OAI211_X1 U10834 ( .C1(n9897), .C2(n10810), .A(n9896), .B(n9895), .ZN(n9898)
         );
  INV_X1 U10835 ( .A(n9898), .ZN(n9958) );
  MUX2_X1 U10836 ( .A(n9899), .B(n9958), .S(n10819), .Z(n9900) );
  OAI21_X1 U10837 ( .B1(n9961), .B2(n9928), .A(n9900), .ZN(P1_U3544) );
  AOI211_X1 U10838 ( .C1(n9903), .C2(n10806), .A(n9902), .B(n9901), .ZN(n9962)
         );
  MUX2_X1 U10839 ( .A(n9904), .B(n9962), .S(n10819), .Z(n9905) );
  OAI21_X1 U10840 ( .B1(n9965), .B2(n9928), .A(n9905), .ZN(P1_U3543) );
  INV_X1 U10841 ( .A(n9906), .ZN(n9969) );
  AOI211_X1 U10842 ( .C1(n10806), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9966)
         );
  MUX2_X1 U10843 ( .A(n9910), .B(n9966), .S(n10819), .Z(n9911) );
  OAI21_X1 U10844 ( .B1(n9969), .B2(n9928), .A(n9911), .ZN(P1_U3542) );
  INV_X1 U10845 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9916) );
  INV_X1 U10846 ( .A(n9912), .ZN(n9913) );
  AOI211_X1 U10847 ( .C1(n9915), .C2(n10806), .A(n9914), .B(n9913), .ZN(n9970)
         );
  MUX2_X1 U10848 ( .A(n9916), .B(n9970), .S(n10819), .Z(n9917) );
  OAI21_X1 U10849 ( .B1(n9558), .B2(n9928), .A(n9917), .ZN(P1_U3541) );
  AOI21_X1 U10850 ( .B1(n9931), .B2(n9919), .A(n9918), .ZN(n9920) );
  OAI211_X1 U10851 ( .C1(n9922), .C2(n10810), .A(n9921), .B(n9920), .ZN(n9973)
         );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9973), .S(n10819), .Z(
        P1_U3540) );
  AOI211_X1 U10853 ( .C1(n10806), .C2(n9925), .A(n9924), .B(n9923), .ZN(n9974)
         );
  MUX2_X1 U10854 ( .A(n9926), .B(n9974), .S(n10819), .Z(n9927) );
  OAI21_X1 U10855 ( .B1(n9978), .B2(n9928), .A(n9927), .ZN(P1_U3539) );
  AOI21_X1 U10856 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9932) );
  OAI211_X1 U10857 ( .C1(n9934), .C2(n10810), .A(n9933), .B(n9932), .ZN(n9979)
         );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9979), .S(n10819), .Z(
        P1_U3538) );
  MUX2_X1 U10859 ( .A(n9938), .B(n9937), .S(n10823), .Z(n9939) );
  OAI21_X1 U10860 ( .B1(n9940), .B2(n9977), .A(n9939), .ZN(P1_U3520) );
  MUX2_X1 U10861 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9941), .S(n10823), .Z(
        P1_U3519) );
  MUX2_X1 U10862 ( .A(n9946), .B(n9945), .S(n10823), .Z(n9947) );
  OAI21_X1 U10863 ( .B1(n9948), .B2(n9977), .A(n9947), .ZN(P1_U3517) );
  MUX2_X1 U10864 ( .A(n9950), .B(n9949), .S(n10823), .Z(n9951) );
  OAI21_X1 U10865 ( .B1(n9952), .B2(n9977), .A(n9951), .ZN(P1_U3516) );
  MUX2_X1 U10866 ( .A(n9953), .B(P1_REG0_REG_25__SCAN_IN), .S(n10820), .Z(
        P1_U3515) );
  MUX2_X1 U10867 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9954), .S(n10823), .Z(
        P1_U3514) );
  MUX2_X1 U10868 ( .A(n9956), .B(n9955), .S(n10823), .Z(n9957) );
  OAI21_X1 U10869 ( .B1(n9559), .B2(n9977), .A(n9957), .ZN(P1_U3513) );
  MUX2_X1 U10870 ( .A(n9959), .B(n9958), .S(n10823), .Z(n9960) );
  OAI21_X1 U10871 ( .B1(n9961), .B2(n9977), .A(n9960), .ZN(P1_U3512) );
  MUX2_X1 U10872 ( .A(n9963), .B(n9962), .S(n10823), .Z(n9964) );
  OAI21_X1 U10873 ( .B1(n9965), .B2(n9977), .A(n9964), .ZN(P1_U3511) );
  MUX2_X1 U10874 ( .A(n9967), .B(n9966), .S(n10823), .Z(n9968) );
  OAI21_X1 U10875 ( .B1(n9969), .B2(n9977), .A(n9968), .ZN(P1_U3510) );
  INV_X1 U10876 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9971) );
  MUX2_X1 U10877 ( .A(n9971), .B(n9970), .S(n10823), .Z(n9972) );
  OAI21_X1 U10878 ( .B1(n9558), .B2(n9977), .A(n9972), .ZN(P1_U3509) );
  MUX2_X1 U10879 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9973), .S(n10823), .Z(
        P1_U3507) );
  INV_X1 U10880 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9975) );
  MUX2_X1 U10881 ( .A(n9975), .B(n9974), .S(n10823), .Z(n9976) );
  OAI21_X1 U10882 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(P1_U3504) );
  MUX2_X1 U10883 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9979), .S(n10823), .Z(
        P1_U3501) );
  INV_X1 U10884 ( .A(n9983), .ZN(n9981) );
  MUX2_X1 U10885 ( .A(n9982), .B(P1_D_REG_1__SCAN_IN), .S(n10003), .Z(P1_U3440) );
  MUX2_X1 U10886 ( .A(n9984), .B(P1_D_REG_0__SCAN_IN), .S(n9983), .Z(P1_U3439)
         );
  NOR4_X1 U10887 ( .A1(n9987), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9985), .ZN(n9988) );
  AOI21_X1 U10888 ( .B1(n9997), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9988), .ZN(
        n9989) );
  OAI21_X1 U10889 ( .B1(n9990), .B2(n8027), .A(n9989), .ZN(P1_U3324) );
  AOI22_X1 U10890 ( .A1(n9991), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9997), .ZN(n9992) );
  OAI21_X1 U10891 ( .B1(n9993), .B2(n10000), .A(n9992), .ZN(P1_U3325) );
  AOI22_X1 U10892 ( .A1(n5034), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9997), .ZN(n9994) );
  OAI21_X1 U10893 ( .B1(n9995), .B2(n10000), .A(n9994), .ZN(P1_U3326) );
  INV_X1 U10894 ( .A(n9996), .ZN(n10001) );
  AOI22_X1 U10895 ( .A1(n9998), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9997), .ZN(n9999) );
  OAI21_X1 U10896 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(P1_U3327) );
  MUX2_X1 U10897 ( .A(n10002), .B(n10302), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  AND2_X1 U10898 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10003), .ZN(P1_U3323) );
  AND2_X1 U10899 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10003), .ZN(P1_U3322) );
  AND2_X1 U10900 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10003), .ZN(P1_U3321) );
  AND2_X1 U10901 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10003), .ZN(P1_U3320) );
  AND2_X1 U10902 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10003), .ZN(P1_U3319) );
  AND2_X1 U10903 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10003), .ZN(P1_U3318) );
  AND2_X1 U10904 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10003), .ZN(P1_U3317) );
  AND2_X1 U10905 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10003), .ZN(P1_U3316) );
  AND2_X1 U10906 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10003), .ZN(P1_U3315) );
  AND2_X1 U10907 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10003), .ZN(P1_U3314) );
  AND2_X1 U10908 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10003), .ZN(P1_U3313) );
  AND2_X1 U10909 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10003), .ZN(P1_U3312) );
  AND2_X1 U10910 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10003), .ZN(P1_U3311) );
  AND2_X1 U10911 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10003), .ZN(P1_U3310) );
  AND2_X1 U10912 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10003), .ZN(P1_U3309) );
  AND2_X1 U10913 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10003), .ZN(P1_U3308) );
  AND2_X1 U10914 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10003), .ZN(P1_U3307) );
  AND2_X1 U10915 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10003), .ZN(P1_U3306) );
  AND2_X1 U10916 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10003), .ZN(P1_U3305) );
  AND2_X1 U10917 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10003), .ZN(P1_U3304) );
  AND2_X1 U10918 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10003), .ZN(P1_U3303) );
  AND2_X1 U10919 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10003), .ZN(P1_U3302) );
  AND2_X1 U10920 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10003), .ZN(P1_U3301) );
  AND2_X1 U10921 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10003), .ZN(P1_U3300) );
  AND2_X1 U10922 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10003), .ZN(P1_U3299) );
  AND2_X1 U10923 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10003), .ZN(P1_U3298) );
  AND2_X1 U10924 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10003), .ZN(P1_U3297) );
  AND2_X1 U10925 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10003), .ZN(P1_U3296) );
  AND2_X1 U10926 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10003), .ZN(P1_U3295) );
  AND2_X1 U10927 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10003), .ZN(P1_U3294) );
  INV_X1 U10928 ( .A(keyinput_114), .ZN(n10083) );
  OAI22_X1 U10929 ( .A1(n5783), .A2(keyinput_113), .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .ZN(n10004) );
  AOI221_X1 U10930 ( .B1(n5783), .B2(keyinput_113), .C1(keyinput_111), .C2(
        P2_REG3_REG_25__SCAN_IN), .A(n10004), .ZN(n10079) );
  INV_X1 U10931 ( .A(keyinput_107), .ZN(n10073) );
  INV_X1 U10932 ( .A(keyinput_106), .ZN(n10071) );
  OAI22_X1 U10933 ( .A1(n10179), .A2(keyinput_105), .B1(keyinput_103), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n10005) );
  AOI221_X1 U10934 ( .B1(n10179), .B2(keyinput_105), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_103), .A(n10005), .ZN(n10068)
         );
  OAI22_X1 U10935 ( .A1(n10007), .A2(keyinput_100), .B1(n10110), .B2(
        keyinput_101), .ZN(n10006) );
  AOI221_X1 U10936 ( .B1(n10007), .B2(keyinput_100), .C1(keyinput_101), .C2(
        n10110), .A(n10006), .ZN(n10064) );
  INV_X1 U10937 ( .A(keyinput_96), .ZN(n10058) );
  INV_X1 U10938 ( .A(SI_0_), .ZN(n10170) );
  OAI22_X1 U10939 ( .A1(n10114), .A2(keyinput_83), .B1(keyinput_82), .B2(
        SI_14_), .ZN(n10008) );
  AOI221_X1 U10940 ( .B1(n10114), .B2(keyinput_83), .C1(SI_14_), .C2(
        keyinput_82), .A(n10008), .ZN(n10037) );
  INV_X1 U10941 ( .A(keyinput_80), .ZN(n10035) );
  INV_X1 U10942 ( .A(SI_21_), .ZN(n10010) );
  OAI22_X1 U10943 ( .A1(n10010), .A2(keyinput_75), .B1(n10116), .B2(
        keyinput_76), .ZN(n10009) );
  AOI221_X1 U10944 ( .B1(n10010), .B2(keyinput_75), .C1(keyinput_76), .C2(
        n10116), .A(n10009), .ZN(n10027) );
  INV_X1 U10945 ( .A(SI_25_), .ZN(n10118) );
  AOI22_X1 U10946 ( .A1(n10118), .A2(keyinput_71), .B1(keyinput_72), .B2(
        n10012), .ZN(n10011) );
  OAI221_X1 U10947 ( .B1(n10118), .B2(keyinput_71), .C1(n10012), .C2(
        keyinput_72), .A(n10011), .ZN(n10025) );
  INV_X1 U10948 ( .A(SI_26_), .ZN(n10127) );
  INV_X1 U10949 ( .A(keyinput_70), .ZN(n10022) );
  OAI22_X1 U10950 ( .A1(n10014), .A2(keyinput_66), .B1(SI_29_), .B2(
        keyinput_67), .ZN(n10013) );
  AOI221_X1 U10951 ( .B1(n10014), .B2(keyinput_66), .C1(keyinput_67), .C2(
        SI_29_), .A(n10013), .ZN(n10020) );
  AOI22_X1 U10952 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n10015) );
  OAI221_X1 U10953 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n10015), .ZN(n10019) );
  AOI22_X1 U10954 ( .A1(n10017), .A2(keyinput_68), .B1(n10122), .B2(
        keyinput_69), .ZN(n10016) );
  OAI221_X1 U10955 ( .B1(n10017), .B2(keyinput_68), .C1(n10122), .C2(
        keyinput_69), .A(n10016), .ZN(n10018) );
  AOI21_X1 U10956 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10021) );
  AOI221_X1 U10957 ( .B1(SI_26_), .B2(keyinput_70), .C1(n10127), .C2(n10022), 
        .A(n10021), .ZN(n10024) );
  NAND2_X1 U10958 ( .A1(SI_23_), .A2(keyinput_73), .ZN(n10023) );
  OAI221_X1 U10959 ( .B1(n10025), .B2(n10024), .C1(SI_23_), .C2(keyinput_73), 
        .A(n10023), .ZN(n10026) );
  OAI211_X1 U10960 ( .C1(SI_22_), .C2(keyinput_74), .A(n10027), .B(n10026), 
        .ZN(n10028) );
  AOI21_X1 U10961 ( .B1(SI_22_), .B2(keyinput_74), .A(n10028), .ZN(n10032) );
  AOI22_X1 U10962 ( .A1(SI_18_), .A2(keyinput_78), .B1(n10030), .B2(
        keyinput_77), .ZN(n10029) );
  OAI221_X1 U10963 ( .B1(SI_18_), .B2(keyinput_78), .C1(n10030), .C2(
        keyinput_77), .A(n10029), .ZN(n10031) );
  AOI211_X1 U10964 ( .C1(n10137), .C2(keyinput_79), .A(n10032), .B(n10031), 
        .ZN(n10033) );
  OAI21_X1 U10965 ( .B1(n10137), .B2(keyinput_79), .A(n10033), .ZN(n10034) );
  OAI221_X1 U10966 ( .B1(SI_16_), .B2(n10035), .C1(n10143), .C2(keyinput_80), 
        .A(n10034), .ZN(n10036) );
  OAI211_X1 U10967 ( .C1(SI_15_), .C2(keyinput_81), .A(n10037), .B(n10036), 
        .ZN(n10038) );
  AOI21_X1 U10968 ( .B1(SI_15_), .B2(keyinput_81), .A(n10038), .ZN(n10051) );
  INV_X1 U10969 ( .A(SI_12_), .ZN(n10150) );
  XOR2_X1 U10970 ( .A(n10150), .B(keyinput_84), .Z(n10050) );
  OAI22_X1 U10971 ( .A1(n10040), .A2(keyinput_88), .B1(keyinput_85), .B2(
        SI_11_), .ZN(n10039) );
  AOI221_X1 U10972 ( .B1(n10040), .B2(keyinput_88), .C1(SI_11_), .C2(
        keyinput_85), .A(n10039), .ZN(n10049) );
  OAI22_X1 U10973 ( .A1(SI_7_), .A2(keyinput_89), .B1(keyinput_91), .B2(SI_5_), 
        .ZN(n10041) );
  AOI221_X1 U10974 ( .B1(SI_7_), .B2(keyinput_89), .C1(SI_5_), .C2(keyinput_91), .A(n10041), .ZN(n10045) );
  INV_X1 U10975 ( .A(SI_6_), .ZN(n10152) );
  OAI22_X1 U10976 ( .A1(n10043), .A2(keyinput_86), .B1(n10152), .B2(
        keyinput_90), .ZN(n10042) );
  AOI221_X1 U10977 ( .B1(n10043), .B2(keyinput_86), .C1(keyinput_90), .C2(
        n10152), .A(n10042), .ZN(n10044) );
  OAI211_X1 U10978 ( .C1(n10047), .C2(keyinput_87), .A(n10045), .B(n10044), 
        .ZN(n10046) );
  AOI21_X1 U10979 ( .B1(n10047), .B2(keyinput_87), .A(n10046), .ZN(n10048) );
  OAI211_X1 U10980 ( .C1(n10051), .C2(n10050), .A(n10049), .B(n10048), .ZN(
        n10056) );
  OAI22_X1 U10981 ( .A1(SI_4_), .A2(keyinput_92), .B1(SI_3_), .B2(keyinput_93), 
        .ZN(n10052) );
  AOI221_X1 U10982 ( .B1(SI_4_), .B2(keyinput_92), .C1(keyinput_93), .C2(SI_3_), .A(n10052), .ZN(n10055) );
  XNOR2_X1 U10983 ( .A(n10164), .B(keyinput_95), .ZN(n10054) );
  XNOR2_X1 U10984 ( .A(SI_2_), .B(keyinput_94), .ZN(n10053) );
  AOI211_X1 U10985 ( .C1(n10056), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10057) );
  AOI221_X1 U10986 ( .B1(SI_0_), .B2(n10058), .C1(n10170), .C2(keyinput_96), 
        .A(n10057), .ZN(n10061) );
  AOI22_X1 U10987 ( .A1(n5060), .A2(keyinput_97), .B1(keyinput_98), .B2(
        P2_U3151), .ZN(n10059) );
  OAI221_X1 U10988 ( .B1(n5060), .B2(keyinput_97), .C1(P2_U3151), .C2(
        keyinput_98), .A(n10059), .ZN(n10060) );
  AOI211_X1 U10989 ( .C1(P2_REG3_REG_7__SCAN_IN), .C2(keyinput_99), .A(n10061), 
        .B(n10060), .ZN(n10062) );
  OAI21_X1 U10990 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .A(n10062), 
        .ZN(n10063) );
  AOI22_X1 U10991 ( .A1(keyinput_102), .A2(n10066), .B1(n10064), .B2(n10063), 
        .ZN(n10065) );
  OAI21_X1 U10992 ( .B1(n10066), .B2(keyinput_102), .A(n10065), .ZN(n10067) );
  OAI211_X1 U10993 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(keyinput_104), .A(n10068), .B(n10067), .ZN(n10069) );
  AOI21_X1 U10994 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .A(n10069), 
        .ZN(n10070) );
  AOI221_X1 U10995 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .C1(
        n6092), .C2(n10071), .A(n10070), .ZN(n10072) );
  AOI221_X1 U10996 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n10187), .C2(n10073), .A(n10072), .ZN(n10076) );
  AOI22_X1 U10997 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_108), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .ZN(n10074) );
  OAI221_X1 U10998 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_109), .A(n10074), .ZN(n10075)
         );
  AOI211_X1 U10999 ( .C1(P2_REG3_REG_12__SCAN_IN), .C2(keyinput_110), .A(
        n10076), .B(n10075), .ZN(n10077) );
  OAI21_X1 U11000 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .A(n10077), .ZN(n10078) );
  OAI211_X1 U11001 ( .C1(n10081), .C2(keyinput_112), .A(n10079), .B(n10078), 
        .ZN(n10080) );
  AOI21_X1 U11002 ( .B1(n10081), .B2(keyinput_112), .A(n10080), .ZN(n10082) );
  AOI221_X1 U11003 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n10083), .C1(n5965), 
        .C2(keyinput_114), .A(n10082), .ZN(n10087) );
  AOI22_X1 U11004 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_117), .B1(n10085), .B2(keyinput_115), .ZN(n10084) );
  OAI221_X1 U11005 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .C1(
        n10085), .C2(keyinput_115), .A(n10084), .ZN(n10086) );
  AOI211_X1 U11006 ( .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_116), .A(n10087), .B(n10086), .ZN(n10088) );
  OAI21_X1 U11007 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .A(n10088), 
        .ZN(n10092) );
  XOR2_X1 U11008 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_118), .Z(n10090) );
  XNOR2_X1 U11009 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_119), .ZN(n10089)
         );
  NOR2_X1 U11010 ( .A1(n10090), .A2(n10089), .ZN(n10091) );
  AOI22_X1 U11011 ( .A1(n10092), .A2(n10091), .B1(keyinput_121), .B2(n10206), 
        .ZN(n10093) );
  OAI21_X1 U11012 ( .B1(keyinput_121), .B2(n10206), .A(n10093), .ZN(n10101) );
  INV_X1 U11013 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11014 ( .A1(n10208), .A2(keyinput_122), .B1(n5918), .B2(
        keyinput_120), .ZN(n10094) );
  OAI221_X1 U11015 ( .B1(n10208), .B2(keyinput_122), .C1(n5918), .C2(
        keyinput_120), .A(n10094), .ZN(n10100) );
  OAI22_X1 U11016 ( .A1(n10096), .A2(keyinput_124), .B1(n10211), .B2(
        keyinput_123), .ZN(n10095) );
  AOI221_X1 U11017 ( .B1(n10096), .B2(keyinput_124), .C1(keyinput_123), .C2(
        n10211), .A(n10095), .ZN(n10099) );
  OAI22_X1 U11018 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_126), .B1(
        keyinput_125), .B2(P2_REG3_REG_6__SCAN_IN), .ZN(n10097) );
  AOI221_X1 U11019 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_125), .A(n10097), .ZN(n10098) );
  OAI211_X1 U11020 ( .C1(n10101), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10103) );
  AOI21_X1 U11021 ( .B1(keyinput_127), .B2(n10103), .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10105) );
  INV_X1 U11022 ( .A(keyinput_127), .ZN(n10102) );
  AOI21_X1 U11023 ( .B1(n10103), .B2(n10102), .A(keyinput_63), .ZN(n10104) );
  AOI22_X1 U11024 ( .A1(keyinput_63), .A2(n10105), .B1(P2_REG3_REG_15__SCAN_IN), .B2(n10104), .ZN(n10218) );
  OAI22_X1 U11025 ( .A1(n5837), .A2(keyinput_53), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(keyinput_51), .ZN(n10106) );
  AOI221_X1 U11026 ( .B1(n5837), .B2(keyinput_53), .C1(keyinput_51), .C2(
        P2_REG3_REG_24__SCAN_IN), .A(n10106), .ZN(n10199) );
  INV_X1 U11027 ( .A(keyinput_50), .ZN(n10197) );
  INV_X1 U11028 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10108) );
  OAI22_X1 U11029 ( .A1(n10108), .A2(keyinput_46), .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .ZN(n10107) );
  AOI221_X1 U11030 ( .B1(n10108), .B2(keyinput_46), .C1(keyinput_45), .C2(
        P2_REG3_REG_21__SCAN_IN), .A(n10107), .ZN(n10189) );
  INV_X1 U11031 ( .A(keyinput_43), .ZN(n10186) );
  INV_X1 U11032 ( .A(keyinput_42), .ZN(n10184) );
  AOI22_X1 U11033 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .B1(n10110), .B2(keyinput_37), .ZN(n10109) );
  OAI221_X1 U11034 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        n10110), .C2(keyinput_37), .A(n10109), .ZN(n10175) );
  INV_X1 U11035 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10112) );
  OAI22_X1 U11036 ( .A1(n10112), .A2(keyinput_35), .B1(keyinput_33), .B2(
        P2_RD_REG_SCAN_IN), .ZN(n10111) );
  AOI221_X1 U11037 ( .B1(n10112), .B2(keyinput_35), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_33), .A(n10111), .ZN(n10172) );
  INV_X1 U11038 ( .A(keyinput_20), .ZN(n10149) );
  OAI22_X1 U11039 ( .A1(n10114), .A2(keyinput_19), .B1(SI_14_), .B2(
        keyinput_18), .ZN(n10113) );
  AOI221_X1 U11040 ( .B1(n10114), .B2(keyinput_19), .C1(keyinput_18), .C2(
        SI_14_), .A(n10113), .ZN(n10145) );
  INV_X1 U11041 ( .A(keyinput_16), .ZN(n10142) );
  OAI22_X1 U11042 ( .A1(n10116), .A2(keyinput_12), .B1(SI_21_), .B2(
        keyinput_11), .ZN(n10115) );
  AOI221_X1 U11043 ( .B1(n10116), .B2(keyinput_12), .C1(keyinput_11), .C2(
        SI_21_), .A(n10115), .ZN(n10134) );
  OAI22_X1 U11044 ( .A1(n10118), .A2(keyinput_7), .B1(keyinput_8), .B2(SI_24_), 
        .ZN(n10117) );
  AOI221_X1 U11045 ( .B1(n10118), .B2(keyinput_7), .C1(SI_24_), .C2(keyinput_8), .A(n10117), .ZN(n10130) );
  INV_X1 U11046 ( .A(keyinput_6), .ZN(n10128) );
  OAI22_X1 U11047 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10119) );
  AOI221_X1 U11048 ( .B1(SI_31_), .B2(keyinput_1), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n10119), .ZN(n10125) );
  AOI22_X1 U11049 ( .A1(SI_30_), .A2(keyinput_2), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n10120) );
  OAI221_X1 U11050 ( .B1(SI_30_), .B2(keyinput_2), .C1(SI_29_), .C2(keyinput_3), .A(n10120), .ZN(n10124) );
  OAI22_X1 U11051 ( .A1(n10122), .A2(keyinput_5), .B1(SI_28_), .B2(keyinput_4), 
        .ZN(n10121) );
  AOI221_X1 U11052 ( .B1(n10122), .B2(keyinput_5), .C1(keyinput_4), .C2(SI_28_), .A(n10121), .ZN(n10123) );
  OAI21_X1 U11053 ( .B1(n10125), .B2(n10124), .A(n10123), .ZN(n10126) );
  OAI221_X1 U11054 ( .B1(SI_26_), .B2(n10128), .C1(n10127), .C2(keyinput_6), 
        .A(n10126), .ZN(n10129) );
  AOI22_X1 U11055 ( .A1(keyinput_9), .A2(n10132), .B1(n10130), .B2(n10129), 
        .ZN(n10131) );
  OAI21_X1 U11056 ( .B1(n10132), .B2(keyinput_9), .A(n10131), .ZN(n10133) );
  OAI211_X1 U11057 ( .C1(SI_22_), .C2(keyinput_10), .A(n10134), .B(n10133), 
        .ZN(n10135) );
  AOI21_X1 U11058 ( .B1(SI_22_), .B2(keyinput_10), .A(n10135), .ZN(n10139) );
  AOI22_X1 U11059 ( .A1(SI_19_), .A2(keyinput_13), .B1(n10137), .B2(
        keyinput_15), .ZN(n10136) );
  OAI221_X1 U11060 ( .B1(SI_19_), .B2(keyinput_13), .C1(n10137), .C2(
        keyinput_15), .A(n10136), .ZN(n10138) );
  AOI211_X1 U11061 ( .C1(SI_18_), .C2(keyinput_14), .A(n10139), .B(n10138), 
        .ZN(n10140) );
  OAI21_X1 U11062 ( .B1(SI_18_), .B2(keyinput_14), .A(n10140), .ZN(n10141) );
  OAI221_X1 U11063 ( .B1(SI_16_), .B2(keyinput_16), .C1(n10143), .C2(n10142), 
        .A(n10141), .ZN(n10144) );
  OAI211_X1 U11064 ( .C1(n10147), .C2(keyinput_17), .A(n10145), .B(n10144), 
        .ZN(n10146) );
  AOI21_X1 U11065 ( .B1(n10147), .B2(keyinput_17), .A(n10146), .ZN(n10148) );
  AOI221_X1 U11066 ( .B1(SI_12_), .B2(keyinput_20), .C1(n10150), .C2(n10149), 
        .A(n10148), .ZN(n10163) );
  INV_X1 U11067 ( .A(SI_11_), .ZN(n10153) );
  OAI22_X1 U11068 ( .A1(n10153), .A2(keyinput_21), .B1(n10152), .B2(
        keyinput_26), .ZN(n10151) );
  AOI221_X1 U11069 ( .B1(n10153), .B2(keyinput_21), .C1(keyinput_26), .C2(
        n10152), .A(n10151), .ZN(n10159) );
  OAI22_X1 U11070 ( .A1(SI_8_), .A2(keyinput_24), .B1(keyinput_25), .B2(SI_7_), 
        .ZN(n10154) );
  AOI221_X1 U11071 ( .B1(SI_8_), .B2(keyinput_24), .C1(SI_7_), .C2(keyinput_25), .A(n10154), .ZN(n10158) );
  OAI22_X1 U11072 ( .A1(SI_10_), .A2(keyinput_22), .B1(keyinput_23), .B2(SI_9_), .ZN(n10155) );
  AOI221_X1 U11073 ( .B1(SI_10_), .B2(keyinput_22), .C1(SI_9_), .C2(
        keyinput_23), .A(n10155), .ZN(n10157) );
  XNOR2_X1 U11074 ( .A(SI_5_), .B(keyinput_27), .ZN(n10156) );
  NAND4_X1 U11075 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10162) );
  OAI22_X1 U11076 ( .A1(SI_4_), .A2(keyinput_28), .B1(keyinput_29), .B2(SI_3_), 
        .ZN(n10160) );
  AOI221_X1 U11077 ( .B1(SI_4_), .B2(keyinput_28), .C1(SI_3_), .C2(keyinput_29), .A(n10160), .ZN(n10161) );
  OAI21_X1 U11078 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(n10168) );
  XNOR2_X1 U11079 ( .A(n10164), .B(keyinput_31), .ZN(n10166) );
  XNOR2_X1 U11080 ( .A(SI_2_), .B(keyinput_30), .ZN(n10165) );
  NOR2_X1 U11081 ( .A1(n10166), .A2(n10165), .ZN(n10167) );
  AOI22_X1 U11082 ( .A1(n10168), .A2(n10167), .B1(keyinput_32), .B2(n10170), 
        .ZN(n10169) );
  OAI21_X1 U11083 ( .B1(n10170), .B2(keyinput_32), .A(n10169), .ZN(n10171) );
  OAI211_X1 U11084 ( .C1(P2_STATE_REG_SCAN_IN), .C2(keyinput_34), .A(n10172), 
        .B(n10171), .ZN(n10173) );
  AOI21_X1 U11085 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .A(n10173), 
        .ZN(n10174) );
  OAI22_X1 U11086 ( .A1(n10175), .A2(n10174), .B1(keyinput_38), .B2(
        P2_REG3_REG_23__SCAN_IN), .ZN(n10176) );
  AOI21_X1 U11087 ( .B1(keyinput_38), .B2(P2_REG3_REG_23__SCAN_IN), .A(n10176), 
        .ZN(n10181) );
  AOI22_X1 U11088 ( .A1(n10179), .A2(keyinput_41), .B1(keyinput_40), .B2(
        n10178), .ZN(n10177) );
  OAI221_X1 U11089 ( .B1(n10179), .B2(keyinput_41), .C1(n10178), .C2(
        keyinput_40), .A(n10177), .ZN(n10180) );
  AOI211_X1 U11090 ( .C1(P2_REG3_REG_10__SCAN_IN), .C2(keyinput_39), .A(n10181), .B(n10180), .ZN(n10182) );
  OAI21_X1 U11091 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .A(n10182), 
        .ZN(n10183) );
  OAI221_X1 U11092 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(n10184), .C1(n6092), 
        .C2(keyinput_42), .A(n10183), .ZN(n10185) );
  OAI221_X1 U11093 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(n10187), .C2(n10186), .A(n10185), .ZN(n10188) );
  OAI211_X1 U11094 ( .C1(n7333), .C2(keyinput_44), .A(n10189), .B(n10188), 
        .ZN(n10190) );
  AOI21_X1 U11095 ( .B1(n7333), .B2(keyinput_44), .A(n10190), .ZN(n10194) );
  AOI22_X1 U11096 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(n10192), 
        .B2(keyinput_47), .ZN(n10191) );
  OAI221_X1 U11097 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(n10192), .C2(keyinput_47), .A(n10191), .ZN(n10193) );
  AOI211_X1 U11098 ( .C1(P2_REG3_REG_16__SCAN_IN), .C2(keyinput_48), .A(n10194), .B(n10193), .ZN(n10195) );
  OAI21_X1 U11099 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .A(n10195), 
        .ZN(n10196) );
  OAI221_X1 U11100 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n10197), .C1(n5965), 
        .C2(keyinput_50), .A(n10196), .ZN(n10198) );
  OAI211_X1 U11101 ( .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_52), .A(n10199), 
        .B(n10198), .ZN(n10200) );
  AOI21_X1 U11102 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .A(n10200), 
        .ZN(n10204) );
  XOR2_X1 U11103 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .Z(n10202) );
  XNOR2_X1 U11104 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n10201)
         );
  NAND2_X1 U11105 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  OAI22_X1 U11106 ( .A1(n10204), .A2(n10203), .B1(keyinput_57), .B2(n10206), 
        .ZN(n10205) );
  AOI21_X1 U11107 ( .B1(n10206), .B2(keyinput_57), .A(n10205), .ZN(n10216) );
  OAI22_X1 U11108 ( .A1(n5918), .A2(keyinput_56), .B1(n10208), .B2(keyinput_58), .ZN(n10207) );
  AOI221_X1 U11109 ( .B1(n5918), .B2(keyinput_56), .C1(keyinput_58), .C2(
        n10208), .A(n10207), .ZN(n10215) );
  AOI22_X1 U11110 ( .A1(n10211), .A2(keyinput_59), .B1(n10210), .B2(
        keyinput_61), .ZN(n10209) );
  OAI221_X1 U11111 ( .B1(n10211), .B2(keyinput_59), .C1(n10210), .C2(
        keyinput_61), .A(n10209), .ZN(n10214) );
  AOI22_X1 U11112 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .ZN(n10212) );
  OAI221_X1 U11113 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_62), .A(n10212), .ZN(n10213) );
  AOI211_X1 U11114 ( .C1(n10216), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n10217) );
  NOR2_X1 U11115 ( .A1(n10218), .A2(n10217), .ZN(n10241) );
  XNOR2_X1 U11116 ( .A(n10219), .B(n10223), .ZN(n10732) );
  INV_X1 U11117 ( .A(n10732), .ZN(n10739) );
  OAI211_X1 U11118 ( .C1(n10221), .C2(n10735), .A(n10220), .B(n9562), .ZN(
        n10733) );
  OAI22_X1 U11119 ( .A1(n10733), .A2(n10222), .B1(n6328), .B2(n10709), .ZN(
        n10232) );
  XNOR2_X1 U11120 ( .A(n10224), .B(n10223), .ZN(n10229) );
  AOI222_X1 U11121 ( .A1(n10230), .A2(n10229), .B1(n10228), .B2(n10227), .C1(
        n10226), .C2(n10225), .ZN(n10734) );
  INV_X1 U11122 ( .A(n10734), .ZN(n10231) );
  AOI211_X1 U11123 ( .C1(n10739), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n10234) );
  NOR2_X1 U11124 ( .A1(n10234), .A2(n4932), .ZN(n10239) );
  OAI22_X1 U11125 ( .A1(n10237), .A2(n10735), .B1(n10236), .B2(n10235), .ZN(
        n10238) );
  NOR2_X1 U11126 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  XNOR2_X1 U11127 ( .A(n10241), .B(n10240), .ZN(P1_U3291) );
  OAI21_X1 U11128 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10244), .ZN(n10242) );
  INV_X1 U11129 ( .A(n10242), .ZN(ADD_1068_U46) );
  OAI21_X1 U11130 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(n10246) );
  XNOR2_X1 U11131 ( .A(n10246), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  AOI21_X1 U11132 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(ADD_1068_U54) );
  AOI21_X1 U11133 ( .B1(n10252), .B2(n10251), .A(n10250), .ZN(ADD_1068_U53) );
  OAI21_X1 U11134 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(ADD_1068_U52) );
  OAI21_X1 U11135 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(ADD_1068_U51) );
  OAI21_X1 U11136 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(ADD_1068_U50) );
  OAI21_X1 U11137 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(ADD_1068_U49) );
  OAI21_X1 U11138 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(ADD_1068_U48) );
  OAI21_X1 U11139 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(ADD_1068_U47) );
  OAI21_X1 U11140 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(ADD_1068_U63) );
  OAI21_X1 U11141 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(ADD_1068_U62) );
  OAI21_X1 U11142 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(ADD_1068_U61) );
  OAI21_X1 U11143 ( .B1(n10282), .B2(n10281), .A(n10280), .ZN(ADD_1068_U60) );
  OAI21_X1 U11144 ( .B1(n10285), .B2(n10284), .A(n10283), .ZN(ADD_1068_U59) );
  OAI21_X1 U11145 ( .B1(n10288), .B2(n10287), .A(n10286), .ZN(ADD_1068_U58) );
  OAI21_X1 U11146 ( .B1(n10291), .B2(n10290), .A(n10289), .ZN(ADD_1068_U57) );
  OAI21_X1 U11147 ( .B1(n10294), .B2(n10293), .A(n10292), .ZN(ADD_1068_U56) );
  OAI21_X1 U11148 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(ADD_1068_U55) );
  AOI22_X1 U11149 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n10300), .B1(n10299), 
        .B2(n10298), .ZN(n10301) );
  XOR2_X1 U11150 ( .A(n10302), .B(n10301), .Z(n10305) );
  AOI22_X1 U11151 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10683), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10303) );
  OAI21_X1 U11152 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(P1_U3243) );
  INV_X1 U11153 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10319) );
  INV_X1 U11154 ( .A(n10306), .ZN(n10307) );
  OAI211_X1 U11155 ( .C1(n10309), .C2(n10308), .A(n10685), .B(n10307), .ZN(
        n10316) );
  OAI211_X1 U11156 ( .C1(n10312), .C2(n10311), .A(n10689), .B(n10310), .ZN(
        n10315) );
  NAND2_X1 U11157 ( .A1(n10693), .A2(n10313), .ZN(n10314) );
  AND3_X1 U11158 ( .A1(n10316), .A2(n10315), .A3(n10314), .ZN(n10318) );
  OAI211_X1 U11159 ( .C1(n10480), .C2(n10319), .A(n10318), .B(n10317), .ZN(
        P1_U3249) );
  INV_X1 U11160 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U11161 ( .A1(n10321), .A2(n10320), .ZN(n10324) );
  INV_X1 U11162 ( .A(n10322), .ZN(n10323) );
  NAND3_X1 U11163 ( .A1(n10689), .A2(n10324), .A3(n10323), .ZN(n10332) );
  NAND2_X1 U11164 ( .A1(n10693), .A2(n10325), .ZN(n10331) );
  AOI21_X1 U11165 ( .B1(n10328), .B2(n10327), .A(n10326), .ZN(n10329) );
  NAND2_X1 U11166 ( .A1(n10685), .A2(n10329), .ZN(n10330) );
  AND3_X1 U11167 ( .A1(n10332), .A2(n10331), .A3(n10330), .ZN(n10334) );
  OAI211_X1 U11168 ( .C1(n10480), .C2(n10335), .A(n10334), .B(n10333), .ZN(
        P1_U3250) );
  INV_X1 U11169 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10351) );
  INV_X1 U11170 ( .A(n10336), .ZN(n10347) );
  AOI21_X1 U11171 ( .B1(n10339), .B2(n10338), .A(n10337), .ZN(n10340) );
  NAND2_X1 U11172 ( .A1(n10685), .A2(n10340), .ZN(n10346) );
  AOI21_X1 U11173 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(n10344) );
  NAND2_X1 U11174 ( .A1(n10689), .A2(n10344), .ZN(n10345) );
  OAI211_X1 U11175 ( .C1(n10461), .C2(n10347), .A(n10346), .B(n10345), .ZN(
        n10348) );
  INV_X1 U11176 ( .A(n10348), .ZN(n10350) );
  OAI211_X1 U11177 ( .C1(n10480), .C2(n10351), .A(n10350), .B(n10349), .ZN(
        P1_U3251) );
  INV_X1 U11178 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10363) );
  AOI211_X1 U11179 ( .C1(n10354), .C2(n10353), .A(n10352), .B(n10470), .ZN(
        n10359) );
  AOI211_X1 U11180 ( .C1(n10357), .C2(n10356), .A(n10355), .B(n10466), .ZN(
        n10358) );
  AOI211_X1 U11181 ( .C1(n10693), .C2(n10360), .A(n10359), .B(n10358), .ZN(
        n10362) );
  OAI211_X1 U11182 ( .C1(n10480), .C2(n10363), .A(n10362), .B(n10361), .ZN(
        P1_U3254) );
  INV_X1 U11183 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10379) );
  INV_X1 U11184 ( .A(n10364), .ZN(n10375) );
  AOI21_X1 U11185 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10368) );
  NAND2_X1 U11186 ( .A1(n10689), .A2(n10368), .ZN(n10374) );
  AOI21_X1 U11187 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(n10372) );
  NAND2_X1 U11188 ( .A1(n10685), .A2(n10372), .ZN(n10373) );
  OAI211_X1 U11189 ( .C1(n10461), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        n10376) );
  INV_X1 U11190 ( .A(n10376), .ZN(n10378) );
  OAI211_X1 U11191 ( .C1(n10480), .C2(n10379), .A(n10378), .B(n10377), .ZN(
        P1_U3257) );
  INV_X1 U11192 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10391) );
  AOI211_X1 U11193 ( .C1(n10382), .C2(n10381), .A(n10380), .B(n10466), .ZN(
        n10387) );
  AOI211_X1 U11194 ( .C1(n10385), .C2(n10384), .A(n10383), .B(n10470), .ZN(
        n10386) );
  AOI211_X1 U11195 ( .C1(n10693), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        n10390) );
  OAI211_X1 U11196 ( .C1(n10480), .C2(n10391), .A(n10390), .B(n10389), .ZN(
        P1_U3258) );
  INV_X1 U11197 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10403) );
  OAI21_X1 U11198 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(n10400) );
  OAI21_X1 U11199 ( .B1(n10397), .B2(n10396), .A(n10395), .ZN(n10398) );
  AOI222_X1 U11200 ( .A1(n10400), .A2(n10685), .B1(n10399), .B2(n10693), .C1(
        n10398), .C2(n10689), .ZN(n10402) );
  OAI211_X1 U11201 ( .C1(n10480), .C2(n10403), .A(n10402), .B(n10401), .ZN(
        P1_U3260) );
  INV_X1 U11202 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10419) );
  INV_X1 U11203 ( .A(n10404), .ZN(n10406) );
  NAND2_X1 U11204 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  NAND3_X1 U11205 ( .A1(n10689), .A2(n10408), .A3(n10407), .ZN(n10416) );
  NAND2_X1 U11206 ( .A1(n10410), .A2(n10409), .ZN(n10411) );
  NAND3_X1 U11207 ( .A1(n10685), .A2(n10412), .A3(n10411), .ZN(n10415) );
  NAND2_X1 U11208 ( .A1(n10693), .A2(n10413), .ZN(n10414) );
  OAI211_X1 U11209 ( .C1(n10480), .C2(n10419), .A(n10418), .B(n10417), .ZN(
        P1_U3261) );
  INV_X1 U11210 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10432) );
  OAI21_X1 U11211 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(n10429) );
  NOR2_X1 U11212 ( .A1(n10461), .A2(n10423), .ZN(n10428) );
  AOI211_X1 U11213 ( .C1(n10426), .C2(n10425), .A(n10424), .B(n10470), .ZN(
        n10427) );
  AOI211_X1 U11214 ( .C1(n10689), .C2(n10429), .A(n10428), .B(n10427), .ZN(
        n10431) );
  OAI211_X1 U11215 ( .C1(n10480), .C2(n10432), .A(n10431), .B(n10430), .ZN(
        P1_U3259) );
  INV_X1 U11216 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10448) );
  INV_X1 U11217 ( .A(n10433), .ZN(n10444) );
  AOI21_X1 U11218 ( .B1(n10436), .B2(n10435), .A(n10434), .ZN(n10437) );
  NAND2_X1 U11219 ( .A1(n10685), .A2(n10437), .ZN(n10443) );
  AOI21_X1 U11220 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(n10441) );
  NAND2_X1 U11221 ( .A1(n10689), .A2(n10441), .ZN(n10442) );
  OAI211_X1 U11222 ( .C1(n10461), .C2(n10444), .A(n10443), .B(n10442), .ZN(
        n10445) );
  INV_X1 U11223 ( .A(n10445), .ZN(n10447) );
  OAI211_X1 U11224 ( .C1(n10480), .C2(n10448), .A(n10447), .B(n10446), .ZN(
        P1_U3256) );
  INV_X1 U11225 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10465) );
  INV_X1 U11226 ( .A(n10449), .ZN(n10460) );
  OAI21_X1 U11227 ( .B1(n10452), .B2(n10451), .A(n10450), .ZN(n10453) );
  NAND2_X1 U11228 ( .A1(n10689), .A2(n10453), .ZN(n10459) );
  OAI21_X1 U11229 ( .B1(n10456), .B2(n10455), .A(n10454), .ZN(n10457) );
  NAND2_X1 U11230 ( .A1(n10685), .A2(n10457), .ZN(n10458) );
  OAI211_X1 U11231 ( .C1(n10461), .C2(n10460), .A(n10459), .B(n10458), .ZN(
        n10462) );
  INV_X1 U11232 ( .A(n10462), .ZN(n10464) );
  OAI211_X1 U11233 ( .C1(n10480), .C2(n10465), .A(n10464), .B(n10463), .ZN(
        P1_U3255) );
  INV_X1 U11234 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10479) );
  AOI211_X1 U11235 ( .C1(n10469), .C2(n10468), .A(n10467), .B(n10466), .ZN(
        n10475) );
  AOI211_X1 U11236 ( .C1(n10473), .C2(n10472), .A(n10471), .B(n10470), .ZN(
        n10474) );
  AOI211_X1 U11237 ( .C1(n10693), .C2(n10476), .A(n10475), .B(n10474), .ZN(
        n10478) );
  OAI211_X1 U11238 ( .C1(n10480), .C2(n10479), .A(n10478), .B(n10477), .ZN(
        P1_U3253) );
  OAI21_X1 U11239 ( .B1(n10482), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10481), .ZN(
        n10484) );
  AOI22_X1 U11240 ( .A1(n10484), .A2(n10671), .B1(n10483), .B2(n10662), .ZN(
        n10497) );
  OAI21_X1 U11241 ( .B1(n10486), .B2(n10485), .A(n10670), .ZN(n10488) );
  NOR2_X1 U11242 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  AOI21_X1 U11243 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(n10661), .A(n10489), .ZN(
        n10496) );
  OAI21_X1 U11244 ( .B1(n10491), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10490), .ZN(
        n10493) );
  NAND2_X1 U11245 ( .A1(n10493), .A2(n10492), .ZN(n10494) );
  NAND4_X1 U11246 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        P2_U3187) );
  OAI21_X1 U11247 ( .B1(n10499), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10498), .ZN(
        n10501) );
  AOI22_X1 U11248 ( .A1(n10501), .A2(n10671), .B1(n10500), .B2(n10662), .ZN(
        n10513) );
  OAI21_X1 U11249 ( .B1(n10504), .B2(n10503), .A(n10502), .ZN(n10505) );
  AOI22_X1 U11250 ( .A1(n10505), .A2(n10670), .B1(n10661), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n10512) );
  AOI21_X1 U11251 ( .B1(n10508), .B2(n10507), .A(n10506), .ZN(n10509) );
  OR2_X1 U11252 ( .A1(n10509), .A2(n10677), .ZN(n10510) );
  NAND4_X1 U11253 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        P2_U3189) );
  AOI22_X1 U11254 ( .A1(n10514), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n10529) );
  OAI21_X1 U11255 ( .B1(n10517), .B2(n10516), .A(n10515), .ZN(n10522) );
  OAI21_X1 U11256 ( .B1(n10520), .B2(n10519), .A(n10518), .ZN(n10521) );
  AOI22_X1 U11257 ( .A1(n10522), .A2(n10671), .B1(n10670), .B2(n10521), .ZN(
        n10528) );
  AOI21_X1 U11258 ( .B1(n10523), .B2(n10524), .A(n5025), .ZN(n10525) );
  OR2_X1 U11259 ( .A1(n10525), .A2(n10677), .ZN(n10526) );
  NAND4_X1 U11260 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        P2_U3190) );
  AOI22_X1 U11261 ( .A1(n10530), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n10545) );
  OAI21_X1 U11262 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10532), .A(n10531), .ZN(
        n10537) );
  OAI21_X1 U11263 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(n10536) );
  AOI22_X1 U11264 ( .A1(n10537), .A2(n10671), .B1(n10670), .B2(n10536), .ZN(
        n10544) );
  AOI21_X1 U11265 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(n10541) );
  OR2_X1 U11266 ( .A1(n10677), .A2(n10541), .ZN(n10542) );
  NAND4_X1 U11267 ( .A1(n10545), .A2(n10544), .A3(n10543), .A4(n10542), .ZN(
        P2_U3191) );
  AOI22_X1 U11268 ( .A1(n10546), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10562) );
  OAI21_X1 U11269 ( .B1(n10549), .B2(n10548), .A(n10547), .ZN(n10554) );
  OAI21_X1 U11270 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(n10553) );
  AOI22_X1 U11271 ( .A1(n10554), .A2(n10671), .B1(n10670), .B2(n10553), .ZN(
        n10561) );
  AOI21_X1 U11272 ( .B1(n10557), .B2(n10556), .A(n10555), .ZN(n10558) );
  OR2_X1 U11273 ( .A1(n10558), .A2(n10677), .ZN(n10559) );
  NAND4_X1 U11274 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        P2_U3192) );
  AOI22_X1 U11275 ( .A1(n10563), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10578) );
  OAI21_X1 U11276 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10565), .A(n10564), 
        .ZN(n10570) );
  OAI21_X1 U11277 ( .B1(n10568), .B2(n10567), .A(n10566), .ZN(n10569) );
  AOI22_X1 U11278 ( .A1(n10570), .A2(n10671), .B1(n10670), .B2(n10569), .ZN(
        n10577) );
  AOI21_X1 U11279 ( .B1(n10573), .B2(n10572), .A(n10571), .ZN(n10574) );
  OR2_X1 U11280 ( .A1(n10677), .A2(n10574), .ZN(n10575) );
  NAND4_X1 U11281 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        P2_U3193) );
  AOI22_X1 U11282 ( .A1(n10661), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n10579), 
        .B2(n10662), .ZN(n10596) );
  OAI21_X1 U11283 ( .B1(n10582), .B2(n10581), .A(n10580), .ZN(n10587) );
  OAI21_X1 U11284 ( .B1(n10585), .B2(n10584), .A(n10583), .ZN(n10586) );
  AOI22_X1 U11285 ( .A1(n10587), .A2(n10671), .B1(n10670), .B2(n10586), .ZN(
        n10595) );
  INV_X1 U11286 ( .A(n10588), .ZN(n10589) );
  AOI21_X1 U11287 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(n10592) );
  OR2_X1 U11288 ( .A1(n10592), .A2(n10677), .ZN(n10593) );
  NAND4_X1 U11289 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        P2_U3194) );
  AOI22_X1 U11290 ( .A1(n10597), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10612) );
  OAI21_X1 U11291 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10599), .A(n10598), 
        .ZN(n10604) );
  OAI21_X1 U11292 ( .B1(n10602), .B2(n10601), .A(n10600), .ZN(n10603) );
  AOI22_X1 U11293 ( .A1(n10604), .A2(n10671), .B1(n10670), .B2(n10603), .ZN(
        n10611) );
  AOI21_X1 U11294 ( .B1(n10607), .B2(n10606), .A(n10605), .ZN(n10608) );
  OR2_X1 U11295 ( .A1(n10608), .A2(n10677), .ZN(n10609) );
  NAND4_X1 U11296 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        P2_U3195) );
  AOI22_X1 U11297 ( .A1(n10613), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10628) );
  OAI21_X1 U11298 ( .B1(n10616), .B2(n10615), .A(n10614), .ZN(n10621) );
  OAI21_X1 U11299 ( .B1(n10619), .B2(n10618), .A(n10617), .ZN(n10620) );
  AOI22_X1 U11300 ( .A1(n10621), .A2(n10671), .B1(n10670), .B2(n10620), .ZN(
        n10627) );
  NAND2_X1 U11301 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10626)
         );
  AOI21_X1 U11302 ( .B1(n4974), .B2(n10623), .A(n10622), .ZN(n10624) );
  OR2_X1 U11303 ( .A1(n10624), .A2(n10677), .ZN(n10625) );
  NAND4_X1 U11304 ( .A1(n10628), .A2(n10627), .A3(n10626), .A4(n10625), .ZN(
        P2_U3196) );
  AOI22_X1 U11305 ( .A1(n10629), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10644) );
  OAI21_X1 U11306 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10631), .A(n10630), 
        .ZN(n10636) );
  OAI21_X1 U11307 ( .B1(n10634), .B2(n10633), .A(n10632), .ZN(n10635) );
  AOI22_X1 U11308 ( .A1(n10636), .A2(n10671), .B1(n10670), .B2(n10635), .ZN(
        n10643) );
  AOI21_X1 U11309 ( .B1(n10639), .B2(n10638), .A(n10637), .ZN(n10640) );
  OR2_X1 U11310 ( .A1(n10677), .A2(n10640), .ZN(n10641) );
  NAND4_X1 U11311 ( .A1(n10644), .A2(n10643), .A3(n10642), .A4(n10641), .ZN(
        P2_U3197) );
  AOI22_X1 U11312 ( .A1(n10645), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10660) );
  OAI21_X1 U11313 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(n10653) );
  OAI21_X1 U11314 ( .B1(n10651), .B2(n10650), .A(n10649), .ZN(n10652) );
  AOI22_X1 U11315 ( .A1(n10653), .A2(n10671), .B1(n10670), .B2(n10652), .ZN(
        n10659) );
  AOI21_X1 U11316 ( .B1(n10655), .B2(n10654), .A(n4981), .ZN(n10656) );
  OR2_X1 U11317 ( .A1(n10656), .A2(n10677), .ZN(n10657) );
  NAND4_X1 U11318 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        P2_U3198) );
  AOI22_X1 U11319 ( .A1(n10663), .A2(n10662), .B1(n10661), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10681) );
  OAI21_X1 U11320 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10665), .A(n10664), 
        .ZN(n10672) );
  OAI21_X1 U11321 ( .B1(n10668), .B2(n10667), .A(n10666), .ZN(n10669) );
  AOI22_X1 U11322 ( .A1(n10672), .A2(n10671), .B1(n10670), .B2(n10669), .ZN(
        n10680) );
  NAND2_X1 U11323 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10679)
         );
  AOI21_X1 U11324 ( .B1(n10675), .B2(n10674), .A(n10673), .ZN(n10676) );
  OR2_X1 U11325 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  NAND4_X1 U11326 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        P2_U3199) );
  XOR2_X1 U11327 ( .A(P1_RD_REG_SCAN_IN), .B(n5060), .Z(U126) );
  AOI21_X1 U11328 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n10683), .A(n10682), .ZN(
        n10699) );
  OAI211_X1 U11329 ( .C1(n10687), .C2(n10686), .A(n10685), .B(n10684), .ZN(
        n10696) );
  OAI211_X1 U11330 ( .C1(n10691), .C2(n10690), .A(n10689), .B(n10688), .ZN(
        n10695) );
  NAND2_X1 U11331 ( .A1(n10693), .A2(n10692), .ZN(n10694) );
  AND3_X1 U11332 ( .A1(n10696), .A2(n10695), .A3(n10694), .ZN(n10698) );
  NAND3_X1 U11333 ( .A1(n10699), .A2(n10698), .A3(n10697), .ZN(P1_U3247) );
  INV_X1 U11334 ( .A(n10700), .ZN(n10715) );
  INV_X1 U11335 ( .A(n10701), .ZN(n10703) );
  INV_X1 U11336 ( .A(n10702), .ZN(n10719) );
  NOR3_X1 U11337 ( .A1(n10715), .A2(n10703), .A3(n10719), .ZN(n10711) );
  NOR2_X1 U11338 ( .A1(n10705), .A2(n10704), .ZN(n10718) );
  NAND3_X1 U11339 ( .A1(n7554), .A2(n10719), .A3(n10706), .ZN(n10707) );
  OAI21_X1 U11340 ( .B1(n10709), .B2(n10708), .A(n10707), .ZN(n10710) );
  NOR3_X1 U11341 ( .A1(n10711), .A2(n10718), .A3(n10710), .ZN(n10713) );
  AOI22_X1 U11342 ( .A1(n4932), .A2(n10714), .B1(n10713), .B2(n10712), .ZN(
        P1_U3293) );
  AOI21_X1 U11343 ( .B1(n10810), .B2(n10716), .A(n10715), .ZN(n10717) );
  AOI211_X1 U11344 ( .C1(n10719), .C2(n7554), .A(n10718), .B(n10717), .ZN(
        n10722) );
  INV_X1 U11345 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U11346 ( .A1(n10819), .A2(n10722), .B1(n10720), .B2(n10818), .ZN(
        P1_U3522) );
  INV_X1 U11347 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U11348 ( .A1(n10823), .A2(n10722), .B1(n10721), .B2(n10820), .ZN(
        P1_U3453) );
  INV_X1 U11349 ( .A(n10723), .ZN(n10728) );
  OAI21_X1 U11350 ( .B1(n10725), .B2(n10814), .A(n10724), .ZN(n10727) );
  AOI211_X1 U11351 ( .C1(n10746), .C2(n10728), .A(n10727), .B(n10726), .ZN(
        n10730) );
  AOI22_X1 U11352 ( .A1(n10819), .A2(n10730), .B1(n6349), .B2(n10818), .ZN(
        P1_U3523) );
  INV_X1 U11353 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U11354 ( .A1(n10823), .A2(n10730), .B1(n10729), .B2(n10820), .ZN(
        P1_U3456) );
  NOR2_X1 U11355 ( .A1(n10732), .A2(n10731), .ZN(n10737) );
  OAI211_X1 U11356 ( .C1(n10735), .C2(n10814), .A(n10734), .B(n10733), .ZN(
        n10736) );
  AOI211_X1 U11357 ( .C1(n10739), .C2(n10738), .A(n10737), .B(n10736), .ZN(
        n10740) );
  AOI22_X1 U11358 ( .A1(n10819), .A2(n10740), .B1(n6330), .B2(n10818), .ZN(
        P1_U3524) );
  AOI22_X1 U11359 ( .A1(n10823), .A2(n10740), .B1(n6329), .B2(n10820), .ZN(
        P1_U3459) );
  INV_X1 U11360 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U11361 ( .A1(n10843), .A2(n10742), .B1(n10741), .B2(n10840), .ZN(
        P2_U3396) );
  OAI21_X1 U11362 ( .B1(n10744), .B2(n10814), .A(n10743), .ZN(n10745) );
  AOI21_X1 U11363 ( .B1(n10747), .B2(n10746), .A(n10745), .ZN(n10748) );
  AND2_X1 U11364 ( .A1(n10749), .A2(n10748), .ZN(n10750) );
  AOI22_X1 U11365 ( .A1(n10819), .A2(n10750), .B1(n9463), .B2(n10818), .ZN(
        P1_U3525) );
  AOI22_X1 U11366 ( .A1(n10823), .A2(n10750), .B1(n6366), .B2(n10820), .ZN(
        P1_U3462) );
  INV_X1 U11367 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U11368 ( .A1(n10843), .A2(n10752), .B1(n10751), .B2(n10840), .ZN(
        P2_U3399) );
  INV_X1 U11369 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U11370 ( .A1(n10843), .A2(n10754), .B1(n10753), .B2(n10840), .ZN(
        P2_U3402) );
  OAI211_X1 U11371 ( .C1(n10757), .C2(n10814), .A(n10756), .B(n10755), .ZN(
        n10758) );
  AOI21_X1 U11372 ( .B1(n10806), .B2(n10759), .A(n10758), .ZN(n10760) );
  AOI22_X1 U11373 ( .A1(n10819), .A2(n10760), .B1(n6383), .B2(n10818), .ZN(
        P1_U3526) );
  AOI22_X1 U11374 ( .A1(n10823), .A2(n10760), .B1(n6379), .B2(n10820), .ZN(
        P1_U3465) );
  INV_X1 U11375 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U11376 ( .A1(n10843), .A2(n10762), .B1(n10761), .B2(n10840), .ZN(
        P2_U3405) );
  INV_X1 U11377 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U11378 ( .A1(n10843), .A2(n10764), .B1(n10763), .B2(n10840), .ZN(
        P2_U3408) );
  OAI211_X1 U11379 ( .C1(n10767), .C2(n10814), .A(n10766), .B(n10765), .ZN(
        n10768) );
  AOI21_X1 U11380 ( .B1(n10806), .B2(n10769), .A(n10768), .ZN(n10771) );
  AOI22_X1 U11381 ( .A1(n10819), .A2(n10771), .B1(n10770), .B2(n10818), .ZN(
        P1_U3528) );
  AOI22_X1 U11382 ( .A1(n10823), .A2(n10771), .B1(n6418), .B2(n10820), .ZN(
        P1_U3471) );
  INV_X1 U11383 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U11384 ( .A1(n10843), .A2(n10773), .B1(n10772), .B2(n10840), .ZN(
        P2_U3411) );
  OAI211_X1 U11385 ( .C1(n5342), .C2(n10814), .A(n10775), .B(n10774), .ZN(
        n10776) );
  AOI21_X1 U11386 ( .B1(n10806), .B2(n10777), .A(n10776), .ZN(n10779) );
  AOI22_X1 U11387 ( .A1(n10819), .A2(n10779), .B1(n6438), .B2(n10818), .ZN(
        P1_U3530) );
  INV_X1 U11388 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U11389 ( .A1(n10823), .A2(n10779), .B1(n10778), .B2(n10820), .ZN(
        P1_U3477) );
  INV_X1 U11390 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U11391 ( .A1(n10843), .A2(n10781), .B1(n10780), .B2(n10840), .ZN(
        P2_U3414) );
  OAI211_X1 U11392 ( .C1(n10784), .C2(n10814), .A(n10783), .B(n10782), .ZN(
        n10785) );
  AOI21_X1 U11393 ( .B1(n10806), .B2(n10786), .A(n10785), .ZN(n10788) );
  AOI22_X1 U11394 ( .A1(n10819), .A2(n10788), .B1(n6454), .B2(n10818), .ZN(
        P1_U3531) );
  INV_X1 U11395 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U11396 ( .A1(n10823), .A2(n10788), .B1(n10787), .B2(n10820), .ZN(
        P1_U3480) );
  INV_X1 U11397 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U11398 ( .A1(n10843), .A2(n10790), .B1(n10789), .B2(n10840), .ZN(
        P2_U3417) );
  OAI211_X1 U11399 ( .C1(n10793), .C2(n10814), .A(n10792), .B(n10791), .ZN(
        n10794) );
  AOI21_X1 U11400 ( .B1(n10795), .B2(n10806), .A(n10794), .ZN(n10797) );
  AOI22_X1 U11401 ( .A1(n10819), .A2(n10797), .B1(n9524), .B2(n10818), .ZN(
        P1_U3532) );
  INV_X1 U11402 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U11403 ( .A1(n10823), .A2(n10797), .B1(n10796), .B2(n10820), .ZN(
        P1_U3483) );
  INV_X1 U11404 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U11405 ( .A1(n10843), .A2(n10799), .B1(n10798), .B2(n10840), .ZN(
        P2_U3420) );
  INV_X1 U11406 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U11407 ( .A1(n10843), .A2(n10801), .B1(n10800), .B2(n10840), .ZN(
        P2_U3423) );
  OAI21_X1 U11408 ( .B1(n10803), .B2(n10814), .A(n10802), .ZN(n10804) );
  AOI211_X1 U11409 ( .C1(n10807), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        n10809) );
  AOI22_X1 U11410 ( .A1(n10819), .A2(n10809), .B1(n9522), .B2(n10818), .ZN(
        P1_U3534) );
  INV_X1 U11411 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U11412 ( .A1(n10823), .A2(n10809), .B1(n10808), .B2(n10820), .ZN(
        P1_U3489) );
  NOR2_X1 U11413 ( .A1(n10811), .A2(n10810), .ZN(n10817) );
  OAI211_X1 U11414 ( .C1(n10815), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n10816) );
  AOI21_X1 U11415 ( .B1(n10817), .B2(n8077), .A(n10816), .ZN(n10822) );
  AOI22_X1 U11416 ( .A1(n10819), .A2(n10822), .B1(n9521), .B2(n10818), .ZN(
        P1_U3535) );
  INV_X1 U11417 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U11418 ( .A1(n10823), .A2(n10822), .B1(n10821), .B2(n10820), .ZN(
        P1_U3492) );
  INV_X1 U11419 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U11420 ( .A1(n10843), .A2(n10825), .B1(n10824), .B2(n10840), .ZN(
        P2_U3429) );
  INV_X1 U11421 ( .A(n10826), .ZN(n10836) );
  INV_X1 U11422 ( .A(n10827), .ZN(n10832) );
  INV_X1 U11423 ( .A(n10828), .ZN(n10830) );
  OAI22_X1 U11424 ( .A1(n10832), .A2(n10831), .B1(n10830), .B2(n10829), .ZN(
        n10834) );
  AOI211_X1 U11425 ( .C1(n10836), .C2(n10835), .A(n10834), .B(n10833), .ZN(
        n10838) );
  AOI22_X1 U11426 ( .A1(n10839), .A2(n6936), .B1(n10838), .B2(n10837), .ZN(
        P2_U3219) );
  INV_X1 U11427 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U11428 ( .A1(n10843), .A2(n10842), .B1(n10841), .B2(n10840), .ZN(
        P2_U3432) );
  AOI22_X1 U11429 ( .A1(n10847), .A2(n10846), .B1(n10845), .B2(n10844), .ZN(
        n10859) );
  NAND2_X1 U11430 ( .A1(n10849), .A2(n10848), .ZN(n10850) );
  NAND2_X1 U11431 ( .A1(n10851), .A2(n10850), .ZN(n10855) );
  AOI222_X1 U11432 ( .A1(n10857), .A2(n10856), .B1(n10855), .B2(n10854), .C1(
        n10853), .C2(n10852), .ZN(n10858) );
  OAI211_X1 U11433 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5965), .A(n10859), .B(
        n10858), .ZN(P2_U3168) );
  XNOR2_X1 U11434 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X2 U5046 ( .A(n6666), .Z(n4939) );
  CLKBUF_X1 U5051 ( .A(n5734), .Z(n6112) );
  CLKBUF_X1 U5125 ( .A(n6147), .Z(n4941) );
  NAND2_X1 U5231 ( .A1(n7345), .A2(n7383), .ZN(n7350) );
  CLKBUF_X1 U8422 ( .A(n5376), .Z(n4934) );
endmodule

