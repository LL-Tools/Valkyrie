

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677;

  BUF_X1 U2246 ( .A(n2420), .Z(n3842) );
  CLKBUF_X2 U2247 ( .A(n2414), .Z(n2611) );
  CLKBUF_X2 U2248 ( .A(n2652), .Z(n3838) );
  INV_X2 U2249 ( .A(n3523), .ZN(n3530) );
  INV_X1 U2250 ( .A(n3531), .ZN(n2865) );
  NAND2_X1 U2251 ( .A1(n2722), .A2(n4334), .ZN(n2986) );
  NOR2_X2 U2252 ( .A1(n3276), .A2(n3698), .ZN(n3305) );
  AND2_X1 U2253 ( .A1(n2722), .A2(n2850), .ZN(n4504) );
  OR2_X2 U2254 ( .A1(n2830), .A2(n2829), .ZN(n2833) );
  NAND2_X2 U2255 ( .A1(n2665), .A2(n3874), .ZN(n3008) );
  XNOR2_X2 U2256 ( .A(n2384), .B(IR_REG_30__SCAN_IN), .ZN(n2391) );
  NAND2_X2 U2257 ( .A1(n2736), .A2(IR_REG_31__SCAN_IN), .ZN(n2384) );
  AOI21_X2 U2258 ( .B1(n3705), .B2(n3707), .A(n3704), .ZN(n3676) );
  XNOR2_X2 U2259 ( .A(n2202), .B(n2209), .ZN(n4028) );
  OAI21_X1 U2260 ( .B1(n4146), .B2(n2651), .A(n2600), .ZN(n4228) );
  NAND2_X1 U2261 ( .A1(n2878), .A2(n4145), .ZN(n3827) );
  NAND2_X1 U2262 ( .A1(n3014), .A2(n3376), .ZN(n3104) );
  NAND2_X1 U2263 ( .A1(n2400), .A2(n2399), .ZN(n2661) );
  INV_X2 U2264 ( .A(n2407), .ZN(n2400) );
  CLKBUF_X3 U2265 ( .A(n2417), .Z(n2418) );
  NAND2_X1 U2266 ( .A1(n2311), .A2(n2699), .ZN(n2934) );
  AOI21_X1 U2267 ( .B1(n4504), .B2(n4207), .A(n4206), .ZN(n4208) );
  OAI21_X2 U2268 ( .B1(n3692), .B2(n3693), .A(n3694), .ZN(n3615) );
  NOR2_X2 U2269 ( .A1(n4106), .A2(n4085), .ZN(n4084) );
  OR2_X1 U2270 ( .A1(n4401), .A2(n2269), .ZN(n2274) );
  OAI21_X1 U2271 ( .B1(n3658), .B2(n3659), .A(n3660), .ZN(n3753) );
  NOR2_X1 U2272 ( .A1(n2183), .A2(n2261), .ZN(n2263) );
  NAND2_X1 U2273 ( .A1(n2128), .A2(n2127), .ZN(n3717) );
  AND2_X1 U2274 ( .A1(n2955), .A2(n2950), .ZN(n2127) );
  NAND2_X1 U2275 ( .A1(n2040), .A2(n3115), .ZN(n3106) );
  INV_X1 U2276 ( .A(n3104), .ZN(n2040) );
  INV_X2 U2277 ( .A(n2999), .ZN(n4182) );
  NAND2_X2 U2278 ( .A1(n2979), .A2(n4145), .ZN(n2999) );
  NAND4_X1 U2279 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(n3801)
         );
  NAND4_X2 U2280 ( .A1(n2425), .A2(n2424), .A3(n2423), .A4(n2422), .ZN(n4006)
         );
  NAND4_X1 U2281 ( .A1(n2413), .A2(n2412), .A3(n2411), .A4(n2410), .ZN(n3609)
         );
  NAND2_X2 U2282 ( .A1(n2986), .A2(n2859), .ZN(n3531) );
  NAND4_X1 U2283 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .ZN(n4008)
         );
  INV_X1 U2284 ( .A(n4504), .ZN(n4478) );
  NAND2_X1 U2285 ( .A1(n2646), .A2(IR_REG_31__SCAN_IN), .ZN(n2648) );
  AND2_X1 U2286 ( .A1(n2391), .A2(n2389), .ZN(n2417) );
  INV_X1 U2287 ( .A(n3610), .ZN(n3083) );
  NAND2_X1 U2288 ( .A1(n2646), .A2(n2369), .ZN(n3986) );
  AND2_X1 U2289 ( .A1(n2857), .A2(n2711), .ZN(n2850) );
  AOI22_X1 U2290 ( .A1(n2780), .A2(REG2_REG_3__SCAN_IN), .B1(n2324), .B2(n4339), .ZN(n2325) );
  OAI21_X1 U2291 ( .B1(n2366), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2368) );
  XNOR2_X1 U2292 ( .A(n2307), .B(n2303), .ZN(n2744) );
  OR2_X1 U2293 ( .A1(n2304), .A2(n2225), .ZN(n2305) );
  AND2_X1 U2294 ( .A1(n2293), .A2(n2302), .ZN(n3992) );
  NOR2_X1 U2295 ( .A1(n2302), .A2(n2301), .ZN(n2306) );
  AND2_X1 U2296 ( .A1(n2282), .A2(n2284), .ZN(n2166) );
  AND4_X1 U2297 ( .A1(n2281), .A2(n2280), .A3(n2279), .A4(n2278), .ZN(n2282)
         );
  NOR2_X1 U2298 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2190)
         );
  NOR2_X1 U2299 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2191)
         );
  NOR2_X1 U2300 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2189)
         );
  INV_X1 U2301 ( .A(IR_REG_3__SCAN_IN), .ZN(n2188) );
  NOR2_X1 U2302 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2044)
         );
  NOR2_X2 U2303 ( .A1(n3201), .A2(n3756), .ZN(n2043) );
  OR2_X2 U2304 ( .A1(n3161), .A2(n3664), .ZN(n3201) );
  NOR2_X4 U2305 ( .A1(n2199), .A2(n2193), .ZN(n2283) );
  NAND3_X2 U2306 ( .A1(n2210), .A2(n2044), .A3(n2188), .ZN(n2199) );
  MUX2_X1 U2307 ( .A(n2312), .B(n2313), .S(n2317), .Z(n2004) );
  NOR2_X2 U2308 ( .A1(n2996), .A2(n2906), .ZN(n3084) );
  AND2_X1 U2309 ( .A1(n2905), .A2(n4478), .ZN(n2005) );
  AND2_X1 U2310 ( .A1(n2905), .A2(n4478), .ZN(n2006) );
  AND2_X1 U2311 ( .A1(n2905), .A2(n4478), .ZN(n2946) );
  XNOR2_X2 U2312 ( .A(n2648), .B(n2647), .ZN(n2722) );
  INV_X1 U2313 ( .A(n2986), .ZN(n2125) );
  NAND2_X1 U2314 ( .A1(n2102), .A2(n2104), .ZN(n2100) );
  NAND2_X1 U2315 ( .A1(n3672), .A2(n3673), .ZN(n2147) );
  NOR2_X1 U2316 ( .A1(n2087), .A2(n2084), .ZN(n2083) );
  INV_X1 U2317 ( .A(n2464), .ZN(n2084) );
  INV_X1 U2318 ( .A(n2088), .ZN(n2087) );
  NOR2_X1 U2319 ( .A1(n2288), .A2(IR_REG_27__SCAN_IN), .ZN(n2381) );
  INV_X1 U2320 ( .A(IR_REG_17__SCAN_IN), .ZN(n2196) );
  INV_X1 U2321 ( .A(n2276), .ZN(n2197) );
  INV_X1 U2322 ( .A(n3811), .ZN(n2148) );
  NAND2_X1 U2323 ( .A1(n2140), .A2(n2137), .ZN(n2136) );
  NAND2_X1 U2324 ( .A1(n2142), .A2(n2138), .ZN(n2137) );
  NAND2_X1 U2325 ( .A1(n2126), .A2(n2124), .ZN(n2860) );
  NAND2_X1 U2326 ( .A1(n2905), .A2(n2399), .ZN(n2126) );
  BUF_X1 U2327 ( .A(n2419), .Z(n2651) );
  NAND2_X1 U2328 ( .A1(n2391), .A2(n2392), .ZN(n2419) );
  AND2_X1 U2329 ( .A1(n2390), .A2(n2389), .ZN(n2652) );
  XNOR2_X1 U2330 ( .A(n2323), .B(n4339), .ZN(n2780) );
  NAND2_X1 U2331 ( .A1(n2062), .A2(n2061), .ZN(n2060) );
  INV_X1 U2332 ( .A(n4350), .ZN(n2061) );
  NOR2_X1 U2333 ( .A1(n2011), .A2(n2623), .ZN(n2631) );
  AND2_X1 U2334 ( .A1(n2031), .A2(n2103), .ZN(n2102) );
  OR2_X1 U2335 ( .A1(n2104), .A2(n3940), .ZN(n2103) );
  NOR2_X1 U2336 ( .A1(n2117), .A2(n2520), .ZN(n2114) );
  AND2_X1 U2337 ( .A1(n3756), .A2(n3665), .ZN(n2520) );
  NOR2_X1 U2338 ( .A1(n2119), .A2(n2021), .ZN(n2117) );
  NOR2_X1 U2339 ( .A1(n3409), .A2(n2132), .ZN(n2131) );
  NOR2_X1 U2340 ( .A1(n3648), .A2(n2170), .ZN(n2169) );
  INV_X1 U2341 ( .A(n2176), .ZN(n2170) );
  INV_X1 U2342 ( .A(n3596), .ZN(n3403) );
  INV_X1 U2343 ( .A(n3253), .ZN(n2070) );
  INV_X1 U2344 ( .A(n2260), .ZN(n2261) );
  NOR2_X1 U2345 ( .A1(n4406), .A2(n2073), .ZN(n2350) );
  AND2_X1 U2346 ( .A1(n2349), .A2(REG2_REG_15__SCAN_IN), .ZN(n2073) );
  NAND2_X1 U2347 ( .A1(n2025), .A2(n2629), .ZN(n2097) );
  NOR2_X1 U2348 ( .A1(n2089), .A2(n2483), .ZN(n2088) );
  INV_X1 U2349 ( .A(n2474), .ZN(n2089) );
  INV_X1 U2350 ( .A(n2473), .ZN(n2086) );
  NAND2_X1 U2351 ( .A1(n2053), .A2(REG3_REG_7__SCAN_IN), .ZN(n2465) );
  INV_X1 U2352 ( .A(n2455), .ZN(n2053) );
  OR2_X1 U2353 ( .A1(n4004), .A2(n3376), .ZN(n3859) );
  OR2_X1 U2354 ( .A1(n3609), .A2(n2921), .ZN(n3848) );
  INV_X1 U2355 ( .A(n4155), .ZN(n4162) );
  INV_X1 U2356 ( .A(n3992), .ZN(n2857) );
  NAND2_X1 U2357 ( .A1(n2178), .A2(n2286), .ZN(n2288) );
  INV_X1 U2358 ( .A(n2301), .ZN(n2286) );
  INV_X1 U2359 ( .A(IR_REG_26__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2360 ( .A1(n2309), .A2(n2297), .ZN(n2301) );
  INV_X1 U2361 ( .A(IR_REG_23__SCAN_IN), .ZN(n2297) );
  AND3_X1 U2362 ( .A1(n2266), .A2(n2264), .A3(n2271), .ZN(n2195) );
  INV_X1 U2363 ( .A(IR_REG_15__SCAN_IN), .ZN(n2266) );
  INV_X1 U2364 ( .A(IR_REG_6__SCAN_IN), .ZN(n2200) );
  AND2_X1 U2365 ( .A1(n2631), .A2(REG3_REG_27__SCAN_IN), .ZN(n2637) );
  AND2_X1 U2366 ( .A1(n3587), .A2(n3588), .ZN(n3497) );
  INV_X1 U2367 ( .A(n3535), .ZN(n2138) );
  AOI21_X1 U2368 ( .B1(n2143), .B2(n2141), .A(n2026), .ZN(n2140) );
  INV_X1 U2369 ( .A(n2023), .ZN(n2141) );
  AND2_X1 U2370 ( .A1(n2174), .A2(n2035), .ZN(n2172) );
  NAND2_X1 U2371 ( .A1(n2151), .A2(n3450), .ZN(n2150) );
  INV_X1 U2372 ( .A(n2153), .ZN(n2151) );
  NAND2_X1 U2373 ( .A1(n2175), .A2(n3470), .ZN(n2174) );
  NOR2_X1 U2374 ( .A1(n2744), .A2(n2697), .ZN(n2311) );
  NAND2_X1 U2375 ( .A1(n2216), .A2(n2215), .ZN(n2219) );
  NAND2_X1 U2376 ( .A1(n2790), .A2(n2224), .ZN(n2228) );
  OAI21_X1 U2377 ( .B1(n2827), .B2(n2232), .A(n2233), .ZN(n2238) );
  NAND2_X1 U2378 ( .A1(n2833), .A2(n2334), .ZN(n2335) );
  OR2_X1 U2379 ( .A1(n4335), .A2(n2980), .ZN(n2334) );
  NAND2_X1 U2380 ( .A1(n4353), .A2(n2069), .ZN(n2339) );
  OR2_X1 U2381 ( .A1(n4469), .A2(n2338), .ZN(n2069) );
  AND2_X1 U2382 ( .A1(n2060), .A2(n2033), .ZN(n2248) );
  NAND2_X1 U2383 ( .A1(n4372), .A2(n2342), .ZN(n2344) );
  XNOR2_X1 U2384 ( .A(n2350), .B(n2547), .ZN(n4418) );
  NAND2_X1 U2385 ( .A1(n4418), .A2(n4417), .ZN(n4416) );
  NAND2_X1 U2386 ( .A1(n4428), .A2(n2067), .ZN(n2353) );
  NAND2_X1 U2387 ( .A1(n4458), .A2(n2068), .ZN(n2067) );
  INV_X1 U2388 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2068) );
  NOR2_X1 U2389 ( .A1(n2353), .A2(n2354), .ZN(n2365) );
  OR2_X1 U2390 ( .A1(n4036), .A2(n2645), .ZN(n4049) );
  NAND2_X1 U2391 ( .A1(n2094), .A2(n2091), .ZN(n4050) );
  NOR2_X1 U2392 ( .A1(n2093), .A2(n2092), .ZN(n2091) );
  OR2_X1 U2393 ( .A1(n2622), .A2(n2097), .ZN(n2094) );
  NOR2_X1 U2394 ( .A1(n2097), .A2(n2621), .ZN(n2092) );
  AND2_X1 U2395 ( .A1(n4228), .A2(n3488), .ZN(n2601) );
  NAND2_X1 U2396 ( .A1(n2581), .A2(n2685), .ZN(n2106) );
  NAND2_X1 U2397 ( .A1(n2582), .A2(n2105), .ZN(n2104) );
  NAND2_X1 U2398 ( .A1(n3939), .A2(n3940), .ZN(n2105) );
  AOI21_X1 U2399 ( .B1(n4174), .B2(n3940), .A(n2104), .ZN(n2101) );
  AOI21_X1 U2400 ( .B1(n2110), .B2(n2010), .A(n2027), .ZN(n2109) );
  OR2_X1 U2401 ( .A1(n3286), .A2(n2010), .ZN(n2111) );
  AND2_X1 U2402 ( .A1(n3930), .A2(n2029), .ZN(n2110) );
  NAND2_X1 U2403 ( .A1(n4284), .A2(n4278), .ZN(n2538) );
  OR2_X1 U2404 ( .A1(n4278), .A2(n4284), .ZN(n2537) );
  NAND2_X1 U2405 ( .A1(n3146), .A2(n2118), .ZN(n2115) );
  NOR2_X1 U2406 ( .A1(n2120), .A2(n2021), .ZN(n2118) );
  NAND2_X1 U2407 ( .A1(n2121), .A2(n2500), .ZN(n2120) );
  INV_X1 U2408 ( .A(n2510), .ZN(n2121) );
  OR2_X1 U2409 ( .A1(n2510), .A2(n2511), .ZN(n2119) );
  AND2_X1 U2410 ( .A1(n2512), .A2(REG3_REG_13__SCAN_IN), .ZN(n2521) );
  OR2_X1 U2411 ( .A1(n3150), .A2(n3131), .ZN(n2491) );
  OR2_X1 U2412 ( .A1(n3144), .A2(n3143), .ZN(n3146) );
  NOR2_X1 U2413 ( .A1(n2437), .A2(n2789), .ZN(n2446) );
  NAND2_X1 U2414 ( .A1(n2039), .A2(n3031), .ZN(n3067) );
  AND2_X1 U2415 ( .A1(n2990), .A2(n2408), .ZN(n2891) );
  INV_X1 U2416 ( .A(IR_REG_20__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U2417 ( .A1(n2717), .A2(n2755), .ZN(n2976) );
  INV_X1 U2418 ( .A(IR_REG_24__SCAN_IN), .ZN(n2309) );
  INV_X1 U2419 ( .A(IR_REG_19__SCAN_IN), .ZN(n2367) );
  OR2_X1 U2420 ( .A1(n2637), .A2(n2051), .ZN(n4067) );
  NOR2_X1 U2421 ( .A1(n2631), .A2(REG3_REG_27__SCAN_IN), .ZN(n2051) );
  XNOR2_X1 U2422 ( .A(n2912), .B(n2910), .ZN(n2874) );
  AND2_X1 U2423 ( .A1(n2011), .A2(n2615), .ZN(n4107) );
  INV_X1 U2424 ( .A(n3454), .ZN(n3698) );
  INV_X1 U2425 ( .A(n4120), .ZN(n4231) );
  XNOR2_X1 U2426 ( .A(n2940), .B(n2939), .ZN(n2919) );
  OAI21_X1 U2427 ( .B1(n4083), .B2(n2651), .A(n2628), .ZN(n4211) );
  NAND4_X1 U2428 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(n4275)
         );
  NAND4_X1 U2429 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n4005)
         );
  OAI21_X1 U2430 ( .B1(n2798), .B2(n2328), .A(n2327), .ZN(n2329) );
  AND2_X1 U2431 ( .A1(n2329), .A2(n2074), .ZN(n2786) );
  INV_X1 U2432 ( .A(n2787), .ZN(n2074) );
  XNOR2_X1 U2433 ( .A(n2335), .B(n2838), .ZN(n2837) );
  XNOR2_X1 U2434 ( .A(n2248), .B(n4467), .ZN(n4359) );
  NAND2_X1 U2435 ( .A1(n4425), .A2(n2185), .ZN(n2314) );
  NOR2_X1 U2436 ( .A1(n2314), .A2(n2315), .ZN(n2375) );
  NAND2_X1 U2437 ( .A1(n2162), .A2(n3573), .ZN(n2155) );
  AOI21_X1 U2438 ( .B1(n2163), .B2(n2160), .A(n2159), .ZN(n2158) );
  INV_X1 U2439 ( .A(n3821), .ZN(n2159) );
  INV_X1 U2440 ( .A(n3574), .ZN(n2160) );
  NOR2_X1 U2441 ( .A1(n3947), .A2(n3948), .ZN(n2050) );
  INV_X1 U2442 ( .A(n3946), .ZN(n2049) );
  INV_X1 U2443 ( .A(IR_REG_14__SCAN_IN), .ZN(n2264) );
  AOI21_X1 U2444 ( .B1(n2158), .B2(n2161), .A(n2154), .ZN(n2153) );
  NAND2_X1 U2445 ( .A1(n2155), .A2(n2164), .ZN(n2154) );
  INV_X1 U2446 ( .A(n2163), .ZN(n2161) );
  INV_X1 U2447 ( .A(n3685), .ZN(n2164) );
  AND2_X1 U2448 ( .A1(n2156), .A2(n3450), .ZN(n2152) );
  OR2_X1 U2449 ( .A1(n2158), .A2(n2162), .ZN(n2156) );
  NOR2_X1 U2450 ( .A1(n3739), .A2(n2177), .ZN(n2176) );
  INV_X1 U2451 ( .A(n3471), .ZN(n2177) );
  AND2_X1 U2452 ( .A1(n3574), .A2(n2022), .ZN(n2162) );
  AOI21_X1 U2453 ( .B1(n3573), .B2(n3574), .A(n2022), .ZN(n2163) );
  NAND2_X1 U2454 ( .A1(n2054), .A2(REG3_REG_15__SCAN_IN), .ZN(n2541) );
  INV_X1 U2455 ( .A(n2530), .ZN(n2054) );
  NAND2_X1 U2456 ( .A1(n2521), .A2(REG3_REG_14__SCAN_IN), .ZN(n2530) );
  NOR2_X1 U2457 ( .A1(n4023), .A2(n2016), .ZN(n2323) );
  INV_X1 U2458 ( .A(n2095), .ZN(n2093) );
  AOI21_X1 U2459 ( .B1(n2630), .B2(n2096), .A(n2028), .ZN(n2095) );
  INV_X1 U2460 ( .A(n2097), .ZN(n2096) );
  OR2_X1 U2461 ( .A1(n4231), .A2(n4099), .ZN(n2621) );
  OR2_X1 U2462 ( .A1(n3309), .A2(n3308), .ZN(n3347) );
  NOR2_X1 U2463 ( .A1(n2541), .A2(n2540), .ZN(n2549) );
  NOR2_X1 U2464 ( .A1(n2557), .A2(n4619), .ZN(n2055) );
  OR2_X1 U2465 ( .A1(n2493), .A2(n3775), .ZN(n2502) );
  NAND2_X1 U2466 ( .A1(n2484), .A2(REG3_REG_10__SCAN_IN), .ZN(n2493) );
  INV_X1 U2467 ( .A(n2435), .ZN(n2080) );
  OR2_X1 U2468 ( .A1(n4005), .A2(n3031), .ZN(n3854) );
  INV_X1 U2469 ( .A(n2416), .ZN(n2077) );
  NAND2_X1 U2470 ( .A1(n2042), .A2(n2041), .ZN(n3276) );
  INV_X1 U2471 ( .A(n3277), .ZN(n2042) );
  OR2_X1 U2472 ( .A1(n3242), .A2(n3921), .ZN(n3243) );
  INV_X1 U2473 ( .A(n2754), .ZN(n2848) );
  AOI21_X1 U2474 ( .B1(n2015), .B2(n3772), .A(n2131), .ZN(n2130) );
  NAND2_X1 U2475 ( .A1(n2186), .A2(n3469), .ZN(n3470) );
  INV_X1 U2476 ( .A(n3619), .ZN(n3469) );
  NOR2_X1 U2477 ( .A1(n2572), .A2(n3746), .ZN(n2577) );
  NAND2_X1 U2478 ( .A1(n2168), .A2(n2167), .ZN(n3763) );
  OR2_X1 U2479 ( .A1(n2171), .A2(n3648), .ZN(n2167) );
  AND2_X1 U2480 ( .A1(n2172), .A2(n3647), .ZN(n2171) );
  NAND2_X1 U2481 ( .A1(n3404), .A2(n3403), .ZN(n3597) );
  INV_X1 U2482 ( .A(n2883), .ZN(n2872) );
  NAND2_X1 U2483 ( .A1(n2157), .A2(n2163), .ZN(n3820) );
  NAND2_X1 U2484 ( .A1(n3572), .A2(n3574), .ZN(n2157) );
  NOR3_X1 U2485 ( .A1(n4051), .A2(n2048), .A3(n3952), .ZN(n2047) );
  INV_X1 U2486 ( .A(n4049), .ZN(n2046) );
  AND3_X1 U2487 ( .A1(n4018), .A2(IR_REG_0__SCAN_IN), .A3(REG2_REG_0__SCAN_IN), 
        .ZN(n4015) );
  NAND2_X1 U2488 ( .A1(n2056), .A2(n2208), .ZN(n2214) );
  NOR2_X1 U2489 ( .A1(n2786), .A2(n2331), .ZN(n2332) );
  NOR2_X1 U2490 ( .A1(n2795), .A2(n2330), .ZN(n2331) );
  NAND2_X1 U2491 ( .A1(n2840), .A2(n2241), .ZN(n2062) );
  NAND2_X1 U2492 ( .A1(n2240), .A2(n2239), .ZN(n2241) );
  INV_X1 U2493 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3775) );
  NOR2_X1 U2494 ( .A1(n4367), .A2(n2065), .ZN(n2254) );
  INV_X1 U2495 ( .A(IR_REG_13__SCAN_IN), .ZN(n2194) );
  NAND2_X1 U2496 ( .A1(n2072), .A2(n2071), .ZN(n2346) );
  OR2_X1 U2497 ( .A1(n2732), .A2(REG2_REG_13__SCAN_IN), .ZN(n2071) );
  AND2_X1 U2498 ( .A1(n2058), .A2(n2019), .ZN(n4403) );
  NAND2_X1 U2499 ( .A1(n4416), .A2(n2351), .ZN(n4429) );
  AND2_X1 U2500 ( .A1(n2357), .A2(n2356), .ZN(n2772) );
  AND2_X1 U2501 ( .A1(n4035), .A2(n2638), .ZN(n3542) );
  AND2_X1 U2502 ( .A1(n3936), .A2(n3935), .ZN(n4077) );
  AND2_X1 U2503 ( .A1(n2609), .A2(n2608), .ZN(n4100) );
  NOR2_X1 U2504 ( .A1(n2595), .A2(n2594), .ZN(n2603) );
  NAND2_X1 U2505 ( .A1(n2100), .A2(n2593), .ZN(n2099) );
  OR2_X1 U2506 ( .A1(n2584), .A2(n2583), .ZN(n2595) );
  NAND2_X1 U2507 ( .A1(n2577), .A2(REG3_REG_21__SCAN_IN), .ZN(n2584) );
  NOR2_X2 U2508 ( .A1(n4177), .A2(n4245), .ZN(n4163) );
  NAND2_X1 U2509 ( .A1(n2055), .A2(REG3_REG_19__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U2510 ( .A1(n2549), .A2(REG3_REG_17__SCAN_IN), .ZN(n2557) );
  INV_X1 U2511 ( .A(n2055), .ZN(n2565) );
  NAND2_X1 U2512 ( .A1(n3245), .A2(n4284), .ZN(n3277) );
  AND2_X1 U2513 ( .A1(n3958), .A2(n3956), .ZN(n3920) );
  NAND2_X1 U2514 ( .A1(n3230), .A2(n2528), .ZN(n2529) );
  INV_X1 U2515 ( .A(n4291), .ZN(n2528) );
  NOR2_X1 U2516 ( .A1(n2502), .A2(n2501), .ZN(n2512) );
  AOI21_X1 U2517 ( .B1(n2088), .B2(n2086), .A(n2017), .ZN(n2085) );
  NAND2_X1 U2518 ( .A1(n2052), .A2(REG3_REG_8__SCAN_IN), .ZN(n2475) );
  INV_X1 U2519 ( .A(n2465), .ZN(n2052) );
  INV_X1 U2520 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3731) );
  NOR2_X1 U2521 ( .A1(n2475), .A2(n3731), .ZN(n2484) );
  INV_X1 U2522 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U2523 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2437) );
  NAND2_X1 U2524 ( .A1(n3848), .A2(n3851), .ZN(n3926) );
  NAND2_X1 U2525 ( .A1(n2891), .A2(n3926), .ZN(n2890) );
  AND2_X1 U2526 ( .A1(n4008), .A2(n2803), .ZN(n2991) );
  NOR2_X2 U2527 ( .A1(n4053), .A2(n4054), .ZN(n4200) );
  INV_X1 U2528 ( .A(n4099), .ZN(n4104) );
  OR2_X2 U2529 ( .A1(n2012), .A2(n4104), .ZN(n4106) );
  NOR2_X1 U2530 ( .A1(n2611), .A2(n2610), .ZN(n4227) );
  NAND2_X1 U2531 ( .A1(n4241), .A2(n4143), .ZN(n4142) );
  INV_X1 U2532 ( .A(n2685), .ZN(n4245) );
  NAND2_X1 U2533 ( .A1(n3154), .A2(n3153), .ZN(n3161) );
  INV_X1 U2534 ( .A(n3599), .ZN(n3131) );
  INV_X1 U2535 ( .A(n4277), .ZN(n4292) );
  AND2_X1 U2536 ( .A1(n2693), .A2(n2692), .ZN(n4259) );
  INV_X1 U2537 ( .A(n3802), .ZN(n3039) );
  INV_X1 U2538 ( .A(n4286), .ZN(n4274) );
  OR2_X1 U2539 ( .A1(n4341), .A2(n2852), .ZN(n4277) );
  INV_X1 U2540 ( .A(n4502), .ZN(n4490) );
  NAND2_X1 U2541 ( .A1(n2316), .A2(n2291), .ZN(n2313) );
  AOI21_X1 U2542 ( .B1(n2289), .B2(n2287), .A(n2184), .ZN(n2312) );
  NAND2_X1 U2543 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2184) );
  INV_X1 U2544 ( .A(IR_REG_16__SCAN_IN), .ZN(n2271) );
  AND2_X1 U2545 ( .A1(n2270), .A2(n2268), .ZN(n2349) );
  INV_X1 U2546 ( .A(IR_REG_7__SCAN_IN), .ZN(n4535) );
  INV_X1 U2547 ( .A(IR_REG_4__SCAN_IN), .ZN(n2187) );
  INV_X1 U2548 ( .A(IR_REG_2__SCAN_IN), .ZN(n2209) );
  NAND2_X1 U2549 ( .A1(n2144), .A2(n2145), .ZN(n3566) );
  INV_X1 U2550 ( .A(n3466), .ZN(n3624) );
  INV_X1 U2551 ( .A(n2135), .ZN(n2134) );
  OAI21_X1 U2552 ( .B1(n2140), .B2(n3535), .A(n2136), .ZN(n2135) );
  NAND2_X1 U2553 ( .A1(n2143), .A2(n3535), .ZN(n2139) );
  AND2_X1 U2554 ( .A1(n2173), .A2(n2172), .ZN(n3652) );
  INV_X1 U2555 ( .A(n3818), .ZN(n3823) );
  AOI21_X1 U2556 ( .B1(n3615), .B2(n3471), .A(n3470), .ZN(n3741) );
  NAND2_X1 U2557 ( .A1(n2173), .A2(n2174), .ZN(n3742) );
  INV_X1 U2558 ( .A(n3427), .ZN(n3756) );
  NAND2_X1 U2559 ( .A1(n2938), .A2(n2937), .ZN(n3830) );
  OAI21_X1 U2560 ( .B1(n4067), .B2(n2651), .A(n2636), .ZN(n4080) );
  NAND2_X1 U2561 ( .A1(n2620), .A2(n2619), .ZN(n4120) );
  INV_X1 U2562 ( .A(n4100), .ZN(n4139) );
  INV_X1 U2563 ( .A(n4248), .ZN(n3997) );
  NAND4_X1 U2564 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n4179)
         );
  NAND4_X1 U2565 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(n3999)
         );
  NAND4_X1 U2566 ( .A1(n2517), .A2(n2516), .A3(n2515), .A4(n2514), .ZN(n3665)
         );
  NAND4_X1 U2567 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n4004)
         );
  OR2_X1 U2568 ( .A1(n2419), .A2(n2409), .ZN(n2411) );
  NAND2_X1 U2569 ( .A1(n2652), .A2(REG0_REG_1__SCAN_IN), .ZN(n2395) );
  NOR2_X1 U2570 ( .A1(n4025), .A2(n4024), .ZN(n4023) );
  AOI21_X1 U2571 ( .B1(n4009), .B2(REG2_REG_1__SCAN_IN), .A(n4015), .ZN(n4025)
         );
  XNOR2_X1 U2572 ( .A(n2214), .B(n2785), .ZN(n2779) );
  XNOR2_X1 U2573 ( .A(n2332), .B(n4337), .ZN(n2818) );
  NAND2_X1 U2574 ( .A1(n2230), .A2(n2229), .ZN(n2827) );
  NAND2_X1 U2575 ( .A1(n2013), .A2(REG1_REG_8__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U2576 ( .A1(n2337), .A2(n2336), .ZN(n4354) );
  NAND2_X1 U2577 ( .A1(n4354), .A2(n4355), .ZN(n4353) );
  INV_X1 U2578 ( .A(n2060), .ZN(n4349) );
  INV_X1 U2579 ( .A(n2062), .ZN(n2179) );
  XNOR2_X1 U2580 ( .A(n2339), .B(n4467), .ZN(n4364) );
  NAND2_X1 U2581 ( .A1(n4364), .A2(REG2_REG_10__SCAN_IN), .ZN(n4363) );
  INV_X1 U2582 ( .A(n4464), .ZN(n4377) );
  NOR2_X1 U2583 ( .A1(n2249), .A2(n4358), .ZN(n4369) );
  NOR2_X1 U2584 ( .A1(n4369), .A2(n4368), .ZN(n4367) );
  XNOR2_X1 U2585 ( .A(n2344), .B(n2343), .ZN(n4384) );
  NAND2_X1 U2586 ( .A1(n4384), .A2(REG2_REG_12__SCAN_IN), .ZN(n4383) );
  XNOR2_X1 U2587 ( .A(n2254), .B(n2343), .ZN(n4379) );
  NOR2_X1 U2588 ( .A1(n4379), .A2(n4380), .ZN(n4378) );
  NAND2_X1 U2589 ( .A1(n4383), .A2(n2345), .ZN(n3257) );
  XNOR2_X1 U2590 ( .A(n2274), .B(n4459), .ZN(n4415) );
  NAND2_X1 U2591 ( .A1(n4426), .A2(n4427), .ZN(n4425) );
  XNOR2_X1 U2592 ( .A(n2063), .B(n2376), .ZN(n2181) );
  OR2_X1 U2593 ( .A1(n2375), .A2(n2038), .ZN(n2063) );
  AND2_X1 U2594 ( .A1(n2772), .A2(n2806), .ZN(n4434) );
  XNOR2_X1 U2595 ( .A(n2066), .B(n2371), .ZN(n2374) );
  NOR2_X1 U2596 ( .A1(n2365), .A2(n2037), .ZN(n2066) );
  AND2_X1 U2597 ( .A1(n2772), .A2(n3990), .ZN(n4432) );
  AOI21_X1 U2598 ( .B1(n4050), .B2(n4049), .A(n4048), .ZN(n4052) );
  XNOR2_X1 U2599 ( .A(n4050), .B(n4049), .ZN(n3552) );
  AND2_X1 U2600 ( .A1(n4061), .A2(n4159), .ZN(n4217) );
  OR2_X1 U2601 ( .A1(n2624), .A2(n2631), .ZN(n4083) );
  OAI21_X1 U2602 ( .B1(n4174), .B2(n2104), .A(n2102), .ZN(n4151) );
  AND2_X1 U2603 ( .A1(n2107), .A2(n2106), .ZN(n4152) );
  INV_X1 U2604 ( .A(n2101), .ZN(n2107) );
  OAI21_X1 U2605 ( .B1(n4174), .B2(n3939), .A(n3940), .ZN(n3339) );
  NAND2_X1 U2606 ( .A1(n2111), .A2(n2110), .ZN(n3303) );
  NOR2_X1 U2607 ( .A1(n2113), .A2(n2112), .ZN(n3177) );
  INV_X1 U2608 ( .A(n2114), .ZN(n2112) );
  INV_X1 U2609 ( .A(n2115), .ZN(n2113) );
  OAI21_X1 U2610 ( .B1(n2116), .B2(n2120), .A(n2119), .ZN(n3189) );
  INV_X1 U2611 ( .A(n3146), .ZN(n2116) );
  NAND2_X1 U2612 ( .A1(n3103), .A2(n2473), .ZN(n2090) );
  AND2_X1 U2613 ( .A1(n2999), .A2(n2987), .ZN(n4176) );
  INV_X1 U2614 ( .A(n4439), .ZN(n4164) );
  NAND2_X1 U2615 ( .A1(n3021), .A2(n2435), .ZN(n3060) );
  INV_X1 U2616 ( .A(n4448), .ZN(n4145) );
  AND2_X1 U2617 ( .A1(n3317), .A2(n4504), .ZN(n4439) );
  AND2_X1 U2618 ( .A1(n2877), .A2(n2977), .ZN(n4448) );
  OR2_X1 U2619 ( .A1(n2724), .A2(n2976), .ZN(n4519) );
  AND2_X2 U2620 ( .A1(n2725), .A2(n2976), .ZN(n4511) );
  XNOR2_X1 U2621 ( .A(n2386), .B(IR_REG_29__SCAN_IN), .ZN(n2392) );
  AND2_X1 U2622 ( .A1(n2306), .A2(n2303), .ZN(n2304) );
  NAND2_X1 U2623 ( .A1(n2308), .A2(IR_REG_31__SCAN_IN), .ZN(n2310) );
  INV_X1 U2624 ( .A(n2711), .ZN(n4334) );
  XNOR2_X1 U2625 ( .A(n2251), .B(IR_REG_11__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U2626 ( .A1(n2245), .A2(n2244), .ZN(n4469) );
  AND2_X1 U2627 ( .A1(n2217), .A2(n2213), .ZN(n4339) );
  NAND2_X1 U2628 ( .A1(n2064), .A2(IR_REG_31__SCAN_IN), .ZN(n2202) );
  INV_X1 U2629 ( .A(n2210), .ZN(n2064) );
  XNOR2_X1 U2630 ( .A(n2204), .B(n2203), .ZN(n4010) );
  INV_X1 U2631 ( .A(n2329), .ZN(n2788) );
  INV_X1 U2632 ( .A(IR_REG_31__SCAN_IN), .ZN(n2225) );
  INV_X1 U2633 ( .A(n2905), .ZN(n3521) );
  AND2_X2 U2634 ( .A1(n2934), .A2(n2125), .ZN(n2908) );
  OR2_X1 U2635 ( .A1(n3753), .A2(n3750), .ZN(n2007) );
  INV_X1 U2636 ( .A(n3031), .ZN(n3721) );
  AND2_X1 U2637 ( .A1(n2114), .A2(n3929), .ZN(n2008) );
  AND2_X1 U2638 ( .A1(n3403), .A2(n2024), .ZN(n2009) );
  AND2_X1 U2639 ( .A1(n3312), .A2(n3454), .ZN(n2010) );
  NAND4_X1 U2640 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .ZN(n4000)
         );
  NAND2_X1 U2641 ( .A1(n3859), .A2(n3865), .ZN(n2985) );
  OR2_X1 U2642 ( .A1(n2614), .A2(n4623), .ZN(n2011) );
  OR2_X1 U2643 ( .A1(n4142), .A2(n4227), .ZN(n2012) );
  XOR2_X1 U2644 ( .A(n2238), .B(n2838), .Z(n2013) );
  INV_X1 U2645 ( .A(n2908), .ZN(n3523) );
  NAND2_X1 U2646 ( .A1(n2390), .A2(n2392), .ZN(n2420) );
  INV_X1 U2647 ( .A(n2414), .ZN(n3906) );
  OAI21_X1 U2648 ( .B1(n4073), .B2(n2630), .A(n2629), .ZN(n4058) );
  OAI21_X1 U2649 ( .B1(n2414), .B2(DATAI_1_), .A(n2398), .ZN(n2997) );
  INV_X1 U2650 ( .A(n2997), .ZN(n2399) );
  INV_X1 U2651 ( .A(n3115), .ZN(n3640) );
  INV_X1 U2652 ( .A(n2946), .ZN(n3524) );
  NOR2_X1 U2653 ( .A1(n3368), .A2(n3367), .ZN(n2014) );
  NAND2_X1 U2654 ( .A1(n3409), .A2(n2132), .ZN(n2015) );
  INV_X1 U2655 ( .A(n2146), .ZN(n2145) );
  OAI21_X1 U2656 ( .B1(n3811), .B2(n2147), .A(n3809), .ZN(n2146) );
  AND2_X1 U2657 ( .A1(n2322), .A2(REG2_REG_2__SCAN_IN), .ZN(n2016) );
  AND2_X1 U2658 ( .A1(n3116), .A2(n3050), .ZN(n2017) );
  NAND2_X1 U2659 ( .A1(n2283), .A2(n2282), .ZN(n2018) );
  OR2_X1 U2660 ( .A1(n2263), .A2(n4462), .ZN(n2019) );
  INV_X1 U2661 ( .A(IR_REG_28__SCAN_IN), .ZN(n2317) );
  AND2_X1 U2662 ( .A1(n2345), .A2(n2070), .ZN(n2020) );
  NAND2_X1 U2663 ( .A1(n3615), .A2(n2176), .ZN(n2173) );
  AND2_X1 U2664 ( .A1(n2283), .A2(n2194), .ZN(n2257) );
  INV_X1 U2665 ( .A(n4272), .ZN(n2041) );
  AND2_X1 U2666 ( .A1(n2519), .A2(n3427), .ZN(n2021) );
  OAI21_X1 U2667 ( .B1(n3320), .B2(n3322), .A(n3321), .ZN(n4174) );
  XOR2_X1 U2668 ( .A(n3442), .B(n2865), .Z(n2022) );
  AND2_X1 U2669 ( .A1(n2148), .A2(n3673), .ZN(n2023) );
  NAND2_X1 U2670 ( .A1(n2129), .A2(n2130), .ZN(n3658) );
  NAND2_X1 U2671 ( .A1(n3597), .A2(n3409), .ZN(n3770) );
  INV_X1 U2672 ( .A(n3771), .ZN(n2132) );
  INV_X1 U2673 ( .A(IR_REG_25__SCAN_IN), .ZN(n2303) );
  OR2_X1 U2674 ( .A1(n3772), .A2(n3771), .ZN(n2024) );
  OR2_X1 U2675 ( .A1(n4080), .A2(n4210), .ZN(n2025) );
  INV_X1 U2676 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4657) );
  INV_X1 U2677 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2454) );
  OAI21_X1 U2678 ( .B1(n3572), .B2(n3573), .A(n2162), .ZN(n2165) );
  NOR2_X1 U2679 ( .A1(n3528), .A2(n3529), .ZN(n2026) );
  AND2_X1 U2680 ( .A1(n3627), .A2(n2719), .ZN(n2027) );
  INV_X1 U2681 ( .A(n2143), .ZN(n2142) );
  NOR2_X1 U2682 ( .A1(n3565), .A2(n2146), .ZN(n2143) );
  NOR2_X1 U2683 ( .A1(n3525), .A2(n4062), .ZN(n2028) );
  NAND2_X1 U2684 ( .A1(n4275), .A2(n3698), .ZN(n2029) );
  AND2_X1 U2685 ( .A1(n2140), .A2(n2138), .ZN(n2030) );
  AND2_X1 U2686 ( .A1(n4153), .A2(n2106), .ZN(n2031) );
  OR2_X1 U2687 ( .A1(n4120), .A2(n4104), .ZN(n2032) );
  NAND2_X1 U2688 ( .A1(n2482), .A2(REG1_REG_9__SCAN_IN), .ZN(n2033) );
  INV_X1 U2689 ( .A(IR_REG_8__SCAN_IN), .ZN(n2236) );
  AND2_X1 U2690 ( .A1(n2111), .A2(n2029), .ZN(n2034) );
  NAND2_X1 U2691 ( .A1(n3477), .A2(n3476), .ZN(n2035) );
  INV_X1 U2692 ( .A(n3739), .ZN(n2175) );
  OAI21_X1 U2693 ( .B1(n3633), .B2(n3634), .A(n3635), .ZN(n3728) );
  NAND2_X1 U2694 ( .A1(n2983), .A2(n2464), .ZN(n3103) );
  NAND2_X1 U2695 ( .A1(n2090), .A2(n2474), .ZN(n3055) );
  NAND2_X1 U2696 ( .A1(n3146), .A2(n2500), .ZN(n3160) );
  XNOR2_X1 U2697 ( .A(n2305), .B(IR_REG_26__SCAN_IN), .ZN(n2699) );
  AND4_X1 U2698 ( .A1(n3951), .A2(n3949), .A3(n2050), .A4(n2049), .ZN(n2036)
         );
  NAND2_X1 U2699 ( .A1(n2128), .A2(n2950), .ZN(n3715) );
  NAND2_X1 U2700 ( .A1(n2434), .A2(n3932), .ZN(n3021) );
  INV_X1 U2701 ( .A(n2043), .ZN(n3202) );
  INV_X1 U2702 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U2703 ( .A1(n2890), .A2(n2416), .ZN(n3074) );
  INV_X1 U2704 ( .A(n3082), .ZN(n2039) );
  AND2_X1 U2705 ( .A1(n2563), .A2(REG2_REG_18__SCAN_IN), .ZN(n2037) );
  AND2_X1 U2706 ( .A1(n2563), .A2(REG1_REG_18__SCAN_IN), .ZN(n2038) );
  AND2_X2 U2707 ( .A1(n3069), .A2(n3039), .ZN(n3014) );
  NOR2_X2 U2708 ( .A1(n3067), .A2(n3066), .ZN(n3069) );
  NAND2_X1 U2709 ( .A1(n3084), .A2(n3083), .ZN(n3082) );
  NAND2_X1 U2710 ( .A1(n2289), .A2(n2381), .ZN(n2316) );
  NOR2_X2 U2711 ( .A1(n2295), .A2(IR_REG_22__SCAN_IN), .ZN(n2289) );
  NAND2_X2 U2712 ( .A1(n2166), .A2(n2283), .ZN(n2295) );
  AND2_X2 U2713 ( .A1(n3093), .A2(n3131), .ZN(n3154) );
  NOR2_X2 U2714 ( .A1(n3106), .A2(n3732), .ZN(n3093) );
  NOR2_X2 U2715 ( .A1(n3202), .A2(n3579), .ZN(n3245) );
  AND2_X2 U2716 ( .A1(n2203), .A2(n2045), .ZN(n2210) );
  INV_X2 U2717 ( .A(IR_REG_0__SCAN_IN), .ZN(n2045) );
  AND2_X2 U2718 ( .A1(n4163), .A2(n4162), .ZN(n4241) );
  NAND3_X1 U2719 ( .A1(n3945), .A2(n2047), .A3(n2046), .ZN(n3982) );
  NAND3_X1 U2720 ( .A1(n3944), .A2(n3950), .A3(n2036), .ZN(n2048) );
  XNOR2_X1 U2721 ( .A(n4028), .B(REG1_REG_2__SCAN_IN), .ZN(n4027) );
  NAND2_X1 U2722 ( .A1(n4026), .A2(n4027), .ZN(n2056) );
  NAND2_X1 U2723 ( .A1(n4014), .A2(n2207), .ZN(n4026) );
  AND2_X1 U2724 ( .A1(n2058), .A2(n2057), .ZN(n4394) );
  AOI21_X1 U2725 ( .B1(n4387), .B2(n4388), .A(n4400), .ZN(n2057) );
  NAND2_X1 U2726 ( .A1(n2059), .A2(REG1_REG_14__SCAN_IN), .ZN(n2058) );
  INV_X1 U2727 ( .A(n4387), .ZN(n2059) );
  AND2_X1 U2728 ( .A1(n4464), .A2(REG1_REG_11__SCAN_IN), .ZN(n2065) );
  NAND2_X1 U2729 ( .A1(n3333), .A2(n3624), .ZN(n3332) );
  XNOR2_X1 U2730 ( .A(n2263), .B(n4462), .ZN(n4387) );
  NAND2_X1 U2731 ( .A1(n2181), .A2(n4434), .ZN(n2377) );
  NAND2_X1 U2732 ( .A1(n4383), .A2(n2020), .ZN(n2072) );
  NAND3_X1 U2733 ( .A1(n2427), .A2(n2076), .A3(n2075), .ZN(n3022) );
  NAND2_X1 U2734 ( .A1(n2426), .A2(n2077), .ZN(n2075) );
  NAND3_X1 U2735 ( .A1(n2426), .A2(n3926), .A3(n2891), .ZN(n2076) );
  OAI21_X1 U2736 ( .B1(n2434), .B2(n2080), .A(n2078), .ZN(n2081) );
  INV_X1 U2737 ( .A(n2079), .ZN(n2078) );
  OAI21_X1 U2738 ( .B1(n3932), .B2(n2080), .A(n2444), .ZN(n2079) );
  NAND2_X1 U2739 ( .A1(n2081), .A2(n2445), .ZN(n3006) );
  NAND2_X1 U2740 ( .A1(n2983), .A2(n2083), .ZN(n2082) );
  NAND2_X1 U2741 ( .A1(n2082), .A2(n2085), .ZN(n3099) );
  NAND2_X1 U2742 ( .A1(n2622), .A2(n2621), .ZN(n4073) );
  AOI21_X1 U2743 ( .B1(n4174), .B2(n2102), .A(n2099), .ZN(n2098) );
  INV_X1 U2744 ( .A(n2098), .ZN(n4130) );
  NAND2_X1 U2745 ( .A1(n3286), .A2(n2110), .ZN(n2108) );
  NAND2_X1 U2746 ( .A1(n2108), .A2(n2109), .ZN(n3320) );
  NAND2_X1 U2747 ( .A1(n2115), .A2(n2008), .ZN(n3176) );
  XNOR2_X1 U2748 ( .A(n2122), .B(n2865), .ZN(n2940) );
  NAND2_X1 U2749 ( .A1(n2123), .A2(n2907), .ZN(n2122) );
  NAND2_X1 U2750 ( .A1(n2908), .A2(n3609), .ZN(n2123) );
  NAND2_X1 U2751 ( .A1(n2908), .A2(n2407), .ZN(n2124) );
  AND2_X4 U2752 ( .A1(n2934), .A2(n2986), .ZN(n2905) );
  NAND2_X1 U2753 ( .A1(n3605), .A2(n3606), .ZN(n2128) );
  NAND2_X1 U2754 ( .A1(n3404), .A2(n2009), .ZN(n2129) );
  AOI21_X1 U2755 ( .B1(n3676), .B2(n2030), .A(n2134), .ZN(n2133) );
  OAI21_X1 U2756 ( .B1(n3676), .B2(n2139), .A(n2133), .ZN(n3541) );
  NAND2_X1 U2757 ( .A1(n3676), .A2(n2023), .ZN(n2144) );
  OAI21_X1 U2758 ( .B1(n3676), .B2(n3672), .A(n3673), .ZN(n3808) );
  NAND2_X1 U2759 ( .A1(n3572), .A2(n2152), .ZN(n2149) );
  NAND2_X1 U2760 ( .A1(n2149), .A2(n2150), .ZN(n3692) );
  INV_X1 U2761 ( .A(n2165), .ZN(n3683) );
  OR2_X1 U2762 ( .A1(n2295), .A2(IR_REG_22__SCAN_IN), .ZN(n2302) );
  NAND2_X1 U2763 ( .A1(n3615), .A2(n2169), .ZN(n2168) );
  OAI21_X1 U2764 ( .B1(n2004), .B2(n2406), .A(n2405), .ZN(n2803) );
  NAND2_X1 U2765 ( .A1(n2414), .A2(IR_REG_0__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U2766 ( .A1(n2004), .A2(n4010), .ZN(n2398) );
  AND2_X1 U2767 ( .A1(n2399), .A2(n2908), .ZN(n2861) );
  OR2_X1 U2768 ( .A1(n2385), .A2(n2225), .ZN(n2386) );
  OR2_X1 U2769 ( .A1(n2934), .A2(n2729), .ZN(n4007) );
  MUX2_X2 U2770 ( .A(REG0_REG_28__SCAN_IN), .B(n2726), .S(n4511), .Z(n2727) );
  MUX2_X2 U2771 ( .A(REG1_REG_28__SCAN_IN), .B(n2726), .S(n4521), .Z(n2718) );
  NAND2_X1 U2772 ( .A1(n3585), .A2(n3502), .ZN(n3705) );
  INV_X1 U2773 ( .A(n2391), .ZN(n2390) );
  AND2_X1 U2774 ( .A1(n2285), .A2(n2303), .ZN(n2178) );
  INV_X1 U2775 ( .A(n3716), .ZN(n2955) );
  OR2_X1 U2776 ( .A1(n3547), .A2(n4329), .ZN(n2180) );
  OR2_X1 U2777 ( .A1(n3547), .A2(n4268), .ZN(n2182) );
  INV_X1 U2778 ( .A(n2838), .ZN(n2239) );
  INV_X1 U2779 ( .A(DATAI_0_), .ZN(n2406) );
  NOR2_X1 U2780 ( .A1(n3260), .A2(n3259), .ZN(n2183) );
  OR2_X1 U2781 ( .A1(n2352), .A2(REG1_REG_17__SCAN_IN), .ZN(n2185) );
  INV_X1 U2782 ( .A(n4395), .ZN(n4462) );
  INV_X1 U2783 ( .A(n3928), .ZN(n3143) );
  OR3_X1 U2784 ( .A1(n3620), .A2(n3617), .A3(n3784), .ZN(n2186) );
  INV_X1 U2785 ( .A(n2985), .ZN(n2462) );
  AOI21_X1 U2786 ( .B1(n3370), .B2(n3369), .A(n2014), .ZN(n3371) );
  INV_X1 U2787 ( .A(IR_REG_22__SCAN_IN), .ZN(n2379) );
  INV_X1 U2788 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2501) );
  INV_X1 U2789 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2540) );
  INV_X1 U2790 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2330) );
  INV_X1 U2791 ( .A(n2274), .ZN(n2273) );
  OR2_X1 U2792 ( .A1(n4248), .A2(n4162), .ZN(n2593) );
  AND2_X1 U2793 ( .A1(n2379), .A2(n2317), .ZN(n2380) );
  INV_X1 U2794 ( .A(IR_REG_21__SCAN_IN), .ZN(n2284) );
  INV_X1 U2795 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4619) );
  NOR2_X1 U2796 ( .A1(n3501), .A2(n3505), .ZN(n3502) );
  NAND2_X1 U2797 ( .A1(n2446), .A2(REG3_REG_6__SCAN_IN), .ZN(n2455) );
  OR3_X1 U2798 ( .A1(n3523), .A2(n2857), .A3(n2856), .ZN(n2881) );
  NAND2_X1 U2799 ( .A1(n2326), .A2(n4338), .ZN(n2327) );
  AND2_X1 U2800 ( .A1(n4212), .A2(n4047), .ZN(n4048) );
  AND2_X1 U2801 ( .A1(n2691), .A2(n3911), .ZN(n3974) );
  AND2_X1 U2802 ( .A1(n3999), .A2(n4272), .ZN(n2548) );
  OR2_X1 U2803 ( .A1(n3047), .A2(n3875), .ZN(n2668) );
  INV_X1 U2804 ( .A(n4000), .ZN(n4278) );
  INV_X1 U2805 ( .A(n2965), .ZN(n3066) );
  NAND2_X1 U2806 ( .A1(n2381), .A2(n2380), .ZN(n2382) );
  OR3_X1 U2807 ( .A1(n2231), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2242) );
  XNOR2_X1 U2808 ( .A(n3380), .B(n3378), .ZN(n3554) );
  AND2_X1 U2809 ( .A1(n2849), .A2(n2978), .ZN(n2883) );
  INV_X1 U2810 ( .A(n4469), .ZN(n2482) );
  INV_X1 U2811 ( .A(n2509), .ZN(n2343) );
  INV_X1 U2812 ( .A(n3974), .ZN(n4059) );
  OR2_X1 U2813 ( .A1(n3347), .A2(n3346), .ZN(n4172) );
  INV_X1 U2814 ( .A(n4273), .ZN(n4285) );
  NOR2_X1 U2815 ( .A1(n2611), .A2(n2576), .ZN(n3743) );
  NOR2_X1 U2816 ( .A1(n2242), .A2(IR_REG_9__SCAN_IN), .ZN(n2246) );
  NOR2_X1 U2817 ( .A1(n2199), .A2(IR_REG_5__SCAN_IN), .ZN(n2226) );
  INV_X1 U2818 ( .A(n3230), .ZN(n3579) );
  AND2_X1 U2819 ( .A1(n2591), .A2(n2590), .ZN(n4248) );
  XNOR2_X1 U2820 ( .A(n2325), .B(n2812), .ZN(n2798) );
  AND2_X1 U2821 ( .A1(n2772), .A2(n4341), .ZN(n4396) );
  AND2_X1 U2822 ( .A1(n3983), .A2(n2850), .ZN(n4273) );
  AND2_X1 U2823 ( .A1(n3898), .A2(n4131), .ZN(n4133) );
  INV_X1 U2824 ( .A(n4259), .ZN(n4159) );
  AND2_X1 U2825 ( .A1(n2722), .A2(n2650), .ZN(n4487) );
  AND2_X1 U2826 ( .A1(n2934), .A2(n4455), .ZN(n2977) );
  XNOR2_X1 U2827 ( .A(n2234), .B(n4535), .ZN(n4335) );
  OR2_X1 U2828 ( .A1(n2872), .A2(n2871), .ZN(n3818) );
  NAND2_X1 U2829 ( .A1(n2644), .A2(n2643), .ZN(n4212) );
  INV_X1 U2830 ( .A(n4434), .ZN(n4400) );
  INV_X1 U2831 ( .A(n4432), .ZN(n4389) );
  INV_X1 U2832 ( .A(n4396), .ZN(n4437) );
  INV_X1 U2833 ( .A(n4176), .ZN(n4169) );
  INV_X1 U2834 ( .A(n4519), .ZN(n4521) );
  INV_X1 U2835 ( .A(n4519), .ZN(n4518) );
  INV_X1 U2836 ( .A(n4511), .ZN(n4509) );
  NAND2_X1 U2837 ( .A1(n2977), .A2(n2754), .ZN(n4634) );
  AND2_X1 U2838 ( .A1(n2933), .A2(STATE_REG_SCAN_IN), .ZN(n4455) );
  INV_X1 U2839 ( .A(n2349), .ZN(n4461) );
  OR2_X1 U2840 ( .A1(n2364), .A2(n2363), .ZN(U3258) );
  INV_X2 U2841 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U2842 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2192)
         );
  NAND4_X1 U2843 ( .A1(n2192), .A2(n2191), .A3(n2190), .A4(n2189), .ZN(n2193)
         );
  NAND2_X1 U2844 ( .A1(n2257), .A2(n2195), .ZN(n2276) );
  NAND2_X1 U2845 ( .A1(n2197), .A2(n2196), .ZN(n2366) );
  NAND2_X1 U2846 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2198) );
  XNOR2_X1 U2847 ( .A(n2198), .B(IR_REG_18__SCAN_IN), .ZN(n2563) );
  INV_X1 U2848 ( .A(n2563), .ZN(n4457) );
  INV_X1 U2849 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2556) );
  AOI22_X1 U2850 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4457), .B1(n2563), .B2(
        n2556), .ZN(n2315) );
  NAND2_X1 U2851 ( .A1(n2226), .A2(n2200), .ZN(n2231) );
  INV_X1 U2852 ( .A(IR_REG_10__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U2853 ( .A1(n2246), .A2(n4640), .ZN(n2201) );
  NAND2_X1 U2854 ( .A1(n2201), .A2(IR_REG_31__SCAN_IN), .ZN(n2251) );
  NAND2_X1 U2855 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2204)
         );
  INV_X1 U2856 ( .A(IR_REG_1__SCAN_IN), .ZN(n2203) );
  INV_X1 U2857 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U2858 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2205) );
  AOI21_X1 U2859 ( .B1(n4010), .B2(n4512), .A(n2205), .ZN(n2206) );
  OR2_X1 U2860 ( .A1(n4010), .A2(n4512), .ZN(n2207) );
  NAND2_X1 U2861 ( .A1(n2206), .A2(n2207), .ZN(n4014) );
  INV_X1 U2862 ( .A(n4028), .ZN(n2322) );
  NAND2_X1 U2863 ( .A1(n2322), .A2(REG1_REG_2__SCAN_IN), .ZN(n2208) );
  NAND2_X1 U2864 ( .A1(n2210), .A2(n2209), .ZN(n2211) );
  NAND2_X1 U2865 ( .A1(n2211), .A2(IR_REG_31__SCAN_IN), .ZN(n2212) );
  NAND2_X1 U2866 ( .A1(n2212), .A2(n2188), .ZN(n2217) );
  OR2_X1 U2867 ( .A1(n2212), .A2(n2188), .ZN(n2213) );
  INV_X1 U2868 ( .A(n4339), .ZN(n2785) );
  NAND2_X1 U2869 ( .A1(n2779), .A2(REG1_REG_3__SCAN_IN), .ZN(n2216) );
  NAND2_X1 U2870 ( .A1(n2214), .A2(n4339), .ZN(n2215) );
  NAND2_X1 U2871 ( .A1(n2217), .A2(IR_REG_31__SCAN_IN), .ZN(n2218) );
  XNOR2_X1 U2872 ( .A(n2218), .B(n2187), .ZN(n2812) );
  XNOR2_X1 U2873 ( .A(n2219), .B(n2812), .ZN(n2810) );
  NAND2_X1 U2874 ( .A1(n2810), .A2(REG1_REG_4__SCAN_IN), .ZN(n2221) );
  INV_X1 U2875 ( .A(n2812), .ZN(n4338) );
  NAND2_X1 U2876 ( .A1(n2219), .A2(n4338), .ZN(n2220) );
  NAND2_X1 U2877 ( .A1(n2221), .A2(n2220), .ZN(n2791) );
  INV_X1 U2878 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U2879 ( .A1(n2199), .A2(IR_REG_31__SCAN_IN), .ZN(n2223) );
  INV_X1 U2880 ( .A(IR_REG_5__SCAN_IN), .ZN(n2222) );
  XNOR2_X1 U2881 ( .A(n2223), .B(n2222), .ZN(n2795) );
  MUX2_X1 U2882 ( .A(n2436), .B(REG1_REG_5__SCAN_IN), .S(n2795), .Z(n2792) );
  NAND2_X1 U2883 ( .A1(n2791), .A2(n2792), .ZN(n2790) );
  OR2_X1 U2884 ( .A1(n2795), .A2(n2436), .ZN(n2224) );
  OR2_X1 U2885 ( .A1(n2226), .A2(n2225), .ZN(n2227) );
  XNOR2_X1 U2886 ( .A(n2227), .B(IR_REG_6__SCAN_IN), .ZN(n4337) );
  INV_X1 U2887 ( .A(n4337), .ZN(n2822) );
  XNOR2_X1 U2888 ( .A(n2228), .B(n2822), .ZN(n2819) );
  NAND2_X1 U2889 ( .A1(n2819), .A2(REG1_REG_6__SCAN_IN), .ZN(n2230) );
  NAND2_X1 U2890 ( .A1(n2228), .A2(n4337), .ZN(n2229) );
  NAND2_X1 U2891 ( .A1(n2231), .A2(IR_REG_31__SCAN_IN), .ZN(n2234) );
  INV_X1 U2892 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2457) );
  NOR2_X1 U2893 ( .A1(n4335), .A2(n2457), .ZN(n2232) );
  NAND2_X1 U2894 ( .A1(n4335), .A2(n2457), .ZN(n2233) );
  NAND2_X1 U2895 ( .A1(n2234), .A2(n4535), .ZN(n2235) );
  NAND2_X1 U2896 ( .A1(n2235), .A2(IR_REG_31__SCAN_IN), .ZN(n2237) );
  XNOR2_X1 U2897 ( .A(n2237), .B(n2236), .ZN(n2838) );
  INV_X1 U2898 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3122) );
  INV_X1 U2899 ( .A(n2238), .ZN(n2240) );
  NAND2_X1 U2900 ( .A1(n2242), .A2(IR_REG_31__SCAN_IN), .ZN(n2243) );
  MUX2_X1 U2901 ( .A(IR_REG_31__SCAN_IN), .B(n2243), .S(IR_REG_9__SCAN_IN), 
        .Z(n2245) );
  INV_X1 U2902 ( .A(n2246), .ZN(n2244) );
  INV_X1 U2903 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U2904 ( .A1(n2482), .A2(n4644), .B1(REG1_REG_9__SCAN_IN), .B2(n4469), .ZN(n4350) );
  OR2_X1 U2905 ( .A1(n2246), .A2(n2225), .ZN(n2247) );
  XNOR2_X1 U2906 ( .A(n2247), .B(IR_REG_10__SCAN_IN), .ZN(n2490) );
  INV_X1 U2907 ( .A(n2490), .ZN(n4467) );
  NOR2_X1 U2908 ( .A1(n2248), .A2(n4467), .ZN(n2249) );
  INV_X1 U2909 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4360) );
  NOR2_X1 U2910 ( .A1(n4360), .A2(n4359), .ZN(n4358) );
  INV_X1 U2911 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U2912 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4377), .B1(n4464), .B2(
        n4576), .ZN(n4368) );
  INV_X1 U2913 ( .A(IR_REG_11__SCAN_IN), .ZN(n2250) );
  NAND2_X1 U2914 ( .A1(n2251), .A2(n2250), .ZN(n2252) );
  NAND2_X1 U2915 ( .A1(n2252), .A2(IR_REG_31__SCAN_IN), .ZN(n2253) );
  XNOR2_X1 U2916 ( .A(n2253), .B(IR_REG_12__SCAN_IN), .ZN(n2509) );
  NOR2_X1 U2917 ( .A1(n2254), .A2(n2343), .ZN(n2255) );
  INV_X1 U2918 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4380) );
  NOR2_X1 U2919 ( .A1(n2255), .A2(n4378), .ZN(n3260) );
  NOR2_X1 U2920 ( .A1(n2283), .A2(n2225), .ZN(n2256) );
  MUX2_X1 U2921 ( .A(n2225), .B(n2256), .S(IR_REG_13__SCAN_IN), .Z(n2258) );
  OR2_X1 U2922 ( .A1(n2258), .A2(n2257), .ZN(n3264) );
  INV_X1 U2923 ( .A(n3264), .ZN(n2732) );
  NAND2_X1 U2924 ( .A1(n2732), .A2(REG1_REG_13__SCAN_IN), .ZN(n2260) );
  INV_X1 U2925 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U2926 ( .A1(n3264), .A2(n3268), .ZN(n2259) );
  NAND2_X1 U2927 ( .A1(n2260), .A2(n2259), .ZN(n3259) );
  OR2_X1 U2928 ( .A1(n2257), .A2(n2225), .ZN(n2262) );
  XNOR2_X1 U2929 ( .A(n2262), .B(IR_REG_14__SCAN_IN), .ZN(n4395) );
  INV_X1 U2930 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U2931 ( .A1(n2257), .A2(n2264), .ZN(n2265) );
  NAND2_X1 U2932 ( .A1(n2265), .A2(IR_REG_31__SCAN_IN), .ZN(n2267) );
  NAND2_X1 U2933 ( .A1(n2267), .A2(n2266), .ZN(n2270) );
  OR2_X1 U2934 ( .A1(n2267), .A2(n2266), .ZN(n2268) );
  INV_X1 U2935 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2532) );
  AOI22_X1 U2936 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4461), .B1(n2349), .B2(
        n2532), .ZN(n4402) );
  NOR2_X1 U2937 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  AND2_X1 U2938 ( .A1(n2349), .A2(REG1_REG_15__SCAN_IN), .ZN(n2269) );
  NAND2_X1 U2939 ( .A1(n2270), .A2(IR_REG_31__SCAN_IN), .ZN(n2272) );
  XNOR2_X1 U2940 ( .A(n2272), .B(n2271), .ZN(n4459) );
  NAND2_X1 U2941 ( .A1(n2273), .A2(n4459), .ZN(n2275) );
  INV_X1 U2942 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U2943 ( .A1(n4415), .A2(n4414), .ZN(n4413) );
  NAND2_X1 U2944 ( .A1(n2275), .A2(n4413), .ZN(n4426) );
  NAND2_X1 U2945 ( .A1(n2276), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  XNOR2_X1 U2946 ( .A(n2277), .B(IR_REG_17__SCAN_IN), .ZN(n2352) );
  INV_X1 U2947 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4645) );
  INV_X1 U2948 ( .A(n2352), .ZN(n4458) );
  AOI22_X1 U2949 ( .A1(n2352), .A2(REG1_REG_17__SCAN_IN), .B1(n4645), .B2(
        n4458), .ZN(n4427) );
  NOR2_X1 U2950 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2281)
         );
  NOR2_X1 U2951 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2280)
         );
  NOR2_X1 U2952 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2279)
         );
  NOR2_X1 U2953 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2278)
         );
  INV_X1 U2954 ( .A(n2288), .ZN(n2287) );
  INV_X1 U2955 ( .A(IR_REG_27__SCAN_IN), .ZN(n2290) );
  NAND2_X1 U2956 ( .A1(n2225), .A2(n2290), .ZN(n2291) );
  MUX2_X2 U2957 ( .A(n2312), .B(n2313), .S(n2317), .Z(n2414) );
  NAND2_X1 U2958 ( .A1(n2295), .A2(IR_REG_31__SCAN_IN), .ZN(n2292) );
  MUX2_X1 U2959 ( .A(IR_REG_31__SCAN_IN), .B(n2292), .S(IR_REG_22__SCAN_IN), 
        .Z(n2293) );
  NAND2_X1 U2960 ( .A1(n2018), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  MUX2_X1 U2961 ( .A(IR_REG_31__SCAN_IN), .B(n2294), .S(IR_REG_21__SCAN_IN), 
        .Z(n2296) );
  NAND2_X1 U2962 ( .A1(n2296), .A2(n2295), .ZN(n2711) );
  AND2_X1 U2963 ( .A1(n3992), .A2(n4334), .ZN(n2712) );
  NAND2_X1 U2964 ( .A1(n2302), .A2(IR_REG_31__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2965 ( .A1(n2298), .A2(n2297), .ZN(n2308) );
  OR2_X1 U2966 ( .A1(n2298), .A2(n2297), .ZN(n2299) );
  NAND2_X1 U2967 ( .A1(n2308), .A2(n2299), .ZN(n2933) );
  AND2_X1 U2968 ( .A1(n2712), .A2(n2933), .ZN(n2300) );
  NOR2_X1 U2969 ( .A1(n2611), .A2(n2300), .ZN(n2357) );
  OR2_X1 U2970 ( .A1(n2306), .A2(n2225), .ZN(n2307) );
  XNOR2_X1 U2971 ( .A(n2310), .B(n2309), .ZN(n2697) );
  NOR2_X1 U2972 ( .A1(n2933), .A2(U3149), .ZN(n3988) );
  OR2_X1 U2973 ( .A1(n2977), .A2(n3988), .ZN(n2356) );
  NOR2_X1 U2974 ( .A1(n2313), .A2(n2312), .ZN(n4040) );
  INV_X1 U2975 ( .A(n4040), .ZN(n2806) );
  AOI211_X1 U2976 ( .C1(n2315), .C2(n2314), .A(n2375), .B(n4400), .ZN(n2364)
         );
  NAND2_X1 U2977 ( .A1(n2316), .A2(IR_REG_31__SCAN_IN), .ZN(n2318) );
  XNOR2_X1 U2978 ( .A(n2318), .B(n2317), .ZN(n4341) );
  INV_X1 U2979 ( .A(n4341), .ZN(n2880) );
  AND2_X1 U2980 ( .A1(n2880), .A2(n4040), .ZN(n3990) );
  NAND2_X1 U2981 ( .A1(REG2_REG_18__SCAN_IN), .A2(n2563), .ZN(n2319) );
  OAI21_X1 U2982 ( .B1(REG2_REG_18__SCAN_IN), .B2(n2563), .A(n2319), .ZN(n2354) );
  NOR2_X1 U2983 ( .A1(n2352), .A2(REG2_REG_17__SCAN_IN), .ZN(n2320) );
  AOI21_X1 U2984 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2352), .A(n2320), .ZN(n4430) );
  INV_X1 U2985 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2338) );
  INV_X1 U2986 ( .A(n4010), .ZN(n4009) );
  XNOR2_X1 U2987 ( .A(n4010), .B(REG2_REG_1__SCAN_IN), .ZN(n4018) );
  INV_X1 U2988 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2321) );
  MUX2_X1 U2989 ( .A(REG2_REG_2__SCAN_IN), .B(n2321), .S(n4028), .Z(n4024) );
  INV_X1 U2990 ( .A(n2323), .ZN(n2324) );
  INV_X1 U2991 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2328) );
  INV_X1 U2992 ( .A(n2325), .ZN(n2326) );
  MUX2_X1 U2993 ( .A(REG2_REG_5__SCAN_IN), .B(n2330), .S(n2795), .Z(n2787) );
  INV_X1 U2994 ( .A(n2332), .ZN(n2333) );
  AOI22_X1 U2995 ( .A1(n2818), .A2(REG2_REG_6__SCAN_IN), .B1(n4337), .B2(n2333), .ZN(n2830) );
  INV_X1 U2996 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2980) );
  MUX2_X1 U2997 ( .A(REG2_REG_7__SCAN_IN), .B(n2980), .S(n4335), .Z(n2829) );
  NAND2_X1 U2998 ( .A1(n2837), .A2(REG2_REG_8__SCAN_IN), .ZN(n2337) );
  NAND2_X1 U2999 ( .A1(n2335), .A2(n2239), .ZN(n2336) );
  AOI22_X1 U3000 ( .A1(n2482), .A2(REG2_REG_9__SCAN_IN), .B1(n2338), .B2(n4469), .ZN(n4355) );
  NAND2_X1 U3001 ( .A1(n2490), .A2(n2339), .ZN(n2340) );
  NAND2_X1 U3002 ( .A1(n2340), .A2(n4363), .ZN(n4373) );
  INV_X1 U3003 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2341) );
  AOI22_X1 U3004 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4464), .B1(n4377), .B2(
        n2341), .ZN(n4374) );
  NAND2_X1 U3005 ( .A1(n4373), .A2(n4374), .ZN(n4372) );
  NAND2_X1 U3006 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4464), .ZN(n2342) );
  NAND2_X1 U3007 ( .A1(n2509), .A2(n2344), .ZN(n2345) );
  INV_X1 U3008 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3254) );
  NOR2_X1 U3009 ( .A1(n3264), .A2(n3254), .ZN(n3253) );
  NOR2_X1 U3010 ( .A1(n4462), .A2(n2346), .ZN(n2347) );
  INV_X1 U3011 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4392) );
  XOR2_X1 U3012 ( .A(n4395), .B(n2346), .Z(n4391) );
  NOR2_X1 U3013 ( .A1(n4392), .A2(n4391), .ZN(n4390) );
  NOR2_X1 U3014 ( .A1(n2347), .A2(n4390), .ZN(n4407) );
  INV_X1 U3015 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2348) );
  AOI22_X1 U3016 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4461), .B1(n2349), .B2(
        n2348), .ZN(n4408) );
  NOR2_X1 U3017 ( .A1(n4407), .A2(n4408), .ZN(n4406) );
  NAND2_X1 U3018 ( .A1(n2350), .A2(n4459), .ZN(n2351) );
  INV_X1 U3019 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U3020 ( .A1(n4430), .A2(n4429), .ZN(n4428) );
  AOI21_X1 U3021 ( .B1(n2354), .B2(n2353), .A(n2365), .ZN(n2355) );
  NAND2_X1 U3022 ( .A1(n4432), .A2(n2355), .ZN(n2362) );
  INV_X1 U3023 ( .A(n2356), .ZN(n2358) );
  NOR2_X2 U3024 ( .A1(n2358), .A2(n2357), .ZN(n4424) );
  AND2_X1 U3025 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3787) );
  AOI21_X1 U3026 ( .B1(n4424), .B2(ADDR_REG_18__SCAN_IN), .A(n3787), .ZN(n2359) );
  OAI21_X1 U3027 ( .B1(n4437), .B2(n4457), .A(n2359), .ZN(n2360) );
  INV_X1 U3028 ( .A(n2360), .ZN(n2361) );
  NAND2_X1 U3029 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
  INV_X1 U3030 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3031 ( .A1(n2368), .A2(n2367), .ZN(n2646) );
  OR2_X1 U3032 ( .A1(n2368), .A2(n2367), .ZN(n2369) );
  MUX2_X1 U3033 ( .A(n2370), .B(REG2_REG_19__SCAN_IN), .S(n3986), .Z(n2371) );
  INV_X1 U3034 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2564) );
  NOR2_X1 U3035 ( .A1(n2564), .A2(STATE_REG_SCAN_IN), .ZN(n3629) );
  AOI21_X1 U3036 ( .B1(n4424), .B2(ADDR_REG_19__SCAN_IN), .A(n3629), .ZN(n2372) );
  OAI21_X1 U3037 ( .B1(n4437), .B2(n3986), .A(n2372), .ZN(n2373) );
  AOI21_X1 U3038 ( .B1(n2374), .B2(n4432), .A(n2373), .ZN(n2378) );
  INV_X1 U3039 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4266) );
  XNOR2_X1 U3040 ( .A(n3986), .B(n4266), .ZN(n2376) );
  NAND2_X1 U3041 ( .A1(n2378), .A2(n2377), .ZN(U3259) );
  NOR2_X2 U3042 ( .A1(n2295), .A2(n2382), .ZN(n2385) );
  INV_X1 U3043 ( .A(IR_REG_29__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U3044 ( .A1(n2385), .A2(n2383), .ZN(n2736) );
  OR2_X1 U3045 ( .A1(n2420), .A2(n4512), .ZN(n2388) );
  INV_X1 U3046 ( .A(n2392), .ZN(n2389) );
  NAND2_X1 U3047 ( .A1(n2417), .A2(REG2_REG_1__SCAN_IN), .ZN(n2387) );
  AND2_X1 U3048 ( .A1(n2388), .A2(n2387), .ZN(n2396) );
  INV_X1 U3049 ( .A(n2419), .ZN(n2393) );
  NAND2_X1 U3050 ( .A1(n2393), .A2(REG3_REG_1__SCAN_IN), .ZN(n2394) );
  NAND3_X2 U3051 ( .A1(n2396), .A2(n2395), .A3(n2394), .ZN(n2407) );
  INV_X1 U3052 ( .A(DATAI_1_), .ZN(n2397) );
  NAND2_X1 U3053 ( .A1(n2407), .A2(n2997), .ZN(n3845) );
  NAND2_X1 U3054 ( .A1(n2661), .A2(n3845), .ZN(n2660) );
  NAND2_X1 U3055 ( .A1(n2652), .A2(REG0_REG_0__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3056 ( .A1(n2417), .A2(REG2_REG_0__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3057 ( .A1(n2393), .A2(REG3_REG_0__SCAN_IN), .ZN(n2402) );
  INV_X1 U3058 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4012) );
  OR2_X1 U3059 ( .A1(n2420), .A2(n4012), .ZN(n2401) );
  NAND2_X1 U3060 ( .A1(n2660), .A2(n2991), .ZN(n2990) );
  NAND2_X1 U3061 ( .A1(n2407), .A2(n2399), .ZN(n2408) );
  NAND2_X1 U3062 ( .A1(n2652), .A2(REG0_REG_2__SCAN_IN), .ZN(n2413) );
  INV_X1 U3063 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2928) );
  OR2_X1 U3064 ( .A1(n2420), .A2(n2928), .ZN(n2412) );
  INV_X1 U3065 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3066 ( .A1(n2417), .A2(REG2_REG_2__SCAN_IN), .ZN(n2410) );
  INV_X1 U3067 ( .A(DATAI_2_), .ZN(n2415) );
  MUX2_X1 U3068 ( .A(n2415), .B(n4028), .S(n2414), .Z(n2921) );
  NAND2_X1 U3069 ( .A1(n3609), .A2(n2921), .ZN(n3851) );
  INV_X1 U3070 ( .A(n3609), .ZN(n3078) );
  NAND2_X1 U3071 ( .A1(n3078), .A2(n2921), .ZN(n2416) );
  NAND2_X1 U3072 ( .A1(n3838), .A2(REG0_REG_3__SCAN_IN), .ZN(n2425) );
  NAND2_X1 U3073 ( .A1(n2418), .A2(REG2_REG_3__SCAN_IN), .ZN(n2424) );
  OR2_X1 U3074 ( .A1(n2651), .A2(REG3_REG_3__SCAN_IN), .ZN(n2423) );
  INV_X1 U3075 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2421) );
  OR2_X1 U3076 ( .A1(n2420), .A2(n2421), .ZN(n2422) );
  MUX2_X1 U3077 ( .A(DATAI_3_), .B(n4339), .S(n2004), .Z(n3610) );
  NAND2_X1 U3078 ( .A1(n4006), .A2(n3610), .ZN(n2426) );
  INV_X1 U3079 ( .A(n4006), .ZN(n2898) );
  NAND2_X1 U3080 ( .A1(n2898), .A2(n3083), .ZN(n2427) );
  INV_X1 U3081 ( .A(n3022), .ZN(n2434) );
  NAND2_X1 U3082 ( .A1(n2418), .A2(REG2_REG_4__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U3083 ( .A1(n3838), .A2(REG0_REG_4__SCAN_IN), .ZN(n2431) );
  OAI21_X1 U3084 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2437), .ZN(n3722) );
  OR2_X1 U3085 ( .A1(n2651), .A2(n3722), .ZN(n2430) );
  INV_X1 U3086 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2428) );
  OR2_X1 U3087 ( .A1(n2420), .A2(n2428), .ZN(n2429) );
  INV_X1 U3088 ( .A(DATAI_4_), .ZN(n2433) );
  MUX2_X1 U3089 ( .A(n2433), .B(n2812), .S(n2611), .Z(n3031) );
  NAND2_X1 U3090 ( .A1(n4005), .A2(n3031), .ZN(n3856) );
  NAND2_X1 U3091 ( .A1(n3854), .A2(n3856), .ZN(n3932) );
  NAND2_X1 U3092 ( .A1(n4005), .A2(n3721), .ZN(n2435) );
  NAND2_X1 U3093 ( .A1(n3838), .A2(REG0_REG_5__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U3094 ( .A1(n2418), .A2(REG2_REG_5__SCAN_IN), .ZN(n2441) );
  OR2_X1 U3095 ( .A1(n3842), .A2(n2436), .ZN(n2440) );
  AND2_X1 U3096 ( .A1(n2437), .A2(n2789), .ZN(n2438) );
  OR2_X1 U3097 ( .A1(n2438), .A2(n2446), .ZN(n3070) );
  OR2_X1 U3098 ( .A1(n2651), .A2(n3070), .ZN(n2439) );
  INV_X1 U3099 ( .A(n3801), .ZN(n3010) );
  INV_X1 U3100 ( .A(DATAI_5_), .ZN(n2443) );
  MUX2_X1 U3101 ( .A(n2443), .B(n2795), .S(n2611), .Z(n2965) );
  NAND2_X1 U3102 ( .A1(n3010), .A2(n2965), .ZN(n2444) );
  NAND2_X1 U3103 ( .A1(n3801), .A2(n3066), .ZN(n2445) );
  NAND2_X1 U3104 ( .A1(n2418), .A2(REG2_REG_6__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3105 ( .A1(n3838), .A2(REG0_REG_6__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3106 ( .A1(n2446), .A2(REG3_REG_6__SCAN_IN), .ZN(n2447) );
  NAND2_X1 U3107 ( .A1(n2455), .A2(n2447), .ZN(n3036) );
  OR2_X1 U3108 ( .A1(n2651), .A2(n3036), .ZN(n2450) );
  INV_X1 U3109 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2448) );
  OR2_X1 U3110 ( .A1(n2420), .A2(n2448), .ZN(n2449) );
  NAND4_X1 U3111 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n3557)
         );
  MUX2_X1 U3112 ( .A(DATAI_6_), .B(n4337), .S(n2611), .Z(n3802) );
  AND2_X1 U3113 ( .A1(n3557), .A2(n3802), .ZN(n2453) );
  OAI22_X1 U3114 ( .A1(n3006), .A2(n2453), .B1(n3802), .B2(n3557), .ZN(n2984)
         );
  INV_X1 U3115 ( .A(n2984), .ZN(n2463) );
  NAND2_X1 U3116 ( .A1(n2418), .A2(REG2_REG_7__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3117 ( .A1(n3838), .A2(REG0_REG_7__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3118 ( .A1(n2455), .A2(n2454), .ZN(n2456) );
  NAND2_X1 U3119 ( .A1(n2465), .A2(n2456), .ZN(n3559) );
  OR2_X1 U3120 ( .A1(n2651), .A2(n3559), .ZN(n2459) );
  OR2_X1 U3121 ( .A1(n2420), .A2(n2457), .ZN(n2458) );
  INV_X1 U3122 ( .A(DATAI_7_), .ZN(n4526) );
  MUX2_X1 U3123 ( .A(n4526), .B(n4335), .S(n2611), .Z(n3376) );
  NAND2_X1 U3124 ( .A1(n4004), .A2(n3376), .ZN(n3865) );
  NAND2_X1 U3125 ( .A1(n2463), .A2(n2985), .ZN(n2983) );
  INV_X1 U3126 ( .A(n3376), .ZN(n3558) );
  NAND2_X1 U3127 ( .A1(n4004), .A2(n3558), .ZN(n2464) );
  NAND2_X1 U3128 ( .A1(n3838), .A2(REG0_REG_8__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3129 ( .A1(n2418), .A2(REG2_REG_8__SCAN_IN), .ZN(n2469) );
  OR2_X1 U3130 ( .A1(n3842), .A2(n3122), .ZN(n2468) );
  NAND2_X1 U3131 ( .A1(n2465), .A2(n4657), .ZN(n2466) );
  NAND2_X1 U3132 ( .A1(n2475), .A2(n2466), .ZN(n3107) );
  OR2_X1 U3133 ( .A1(n2651), .A2(n3107), .ZN(n2467) );
  NAND4_X1 U3134 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n4003)
         );
  INV_X1 U3135 ( .A(n4003), .ZN(n2472) );
  INV_X1 U3136 ( .A(DATAI_8_), .ZN(n2471) );
  MUX2_X1 U3137 ( .A(n2471), .B(n2838), .S(n2611), .Z(n3115) );
  NAND2_X1 U3138 ( .A1(n2472), .A2(n3115), .ZN(n2473) );
  NAND2_X1 U3139 ( .A1(n4003), .A2(n3640), .ZN(n2474) );
  NAND2_X1 U3140 ( .A1(n2418), .A2(REG2_REG_9__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3141 ( .A1(n3838), .A2(REG0_REG_9__SCAN_IN), .ZN(n2480) );
  INV_X1 U3142 ( .A(n2484), .ZN(n2477) );
  NAND2_X1 U3143 ( .A1(n2475), .A2(n3731), .ZN(n2476) );
  NAND2_X1 U3144 ( .A1(n2477), .A2(n2476), .ZN(n3733) );
  OR2_X1 U3145 ( .A1(n2651), .A2(n3733), .ZN(n2479) );
  OR2_X1 U3146 ( .A1(n3842), .A2(n4644), .ZN(n2478) );
  NAND4_X1 U3147 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n3641)
         );
  MUX2_X1 U31480 ( .A(DATAI_9_), .B(n2482), .S(n2611), .Z(n3732) );
  AND2_X1 U31490 ( .A1(n3641), .A2(n3732), .ZN(n2483) );
  INV_X1 U3150 ( .A(n3641), .ZN(n3116) );
  INV_X1 U3151 ( .A(n3732), .ZN(n3050) );
  NAND2_X1 U3152 ( .A1(n3838), .A2(REG0_REG_10__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3153 ( .A1(n2418), .A2(REG2_REG_10__SCAN_IN), .ZN(n2488) );
  OR2_X1 U3154 ( .A1(n3842), .A2(n4360), .ZN(n2487) );
  OR2_X1 U3155 ( .A1(n2484), .A2(REG3_REG_10__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U3156 ( .A1(n2493), .A2(n2485), .ZN(n3095) );
  OR2_X1 U3157 ( .A1(n2651), .A2(n3095), .ZN(n2486) );
  NAND4_X1 U3158 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n4002)
         );
  MUX2_X1 U3159 ( .A(DATAI_10_), .B(n2490), .S(n2611), .Z(n3599) );
  NOR2_X1 U3160 ( .A1(n4002), .A2(n3599), .ZN(n2492) );
  INV_X1 U3161 ( .A(n4002), .ZN(n3150) );
  OAI21_X1 U3162 ( .B1(n3099), .B2(n2492), .A(n2491), .ZN(n3144) );
  NAND2_X1 U3163 ( .A1(n3838), .A2(REG0_REG_11__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3164 ( .A1(n2418), .A2(REG2_REG_11__SCAN_IN), .ZN(n2497) );
  OR2_X1 U3165 ( .A1(n3842), .A2(n4576), .ZN(n2496) );
  NAND2_X1 U3166 ( .A1(n2493), .A2(n3775), .ZN(n2494) );
  NAND2_X1 U3167 ( .A1(n2502), .A2(n2494), .ZN(n3156) );
  OR2_X1 U3168 ( .A1(n2651), .A2(n3156), .ZN(n2495) );
  NAND4_X1 U3169 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n4001)
         );
  INV_X1 U3170 ( .A(DATAI_11_), .ZN(n2499) );
  MUX2_X1 U3171 ( .A(n2499), .B(n4377), .S(n2611), .Z(n3153) );
  OR2_X1 U3172 ( .A1(n4001), .A2(n3153), .ZN(n3167) );
  NAND2_X1 U3173 ( .A1(n4001), .A2(n3153), .ZN(n3170) );
  NAND2_X1 U3174 ( .A1(n3167), .A2(n3170), .ZN(n3928) );
  INV_X1 U3175 ( .A(n4001), .ZN(n3212) );
  NAND2_X1 U3176 ( .A1(n3212), .A2(n3153), .ZN(n2500) );
  NAND2_X1 U3177 ( .A1(n2418), .A2(REG2_REG_12__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3178 ( .A1(n3838), .A2(REG0_REG_12__SCAN_IN), .ZN(n2507) );
  INV_X1 U3179 ( .A(n2512), .ZN(n2504) );
  NAND2_X1 U3180 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  NAND2_X1 U3181 ( .A1(n2504), .A2(n2503), .ZN(n3666) );
  OR2_X1 U3182 ( .A1(n2651), .A2(n3666), .ZN(n2506) );
  OR2_X1 U3183 ( .A1(n3842), .A2(n4380), .ZN(n2505) );
  NAND4_X1 U3184 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3776)
         );
  MUX2_X1 U3185 ( .A(DATAI_12_), .B(n2509), .S(n2611), .Z(n3664) );
  NAND2_X1 U3186 ( .A1(n3776), .A2(n3664), .ZN(n2511) );
  NOR2_X1 U3187 ( .A1(n3776), .A2(n3664), .ZN(n2510) );
  NAND2_X1 U3188 ( .A1(n2418), .A2(REG2_REG_13__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3189 ( .A1(n3838), .A2(REG0_REG_13__SCAN_IN), .ZN(n2516) );
  NOR2_X1 U3190 ( .A1(n2512), .A2(REG3_REG_13__SCAN_IN), .ZN(n2513) );
  OR2_X1 U3191 ( .A1(n2521), .A2(n2513), .ZN(n3757) );
  OR2_X1 U3192 ( .A1(n2651), .A2(n3757), .ZN(n2515) );
  OR2_X1 U3193 ( .A1(n3842), .A2(n3268), .ZN(n2514) );
  INV_X1 U3194 ( .A(n3665), .ZN(n2519) );
  INV_X1 U3195 ( .A(DATAI_13_), .ZN(n2518) );
  MUX2_X1 U3196 ( .A(n2518), .B(n3264), .S(n2611), .Z(n3427) );
  NAND2_X1 U3197 ( .A1(n3838), .A2(REG0_REG_14__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U3198 ( .A1(n2418), .A2(REG2_REG_14__SCAN_IN), .ZN(n2525) );
  OR2_X1 U3199 ( .A1(n3842), .A2(n4388), .ZN(n2524) );
  OR2_X1 U3200 ( .A1(n2521), .A2(REG3_REG_14__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3201 ( .A1(n2530), .A2(n2522), .ZN(n3179) );
  OR2_X1 U3202 ( .A1(n2651), .A2(n3179), .ZN(n2523) );
  NAND4_X1 U3203 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n4291)
         );
  INV_X1 U3204 ( .A(DATAI_14_), .ZN(n2527) );
  MUX2_X1 U3205 ( .A(n2527), .B(n4462), .S(n2611), .Z(n3230) );
  OR2_X1 U3206 ( .A1(n4291), .A2(n3230), .ZN(n3889) );
  NAND2_X1 U3207 ( .A1(n4291), .A2(n3230), .ZN(n3869) );
  NAND2_X1 U3208 ( .A1(n3889), .A2(n3869), .ZN(n3929) );
  NAND2_X1 U3209 ( .A1(n3176), .A2(n2529), .ZN(n3241) );
  NAND2_X1 U32100 ( .A1(n2418), .A2(REG2_REG_15__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32110 ( .A1(n3838), .A2(REG0_REG_15__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32120 ( .A1(n2530), .A2(n4617), .ZN(n2531) );
  NAND2_X1 U32130 ( .A1(n2541), .A2(n2531), .ZN(n3246) );
  OR2_X1 U32140 ( .A1(n2651), .A2(n3246), .ZN(n2534) );
  OR2_X1 U32150 ( .A1(n3842), .A2(n2532), .ZN(n2533) );
  INV_X1 U32160 ( .A(DATAI_15_), .ZN(n4460) );
  MUX2_X1 U32170 ( .A(n4460), .B(n4461), .S(n2611), .Z(n4284) );
  NAND2_X1 U32180 ( .A1(n3241), .A2(n2537), .ZN(n2539) );
  INV_X1 U32190 ( .A(n4284), .ZN(n3826) );
  NAND2_X1 U32200 ( .A1(n2539), .A2(n2538), .ZN(n3273) );
  NAND2_X1 U32210 ( .A1(n2418), .A2(REG2_REG_16__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32220 ( .A1(n3838), .A2(REG0_REG_16__SCAN_IN), .ZN(n2545) );
  AND2_X1 U32230 ( .A1(n2541), .A2(n2540), .ZN(n2542) );
  OR2_X1 U32240 ( .A1(n2542), .A2(n2549), .ZN(n3278) );
  OR2_X1 U32250 ( .A1(n2651), .A2(n3278), .ZN(n2544) );
  OR2_X1 U32260 ( .A1(n3842), .A2(n4414), .ZN(n2543) );
  INV_X1 U32270 ( .A(n3999), .ZN(n4287) );
  INV_X1 U32280 ( .A(n4459), .ZN(n2547) );
  MUX2_X1 U32290 ( .A(DATAI_16_), .B(n2547), .S(n2611), .Z(n4272) );
  NAND2_X1 U32300 ( .A1(n4287), .A2(n4272), .ZN(n3958) );
  NAND2_X1 U32310 ( .A1(n3999), .A2(n2041), .ZN(n3956) );
  NOR2_X1 U32320 ( .A1(n3273), .A2(n3920), .ZN(n3274) );
  NOR2_X1 U32330 ( .A1(n3274), .A2(n2548), .ZN(n3286) );
  NAND2_X1 U32340 ( .A1(n3838), .A2(REG0_REG_17__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U32350 ( .A1(n2418), .A2(REG2_REG_17__SCAN_IN), .ZN(n2553) );
  OR2_X1 U32360 ( .A1(n3842), .A2(n4645), .ZN(n2552) );
  OR2_X1 U32370 ( .A1(n2549), .A2(REG3_REG_17__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32380 ( .A1(n2557), .A2(n2550), .ZN(n3292) );
  OR2_X1 U32390 ( .A1(n2651), .A2(n3292), .ZN(n2551) );
  INV_X1 U32400 ( .A(n4275), .ZN(n3312) );
  INV_X1 U32410 ( .A(DATAI_17_), .ZN(n2555) );
  MUX2_X1 U32420 ( .A(n2555), .B(n4458), .S(n2611), .Z(n3454) );
  NAND2_X1 U32430 ( .A1(n3838), .A2(REG0_REG_18__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32440 ( .A1(n2418), .A2(REG2_REG_18__SCAN_IN), .ZN(n2561) );
  OR2_X1 U32450 ( .A1(n3842), .A2(n2556), .ZN(n2560) );
  NAND2_X1 U32460 ( .A1(n2557), .A2(n4619), .ZN(n2558) );
  NAND2_X1 U32470 ( .A1(n2565), .A2(n2558), .ZN(n3789) );
  OR2_X1 U32480 ( .A1(n2651), .A2(n3789), .ZN(n2559) );
  NAND4_X1 U32490 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), .ZN(n3998)
         );
  INV_X1 U32500 ( .A(n3998), .ZN(n3627) );
  MUX2_X1 U32510 ( .A(DATAI_18_), .B(n2563), .S(n2611), .Z(n3788) );
  NAND2_X1 U32520 ( .A1(n3627), .A2(n3788), .ZN(n3324) );
  INV_X1 U32530 ( .A(n3788), .ZN(n2719) );
  NAND2_X1 U32540 ( .A1(n3998), .A2(n2719), .ZN(n3325) );
  NAND2_X1 U32550 ( .A1(n3324), .A2(n3325), .ZN(n3930) );
  NAND2_X1 U32560 ( .A1(n2565), .A2(n2564), .ZN(n2566) );
  NAND2_X1 U32570 ( .A1(n2572), .A2(n2566), .ZN(n3632) );
  INV_X1 U32580 ( .A(n3632), .ZN(n2567) );
  NAND2_X1 U32590 ( .A1(n2567), .A2(n2393), .ZN(n2571) );
  NAND2_X1 U32600 ( .A1(n2418), .A2(REG2_REG_19__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U32610 ( .A1(n3838), .A2(REG0_REG_19__SCAN_IN), .ZN(n2569) );
  OR2_X1 U32620 ( .A1(n3842), .A2(n4266), .ZN(n2568) );
  INV_X1 U32630 ( .A(n3986), .ZN(n4444) );
  MUX2_X1 U32640 ( .A(DATAI_19_), .B(n4444), .S(n2611), .Z(n3466) );
  NOR2_X1 U32650 ( .A1(n4179), .A2(n3466), .ZN(n3322) );
  NAND2_X1 U32660 ( .A1(n4179), .A2(n3466), .ZN(n3321) );
  INV_X1 U32670 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4578) );
  INV_X1 U32680 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3746) );
  AND2_X1 U32690 ( .A1(n2572), .A2(n3746), .ZN(n2573) );
  NOR2_X1 U32700 ( .A1(n2577), .A2(n2573), .ZN(n4183) );
  NAND2_X1 U32710 ( .A1(n4183), .A2(n2393), .ZN(n2575) );
  AOI22_X1 U32720 ( .A1(n2418), .A2(REG2_REG_20__SCAN_IN), .B1(n3838), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2574) );
  OAI211_X1 U32730 ( .C1(n3842), .C2(n4578), .A(n2575), .B(n2574), .ZN(n4246)
         );
  INV_X1 U32740 ( .A(DATAI_20_), .ZN(n2576) );
  AND2_X1 U32750 ( .A1(n4246), .A2(n3743), .ZN(n3939) );
  OR2_X1 U32760 ( .A1(n4246), .A2(n3743), .ZN(n3940) );
  OR2_X1 U32770 ( .A1(n2577), .A2(REG3_REG_21__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32780 ( .A1(n2584), .A2(n2578), .ZN(n3655) );
  AOI22_X1 U32790 ( .A1(n2418), .A2(REG2_REG_21__SCAN_IN), .B1(n3838), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2580) );
  INV_X1 U32800 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4581) );
  OR2_X1 U32810 ( .A1(n3842), .A2(n4581), .ZN(n2579) );
  OAI211_X1 U32820 ( .C1(n3655), .C2(n2651), .A(n2580), .B(n2579), .ZN(n4257)
         );
  NAND2_X1 U32830 ( .A1(n3906), .A2(DATAI_21_), .ZN(n2685) );
  NAND2_X1 U32840 ( .A1(n4257), .A2(n4245), .ZN(n2582) );
  INV_X1 U32850 ( .A(n4257), .ZN(n2581) );
  INV_X1 U32860 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U32870 ( .A1(n2584), .A2(n2583), .ZN(n2585) );
  AND2_X1 U32880 ( .A1(n2595), .A2(n2585), .ZN(n4161) );
  NAND2_X1 U32890 ( .A1(n4161), .A2(n2393), .ZN(n2591) );
  INV_X1 U32900 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U32910 ( .A1(n3838), .A2(REG0_REG_22__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U32920 ( .A1(n2418), .A2(REG2_REG_22__SCAN_IN), .ZN(n2586) );
  OAI211_X1 U32930 ( .C1(n3842), .C2(n2588), .A(n2587), .B(n2586), .ZN(n2589)
         );
  INV_X1 U32940 ( .A(n2589), .ZN(n2590) );
  INV_X1 U32950 ( .A(DATAI_22_), .ZN(n2592) );
  NOR2_X1 U32960 ( .A1(n2611), .A2(n2592), .ZN(n4155) );
  NAND2_X1 U32970 ( .A1(n4248), .A2(n4155), .ZN(n4135) );
  NAND2_X1 U32980 ( .A1(n3997), .A2(n4162), .ZN(n2683) );
  NAND2_X1 U32990 ( .A1(n4135), .A2(n2683), .ZN(n4153) );
  INV_X1 U33000 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2594) );
  AND2_X1 U33010 ( .A1(n2595), .A2(n2594), .ZN(n2596) );
  OR2_X1 U33020 ( .A1(n2596), .A2(n2603), .ZN(n4146) );
  INV_X1 U33030 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U33040 ( .A1(n2418), .A2(REG2_REG_23__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33050 ( .A1(n3838), .A2(REG0_REG_23__SCAN_IN), .ZN(n2597) );
  OAI211_X1 U33060 ( .C1(n4238), .C2(n3842), .A(n2598), .B(n2597), .ZN(n2599)
         );
  INV_X1 U33070 ( .A(n2599), .ZN(n2600) );
  INV_X1 U33080 ( .A(n4228), .ZN(n4125) );
  NAND2_X1 U33090 ( .A1(n3906), .A2(DATAI_23_), .ZN(n4143) );
  NAND2_X1 U33100 ( .A1(n4125), .A2(n4143), .ZN(n2602) );
  INV_X1 U33110 ( .A(n4143), .ZN(n3488) );
  AOI21_X1 U33120 ( .B1(n4130), .B2(n2602), .A(n2601), .ZN(n4116) );
  NAND2_X1 U33130 ( .A1(n2603), .A2(REG3_REG_24__SCAN_IN), .ZN(n2614) );
  OR2_X1 U33140 ( .A1(n2603), .A2(REG3_REG_24__SCAN_IN), .ZN(n2604) );
  AND2_X1 U33150 ( .A1(n2614), .A2(n2604), .ZN(n4121) );
  NAND2_X1 U33160 ( .A1(n4121), .A2(n2393), .ZN(n2609) );
  INV_X1 U33170 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U33180 ( .A1(n2418), .A2(REG2_REG_24__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U33190 ( .A1(n3838), .A2(REG0_REG_24__SCAN_IN), .ZN(n2605) );
  OAI211_X1 U33200 ( .C1(n4234), .C2(n3842), .A(n2606), .B(n2605), .ZN(n2607)
         );
  INV_X1 U33210 ( .A(n2607), .ZN(n2608) );
  INV_X1 U33220 ( .A(DATAI_24_), .ZN(n2610) );
  NAND2_X1 U33230 ( .A1(n4139), .A2(n4227), .ZN(n2613) );
  NOR2_X1 U33240 ( .A1(n4139), .A2(n4227), .ZN(n2612) );
  AOI21_X1 U33250 ( .B1(n4116), .B2(n2613), .A(n2612), .ZN(n4092) );
  INV_X1 U33260 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U33270 ( .A1(n2614), .A2(n4623), .ZN(n2615) );
  NAND2_X1 U33280 ( .A1(n4107), .A2(n2393), .ZN(n2620) );
  INV_X1 U33290 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4225) );
  NAND2_X1 U33300 ( .A1(n2418), .A2(REG2_REG_25__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33310 ( .A1(n3838), .A2(REG0_REG_25__SCAN_IN), .ZN(n2616) );
  OAI211_X1 U33320 ( .C1(n4225), .C2(n3842), .A(n2617), .B(n2616), .ZN(n2618)
         );
  INV_X1 U33330 ( .A(n2618), .ZN(n2619) );
  NAND2_X1 U33340 ( .A1(n3906), .A2(DATAI_25_), .ZN(n4099) );
  NAND2_X1 U33350 ( .A1(n4092), .A2(n2032), .ZN(n2622) );
  INV_X1 U33360 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2623) );
  AND2_X1 U33370 ( .A1(n2011), .A2(n2623), .ZN(n2624) );
  INV_X1 U33380 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4580) );
  NAND2_X1 U33390 ( .A1(n2418), .A2(REG2_REG_26__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U33400 ( .A1(n3838), .A2(REG0_REG_26__SCAN_IN), .ZN(n2625) );
  OAI211_X1 U33410 ( .C1(n4580), .C2(n3842), .A(n2626), .B(n2625), .ZN(n2627)
         );
  INV_X1 U33420 ( .A(n2627), .ZN(n2628) );
  INV_X1 U33430 ( .A(n4211), .ZN(n3679) );
  NAND2_X1 U33440 ( .A1(n3906), .A2(DATAI_26_), .ZN(n4078) );
  NOR2_X1 U33450 ( .A1(n3679), .A2(n4078), .ZN(n2630) );
  NAND2_X1 U33460 ( .A1(n3679), .A2(n4078), .ZN(n2629) );
  INV_X1 U33470 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U33480 ( .A1(n2418), .A2(REG2_REG_27__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U33490 ( .A1(n3838), .A2(REG0_REG_27__SCAN_IN), .ZN(n2632) );
  OAI211_X1 U33500 ( .C1(n2634), .C2(n3842), .A(n2633), .B(n2632), .ZN(n2635)
         );
  INV_X1 U33510 ( .A(n2635), .ZN(n2636) );
  NAND2_X1 U33520 ( .A1(n3906), .A2(DATAI_27_), .ZN(n4062) );
  INV_X1 U3353 ( .A(n4062), .ZN(n4210) );
  INV_X1 U33540 ( .A(n4080), .ZN(n3525) );
  NAND2_X1 U3355 ( .A1(n2637), .A2(REG3_REG_28__SCAN_IN), .ZN(n4035) );
  OR2_X1 U3356 ( .A1(n2637), .A2(REG3_REG_28__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3357 ( .A1(n3542), .A2(n2393), .ZN(n2644) );
  INV_X1 U3358 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3359 ( .A1(n2418), .A2(REG2_REG_28__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3360 ( .A1(n3838), .A2(REG0_REG_28__SCAN_IN), .ZN(n2639) );
  OAI211_X1 U3361 ( .C1(n2641), .C2(n3842), .A(n2640), .B(n2639), .ZN(n2642)
         );
  INV_X1 U3362 ( .A(n2642), .ZN(n2643) );
  NAND2_X1 U3363 ( .A1(n3906), .A2(DATAI_28_), .ZN(n2720) );
  NOR2_X1 U3364 ( .A1(n4212), .A2(n2720), .ZN(n4036) );
  NAND2_X1 U3365 ( .A1(n4212), .A2(n2720), .ZN(n4037) );
  INV_X1 U3366 ( .A(n4037), .ZN(n2645) );
  XNOR2_X1 U3367 ( .A(n2986), .B(n3992), .ZN(n2649) );
  NAND2_X1 U3368 ( .A1(n2649), .A2(n3986), .ZN(n3200) );
  NOR2_X1 U3369 ( .A1(n3986), .A2(n3992), .ZN(n2650) );
  INV_X1 U3370 ( .A(n4487), .ZN(n4479) );
  NAND2_X1 U3371 ( .A1(n3200), .A2(n4479), .ZN(n4502) );
  INV_X1 U3372 ( .A(n2712), .ZN(n2852) );
  OR2_X1 U3373 ( .A1(n4035), .A2(n2651), .ZN(n2658) );
  INV_X1 U3374 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3375 ( .A1(n2418), .A2(REG2_REG_29__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3376 ( .A1(n2652), .A2(REG0_REG_29__SCAN_IN), .ZN(n2653) );
  OAI211_X1 U3377 ( .C1(n2655), .C2(n3842), .A(n2654), .B(n2653), .ZN(n2656)
         );
  INV_X1 U3378 ( .A(n2656), .ZN(n2657) );
  NAND2_X1 U3379 ( .A1(n2658), .A2(n2657), .ZN(n3996) );
  INV_X1 U3380 ( .A(n3996), .ZN(n2659) );
  NAND2_X1 U3381 ( .A1(n4341), .A2(n2712), .ZN(n4286) );
  INV_X1 U3382 ( .A(n2722), .ZN(n3983) );
  OAI22_X1 U3383 ( .A1(n2659), .A2(n4286), .B1(n2720), .B2(n4285), .ZN(n2695)
         );
  INV_X2 U3384 ( .A(n2803), .ZN(n2998) );
  OR2_X1 U3385 ( .A1(n4008), .A2(n2998), .ZN(n3844) );
  OAI21_X1 U3386 ( .B1(n2660), .B2(n3844), .A(n2661), .ZN(n2893) );
  INV_X1 U3387 ( .A(n3926), .ZN(n2894) );
  NAND2_X1 U3388 ( .A1(n2893), .A2(n2894), .ZN(n2892) );
  NAND2_X1 U3389 ( .A1(n2892), .A2(n3848), .ZN(n3076) );
  OR2_X1 U3390 ( .A1(n4006), .A2(n3083), .ZN(n3853) );
  NAND2_X1 U3391 ( .A1(n4006), .A2(n3083), .ZN(n3850) );
  NAND2_X1 U3392 ( .A1(n3853), .A2(n3850), .ZN(n3927) );
  INV_X1 U3393 ( .A(n3927), .ZN(n3075) );
  NAND2_X1 U3394 ( .A1(n3076), .A2(n3075), .ZN(n2662) );
  NAND2_X1 U3395 ( .A1(n2662), .A2(n3853), .ZN(n3025) );
  INV_X1 U3396 ( .A(n3854), .ZN(n2663) );
  OR2_X1 U3397 ( .A1(n3025), .A2(n2663), .ZN(n2664) );
  NAND2_X1 U3398 ( .A1(n2664), .A2(n3856), .ZN(n3061) );
  AND2_X1 U3399 ( .A1(n3801), .A2(n2965), .ZN(n3857) );
  OR2_X1 U3400 ( .A1(n3061), .A2(n3857), .ZN(n2665) );
  OR2_X1 U3401 ( .A1(n3801), .A2(n2965), .ZN(n3874) );
  NAND2_X1 U3402 ( .A1(n3557), .A2(n3039), .ZN(n3007) );
  NOR2_X1 U3403 ( .A1(n3557), .A2(n3039), .ZN(n3860) );
  AOI21_X1 U3404 ( .B1(n3008), .B2(n3007), .A(n3860), .ZN(n2970) );
  NAND2_X1 U3405 ( .A1(n2970), .A2(n3859), .ZN(n2666) );
  NAND2_X1 U3406 ( .A1(n2666), .A2(n3865), .ZN(n3110) );
  OR2_X1 U3407 ( .A1(n4003), .A2(n3115), .ZN(n3866) );
  NAND2_X1 U3408 ( .A1(n3110), .A2(n3866), .ZN(n2667) );
  NAND2_X1 U3409 ( .A1(n4003), .A2(n3115), .ZN(n3864) );
  NAND2_X1 U3410 ( .A1(n2667), .A2(n3864), .ZN(n3047) );
  AND2_X1 U3411 ( .A1(n3641), .A2(n3050), .ZN(n3875) );
  OR2_X1 U3412 ( .A1(n3641), .A2(n3050), .ZN(n3867) );
  NAND2_X1 U3413 ( .A1(n2668), .A2(n3867), .ZN(n3092) );
  NAND2_X1 U3414 ( .A1(n4002), .A2(n3131), .ZN(n3882) );
  NAND2_X1 U3415 ( .A1(n3092), .A2(n3882), .ZN(n2669) );
  OR2_X1 U3416 ( .A1(n4002), .A2(n3131), .ZN(n3878) );
  NAND2_X1 U3417 ( .A1(n2669), .A2(n3878), .ZN(n3169) );
  INV_X1 U3418 ( .A(n3664), .ZN(n2672) );
  NAND2_X1 U3419 ( .A1(n3776), .A2(n2672), .ZN(n3190) );
  NAND2_X1 U3420 ( .A1(n3665), .A2(n3427), .ZN(n3186) );
  NAND2_X1 U3421 ( .A1(n3190), .A2(n3186), .ZN(n2671) );
  INV_X1 U3422 ( .A(n3170), .ZN(n2670) );
  NOR2_X1 U3423 ( .A1(n2671), .A2(n2670), .ZN(n3883) );
  NAND2_X1 U3424 ( .A1(n3169), .A2(n3883), .ZN(n2675) );
  INV_X1 U3425 ( .A(n2671), .ZN(n2674) );
  OR2_X1 U3426 ( .A1(n3776), .A2(n2672), .ZN(n3192) );
  NAND2_X1 U3427 ( .A1(n3167), .A2(n3192), .ZN(n2673) );
  NOR2_X1 U3428 ( .A1(n3665), .A2(n3427), .ZN(n3187) );
  AOI21_X1 U3429 ( .B1(n2674), .B2(n2673), .A(n3187), .ZN(n3892) );
  NAND2_X1 U3430 ( .A1(n2675), .A2(n3892), .ZN(n3955) );
  INV_X1 U3431 ( .A(n3929), .ZN(n2676) );
  NAND2_X1 U3432 ( .A1(n3955), .A2(n2676), .ZN(n2677) );
  NAND2_X1 U3433 ( .A1(n2677), .A2(n3889), .ZN(n3242) );
  OR2_X1 U3434 ( .A1(n4000), .A2(n4284), .ZN(n3888) );
  NAND2_X1 U3435 ( .A1(n4000), .A2(n4284), .ZN(n3870) );
  NAND2_X1 U3436 ( .A1(n3888), .A2(n3870), .ZN(n3921) );
  NAND2_X1 U3437 ( .A1(n3243), .A2(n3870), .ZN(n3282) );
  NAND2_X1 U3438 ( .A1(n3282), .A2(n3920), .ZN(n3281) );
  NAND2_X1 U3439 ( .A1(n3281), .A2(n3956), .ZN(n3309) );
  OR2_X1 U3440 ( .A1(n4257), .A2(n2685), .ZN(n4131) );
  AND2_X1 U3441 ( .A1(n4135), .A2(n4131), .ZN(n3903) );
  NAND2_X1 U3442 ( .A1(n4179), .A2(n3624), .ZN(n2678) );
  AND2_X1 U3443 ( .A1(n2678), .A2(n3325), .ZN(n3345) );
  OR2_X1 U3444 ( .A1(n4275), .A2(n3454), .ZN(n3310) );
  NAND2_X1 U3445 ( .A1(n3324), .A2(n3310), .ZN(n2679) );
  NAND2_X1 U3446 ( .A1(n3345), .A2(n2679), .ZN(n2681) );
  INV_X1 U3447 ( .A(n4179), .ZN(n4255) );
  NAND2_X1 U3448 ( .A1(n4255), .A2(n3466), .ZN(n2680) );
  NAND2_X1 U3449 ( .A1(n2681), .A2(n2680), .ZN(n4170) );
  INV_X1 U3450 ( .A(n3743), .ZN(n4254) );
  NOR2_X1 U3451 ( .A1(n4246), .A2(n4254), .ZN(n2682) );
  NAND2_X1 U3452 ( .A1(n4246), .A2(n4254), .ZN(n3348) );
  OAI21_X1 U3453 ( .B1(n4170), .B2(n2682), .A(n3348), .ZN(n3897) );
  AND2_X1 U3454 ( .A1(n3903), .A2(n3897), .ZN(n3960) );
  NAND2_X1 U3455 ( .A1(n3309), .A2(n3960), .ZN(n2689) );
  NAND2_X1 U3456 ( .A1(n4275), .A2(n3454), .ZN(n3307) );
  NAND3_X1 U3457 ( .A1(n3348), .A2(n3345), .A3(n3307), .ZN(n3895) );
  NAND2_X1 U34580 ( .A1(n3960), .A2(n3895), .ZN(n2688) );
  NAND2_X1 U34590 ( .A1(n4228), .A2(n4143), .ZN(n2684) );
  NAND2_X1 U3460 ( .A1(n2684), .A2(n2683), .ZN(n3901) );
  AND2_X1 U3461 ( .A1(n4257), .A2(n2685), .ZN(n3338) );
  AND2_X1 U3462 ( .A1(n4135), .A2(n3338), .ZN(n2686) );
  NOR2_X1 U3463 ( .A1(n3901), .A2(n2686), .ZN(n2687) );
  AND2_X1 U3464 ( .A1(n2688), .A2(n2687), .ZN(n3961) );
  NAND2_X1 U3465 ( .A1(n2689), .A2(n3961), .ZN(n4113) );
  NAND2_X1 U3466 ( .A1(n4100), .A2(n4227), .ZN(n3942) );
  OR2_X1 U34670 ( .A1(n4228), .A2(n4143), .ZN(n4112) );
  AND2_X1 U3468 ( .A1(n3942), .A2(n4112), .ZN(n3964) );
  NAND2_X1 U34690 ( .A1(n4113), .A2(n3964), .ZN(n4094) );
  INV_X1 U3470 ( .A(n4227), .ZN(n3503) );
  NAND2_X1 U34710 ( .A1(n4139), .A2(n3503), .ZN(n4093) );
  NAND2_X1 U3472 ( .A1(n4120), .A2(n4099), .ZN(n3937) );
  AND2_X1 U34730 ( .A1(n4093), .A2(n3937), .ZN(n3971) );
  NAND2_X1 U3474 ( .A1(n4094), .A2(n3971), .ZN(n4075) );
  OR2_X1 U34750 ( .A1(n4211), .A2(n4078), .ZN(n3935) );
  OR2_X1 U3476 ( .A1(n4120), .A2(n4099), .ZN(n4074) );
  AND2_X1 U34770 ( .A1(n3935), .A2(n4074), .ZN(n3969) );
  NAND2_X1 U3478 ( .A1(n4075), .A2(n3969), .ZN(n2690) );
  AND2_X1 U34790 ( .A1(n4211), .A2(n4078), .ZN(n3907) );
  INV_X1 U3480 ( .A(n3907), .ZN(n3936) );
  NAND2_X1 U34810 ( .A1(n2690), .A2(n3936), .ZN(n4060) );
  AND2_X1 U3482 ( .A1(n4080), .A2(n4062), .ZN(n3909) );
  INV_X1 U34830 ( .A(n3909), .ZN(n2691) );
  OR2_X1 U3484 ( .A1(n4080), .A2(n4062), .ZN(n3911) );
  OAI21_X1 U34850 ( .B1(n4060), .B2(n4059), .A(n3911), .ZN(n4038) );
  XNOR2_X1 U3486 ( .A(n4038), .B(n4049), .ZN(n2694) );
  NAND2_X1 U34870 ( .A1(n3983), .A2(n4334), .ZN(n2693) );
  OR2_X1 U3488 ( .A1(n3986), .A2(n2857), .ZN(n2692) );
  NOR2_X1 U34890 ( .A1(n2694), .A2(n4259), .ZN(n3550) );
  AOI211_X1 U3490 ( .C1(n4292), .C2(n4080), .A(n2695), .B(n3550), .ZN(n2696)
         );
  OAI21_X1 U34910 ( .B1(n3552), .B2(n4490), .A(n2696), .ZN(n2726) );
  NAND2_X1 U3492 ( .A1(n2744), .A2(n2697), .ZN(n2698) );
  MUX2_X1 U34930 ( .A(n2697), .B(n2698), .S(B_REG_SCAN_IN), .Z(n2700) );
  NAND2_X1 U3494 ( .A1(n2700), .A2(n2699), .ZN(n2754) );
  NOR4_X1 U34950 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2704) );
  NOR4_X1 U3496 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2703) );
  NOR4_X1 U34970 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2702) );
  NOR4_X1 U3498 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2701) );
  AND4_X1 U34990 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n2710)
         );
  NOR2_X1 U3500 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_8__SCAN_IN), .ZN(n2708) );
  NOR4_X1 U35010 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2707) );
  NOR4_X1 U3502 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2706) );
  NOR4_X1 U35030 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2705) );
  AND4_X1 U3504 ( .A1(n2708), .A2(n2707), .A3(n2706), .A4(n2705), .ZN(n2709)
         );
  NAND2_X1 U35050 ( .A1(n2710), .A2(n2709), .ZN(n2844) );
  NAND2_X1 U35060 ( .A1(n2848), .A2(n2844), .ZN(n2715) );
  INV_X1 U35070 ( .A(n2699), .ZN(n2716) );
  NAND2_X1 U35080 ( .A1(n2716), .A2(n2744), .ZN(n2758) );
  OAI21_X1 U35090 ( .B1(n2754), .B2(D_REG_1__SCAN_IN), .A(n2758), .ZN(n2714)
         );
  NAND2_X1 U35100 ( .A1(n4487), .A2(n2711), .ZN(n2876) );
  NAND2_X1 U35110 ( .A1(n2722), .A2(n3986), .ZN(n2851) );
  NAND2_X1 U35120 ( .A1(n2851), .A2(n2712), .ZN(n2975) );
  AND2_X1 U35130 ( .A1(n2876), .A2(n2975), .ZN(n2713) );
  NAND4_X1 U35140 ( .A1(n2715), .A2(n2714), .A3(n2713), .A4(n2977), .ZN(n2724)
         );
  INV_X1 U35150 ( .A(D_REG_0__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U35160 ( .A1(n2848), .A2(n2757), .ZN(n2717) );
  NAND2_X1 U35170 ( .A1(n2716), .A2(n2697), .ZN(n2755) );
  INV_X1 U35180 ( .A(n2718), .ZN(n2723) );
  NAND2_X1 U35190 ( .A1(n2997), .A2(n2998), .ZN(n2996) );
  INV_X1 U35200 ( .A(n2921), .ZN(n2906) );
  AND2_X2 U35210 ( .A1(n3305), .A2(n2719), .ZN(n3333) );
  OR2_X2 U35220 ( .A1(n3332), .A2(n3743), .ZN(n4177) );
  INV_X1 U35230 ( .A(n4078), .ZN(n4085) );
  NAND2_X1 U35240 ( .A1(n4084), .A2(n4062), .ZN(n4064) );
  INV_X1 U35250 ( .A(n2720), .ZN(n4047) );
  OR2_X2 U35260 ( .A1(n4064), .A2(n4047), .ZN(n4053) );
  NAND2_X1 U35270 ( .A1(n4064), .A2(n4047), .ZN(n2721) );
  NAND2_X1 U35280 ( .A1(n4053), .A2(n2721), .ZN(n3547) );
  NAND2_X1 U35290 ( .A1(n4518), .A2(n4504), .ZN(n4268) );
  NAND2_X1 U35300 ( .A1(n2723), .A2(n2182), .ZN(U3546) );
  INV_X1 U35310 ( .A(n2724), .ZN(n2725) );
  INV_X1 U35320 ( .A(n2727), .ZN(n2728) );
  NAND2_X1 U35330 ( .A1(n4511), .A2(n4504), .ZN(n4329) );
  NAND2_X1 U35340 ( .A1(n2728), .A2(n2180), .ZN(U3514) );
  INV_X1 U35350 ( .A(n4455), .ZN(n2729) );
  INV_X2 U35360 ( .A(n4007), .ZN(U4043) );
  MUX2_X1 U35370 ( .A(n4010), .B(n2397), .S(U3149), .Z(n2730) );
  INV_X1 U35380 ( .A(n2730), .ZN(U3351) );
  MUX2_X1 U35390 ( .A(n2795), .B(n2443), .S(U3149), .Z(n2731) );
  INV_X1 U35400 ( .A(n2731), .ZN(U3347) );
  NAND2_X1 U35410 ( .A1(n2732), .A2(STATE_REG_SCAN_IN), .ZN(n2733) );
  OAI21_X1 U35420 ( .B1(STATE_REG_SCAN_IN), .B2(n2518), .A(n2733), .ZN(U3339)
         );
  NAND2_X1 U35430 ( .A1(n3992), .A2(STATE_REG_SCAN_IN), .ZN(n2734) );
  OAI21_X1 U35440 ( .B1(STATE_REG_SCAN_IN), .B2(n2592), .A(n2734), .ZN(U3330)
         );
  MUX2_X1 U35450 ( .A(n2471), .B(n2838), .S(STATE_REG_SCAN_IN), .Z(n2735) );
  INV_X1 U35460 ( .A(n2735), .ZN(U3344) );
  INV_X1 U35470 ( .A(DATAI_31_), .ZN(n2738) );
  OR4_X1 U35480 ( .A1(n2736), .A2(IR_REG_30__SCAN_IN), .A3(n2225), .A4(U3149), 
        .ZN(n2737) );
  OAI21_X1 U35490 ( .B1(STATE_REG_SCAN_IN), .B2(n2738), .A(n2737), .ZN(U3321)
         );
  INV_X1 U35500 ( .A(DATAI_30_), .ZN(n2740) );
  NAND2_X1 U35510 ( .A1(n2391), .A2(STATE_REG_SCAN_IN), .ZN(n2739) );
  OAI21_X1 U35520 ( .B1(STATE_REG_SCAN_IN), .B2(n2740), .A(n2739), .ZN(U3322)
         );
  MUX2_X1 U35530 ( .A(n4028), .B(n2415), .S(U3149), .Z(n2741) );
  INV_X1 U35540 ( .A(n2741), .ZN(U3350) );
  INV_X1 U35550 ( .A(DATAI_27_), .ZN(n2743) );
  NAND2_X1 U35560 ( .A1(n4040), .A2(STATE_REG_SCAN_IN), .ZN(n2742) );
  OAI21_X1 U35570 ( .B1(STATE_REG_SCAN_IN), .B2(n2743), .A(n2742), .ZN(U3325)
         );
  INV_X1 U35580 ( .A(DATAI_25_), .ZN(n2747) );
  INV_X1 U35590 ( .A(n2744), .ZN(n2745) );
  NAND2_X1 U35600 ( .A1(n2745), .A2(STATE_REG_SCAN_IN), .ZN(n2746) );
  OAI21_X1 U35610 ( .B1(STATE_REG_SCAN_IN), .B2(n2747), .A(n2746), .ZN(U3327)
         );
  MUX2_X1 U35620 ( .A(n2610), .B(n2697), .S(STATE_REG_SCAN_IN), .Z(n2748) );
  INV_X1 U35630 ( .A(n2748), .ZN(U3328) );
  INV_X1 U35640 ( .A(DATAI_26_), .ZN(n2750) );
  NAND2_X1 U35650 ( .A1(n2699), .A2(STATE_REG_SCAN_IN), .ZN(n2749) );
  OAI21_X1 U35660 ( .B1(STATE_REG_SCAN_IN), .B2(n2750), .A(n2749), .ZN(U3326)
         );
  INV_X1 U35670 ( .A(DATAI_19_), .ZN(n2751) );
  MUX2_X1 U35680 ( .A(n3986), .B(n2751), .S(U3149), .Z(n2752) );
  INV_X1 U35690 ( .A(n2752), .ZN(U3333) );
  NAND2_X1 U35700 ( .A1(n3983), .A2(STATE_REG_SCAN_IN), .ZN(n2753) );
  OAI21_X1 U35710 ( .B1(STATE_REG_SCAN_IN), .B2(n2576), .A(n2753), .ZN(U3332)
         );
  INV_X1 U35720 ( .A(n2755), .ZN(n2756) );
  AOI22_X1 U35730 ( .A1(n4634), .A2(n2757), .B1(n2756), .B2(n4455), .ZN(U3458)
         );
  INV_X1 U35740 ( .A(D_REG_1__SCAN_IN), .ZN(n2759) );
  INV_X1 U35750 ( .A(n2758), .ZN(n2846) );
  AOI22_X1 U35760 ( .A1(n4634), .A2(n2759), .B1(n2846), .B2(n4455), .ZN(U3459)
         );
  INV_X1 U35770 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U35780 ( .A1(n4291), .A2(U4043), .ZN(n2760) );
  OAI21_X1 U35790 ( .B1(U4043), .B2(n4613), .A(n2760), .ZN(U3564) );
  INV_X1 U35800 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U35810 ( .A1(n3609), .A2(U4043), .ZN(n2761) );
  OAI21_X1 U3582 ( .B1(U4043), .B2(n4604), .A(n2761), .ZN(U3552) );
  INV_X1 U3583 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U3584 ( .A1(n3557), .A2(U4043), .ZN(n2762) );
  OAI21_X1 U3585 ( .B1(U4043), .B2(n4655), .A(n2762), .ZN(U3556) );
  INV_X1 U3586 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U3587 ( .A1(n3776), .A2(U4043), .ZN(n2763) );
  OAI21_X1 U3588 ( .B1(U4043), .B2(n4607), .A(n2763), .ZN(U3562) );
  INV_X1 U3589 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U3590 ( .A1(n3641), .A2(U4043), .ZN(n2764) );
  OAI21_X1 U3591 ( .B1(U4043), .B2(n4653), .A(n2764), .ZN(U3559) );
  INV_X1 U3592 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U3593 ( .A1(n3665), .A2(U4043), .ZN(n2765) );
  OAI21_X1 U3594 ( .B1(U4043), .B2(n4614), .A(n2765), .ZN(U3563) );
  INV_X1 U3595 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U3596 ( .A1(n3801), .A2(U4043), .ZN(n2766) );
  OAI21_X1 U3597 ( .B1(U4043), .B2(n4654), .A(n2766), .ZN(U3555) );
  NAND2_X1 U3598 ( .A1(n4008), .A2(n2998), .ZN(n3846) );
  NAND2_X1 U3599 ( .A1(n3844), .A2(n3846), .ZN(n4450) );
  INV_X1 U3600 ( .A(n2850), .ZN(n2767) );
  NOR2_X1 U3601 ( .A1(n2998), .A2(n2767), .ZN(n4447) );
  INV_X1 U3602 ( .A(n3200), .ZN(n3147) );
  OAI21_X1 U3603 ( .B1(n3147), .B2(n4159), .A(n4450), .ZN(n2768) );
  OAI21_X1 U3604 ( .B1(n2400), .B2(n4286), .A(n2768), .ZN(n4445) );
  AOI211_X1 U3605 ( .C1(n4487), .C2(n4450), .A(n4447), .B(n4445), .ZN(n4470)
         );
  NAND2_X1 U3606 ( .A1(n4519), .A2(REG1_REG_0__SCAN_IN), .ZN(n2769) );
  OAI21_X1 U3607 ( .B1(n4470), .B2(n4519), .A(n2769), .ZN(U3518) );
  NOR2_X1 U3608 ( .A1(n4424), .A2(U4043), .ZN(U3148) );
  INV_X1 U3609 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2775) );
  INV_X1 U3610 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U3611 ( .A1(n4040), .A2(n4452), .ZN(n2770) );
  AND2_X1 U3612 ( .A1(n2880), .A2(n2770), .ZN(n2809) );
  NOR2_X1 U3613 ( .A1(n4040), .A2(REG1_REG_0__SCAN_IN), .ZN(n2771) );
  OAI21_X1 U3614 ( .B1(IR_REG_0__SCAN_IN), .B2(n2771), .A(n2809), .ZN(n2773)
         );
  OAI211_X1 U3615 ( .C1(n2809), .C2(IR_REG_0__SCAN_IN), .A(n2773), .B(n2772), 
        .ZN(n2774) );
  OAI21_X1 U3616 ( .B1(STATE_REG_SCAN_IN), .B2(n2775), .A(n2774), .ZN(n2777)
         );
  NOR3_X1 U3617 ( .A1(n4400), .A2(REG1_REG_0__SCAN_IN), .A3(n2045), .ZN(n2776)
         );
  AOI211_X1 U3618 ( .C1(n4424), .C2(ADDR_REG_0__SCAN_IN), .A(n2777), .B(n2776), 
        .ZN(n2778) );
  INV_X1 U3619 ( .A(n2778), .ZN(U3240) );
  XOR2_X1 U3620 ( .A(n2779), .B(REG1_REG_3__SCAN_IN), .Z(n2782) );
  XOR2_X1 U3621 ( .A(REG2_REG_3__SCAN_IN), .B(n2780), .Z(n2781) );
  AOI22_X1 U3622 ( .A1(n4434), .A2(n2782), .B1(n4432), .B2(n2781), .ZN(n2784)
         );
  INV_X1 U3623 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3085) );
  NOR2_X1 U3624 ( .A1(STATE_REG_SCAN_IN), .A2(n3085), .ZN(n3608) );
  AOI21_X1 U3625 ( .B1(n4424), .B2(ADDR_REG_3__SCAN_IN), .A(n3608), .ZN(n2783)
         );
  OAI211_X1 U3626 ( .C1(n2785), .C2(n4437), .A(n2784), .B(n2783), .ZN(U3243)
         );
  AOI211_X1 U3627 ( .C1(n2788), .C2(n2787), .A(n4389), .B(n2786), .ZN(n2797)
         );
  NOR2_X1 U3628 ( .A1(n2789), .A2(STATE_REG_SCAN_IN), .ZN(n2967) );
  AOI21_X1 U3629 ( .B1(n4424), .B2(ADDR_REG_5__SCAN_IN), .A(n2967), .ZN(n2794)
         );
  OAI211_X1 U3630 ( .C1(n2792), .C2(n2791), .A(n4434), .B(n2790), .ZN(n2793)
         );
  OAI211_X1 U3631 ( .C1(n4437), .C2(n2795), .A(n2794), .B(n2793), .ZN(n2796)
         );
  OR2_X1 U3632 ( .A1(n2797), .A2(n2796), .ZN(U3245) );
  XOR2_X1 U3633 ( .A(REG2_REG_4__SCAN_IN), .B(n2798), .Z(n2817) );
  NAND2_X1 U3634 ( .A1(n4008), .A2(n2908), .ZN(n2800) );
  NAND2_X1 U3635 ( .A1(n2803), .A2(n2905), .ZN(n2799) );
  NAND2_X1 U3636 ( .A1(n2800), .A2(n2799), .ZN(n2864) );
  NOR2_X1 U3637 ( .A1(n2934), .A2(n4012), .ZN(n2801) );
  OR2_X1 U3638 ( .A1(n2864), .A2(n2801), .ZN(n2863) );
  NAND2_X1 U3639 ( .A1(n4008), .A2(n2005), .ZN(n2805) );
  INV_X1 U3640 ( .A(n2934), .ZN(n2802) );
  AOI22_X1 U3641 ( .A1(n2803), .A2(n2908), .B1(n2802), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2804) );
  NAND2_X1 U3642 ( .A1(n2805), .A2(n2804), .ZN(n2862) );
  XNOR2_X1 U3643 ( .A(n2863), .B(n2862), .ZN(n2932) );
  NAND3_X1 U3644 ( .A1(n2932), .A2(n2880), .A3(n2806), .ZN(n2808) );
  NOR2_X1 U3645 ( .A1(n2045), .A2(n4452), .ZN(n4017) );
  AOI21_X1 U3646 ( .B1(n3990), .B2(n4017), .A(n4007), .ZN(n2807) );
  OAI211_X1 U3647 ( .C1(IR_REG_0__SCAN_IN), .C2(n2809), .A(n2808), .B(n2807), 
        .ZN(n4034) );
  XOR2_X1 U3648 ( .A(n2810), .B(REG1_REG_4__SCAN_IN), .Z(n2815) );
  INV_X1 U3649 ( .A(n4424), .ZN(n2811) );
  INV_X1 U3650 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U3651 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3719) );
  OAI21_X1 U3652 ( .B1(n2811), .B2(n4652), .A(n3719), .ZN(n2814) );
  NOR2_X1 U3653 ( .A1(n4437), .A2(n2812), .ZN(n2813) );
  AOI211_X1 U3654 ( .C1(n4434), .C2(n2815), .A(n2814), .B(n2813), .ZN(n2816)
         );
  OAI211_X1 U3655 ( .C1(n2817), .C2(n4389), .A(n4034), .B(n2816), .ZN(U3244)
         );
  XNOR2_X1 U3656 ( .A(n2818), .B(REG2_REG_6__SCAN_IN), .ZN(n2826) );
  XOR2_X1 U3657 ( .A(n2819), .B(REG1_REG_6__SCAN_IN), .Z(n2824) );
  INV_X1 U3658 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2820) );
  NOR2_X1 U3659 ( .A1(STATE_REG_SCAN_IN), .A2(n2820), .ZN(n3800) );
  AOI21_X1 U3660 ( .B1(n4424), .B2(ADDR_REG_6__SCAN_IN), .A(n3800), .ZN(n2821)
         );
  OAI21_X1 U3661 ( .B1(n4437), .B2(n2822), .A(n2821), .ZN(n2823) );
  AOI21_X1 U3662 ( .B1(n4434), .B2(n2824), .A(n2823), .ZN(n2825) );
  OAI21_X1 U3663 ( .B1(n2826), .B2(n4389), .A(n2825), .ZN(U3246) );
  MUX2_X1 U3664 ( .A(REG1_REG_7__SCAN_IN), .B(n2457), .S(n4335), .Z(n2828) );
  XOR2_X1 U3665 ( .A(n2828), .B(n2827), .Z(n2836) );
  AOI21_X1 U3666 ( .B1(n2830), .B2(n2829), .A(n4389), .ZN(n2834) );
  AND2_X1 U3667 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3556) );
  AOI21_X1 U3668 ( .B1(n4424), .B2(ADDR_REG_7__SCAN_IN), .A(n3556), .ZN(n2831)
         );
  OAI21_X1 U3669 ( .B1(n4437), .B2(n4335), .A(n2831), .ZN(n2832) );
  AOI21_X1 U3670 ( .B1(n2834), .B2(n2833), .A(n2832), .ZN(n2835) );
  OAI21_X1 U3671 ( .B1(n4400), .B2(n2836), .A(n2835), .ZN(U3247) );
  XNOR2_X1 U3672 ( .A(n2837), .B(REG2_REG_8__SCAN_IN), .ZN(n2843) );
  AND2_X1 U3673 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3639) );
  NOR2_X1 U3674 ( .A1(n4437), .A2(n2838), .ZN(n2839) );
  AOI211_X1 U3675 ( .C1(n4424), .C2(ADDR_REG_8__SCAN_IN), .A(n3639), .B(n2839), 
        .ZN(n2842) );
  OAI211_X1 U3676 ( .C1(n2013), .C2(REG1_REG_8__SCAN_IN), .A(n2840), .B(n4434), 
        .ZN(n2841) );
  OAI211_X1 U3677 ( .C1(n2843), .C2(n4389), .A(n2842), .B(n2841), .ZN(U3248)
         );
  INV_X1 U3678 ( .A(n2976), .ZN(n2849) );
  INV_X1 U3679 ( .A(n2844), .ZN(n2845) );
  NAND2_X1 U3680 ( .A1(n2845), .A2(D_REG_1__SCAN_IN), .ZN(n2847) );
  AOI21_X1 U3681 ( .B1(n2848), .B2(n2847), .A(n2846), .ZN(n2978) );
  NAND2_X1 U3682 ( .A1(n2851), .A2(n2850), .ZN(n2853) );
  NAND2_X1 U3683 ( .A1(n2853), .A2(n2852), .ZN(n2869) );
  NAND2_X1 U3684 ( .A1(n2869), .A2(n4285), .ZN(n2854) );
  NAND2_X1 U3685 ( .A1(n2872), .A2(n2854), .ZN(n2855) );
  NAND2_X1 U3686 ( .A1(n2855), .A2(n2975), .ZN(n2936) );
  INV_X1 U3687 ( .A(n2936), .ZN(n2858) );
  NAND2_X1 U3688 ( .A1(n4455), .A2(n3986), .ZN(n2856) );
  INV_X1 U3689 ( .A(n2881), .ZN(n3989) );
  NAND2_X1 U3690 ( .A1(n2872), .A2(n3989), .ZN(n2937) );
  NAND3_X1 U3691 ( .A1(n2858), .A2(n2977), .A3(n2937), .ZN(n2930) );
  INV_X1 U3692 ( .A(n2930), .ZN(n2889) );
  INV_X1 U3693 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2888) );
  NAND2_X1 U3694 ( .A1(n3986), .A2(n3992), .ZN(n2859) );
  XNOR2_X1 U3695 ( .A(n2860), .B(n3531), .ZN(n2912) );
  AOI21_X1 U3696 ( .B1(n2006), .B2(n2407), .A(n2861), .ZN(n2910) );
  NAND2_X1 U3697 ( .A1(n2863), .A2(n2862), .ZN(n2868) );
  INV_X1 U3698 ( .A(n2864), .ZN(n2866) );
  NAND2_X1 U3699 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  NAND2_X1 U3700 ( .A1(n2868), .A2(n2867), .ZN(n2873) );
  NAND2_X1 U3701 ( .A1(n2874), .A2(n2873), .ZN(n2914) );
  INV_X1 U3702 ( .A(n2869), .ZN(n2870) );
  NAND2_X1 U3703 ( .A1(n2870), .A2(n2977), .ZN(n2871) );
  OAI211_X1 U3704 ( .C1(n2874), .C2(n2873), .A(n2914), .B(n3823), .ZN(n2887)
         );
  AND2_X1 U3705 ( .A1(n2977), .A2(n4273), .ZN(n2875) );
  NAND2_X1 U3706 ( .A1(n2883), .A2(n2875), .ZN(n2878) );
  INV_X1 U3707 ( .A(n2876), .ZN(n2877) );
  INV_X1 U3708 ( .A(n4008), .ZN(n2884) );
  NOR2_X1 U3709 ( .A1(n2881), .A2(n4341), .ZN(n2879) );
  AND2_X2 U3710 ( .A1(n2883), .A2(n2879), .ZN(n3828) );
  INV_X1 U3711 ( .A(n3828), .ZN(n3626) );
  NOR2_X1 U3712 ( .A1(n2881), .A2(n2880), .ZN(n2882) );
  AND2_X2 U3713 ( .A1(n2883), .A2(n2882), .ZN(n3825) );
  INV_X1 U3714 ( .A(n3825), .ZN(n3711) );
  OAI22_X1 U3715 ( .A1(n2884), .A2(n3626), .B1(n3078), .B2(n3711), .ZN(n2885)
         );
  AOI21_X1 U3716 ( .B1(n2399), .B2(n3827), .A(n2885), .ZN(n2886) );
  OAI211_X1 U3717 ( .C1(n2889), .C2(n2888), .A(n2887), .B(n2886), .ZN(U3219)
         );
  INV_X1 U3718 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2904) );
  OAI21_X1 U3719 ( .B1(n2891), .B2(n3926), .A(n2890), .ZN(n4440) );
  INV_X1 U3720 ( .A(n4440), .ZN(n2900) );
  OAI21_X1 U3721 ( .B1(n2894), .B2(n2893), .A(n2892), .ZN(n2895) );
  NAND2_X1 U3722 ( .A1(n2895), .A2(n4159), .ZN(n2897) );
  AOI22_X1 U3723 ( .A1(n2407), .A2(n4292), .B1(n2906), .B2(n4273), .ZN(n2896)
         );
  OAI211_X1 U3724 ( .C1(n2898), .C2(n4286), .A(n2897), .B(n2896), .ZN(n2899)
         );
  AOI21_X1 U3725 ( .B1(n3147), .B2(n4440), .A(n2899), .ZN(n4443) );
  OAI21_X1 U3726 ( .B1(n2900), .B2(n4479), .A(n4443), .ZN(n2925) );
  NAND2_X1 U3727 ( .A1(n2925), .A2(n4511), .ZN(n2903) );
  AND2_X1 U3728 ( .A1(n2996), .A2(n2906), .ZN(n2901) );
  NOR2_X1 U3729 ( .A1(n3084), .A2(n2901), .ZN(n4438) );
  INV_X1 U3730 ( .A(n4329), .ZN(n4296) );
  NAND2_X1 U3731 ( .A1(n4438), .A2(n4296), .ZN(n2902) );
  OAI211_X1 U3732 ( .C1(n4511), .C2(n2904), .A(n2903), .B(n2902), .ZN(U3471)
         );
  NAND2_X1 U3733 ( .A1(n2906), .A2(n2905), .ZN(n2907) );
  NOR2_X1 U3734 ( .A1(n2921), .A2(n3523), .ZN(n2909) );
  AOI21_X1 U3735 ( .B1(n3609), .B2(n2946), .A(n2909), .ZN(n2939) );
  INV_X1 U3736 ( .A(n2910), .ZN(n2911) );
  NAND2_X1 U3737 ( .A1(n2912), .A2(n2911), .ZN(n2913) );
  NAND2_X1 U3738 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  INV_X1 U3739 ( .A(n2915), .ZN(n2917) );
  INV_X1 U3740 ( .A(n2919), .ZN(n2916) );
  NAND2_X1 U3741 ( .A1(n2917), .A2(n2916), .ZN(n2942) );
  INV_X1 U3742 ( .A(n2942), .ZN(n2918) );
  AOI21_X1 U3743 ( .B1(n2919), .B2(n2915), .A(n2918), .ZN(n2924) );
  INV_X1 U3744 ( .A(n3827), .ZN(n3625) );
  AOI22_X1 U3745 ( .A1(n3825), .A2(n4006), .B1(n2407), .B2(n3828), .ZN(n2920)
         );
  OAI21_X1 U3746 ( .B1(n3625), .B2(n2921), .A(n2920), .ZN(n2922) );
  AOI21_X1 U3747 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2930), .A(n2922), .ZN(n2923)
         );
  OAI21_X1 U3748 ( .B1(n2924), .B2(n3818), .A(n2923), .ZN(U3234) );
  NAND2_X1 U3749 ( .A1(n2925), .A2(n4518), .ZN(n2927) );
  INV_X1 U3750 ( .A(n4268), .ZN(n4192) );
  NAND2_X1 U3751 ( .A1(n4438), .A2(n4192), .ZN(n2926) );
  OAI211_X1 U3752 ( .C1(n4518), .C2(n2928), .A(n2927), .B(n2926), .ZN(U3520)
         );
  OAI22_X1 U3753 ( .A1(n2400), .A2(n3711), .B1(n3625), .B2(n2998), .ZN(n2929)
         );
  AOI21_X1 U3754 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2930), .A(n2929), .ZN(n2931)
         );
  OAI21_X1 U3755 ( .B1(n2932), .B2(n3818), .A(n2931), .ZN(U3229) );
  NAND2_X1 U3756 ( .A1(n2934), .A2(n2933), .ZN(n2935) );
  OAI21_X1 U3757 ( .B1(n2936), .B2(n2935), .A(STATE_REG_SCAN_IN), .ZN(n2938)
         );
  INV_X1 U3758 ( .A(n3830), .ZN(n3815) );
  NAND2_X1 U3759 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  NAND2_X1 U3760 ( .A1(n2942), .A2(n2941), .ZN(n3605) );
  NAND2_X1 U3761 ( .A1(n4006), .A2(n2908), .ZN(n2944) );
  NAND2_X1 U3762 ( .A1(n3610), .A2(n2905), .ZN(n2943) );
  NAND2_X1 U3763 ( .A1(n2944), .A2(n2943), .ZN(n2945) );
  XNOR2_X1 U3764 ( .A(n2945), .B(n3531), .ZN(n2947) );
  AOI22_X1 U3765 ( .A1(n4006), .A2(n2946), .B1(n2908), .B2(n3610), .ZN(n2948)
         );
  XNOR2_X1 U3766 ( .A(n2947), .B(n2948), .ZN(n3606) );
  INV_X1 U3767 ( .A(n2947), .ZN(n2949) );
  NAND2_X1 U3768 ( .A1(n2949), .A2(n2948), .ZN(n2950) );
  NAND2_X1 U3769 ( .A1(n4005), .A2(n2908), .ZN(n2952) );
  NAND2_X1 U3770 ( .A1(n3721), .A2(n2905), .ZN(n2951) );
  NAND2_X1 U3771 ( .A1(n2952), .A2(n2951), .ZN(n2953) );
  XNOR2_X1 U3772 ( .A(n2953), .B(n2865), .ZN(n2956) );
  NOR2_X1 U3773 ( .A1(n3031), .A2(n3523), .ZN(n2954) );
  AOI21_X1 U3774 ( .B1(n4005), .B2(n2946), .A(n2954), .ZN(n2957) );
  XNOR2_X1 U3775 ( .A(n2956), .B(n2957), .ZN(n3716) );
  INV_X1 U3776 ( .A(n2956), .ZN(n2959) );
  INV_X1 U3777 ( .A(n2957), .ZN(n2958) );
  NAND2_X1 U3778 ( .A1(n2959), .A2(n2958), .ZN(n3357) );
  NAND2_X1 U3779 ( .A1(n3717), .A2(n3357), .ZN(n3370) );
  NAND2_X1 U3780 ( .A1(n3801), .A2(n2908), .ZN(n2961) );
  NAND2_X1 U3781 ( .A1(n3066), .A2(n2905), .ZN(n2960) );
  NAND2_X1 U3782 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
  XNOR2_X1 U3783 ( .A(n2962), .B(n3531), .ZN(n3356) );
  NOR2_X1 U3784 ( .A1(n2965), .A2(n3523), .ZN(n2963) );
  AOI21_X1 U3785 ( .B1(n3801), .B2(n2946), .A(n2963), .ZN(n3354) );
  XNOR2_X1 U3786 ( .A(n3356), .B(n3354), .ZN(n3366) );
  NAND2_X1 U3787 ( .A1(n3370), .A2(n3366), .ZN(n2964) );
  OAI211_X1 U3788 ( .C1(n3370), .C2(n3366), .A(n2964), .B(n3823), .ZN(n2969)
         );
  INV_X1 U3789 ( .A(n4005), .ZN(n3063) );
  OAI22_X1 U3790 ( .A1(n3063), .A2(n3626), .B1(n3625), .B2(n2965), .ZN(n2966)
         );
  AOI211_X1 U3791 ( .C1(n3825), .C2(n3557), .A(n2967), .B(n2966), .ZN(n2968)
         );
  OAI211_X1 U3792 ( .C1(n3815), .C2(n3070), .A(n2969), .B(n2968), .ZN(U3224)
         );
  XNOR2_X1 U3793 ( .A(n2970), .B(n2985), .ZN(n2974) );
  NAND2_X1 U3794 ( .A1(n3557), .A2(n4292), .ZN(n2972) );
  NAND2_X1 U3795 ( .A1(n4003), .A2(n4274), .ZN(n2971) );
  OAI211_X1 U3796 ( .C1(n4285), .C2(n3376), .A(n2972), .B(n2971), .ZN(n2973)
         );
  AOI21_X1 U3797 ( .B1(n2974), .B2(n4159), .A(n2973), .ZN(n4500) );
  NAND4_X1 U3798 ( .A1(n2978), .A2(n2977), .A3(n2976), .A4(n2975), .ZN(n2979)
         );
  OAI211_X1 U3799 ( .C1(n3014), .C2(n3376), .A(n4504), .B(n3104), .ZN(n4497)
         );
  INV_X1 U3800 ( .A(n4497), .ZN(n2982) );
  AND2_X1 U3801 ( .A1(n2999), .A2(n3986), .ZN(n3317) );
  OAI22_X1 U3802 ( .A1(n2999), .A2(n2980), .B1(n3559), .B2(n4145), .ZN(n2981)
         );
  AOI21_X1 U3803 ( .B1(n2982), .B2(n3317), .A(n2981), .ZN(n2989) );
  NAND2_X1 U3804 ( .A1(n2984), .A2(n2462), .ZN(n4496) );
  OR2_X1 U3805 ( .A1(n2986), .A2(n3986), .ZN(n3000) );
  NAND2_X1 U3806 ( .A1(n3200), .A2(n3000), .ZN(n2987) );
  NAND3_X1 U3807 ( .A1(n2983), .A2(n4496), .A3(n4176), .ZN(n2988) );
  OAI211_X1 U3808 ( .C1(n4500), .C2(n4182), .A(n2989), .B(n2988), .ZN(U3283)
         );
  XNOR2_X1 U3809 ( .A(n2660), .B(n3844), .ZN(n2995) );
  OAI21_X1 U3810 ( .B1(n2660), .B2(n2991), .A(n2990), .ZN(n4473) );
  AOI22_X1 U3811 ( .A1(n3609), .A2(n4274), .B1(n4273), .B2(n2399), .ZN(n2993)
         );
  NAND2_X1 U3812 ( .A1(n4008), .A2(n4292), .ZN(n2992) );
  OAI211_X1 U3813 ( .C1(n4473), .C2(n3200), .A(n2993), .B(n2992), .ZN(n2994)
         );
  AOI21_X1 U3814 ( .B1(n4159), .B2(n2995), .A(n2994), .ZN(n4471) );
  OAI21_X1 U3815 ( .B1(n2998), .B2(n2997), .A(n2996), .ZN(n4472) );
  INV_X1 U3816 ( .A(n4472), .ZN(n3004) );
  INV_X1 U3817 ( .A(n3000), .ZN(n3001) );
  NAND2_X1 U3818 ( .A1(n2999), .A2(n3001), .ZN(n3208) );
  AOI22_X1 U3819 ( .A1(n4182), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4448), .ZN(n3002) );
  OAI21_X1 U3820 ( .B1(n4473), .B2(n3208), .A(n3002), .ZN(n3003) );
  AOI21_X1 U3821 ( .B1(n4439), .B2(n3004), .A(n3003), .ZN(n3005) );
  OAI21_X1 U3822 ( .B1(n4471), .B2(n4182), .A(n3005), .ZN(U3289) );
  INV_X1 U3823 ( .A(n3007), .ZN(n3877) );
  OR2_X1 U3824 ( .A1(n3877), .A2(n3860), .ZN(n3933) );
  XNOR2_X1 U3825 ( .A(n3006), .B(n3933), .ZN(n3045) );
  XOR2_X1 U3826 ( .A(n3933), .B(n3008), .Z(n3043) );
  AOI22_X1 U3827 ( .A1(n4004), .A2(n4274), .B1(n3802), .B2(n4273), .ZN(n3009)
         );
  OAI21_X1 U3828 ( .B1(n3010), .B2(n4277), .A(n3009), .ZN(n3011) );
  AOI21_X1 U3829 ( .B1(n3043), .B2(n4159), .A(n3011), .ZN(n3012) );
  OAI21_X1 U3830 ( .B1(n4490), .B2(n3045), .A(n3012), .ZN(n3019) );
  NOR2_X1 U3831 ( .A1(n3069), .A2(n3039), .ZN(n3013) );
  OR2_X1 U3832 ( .A1(n3014), .A2(n3013), .ZN(n3035) );
  OAI22_X1 U3833 ( .A1(n3035), .A2(n4268), .B1(n4518), .B2(n2448), .ZN(n3015)
         );
  AOI21_X1 U3834 ( .B1(n3019), .B2(n4518), .A(n3015), .ZN(n3016) );
  INV_X1 U3835 ( .A(n3016), .ZN(U3524) );
  INV_X1 U3836 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3017) );
  OAI22_X1 U3837 ( .A1(n3035), .A2(n4329), .B1(n4511), .B2(n3017), .ZN(n3018)
         );
  AOI21_X1 U3838 ( .B1(n3019), .B2(n4511), .A(n3018), .ZN(n3020) );
  INV_X1 U3839 ( .A(n3020), .ZN(U3479) );
  INV_X1 U3840 ( .A(n3932), .ZN(n3024) );
  NAND2_X1 U3841 ( .A1(n3022), .A2(n3024), .ZN(n3023) );
  NAND2_X1 U3842 ( .A1(n3021), .A2(n3023), .ZN(n4483) );
  XNOR2_X1 U3843 ( .A(n3025), .B(n3024), .ZN(n3029) );
  AOI22_X1 U3844 ( .A1(n4006), .A2(n4292), .B1(n3721), .B2(n4273), .ZN(n3027)
         );
  NAND2_X1 U3845 ( .A1(n3801), .A2(n4274), .ZN(n3026) );
  OAI211_X1 U3846 ( .C1(n4483), .C2(n3200), .A(n3027), .B(n3026), .ZN(n3028)
         );
  AOI21_X1 U3847 ( .B1(n3029), .B2(n4159), .A(n3028), .ZN(n3030) );
  INV_X1 U3848 ( .A(n3030), .ZN(n4485) );
  OAI211_X1 U3849 ( .C1(n2039), .C2(n3031), .A(n4504), .B(n3067), .ZN(n4484)
         );
  OAI22_X1 U3850 ( .A1(n4484), .A2(n4444), .B1(n4145), .B2(n3722), .ZN(n3032)
         );
  OAI21_X1 U3851 ( .B1(n4485), .B2(n3032), .A(n2999), .ZN(n3034) );
  NAND2_X1 U3852 ( .A1(n4182), .A2(REG2_REG_4__SCAN_IN), .ZN(n3033) );
  OAI211_X1 U3853 ( .C1(n4483), .C2(n3208), .A(n3034), .B(n3033), .ZN(U3286)
         );
  NAND2_X1 U3854 ( .A1(n2999), .A2(n4159), .ZN(n4191) );
  INV_X1 U3855 ( .A(n4191), .ZN(n3042) );
  NOR2_X1 U3856 ( .A1(n3035), .A2(n4164), .ZN(n3041) );
  AND2_X1 U3857 ( .A1(n2999), .A2(n4273), .ZN(n4119) );
  INV_X1 U3858 ( .A(n4119), .ZN(n4186) );
  AND2_X1 U3859 ( .A1(n2999), .A2(n4274), .ZN(n4181) );
  AND2_X1 U3860 ( .A1(n2999), .A2(n4292), .ZN(n4180) );
  AOI22_X1 U3861 ( .A1(n4181), .A2(n4004), .B1(n3801), .B2(n4180), .ZN(n3038)
         );
  INV_X1 U3862 ( .A(n3036), .ZN(n3803) );
  AOI22_X1 U3863 ( .A1(n4182), .A2(REG2_REG_6__SCAN_IN), .B1(n3803), .B2(n4448), .ZN(n3037) );
  OAI211_X1 U3864 ( .C1(n3039), .C2(n4186), .A(n3038), .B(n3037), .ZN(n3040)
         );
  AOI211_X1 U3865 ( .C1(n3043), .C2(n3042), .A(n3041), .B(n3040), .ZN(n3044)
         );
  OAI21_X1 U3866 ( .B1(n4169), .B2(n3045), .A(n3044), .ZN(U3284) );
  INV_X1 U3867 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U3868 ( .A1(n4120), .A2(U4043), .ZN(n3046) );
  OAI21_X1 U3869 ( .B1(U4043), .B2(n4616), .A(n3046), .ZN(U3575) );
  INV_X1 U3870 ( .A(n3875), .ZN(n3871) );
  NAND2_X1 U3871 ( .A1(n3871), .A2(n3867), .ZN(n3934) );
  XNOR2_X1 U3872 ( .A(n3047), .B(n3934), .ZN(n3052) );
  NAND2_X1 U3873 ( .A1(n4003), .A2(n4292), .ZN(n3049) );
  NAND2_X1 U3874 ( .A1(n4002), .A2(n4274), .ZN(n3048) );
  OAI211_X1 U3875 ( .C1(n4285), .C2(n3050), .A(n3049), .B(n3048), .ZN(n3051)
         );
  AOI21_X1 U3876 ( .B1(n3052), .B2(n4159), .A(n3051), .ZN(n4507) );
  AND2_X1 U3877 ( .A1(n3106), .A2(n3732), .ZN(n3053) );
  NOR2_X1 U3878 ( .A1(n3093), .A2(n3053), .ZN(n4505) );
  OAI22_X1 U3879 ( .A1(n2999), .A2(n2338), .B1(n3733), .B2(n4145), .ZN(n3054)
         );
  AOI21_X1 U3880 ( .B1(n4505), .B2(n4439), .A(n3054), .ZN(n3058) );
  INV_X1 U3881 ( .A(n3934), .ZN(n3056) );
  XNOR2_X1 U3882 ( .A(n3055), .B(n3056), .ZN(n4503) );
  NAND2_X1 U3883 ( .A1(n4503), .A2(n4176), .ZN(n3057) );
  OAI211_X1 U3884 ( .C1(n4507), .C2(n4182), .A(n3058), .B(n3057), .ZN(U3281)
         );
  INV_X1 U3885 ( .A(n3857), .ZN(n3059) );
  NAND2_X1 U3886 ( .A1(n3059), .A2(n3874), .ZN(n3948) );
  XNOR2_X1 U3887 ( .A(n3060), .B(n3948), .ZN(n4491) );
  XNOR2_X1 U3888 ( .A(n3061), .B(n3948), .ZN(n3065) );
  AOI22_X1 U3889 ( .A1(n3557), .A2(n4274), .B1(n4273), .B2(n3066), .ZN(n3062)
         );
  OAI21_X1 U3890 ( .B1(n3063), .B2(n4277), .A(n3062), .ZN(n3064) );
  AOI21_X1 U3891 ( .B1(n3065), .B2(n4159), .A(n3064), .ZN(n4492) );
  MUX2_X1 U3892 ( .A(n4492), .B(n2330), .S(n4182), .Z(n3073) );
  AND2_X1 U3893 ( .A1(n3067), .A2(n3066), .ZN(n3068) );
  NOR2_X1 U3894 ( .A1(n3069), .A2(n3068), .ZN(n4495) );
  INV_X1 U3895 ( .A(n3070), .ZN(n3071) );
  AOI22_X1 U3896 ( .A1(n4495), .A2(n4439), .B1(n3071), .B2(n4448), .ZN(n3072)
         );
  OAI211_X1 U3897 ( .C1(n4169), .C2(n4491), .A(n3073), .B(n3072), .ZN(U3285)
         );
  XNOR2_X1 U3898 ( .A(n3074), .B(n3075), .ZN(n4480) );
  XNOR2_X1 U3899 ( .A(n3076), .B(n3075), .ZN(n3080) );
  AOI22_X1 U3900 ( .A1(n4005), .A2(n4274), .B1(n4273), .B2(n3610), .ZN(n3077)
         );
  OAI21_X1 U3901 ( .B1(n3078), .B2(n4277), .A(n3077), .ZN(n3079) );
  AOI21_X1 U3902 ( .B1(n3080), .B2(n4159), .A(n3079), .ZN(n3081) );
  OAI21_X1 U3903 ( .B1(n4480), .B2(n3200), .A(n3081), .ZN(n4482) );
  INV_X1 U3904 ( .A(n4482), .ZN(n3090) );
  INV_X1 U3905 ( .A(n4480), .ZN(n3088) );
  INV_X1 U3906 ( .A(n3208), .ZN(n4449) );
  OAI21_X1 U3907 ( .B1(n3084), .B2(n3083), .A(n3082), .ZN(n4477) );
  AOI22_X1 U3908 ( .A1(n4182), .A2(REG2_REG_3__SCAN_IN), .B1(n4448), .B2(n3085), .ZN(n3086) );
  OAI21_X1 U3909 ( .B1(n4164), .B2(n4477), .A(n3086), .ZN(n3087) );
  AOI21_X1 U3910 ( .B1(n3088), .B2(n4449), .A(n3087), .ZN(n3089) );
  OAI21_X1 U3911 ( .B1(n3090), .B2(n4182), .A(n3089), .ZN(U3287) );
  NAND2_X1 U3912 ( .A1(n3878), .A2(n3882), .ZN(n3925) );
  INV_X1 U3913 ( .A(n3925), .ZN(n3091) );
  XNOR2_X1 U3914 ( .A(n3092), .B(n3091), .ZN(n3133) );
  INV_X1 U3915 ( .A(n3133), .ZN(n3102) );
  INV_X1 U3916 ( .A(n3093), .ZN(n3094) );
  AOI21_X1 U3917 ( .B1(n3599), .B2(n3094), .A(n3154), .ZN(n3141) );
  AOI22_X1 U3918 ( .A1(n4180), .A2(n3641), .B1(n4001), .B2(n4181), .ZN(n3097)
         );
  INV_X1 U3919 ( .A(n3095), .ZN(n3600) );
  AOI22_X1 U3920 ( .A1(n4182), .A2(REG2_REG_10__SCAN_IN), .B1(n3600), .B2(
        n4448), .ZN(n3096) );
  OAI211_X1 U3921 ( .C1(n3131), .C2(n4186), .A(n3097), .B(n3096), .ZN(n3098)
         );
  AOI21_X1 U3922 ( .B1(n3141), .B2(n4439), .A(n3098), .ZN(n3101) );
  XNOR2_X1 U3923 ( .A(n3099), .B(n3925), .ZN(n3134) );
  NAND2_X1 U3924 ( .A1(n3134), .A2(n4176), .ZN(n3100) );
  OAI211_X1 U3925 ( .C1(n3102), .C2(n4191), .A(n3101), .B(n3100), .ZN(U3280)
         );
  NAND2_X1 U3926 ( .A1(n3866), .A2(n3864), .ZN(n3931) );
  XNOR2_X1 U3927 ( .A(n3103), .B(n3931), .ZN(n3121) );
  NAND2_X1 U3928 ( .A1(n3104), .A2(n3640), .ZN(n3105) );
  NAND2_X1 U3929 ( .A1(n3106), .A2(n3105), .ZN(n3125) );
  INV_X1 U3930 ( .A(n3125), .ZN(n3113) );
  AOI22_X1 U3931 ( .A1(n4181), .A2(n3641), .B1(n4004), .B2(n4180), .ZN(n3109)
         );
  INV_X1 U3932 ( .A(n3107), .ZN(n3642) );
  AOI22_X1 U3933 ( .A1(n4182), .A2(REG2_REG_8__SCAN_IN), .B1(n3642), .B2(n4448), .ZN(n3108) );
  OAI211_X1 U3934 ( .C1(n3115), .C2(n4186), .A(n3109), .B(n3108), .ZN(n3112)
         );
  XOR2_X1 U3935 ( .A(n3931), .B(n3110), .Z(n3117) );
  NOR2_X1 U3936 ( .A1(n3117), .A2(n4191), .ZN(n3111) );
  AOI211_X1 U3937 ( .C1(n3113), .C2(n4439), .A(n3112), .B(n3111), .ZN(n3114)
         );
  OAI21_X1 U3938 ( .B1(n4169), .B2(n3121), .A(n3114), .ZN(U3282) );
  OAI22_X1 U3939 ( .A1(n3116), .A2(n4286), .B1(n3115), .B2(n4285), .ZN(n3119)
         );
  NOR2_X1 U3940 ( .A1(n3117), .A2(n4259), .ZN(n3118) );
  AOI211_X1 U3941 ( .C1(n4292), .C2(n4004), .A(n3119), .B(n3118), .ZN(n3120)
         );
  OAI21_X1 U3942 ( .B1(n4490), .B2(n3121), .A(n3120), .ZN(n3127) );
  OAI22_X1 U3943 ( .A1(n3125), .A2(n4268), .B1(n4518), .B2(n3122), .ZN(n3123)
         );
  AOI21_X1 U3944 ( .B1(n3127), .B2(n4518), .A(n3123), .ZN(n3124) );
  INV_X1 U3945 ( .A(n3124), .ZN(U3526) );
  INV_X1 U3946 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4665) );
  OAI22_X1 U3947 ( .A1(n3125), .A2(n4329), .B1(n4511), .B2(n4665), .ZN(n3126)
         );
  AOI21_X1 U3948 ( .B1(n3127), .B2(n4511), .A(n3126), .ZN(n3128) );
  INV_X1 U3949 ( .A(n3128), .ZN(U3483) );
  NAND2_X1 U3950 ( .A1(n3641), .A2(n4292), .ZN(n3130) );
  NAND2_X1 U3951 ( .A1(n4001), .A2(n4274), .ZN(n3129) );
  OAI211_X1 U3952 ( .C1(n4285), .C2(n3131), .A(n3130), .B(n3129), .ZN(n3132)
         );
  AOI21_X1 U3953 ( .B1(n3133), .B2(n4159), .A(n3132), .ZN(n3136) );
  NAND2_X1 U3954 ( .A1(n3134), .A2(n4502), .ZN(n3135) );
  NAND2_X1 U3955 ( .A1(n3136), .A2(n3135), .ZN(n3139) );
  MUX2_X1 U3956 ( .A(REG1_REG_10__SCAN_IN), .B(n3139), .S(n4521), .Z(n3137) );
  AOI21_X1 U3957 ( .B1(n4192), .B2(n3141), .A(n3137), .ZN(n3138) );
  INV_X1 U3958 ( .A(n3138), .ZN(U3528) );
  MUX2_X1 U3959 ( .A(REG0_REG_10__SCAN_IN), .B(n3139), .S(n4511), .Z(n3140) );
  AOI21_X1 U3960 ( .B1(n3141), .B2(n4296), .A(n3140), .ZN(n3142) );
  INV_X1 U3961 ( .A(n3142), .ZN(U3487) );
  XNOR2_X1 U3962 ( .A(n3169), .B(n3143), .ZN(n3152) );
  NAND2_X1 U3963 ( .A1(n3144), .A2(n3143), .ZN(n3145) );
  NAND2_X1 U3964 ( .A1(n3146), .A2(n3145), .ZN(n3224) );
  NAND2_X1 U3965 ( .A1(n3224), .A2(n3147), .ZN(n3149) );
  INV_X1 U3966 ( .A(n3153), .ZN(n3777) );
  AOI22_X1 U3967 ( .A1(n3776), .A2(n4274), .B1(n4273), .B2(n3777), .ZN(n3148)
         );
  OAI211_X1 U3968 ( .C1(n3150), .C2(n4277), .A(n3149), .B(n3148), .ZN(n3151)
         );
  AOI21_X1 U3969 ( .B1(n3152), .B2(n4159), .A(n3151), .ZN(n3222) );
  OR2_X1 U3970 ( .A1(n3154), .A2(n3153), .ZN(n3155) );
  NAND2_X1 U3971 ( .A1(n3161), .A2(n3155), .ZN(n3229) );
  INV_X1 U3972 ( .A(n3156), .ZN(n3778) );
  AOI22_X1 U3973 ( .A1(n4182), .A2(REG2_REG_11__SCAN_IN), .B1(n3778), .B2(
        n4448), .ZN(n3157) );
  OAI21_X1 U3974 ( .B1(n3229), .B2(n4164), .A(n3157), .ZN(n3158) );
  AOI21_X1 U3975 ( .B1(n3224), .B2(n4449), .A(n3158), .ZN(n3159) );
  OAI21_X1 U3976 ( .B1(n3222), .B2(n4182), .A(n3159), .ZN(U3279) );
  NAND2_X1 U3977 ( .A1(n3192), .A2(n3190), .ZN(n3924) );
  XNOR2_X1 U3978 ( .A(n3160), .B(n3924), .ZN(n3209) );
  NAND2_X1 U3979 ( .A1(n3161), .A2(n3664), .ZN(n3162) );
  NAND2_X1 U3980 ( .A1(n3201), .A2(n3162), .ZN(n3221) );
  INV_X1 U3981 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3163) );
  OAI22_X1 U3982 ( .A1(n2999), .A2(n3163), .B1(n3666), .B2(n4145), .ZN(n3164)
         );
  AOI21_X1 U3983 ( .B1(n4181), .B2(n3665), .A(n3164), .ZN(n3166) );
  AOI22_X1 U3984 ( .A1(n4180), .A2(n4001), .B1(n4119), .B2(n3664), .ZN(n3165)
         );
  OAI211_X1 U3985 ( .C1(n3221), .C2(n4164), .A(n3166), .B(n3165), .ZN(n3174)
         );
  INV_X1 U3986 ( .A(n3167), .ZN(n3168) );
  OR2_X1 U3987 ( .A1(n3169), .A2(n3168), .ZN(n3171) );
  NAND2_X1 U3988 ( .A1(n3171), .A2(n3170), .ZN(n3193) );
  XNOR2_X1 U3989 ( .A(n3193), .B(n3924), .ZN(n3172) );
  NAND2_X1 U3990 ( .A1(n3172), .A2(n4159), .ZN(n3211) );
  NOR2_X1 U3991 ( .A1(n3211), .A2(n4182), .ZN(n3173) );
  AOI211_X1 U3992 ( .C1(n4176), .C2(n3209), .A(n3174), .B(n3173), .ZN(n3175)
         );
  INV_X1 U3993 ( .A(n3175), .ZN(U3278) );
  XNOR2_X1 U3994 ( .A(n3955), .B(n3929), .ZN(n3233) );
  OAI21_X1 U3995 ( .B1(n3177), .B2(n3929), .A(n3176), .ZN(n3235) );
  NAND2_X1 U3996 ( .A1(n3235), .A2(n4176), .ZN(n3185) );
  INV_X1 U3997 ( .A(n3245), .ZN(n3178) );
  OAI21_X1 U3998 ( .B1(n2043), .B2(n3230), .A(n3178), .ZN(n3240) );
  INV_X1 U3999 ( .A(n3240), .ZN(n3183) );
  AOI22_X1 U4000 ( .A1(n4180), .A2(n3665), .B1(n4000), .B2(n4181), .ZN(n3181)
         );
  INV_X1 U4001 ( .A(n3179), .ZN(n3580) );
  AOI22_X1 U4002 ( .A1(n4182), .A2(REG2_REG_14__SCAN_IN), .B1(n3580), .B2(
        n4448), .ZN(n3180) );
  OAI211_X1 U4003 ( .C1(n3230), .C2(n4186), .A(n3181), .B(n3180), .ZN(n3182)
         );
  AOI21_X1 U4004 ( .B1(n3183), .B2(n4439), .A(n3182), .ZN(n3184) );
  OAI211_X1 U4005 ( .C1(n3233), .C2(n4191), .A(n3185), .B(n3184), .ZN(U3276)
         );
  INV_X1 U4006 ( .A(n3186), .ZN(n3188) );
  OR2_X1 U4007 ( .A1(n3188), .A2(n3187), .ZN(n3947) );
  XNOR2_X1 U4008 ( .A(n3189), .B(n3947), .ZN(n3265) );
  INV_X1 U4009 ( .A(n3190), .ZN(n3191) );
  AOI21_X1 U4010 ( .B1(n3193), .B2(n3192), .A(n3191), .ZN(n3194) );
  XOR2_X1 U4011 ( .A(n3947), .B(n3194), .Z(n3198) );
  INV_X1 U4012 ( .A(n3776), .ZN(n3196) );
  AOI22_X1 U4013 ( .A1(n4291), .A2(n4274), .B1(n4273), .B2(n3756), .ZN(n3195)
         );
  OAI21_X1 U4014 ( .B1(n3196), .B2(n4277), .A(n3195), .ZN(n3197) );
  AOI21_X1 U4015 ( .B1(n3198), .B2(n4159), .A(n3197), .ZN(n3199) );
  OAI21_X1 U4016 ( .B1(n3265), .B2(n3200), .A(n3199), .ZN(n3266) );
  NAND2_X1 U4017 ( .A1(n3266), .A2(n2999), .ZN(n3207) );
  INV_X1 U4018 ( .A(n3201), .ZN(n3203) );
  OAI21_X1 U4019 ( .B1(n3203), .B2(n3427), .A(n3202), .ZN(n3272) );
  INV_X1 U4020 ( .A(n3272), .ZN(n3205) );
  OAI22_X1 U4021 ( .A1(n2999), .A2(n3254), .B1(n3757), .B2(n4145), .ZN(n3204)
         );
  AOI21_X1 U4022 ( .B1(n3205), .B2(n4439), .A(n3204), .ZN(n3206) );
  OAI211_X1 U4023 ( .C1(n3265), .C2(n3208), .A(n3207), .B(n3206), .ZN(U3277)
         );
  NAND2_X1 U4024 ( .A1(n3209), .A2(n4502), .ZN(n3215) );
  AOI22_X1 U4025 ( .A1(n3665), .A2(n4274), .B1(n4273), .B2(n3664), .ZN(n3210)
         );
  OAI211_X1 U4026 ( .C1(n3212), .C2(n4277), .A(n3211), .B(n3210), .ZN(n3213)
         );
  INV_X1 U4027 ( .A(n3213), .ZN(n3214) );
  NAND2_X1 U4028 ( .A1(n3215), .A2(n3214), .ZN(n3218) );
  MUX2_X1 U4029 ( .A(n3218), .B(REG1_REG_12__SCAN_IN), .S(n4519), .Z(n3216) );
  INV_X1 U4030 ( .A(n3216), .ZN(n3217) );
  OAI21_X1 U4031 ( .B1(n4268), .B2(n3221), .A(n3217), .ZN(U3530) );
  MUX2_X1 U4032 ( .A(n3218), .B(REG0_REG_12__SCAN_IN), .S(n4509), .Z(n3219) );
  INV_X1 U4033 ( .A(n3219), .ZN(n3220) );
  OAI21_X1 U4034 ( .B1(n3221), .B2(n4329), .A(n3220), .ZN(U3491) );
  INV_X1 U4035 ( .A(n3222), .ZN(n3223) );
  AOI21_X1 U4036 ( .B1(n4487), .B2(n3224), .A(n3223), .ZN(n3226) );
  MUX2_X1 U4037 ( .A(n4576), .B(n3226), .S(n4521), .Z(n3225) );
  OAI21_X1 U4038 ( .B1(n4268), .B2(n3229), .A(n3225), .ZN(U3529) );
  INV_X1 U4039 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3227) );
  MUX2_X1 U4040 ( .A(n3227), .B(n3226), .S(n4511), .Z(n3228) );
  OAI21_X1 U4041 ( .B1(n3229), .B2(n4329), .A(n3228), .ZN(U3489) );
  OAI22_X1 U4042 ( .A1(n4278), .A2(n4286), .B1(n4285), .B2(n3230), .ZN(n3231)
         );
  AOI21_X1 U40430 ( .B1(n4292), .B2(n3665), .A(n3231), .ZN(n3232) );
  OAI21_X1 U4044 ( .B1(n3233), .B2(n4259), .A(n3232), .ZN(n3234) );
  AOI21_X1 U4045 ( .B1(n3235), .B2(n4502), .A(n3234), .ZN(n3237) );
  MUX2_X1 U4046 ( .A(n4388), .B(n3237), .S(n4521), .Z(n3236) );
  OAI21_X1 U4047 ( .B1(n4268), .B2(n3240), .A(n3236), .ZN(U3532) );
  INV_X1 U4048 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3238) );
  MUX2_X1 U4049 ( .A(n3238), .B(n3237), .S(n4511), .Z(n3239) );
  OAI21_X1 U4050 ( .B1(n3240), .B2(n4329), .A(n3239), .ZN(U3495) );
  XOR2_X1 U4051 ( .A(n3921), .B(n3241), .Z(n4295) );
  AOI21_X1 U4052 ( .B1(n3242), .B2(n3921), .A(n4259), .ZN(n3244) );
  NAND2_X1 U4053 ( .A1(n3244), .A2(n3243), .ZN(n4293) );
  INV_X1 U4054 ( .A(n4293), .ZN(n3251) );
  XNOR2_X1 U4055 ( .A(n3245), .B(n4284), .ZN(n4288) );
  NOR2_X1 U4056 ( .A1(n4288), .A2(n4164), .ZN(n3250) );
  INV_X1 U4057 ( .A(n4181), .ZN(n3344) );
  AOI22_X1 U4058 ( .A1(n4180), .A2(n4291), .B1(n4119), .B2(n3826), .ZN(n3248)
         );
  INV_X1 U4059 ( .A(n3246), .ZN(n3829) );
  AOI22_X1 U4060 ( .A1(n4182), .A2(REG2_REG_15__SCAN_IN), .B1(n3829), .B2(
        n4448), .ZN(n3247) );
  OAI211_X1 U4061 ( .C1(n4287), .C2(n3344), .A(n3248), .B(n3247), .ZN(n3249)
         );
  AOI211_X1 U4062 ( .C1(n3251), .C2(n2999), .A(n3250), .B(n3249), .ZN(n3252)
         );
  OAI21_X1 U4063 ( .B1(n4295), .B2(n4169), .A(n3252), .ZN(U3275) );
  AOI21_X1 U4064 ( .B1(n3254), .B2(n3264), .A(n3253), .ZN(n3256) );
  AOI21_X1 U4065 ( .B1(n3256), .B2(n3257), .A(n4389), .ZN(n3255) );
  OAI21_X1 U4066 ( .B1(n3257), .B2(n3256), .A(n3255), .ZN(n3263) );
  INV_X1 U4067 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3258) );
  NOR2_X1 U4068 ( .A1(STATE_REG_SCAN_IN), .A2(n3258), .ZN(n3755) );
  AOI211_X1 U4069 ( .C1(n3260), .C2(n3259), .A(n2183), .B(n4400), .ZN(n3261)
         );
  AOI211_X1 U4070 ( .C1(n4424), .C2(ADDR_REG_13__SCAN_IN), .A(n3755), .B(n3261), .ZN(n3262) );
  OAI211_X1 U4071 ( .C1(n4437), .C2(n3264), .A(n3263), .B(n3262), .ZN(U3253)
         );
  INV_X1 U4072 ( .A(n3265), .ZN(n3267) );
  AOI21_X1 U4073 ( .B1(n4487), .B2(n3267), .A(n3266), .ZN(n3270) );
  MUX2_X1 U4074 ( .A(n3268), .B(n3270), .S(n4521), .Z(n3269) );
  OAI21_X1 U4075 ( .B1(n4268), .B2(n3272), .A(n3269), .ZN(U3531) );
  INV_X1 U4076 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4664) );
  MUX2_X1 U4077 ( .A(n4664), .B(n3270), .S(n4511), .Z(n3271) );
  OAI21_X1 U4078 ( .B1(n3272), .B2(n4329), .A(n3271), .ZN(U3493) );
  AOI21_X1 U4079 ( .B1(n3920), .B2(n3273), .A(n3274), .ZN(n3275) );
  INV_X1 U4080 ( .A(n3275), .ZN(n4283) );
  INV_X1 U4081 ( .A(n3276), .ZN(n3291) );
  AOI21_X1 U4082 ( .B1(n4272), .B2(n3277), .A(n3291), .ZN(n4280) );
  AOI22_X1 U4083 ( .A1(n4180), .A2(n4000), .B1(n4119), .B2(n4272), .ZN(n3280)
         );
  INV_X1 U4084 ( .A(n3278), .ZN(n3687) );
  AOI22_X1 U4085 ( .A1(n4182), .A2(REG2_REG_16__SCAN_IN), .B1(n3687), .B2(
        n4448), .ZN(n3279) );
  OAI211_X1 U4086 ( .C1(n3312), .C2(n3344), .A(n3280), .B(n3279), .ZN(n3284)
         );
  OAI211_X1 U4087 ( .C1(n3282), .C2(n3920), .A(n3281), .B(n4159), .ZN(n4281)
         );
  NOR2_X1 U4088 ( .A1(n4281), .A2(n4182), .ZN(n3283) );
  AOI211_X1 U4089 ( .C1(n4280), .C2(n4439), .A(n3284), .B(n3283), .ZN(n3285)
         );
  OAI21_X1 U4090 ( .B1(n4283), .B2(n4169), .A(n3285), .ZN(U3274) );
  NAND2_X1 U4091 ( .A1(n3310), .A2(n3307), .ZN(n3946) );
  XNOR2_X1 U4092 ( .A(n3286), .B(n3946), .ZN(n3298) );
  INV_X1 U4093 ( .A(n3298), .ZN(n3296) );
  XOR2_X1 U4094 ( .A(n3946), .B(n3309), .Z(n3289) );
  OAI22_X1 U4095 ( .A1(n3627), .A2(n4286), .B1(n3454), .B2(n4285), .ZN(n3287)
         );
  AOI21_X1 U4096 ( .B1(n4292), .B2(n3999), .A(n3287), .ZN(n3288) );
  OAI21_X1 U4097 ( .B1(n3289), .B2(n4259), .A(n3288), .ZN(n3297) );
  INV_X1 U4098 ( .A(n3305), .ZN(n3290) );
  OAI21_X1 U4099 ( .B1(n3291), .B2(n3454), .A(n3290), .ZN(n3302) );
  INV_X1 U4100 ( .A(n3292), .ZN(n3699) );
  AOI22_X1 U4101 ( .A1(n4182), .A2(REG2_REG_17__SCAN_IN), .B1(n3699), .B2(
        n4448), .ZN(n3293) );
  OAI21_X1 U4102 ( .B1(n3302), .B2(n4164), .A(n3293), .ZN(n3294) );
  AOI21_X1 U4103 ( .B1(n3297), .B2(n2999), .A(n3294), .ZN(n3295) );
  OAI21_X1 U4104 ( .B1(n3296), .B2(n4169), .A(n3295), .ZN(U3273) );
  INV_X1 U4105 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4565) );
  AOI21_X1 U4106 ( .B1(n3298), .B2(n4502), .A(n3297), .ZN(n3300) );
  MUX2_X1 U4107 ( .A(n4565), .B(n3300), .S(n4511), .Z(n3299) );
  OAI21_X1 U4108 ( .B1(n3302), .B2(n4329), .A(n3299), .ZN(U3501) );
  MUX2_X1 U4109 ( .A(n4645), .B(n3300), .S(n4521), .Z(n3301) );
  OAI21_X1 U4110 ( .B1(n4268), .B2(n3302), .A(n3301), .ZN(U3535) );
  OAI21_X1 U4111 ( .B1(n2034), .B2(n3930), .A(n3303), .ZN(n3304) );
  INV_X1 U4112 ( .A(n3304), .ZN(n4271) );
  XNOR2_X1 U4113 ( .A(n3305), .B(n3788), .ZN(n3306) );
  NAND2_X1 U4114 ( .A1(n3306), .A2(n4504), .ZN(n4269) );
  INV_X1 U4115 ( .A(n4269), .ZN(n3318) );
  OAI22_X1 U4116 ( .A1(n2999), .A2(n4591), .B1(n3789), .B2(n4145), .ZN(n3316)
         );
  INV_X1 U4117 ( .A(n3307), .ZN(n3308) );
  NAND2_X1 U4118 ( .A1(n3347), .A2(n3310), .ZN(n3327) );
  XOR2_X1 U4119 ( .A(n3930), .B(n3327), .Z(n3314) );
  AOI22_X1 U4120 ( .A1(n4179), .A2(n4274), .B1(n4273), .B2(n3788), .ZN(n3311)
         );
  OAI21_X1 U4121 ( .B1(n3312), .B2(n4277), .A(n3311), .ZN(n3313) );
  AOI21_X1 U4122 ( .B1(n3314), .B2(n4159), .A(n3313), .ZN(n4270) );
  NOR2_X1 U4123 ( .A1(n4270), .A2(n4182), .ZN(n3315) );
  AOI211_X1 U4124 ( .C1(n3318), .C2(n3317), .A(n3316), .B(n3315), .ZN(n3319)
         );
  OAI21_X1 U4125 ( .B1(n4271), .B2(n4169), .A(n3319), .ZN(U3272) );
  INV_X1 U4126 ( .A(n3321), .ZN(n3323) );
  NOR2_X1 U4127 ( .A1(n3323), .A2(n3322), .ZN(n3943) );
  XNOR2_X1 U4128 ( .A(n3320), .B(n3943), .ZN(n4265) );
  INV_X1 U4129 ( .A(n4265), .ZN(n3337) );
  INV_X1 U4130 ( .A(n3324), .ZN(n3326) );
  OAI21_X1 U4131 ( .B1(n3327), .B2(n3326), .A(n3325), .ZN(n3328) );
  XNOR2_X1 U4132 ( .A(n3328), .B(n3943), .ZN(n3329) );
  NAND2_X1 U4133 ( .A1(n3329), .A2(n4159), .ZN(n3331) );
  AOI22_X1 U4134 ( .A1(n4246), .A2(n4274), .B1(n4273), .B2(n3466), .ZN(n3330)
         );
  OAI211_X1 U4135 ( .C1(n3627), .C2(n4277), .A(n3331), .B(n3330), .ZN(n4264)
         );
  OAI21_X1 U4136 ( .B1(n3333), .B2(n3624), .A(n3332), .ZN(n4330) );
  NOR2_X1 U4137 ( .A1(n4330), .A2(n4164), .ZN(n3335) );
  OAI22_X1 U4138 ( .A1(n2999), .A2(n2370), .B1(n3632), .B2(n4145), .ZN(n3334)
         );
  AOI211_X1 U4139 ( .C1(n4264), .C2(n2999), .A(n3335), .B(n3334), .ZN(n3336)
         );
  OAI21_X1 U4140 ( .B1(n3337), .B2(n4169), .A(n3336), .ZN(U3271) );
  INV_X1 U4141 ( .A(n3338), .ZN(n3898) );
  XNOR2_X1 U4142 ( .A(n3339), .B(n4133), .ZN(n4253) );
  AND2_X1 U4143 ( .A1(n4177), .A2(n4245), .ZN(n3340) );
  NOR2_X1 U4144 ( .A1(n4163), .A2(n3340), .ZN(n4250) );
  INV_X1 U4145 ( .A(n3655), .ZN(n3341) );
  AOI22_X1 U4146 ( .A1(n3341), .A2(n4448), .B1(REG2_REG_21__SCAN_IN), .B2(
        n4182), .ZN(n3343) );
  AOI22_X1 U4147 ( .A1(n4246), .A2(n4180), .B1(n4245), .B2(n4119), .ZN(n3342)
         );
  OAI211_X1 U4148 ( .C1(n4248), .C2(n3344), .A(n3343), .B(n3342), .ZN(n3352)
         );
  INV_X1 U4149 ( .A(n3345), .ZN(n3346) );
  INV_X1 U4150 ( .A(n3348), .ZN(n3349) );
  OAI21_X1 U4151 ( .B1(n4172), .B2(n3349), .A(n3897), .ZN(n4134) );
  XNOR2_X1 U4152 ( .A(n4134), .B(n4133), .ZN(n3350) );
  NAND2_X1 U4153 ( .A1(n3350), .A2(n4159), .ZN(n4251) );
  NOR2_X1 U4154 ( .A1(n4251), .A2(n4182), .ZN(n3351) );
  AOI211_X1 U4155 ( .C1(n4250), .C2(n4439), .A(n3352), .B(n3351), .ZN(n3353)
         );
  OAI21_X1 U4156 ( .B1(n4253), .B2(n4169), .A(n3353), .ZN(U3269) );
  INV_X1 U4157 ( .A(n3354), .ZN(n3355) );
  NAND2_X1 U4158 ( .A1(n3356), .A2(n3355), .ZN(n3367) );
  AND2_X1 U4159 ( .A1(n3357), .A2(n3367), .ZN(n3360) );
  INV_X1 U4160 ( .A(n3367), .ZN(n3358) );
  NOR2_X1 U4161 ( .A1(n3358), .A2(n3366), .ZN(n3359) );
  AOI21_X1 U4162 ( .B1(n3717), .B2(n3360), .A(n3359), .ZN(n3798) );
  NAND2_X1 U4163 ( .A1(n3557), .A2(n2946), .ZN(n3362) );
  NAND2_X1 U4164 ( .A1(n3802), .A2(n3530), .ZN(n3361) );
  NAND2_X1 U4165 ( .A1(n3362), .A2(n3361), .ZN(n3795) );
  NAND2_X1 U4166 ( .A1(n3557), .A2(n3530), .ZN(n3364) );
  NAND2_X1 U4167 ( .A1(n3802), .A2(n2905), .ZN(n3363) );
  NAND2_X1 U4168 ( .A1(n3364), .A2(n3363), .ZN(n3365) );
  XNOR2_X1 U4169 ( .A(n3365), .B(n3531), .ZN(n3796) );
  OAI21_X1 U4170 ( .B1(n3798), .B2(n3795), .A(n3796), .ZN(n3372) );
  AND2_X1 U4171 ( .A1(n3366), .A2(n3795), .ZN(n3369) );
  INV_X1 U4172 ( .A(n3795), .ZN(n3368) );
  NAND2_X1 U4173 ( .A1(n3372), .A2(n3371), .ZN(n3553) );
  NAND2_X1 U4174 ( .A1(n4004), .A2(n3530), .ZN(n3374) );
  NAND2_X1 U4175 ( .A1(n3558), .A2(n2905), .ZN(n3373) );
  NAND2_X1 U4176 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  XNOR2_X1 U4177 ( .A(n3375), .B(n3531), .ZN(n3380) );
  NOR2_X1 U4178 ( .A1(n3376), .A2(n3523), .ZN(n3377) );
  AOI21_X1 U4179 ( .B1(n4004), .B2(n2946), .A(n3377), .ZN(n3378) );
  NAND2_X1 U4180 ( .A1(n3553), .A2(n3554), .ZN(n3382) );
  INV_X1 U4181 ( .A(n3378), .ZN(n3379) );
  NAND2_X1 U4182 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  NAND2_X1 U4183 ( .A1(n3382), .A2(n3381), .ZN(n3633) );
  NAND2_X1 U4184 ( .A1(n4003), .A2(n3530), .ZN(n3384) );
  NAND2_X1 U4185 ( .A1(n3640), .A2(n2905), .ZN(n3383) );
  NAND2_X1 U4186 ( .A1(n3384), .A2(n3383), .ZN(n3385) );
  XNOR2_X1 U4187 ( .A(n3385), .B(n3531), .ZN(n3388) );
  NAND2_X1 U4188 ( .A1(n4003), .A2(n2005), .ZN(n3387) );
  NAND2_X1 U4189 ( .A1(n3640), .A2(n3530), .ZN(n3386) );
  NAND2_X1 U4190 ( .A1(n3387), .A2(n3386), .ZN(n3389) );
  AND2_X1 U4191 ( .A1(n3388), .A2(n3389), .ZN(n3634) );
  INV_X1 U4192 ( .A(n3388), .ZN(n3391) );
  INV_X1 U4193 ( .A(n3389), .ZN(n3390) );
  NAND2_X1 U4194 ( .A1(n3391), .A2(n3390), .ZN(n3635) );
  NAND2_X1 U4195 ( .A1(n3641), .A2(n3530), .ZN(n3393) );
  NAND2_X1 U4196 ( .A1(n3732), .A2(n2905), .ZN(n3392) );
  NAND2_X1 U4197 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  XNOR2_X1 U4198 ( .A(n3394), .B(n3531), .ZN(n3395) );
  AOI22_X1 U4199 ( .A1(n3641), .A2(n2946), .B1(n3530), .B2(n3732), .ZN(n3396)
         );
  XNOR2_X1 U4200 ( .A(n3395), .B(n3396), .ZN(n3729) );
  NAND2_X1 U4201 ( .A1(n3728), .A2(n3729), .ZN(n3399) );
  INV_X1 U4202 ( .A(n3395), .ZN(n3397) );
  NAND2_X1 U4203 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  NAND2_X1 U4204 ( .A1(n3399), .A2(n3398), .ZN(n3595) );
  INV_X1 U4205 ( .A(n3595), .ZN(n3404) );
  NAND2_X1 U4206 ( .A1(n4002), .A2(n3530), .ZN(n3401) );
  NAND2_X1 U4207 ( .A1(n3599), .A2(n2905), .ZN(n3400) );
  NAND2_X1 U4208 ( .A1(n3401), .A2(n3400), .ZN(n3402) );
  XNOR2_X1 U4209 ( .A(n3402), .B(n2865), .ZN(n3405) );
  AOI22_X1 U4210 ( .A1(n4002), .A2(n2005), .B1(n3530), .B2(n3599), .ZN(n3406)
         );
  XNOR2_X1 U4211 ( .A(n3405), .B(n3406), .ZN(n3596) );
  INV_X1 U4212 ( .A(n3405), .ZN(n3408) );
  INV_X1 U4213 ( .A(n3406), .ZN(n3407) );
  NAND2_X1 U4214 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  NAND2_X1 U4215 ( .A1(n4001), .A2(n2946), .ZN(n3411) );
  NAND2_X1 U4216 ( .A1(n3777), .A2(n3530), .ZN(n3410) );
  NAND2_X1 U4217 ( .A1(n3411), .A2(n3410), .ZN(n3771) );
  NAND2_X1 U4218 ( .A1(n4001), .A2(n3530), .ZN(n3413) );
  NAND2_X1 U4219 ( .A1(n3777), .A2(n2905), .ZN(n3412) );
  NAND2_X1 U4220 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  XNOR2_X1 U4221 ( .A(n3414), .B(n3531), .ZN(n3772) );
  NAND2_X1 U4222 ( .A1(n3776), .A2(n3530), .ZN(n3416) );
  NAND2_X1 U4223 ( .A1(n3664), .A2(n2905), .ZN(n3415) );
  NAND2_X1 U4224 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  XNOR2_X1 U4225 ( .A(n3417), .B(n3531), .ZN(n3420) );
  NAND2_X1 U4226 ( .A1(n3776), .A2(n2005), .ZN(n3419) );
  NAND2_X1 U4227 ( .A1(n3664), .A2(n2908), .ZN(n3418) );
  NAND2_X1 U4228 ( .A1(n3419), .A2(n3418), .ZN(n3421) );
  AND2_X1 U4229 ( .A1(n3420), .A2(n3421), .ZN(n3659) );
  INV_X1 U4230 ( .A(n3420), .ZN(n3423) );
  INV_X1 U4231 ( .A(n3421), .ZN(n3422) );
  NAND2_X1 U4232 ( .A1(n3423), .A2(n3422), .ZN(n3660) );
  NAND2_X1 U4233 ( .A1(n3665), .A2(n2908), .ZN(n3425) );
  NAND2_X1 U4234 ( .A1(n3756), .A2(n2905), .ZN(n3424) );
  NAND2_X1 U4235 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  XNOR2_X1 U4236 ( .A(n3426), .B(n2865), .ZN(n3750) );
  NOR2_X1 U4237 ( .A1(n3427), .A2(n3523), .ZN(n3428) );
  AOI21_X1 U4238 ( .B1(n3665), .B2(n2005), .A(n3428), .ZN(n3751) );
  AOI21_X1 U4239 ( .B1(n3753), .B2(n3750), .A(n3751), .ZN(n3429) );
  INV_X1 U4240 ( .A(n3429), .ZN(n3430) );
  NAND2_X1 U4241 ( .A1(n3430), .A2(n2007), .ZN(n3572) );
  NAND2_X1 U4242 ( .A1(n4291), .A2(n3530), .ZN(n3432) );
  NAND2_X1 U4243 ( .A1(n3579), .A2(n2905), .ZN(n3431) );
  NAND2_X1 U4244 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  XNOR2_X1 U4245 ( .A(n3433), .B(n3531), .ZN(n3436) );
  NAND2_X1 U4246 ( .A1(n4291), .A2(n2005), .ZN(n3435) );
  NAND2_X1 U4247 ( .A1(n3579), .A2(n3530), .ZN(n3434) );
  NAND2_X1 U4248 ( .A1(n3435), .A2(n3434), .ZN(n3437) );
  AND2_X1 U4249 ( .A1(n3436), .A2(n3437), .ZN(n3573) );
  INV_X1 U4250 ( .A(n3436), .ZN(n3439) );
  INV_X1 U4251 ( .A(n3437), .ZN(n3438) );
  NAND2_X1 U4252 ( .A1(n3439), .A2(n3438), .ZN(n3574) );
  NAND2_X1 U4253 ( .A1(n4000), .A2(n3530), .ZN(n3441) );
  NAND2_X1 U4254 ( .A1(n3826), .A2(n2905), .ZN(n3440) );
  NAND2_X1 U4255 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  NAND2_X1 U4256 ( .A1(n3999), .A2(n3530), .ZN(n3444) );
  NAND2_X1 U4257 ( .A1(n4272), .A2(n2905), .ZN(n3443) );
  NAND2_X1 U4258 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  XNOR2_X1 U4259 ( .A(n3445), .B(n2865), .ZN(n3447) );
  AOI22_X1 U4260 ( .A1(n3999), .A2(n2946), .B1(n2908), .B2(n4272), .ZN(n3446)
         );
  NAND2_X1 U4261 ( .A1(n3447), .A2(n3446), .ZN(n3450) );
  OAI21_X1 U4262 ( .B1(n3447), .B2(n3446), .A(n3450), .ZN(n3685) );
  NAND2_X1 U4263 ( .A1(n4000), .A2(n2005), .ZN(n3449) );
  NAND2_X1 U4264 ( .A1(n3826), .A2(n3530), .ZN(n3448) );
  NAND2_X1 U4265 ( .A1(n3449), .A2(n3448), .ZN(n3821) );
  NAND2_X1 U4266 ( .A1(n4275), .A2(n2908), .ZN(n3452) );
  NAND2_X1 U4267 ( .A1(n3698), .A2(n2905), .ZN(n3451) );
  NAND2_X1 U4268 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  XNOR2_X1 U4269 ( .A(n3453), .B(n2865), .ZN(n3457) );
  NOR2_X1 U4270 ( .A1(n3454), .A2(n3523), .ZN(n3455) );
  AOI21_X1 U4271 ( .B1(n4275), .B2(n2005), .A(n3455), .ZN(n3456) );
  NOR2_X1 U4272 ( .A1(n3457), .A2(n3456), .ZN(n3693) );
  NAND2_X1 U4273 ( .A1(n3457), .A2(n3456), .ZN(n3694) );
  NAND2_X1 U4274 ( .A1(n3998), .A2(n2005), .ZN(n3459) );
  NAND2_X1 U4275 ( .A1(n3788), .A2(n2908), .ZN(n3458) );
  NAND2_X1 U4276 ( .A1(n3459), .A2(n3458), .ZN(n3617) );
  NAND2_X1 U4277 ( .A1(n3998), .A2(n3530), .ZN(n3461) );
  NAND2_X1 U4278 ( .A1(n3788), .A2(n2905), .ZN(n3460) );
  NAND2_X1 U4279 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  XNOR2_X1 U4280 ( .A(n3462), .B(n3531), .ZN(n3784) );
  NAND2_X1 U4281 ( .A1(n4179), .A2(n3530), .ZN(n3464) );
  NAND2_X1 U4282 ( .A1(n3466), .A2(n2905), .ZN(n3463) );
  NAND2_X1 U4283 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  XNOR2_X1 U4284 ( .A(n3465), .B(n2865), .ZN(n3468) );
  AOI22_X1 U4285 ( .A1(n4179), .A2(n2946), .B1(n2908), .B2(n3466), .ZN(n3467)
         );
  NOR2_X1 U4286 ( .A1(n3468), .A2(n3467), .ZN(n3620) );
  AOI21_X1 U4287 ( .B1(n3617), .B2(n3784), .A(n3620), .ZN(n3471) );
  AND2_X1 U4288 ( .A1(n3468), .A2(n3467), .ZN(n3619) );
  NAND2_X1 U4289 ( .A1(n4246), .A2(n2908), .ZN(n3473) );
  NAND2_X1 U4290 ( .A1(n3743), .A2(n2905), .ZN(n3472) );
  NAND2_X1 U4291 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  XNOR2_X1 U4292 ( .A(n3474), .B(n2865), .ZN(n3477) );
  AND2_X1 U4293 ( .A1(n3743), .A2(n2908), .ZN(n3475) );
  AOI21_X1 U4294 ( .B1(n4246), .B2(n2005), .A(n3475), .ZN(n3476) );
  NOR2_X1 U4295 ( .A1(n3477), .A2(n3476), .ZN(n3739) );
  NAND2_X1 U4296 ( .A1(n4257), .A2(n3530), .ZN(n3479) );
  NAND2_X1 U4297 ( .A1(n4245), .A2(n2905), .ZN(n3478) );
  NAND2_X1 U4298 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  XNOR2_X1 U4299 ( .A(n3480), .B(n3531), .ZN(n3486) );
  INV_X1 U4300 ( .A(n3486), .ZN(n3484) );
  NAND2_X1 U4301 ( .A1(n4257), .A2(n2946), .ZN(n3482) );
  NAND2_X1 U4302 ( .A1(n4245), .A2(n3530), .ZN(n3481) );
  NAND2_X1 U4303 ( .A1(n3482), .A2(n3481), .ZN(n3485) );
  INV_X1 U4304 ( .A(n3485), .ZN(n3483) );
  NAND2_X1 U4305 ( .A1(n3484), .A2(n3483), .ZN(n3647) );
  AND2_X1 U4306 ( .A1(n3486), .A2(n3485), .ZN(n3648) );
  OAI22_X1 U4307 ( .A1(n4248), .A2(n3524), .B1(n3523), .B2(n4162), .ZN(n3494)
         );
  OAI22_X1 U4308 ( .A1(n4248), .A2(n3523), .B1(n3521), .B2(n4162), .ZN(n3487)
         );
  XNOR2_X1 U4309 ( .A(n3487), .B(n3531), .ZN(n3493) );
  XOR2_X1 U4310 ( .A(n3494), .B(n3493), .Z(n3764) );
  NAND2_X1 U4311 ( .A1(n3763), .A2(n3764), .ZN(n3586) );
  NAND2_X1 U4312 ( .A1(n4228), .A2(n3530), .ZN(n3490) );
  NAND2_X1 U4313 ( .A1(n3488), .A2(n2905), .ZN(n3489) );
  NAND2_X1 U4314 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  XNOR2_X1 U4315 ( .A(n3491), .B(n3531), .ZN(n3500) );
  NOR2_X1 U4316 ( .A1(n4143), .A2(n3523), .ZN(n3492) );
  AOI21_X1 U4317 ( .B1(n4228), .B2(n2006), .A(n3492), .ZN(n3498) );
  XNOR2_X1 U4318 ( .A(n3500), .B(n3498), .ZN(n3587) );
  INV_X1 U4319 ( .A(n3493), .ZN(n3496) );
  INV_X1 U4320 ( .A(n3494), .ZN(n3495) );
  NAND2_X1 U4321 ( .A1(n3496), .A2(n3495), .ZN(n3588) );
  NAND2_X1 U4322 ( .A1(n3586), .A2(n3497), .ZN(n3585) );
  INV_X1 U4323 ( .A(n3498), .ZN(n3499) );
  NAND2_X1 U4324 ( .A1(n3500), .A2(n3499), .ZN(n3507) );
  INV_X1 U4325 ( .A(n3507), .ZN(n3501) );
  OAI22_X1 U4326 ( .A1(n4100), .A2(n3524), .B1(n3523), .B2(n3503), .ZN(n3505)
         );
  OAI22_X1 U4327 ( .A1(n4100), .A2(n3523), .B1(n3521), .B2(n3503), .ZN(n3504)
         );
  XNOR2_X1 U4328 ( .A(n3504), .B(n3531), .ZN(n3707) );
  INV_X1 U4329 ( .A(n3505), .ZN(n3506) );
  AOI21_X1 U4330 ( .B1(n3585), .B2(n3507), .A(n3506), .ZN(n3704) );
  NAND2_X1 U4331 ( .A1(n4120), .A2(n3530), .ZN(n3509) );
  NAND2_X1 U4332 ( .A1(n4104), .A2(n2905), .ZN(n3508) );
  NAND2_X1 U4333 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  XNOR2_X1 U4334 ( .A(n3510), .B(n3531), .ZN(n3514) );
  NAND2_X1 U4335 ( .A1(n4120), .A2(n2005), .ZN(n3512) );
  NAND2_X1 U4336 ( .A1(n4104), .A2(n2908), .ZN(n3511) );
  NAND2_X1 U4337 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  NOR2_X1 U4338 ( .A1(n3514), .A2(n3513), .ZN(n3672) );
  NAND2_X1 U4339 ( .A1(n3514), .A2(n3513), .ZN(n3673) );
  NAND2_X1 U4340 ( .A1(n4211), .A2(n3530), .ZN(n3516) );
  NAND2_X1 U4341 ( .A1(n4085), .A2(n2905), .ZN(n3515) );
  NAND2_X1 U4342 ( .A1(n3516), .A2(n3515), .ZN(n3517) );
  XNOR2_X1 U4343 ( .A(n3517), .B(n2865), .ZN(n3520) );
  NOR2_X1 U4344 ( .A1(n4078), .A2(n3523), .ZN(n3518) );
  AOI21_X1 U4345 ( .B1(n4211), .B2(n2005), .A(n3518), .ZN(n3519) );
  NOR2_X1 U4346 ( .A1(n3520), .A2(n3519), .ZN(n3811) );
  NAND2_X1 U4347 ( .A1(n3520), .A2(n3519), .ZN(n3809) );
  OAI22_X1 U4348 ( .A1(n3525), .A2(n3523), .B1(n4062), .B2(n3521), .ZN(n3522)
         );
  XNOR2_X1 U4349 ( .A(n3522), .B(n3531), .ZN(n3527) );
  OAI22_X1 U4350 ( .A1(n3525), .A2(n3524), .B1(n4062), .B2(n3523), .ZN(n3526)
         );
  XNOR2_X1 U4351 ( .A(n3527), .B(n3526), .ZN(n3565) );
  INV_X1 U4352 ( .A(n3526), .ZN(n3529) );
  INV_X1 U4353 ( .A(n3527), .ZN(n3528) );
  AOI22_X1 U4354 ( .A1(n4212), .A2(n3530), .B1(n2905), .B2(n4047), .ZN(n3534)
         );
  AOI22_X1 U4355 ( .A1(n4212), .A2(n2005), .B1(n3530), .B2(n4047), .ZN(n3532)
         );
  XNOR2_X1 U4356 ( .A(n3532), .B(n3531), .ZN(n3533) );
  XOR2_X1 U4357 ( .A(n3534), .B(n3533), .Z(n3535) );
  NAND2_X1 U4358 ( .A1(n3996), .A2(n3825), .ZN(n3538) );
  AOI22_X1 U4359 ( .A1(n3827), .A2(n4047), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3537) );
  NAND2_X1 U4360 ( .A1(n3542), .A2(n3830), .ZN(n3536) );
  NAND3_X1 U4361 ( .A1(n3538), .A2(n3537), .A3(n3536), .ZN(n3539) );
  AOI21_X1 U4362 ( .B1(n3828), .B2(n4080), .A(n3539), .ZN(n3540) );
  OAI21_X1 U4363 ( .B1(n3541), .B2(n3818), .A(n3540), .ZN(U3217) );
  NAND2_X1 U4364 ( .A1(n4080), .A2(n4180), .ZN(n3546) );
  AOI22_X1 U4365 ( .A1(n4119), .A2(n4047), .B1(n4182), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3545) );
  NAND2_X1 U4366 ( .A1(n3996), .A2(n4181), .ZN(n3544) );
  NAND2_X1 U4367 ( .A1(n3542), .A2(n4448), .ZN(n3543) );
  NAND4_X1 U4368 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3549)
         );
  NOR2_X1 U4369 ( .A1(n3547), .A2(n4164), .ZN(n3548) );
  AOI211_X1 U4370 ( .C1(n3550), .C2(n2999), .A(n3549), .B(n3548), .ZN(n3551)
         );
  OAI21_X1 U4371 ( .B1(n3552), .B2(n4169), .A(n3551), .ZN(U3262) );
  XOR2_X1 U4372 ( .A(n3553), .B(n3554), .Z(n3555) );
  NAND2_X1 U4373 ( .A1(n3555), .A2(n3823), .ZN(n3564) );
  AOI21_X1 U4374 ( .B1(n3557), .B2(n3828), .A(n3556), .ZN(n3563) );
  AOI22_X1 U4375 ( .A1(n4003), .A2(n3825), .B1(n3827), .B2(n3558), .ZN(n3562)
         );
  INV_X1 U4376 ( .A(n3559), .ZN(n3560) );
  NAND2_X1 U4377 ( .A1(n3830), .A2(n3560), .ZN(n3561) );
  NAND4_X1 U4378 ( .A1(n3564), .A2(n3563), .A3(n3562), .A4(n3561), .ZN(U3210)
         );
  XNOR2_X1 U4379 ( .A(n3566), .B(n3565), .ZN(n3571) );
  NAND2_X1 U4380 ( .A1(n4211), .A2(n3828), .ZN(n3568) );
  AOI22_X1 U4381 ( .A1(n3827), .A2(n4210), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3567) );
  OAI211_X1 U4382 ( .C1(n3815), .C2(n4067), .A(n3568), .B(n3567), .ZN(n3569)
         );
  AOI21_X1 U4383 ( .B1(n3825), .B2(n4212), .A(n3569), .ZN(n3570) );
  OAI21_X1 U4384 ( .B1(n3571), .B2(n3818), .A(n3570), .ZN(U3211) );
  INV_X1 U4385 ( .A(n3573), .ZN(n3575) );
  NAND2_X1 U4386 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  XNOR2_X1 U4387 ( .A(n3572), .B(n3576), .ZN(n3577) );
  NAND2_X1 U4388 ( .A1(n3577), .A2(n3823), .ZN(n3584) );
  NAND2_X1 U4389 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4397) );
  INV_X1 U4390 ( .A(n4397), .ZN(n3578) );
  AOI21_X1 U4391 ( .B1(n3665), .B2(n3828), .A(n3578), .ZN(n3583) );
  AOI22_X1 U4392 ( .A1(n4000), .A2(n3825), .B1(n3827), .B2(n3579), .ZN(n3582)
         );
  NAND2_X1 U4393 ( .A1(n3830), .A2(n3580), .ZN(n3581) );
  NAND4_X1 U4394 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(U3212)
         );
  INV_X1 U4395 ( .A(n3585), .ZN(n3590) );
  AOI21_X1 U4396 ( .B1(n3586), .B2(n3588), .A(n3587), .ZN(n3589) );
  OR3_X1 U4397 ( .A1(n3590), .A2(n3589), .A3(n3818), .ZN(n3594) );
  AOI22_X1 U4398 ( .A1(n3997), .A2(n3828), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3591) );
  OAI21_X1 U4399 ( .B1(n3625), .B2(n4143), .A(n3591), .ZN(n3592) );
  AOI21_X1 U4400 ( .B1(n3825), .B2(n4139), .A(n3592), .ZN(n3593) );
  OAI211_X1 U4401 ( .C1(n3815), .C2(n4146), .A(n3594), .B(n3593), .ZN(U3213)
         );
  AOI21_X1 U4402 ( .B1(n3595), .B2(n3596), .A(n3818), .ZN(n3598) );
  NAND2_X1 U4403 ( .A1(n3598), .A2(n3597), .ZN(n3604) );
  AND2_X1 U4404 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4361) );
  AOI21_X1 U4405 ( .B1(n3641), .B2(n3828), .A(n4361), .ZN(n3603) );
  AOI22_X1 U4406 ( .A1(n4001), .A2(n3825), .B1(n3827), .B2(n3599), .ZN(n3602)
         );
  NAND2_X1 U4407 ( .A1(n3830), .A2(n3600), .ZN(n3601) );
  NAND4_X1 U4408 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(U3214)
         );
  XNOR2_X1 U4409 ( .A(n3605), .B(n3606), .ZN(n3607) );
  NAND2_X1 U4410 ( .A1(n3607), .A2(n3823), .ZN(n3614) );
  AOI21_X1 U4411 ( .B1(n3609), .B2(n3828), .A(n3608), .ZN(n3613) );
  AOI22_X1 U4412 ( .A1(n4005), .A2(n3825), .B1(n3827), .B2(n3610), .ZN(n3612)
         );
  NAND2_X1 U4413 ( .A1(n3830), .A2(n3085), .ZN(n3611) );
  NAND4_X1 U4414 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(U3215)
         );
  INV_X1 U4415 ( .A(n3615), .ZN(n3618) );
  INV_X1 U4416 ( .A(n3617), .ZN(n3783) );
  NAND2_X1 U4417 ( .A1(n3615), .A2(n3783), .ZN(n3616) );
  AOI22_X1 U4418 ( .A1(n3618), .A2(n3617), .B1(n3616), .B2(n3784), .ZN(n3622)
         );
  NOR2_X1 U4419 ( .A1(n3620), .A2(n3619), .ZN(n3621) );
  XNOR2_X1 U4420 ( .A(n3622), .B(n3621), .ZN(n3623) );
  NAND2_X1 U4421 ( .A1(n3623), .A2(n3823), .ZN(n3631) );
  OAI22_X1 U4422 ( .A1(n3627), .A2(n3626), .B1(n3625), .B2(n3624), .ZN(n3628)
         );
  AOI211_X1 U4423 ( .C1(n3825), .C2(n4246), .A(n3629), .B(n3628), .ZN(n3630)
         );
  OAI211_X1 U4424 ( .C1(n3815), .C2(n3632), .A(n3631), .B(n3630), .ZN(U3216)
         );
  INV_X1 U4425 ( .A(n3634), .ZN(n3636) );
  NAND2_X1 U4426 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  XNOR2_X1 U4427 ( .A(n3633), .B(n3637), .ZN(n3638) );
  NAND2_X1 U4428 ( .A1(n3638), .A2(n3823), .ZN(n3646) );
  AOI21_X1 U4429 ( .B1(n4004), .B2(n3828), .A(n3639), .ZN(n3645) );
  AOI22_X1 U4430 ( .A1(n3641), .A2(n3825), .B1(n3827), .B2(n3640), .ZN(n3644)
         );
  NAND2_X1 U4431 ( .A1(n3830), .A2(n3642), .ZN(n3643) );
  NAND4_X1 U4432 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(U3218)
         );
  INV_X1 U4433 ( .A(n3647), .ZN(n3649) );
  NOR2_X1 U4434 ( .A1(n3649), .A2(n3648), .ZN(n3651) );
  AOI211_X1 U4435 ( .C1(n3741), .C2(n2035), .A(n3739), .B(n3651), .ZN(n3650)
         );
  AOI211_X1 U4436 ( .C1(n3652), .C2(n3651), .A(n3818), .B(n3650), .ZN(n3657)
         );
  AOI22_X1 U4437 ( .A1(n3997), .A2(n3825), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3654) );
  AOI22_X1 U4438 ( .A1(n4246), .A2(n3828), .B1(n4245), .B2(n3827), .ZN(n3653)
         );
  OAI211_X1 U4439 ( .C1(n3815), .C2(n3655), .A(n3654), .B(n3653), .ZN(n3656)
         );
  OR2_X1 U4440 ( .A1(n3657), .A2(n3656), .ZN(U3220) );
  INV_X1 U4441 ( .A(n3659), .ZN(n3661) );
  NAND2_X1 U4442 ( .A1(n3661), .A2(n3660), .ZN(n3662) );
  XNOR2_X1 U4443 ( .A(n3658), .B(n3662), .ZN(n3663) );
  NAND2_X1 U4444 ( .A1(n3663), .A2(n3823), .ZN(n3671) );
  AND2_X1 U4445 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4381) );
  AOI21_X1 U4446 ( .B1(n4001), .B2(n3828), .A(n4381), .ZN(n3670) );
  AOI22_X1 U4447 ( .A1(n3665), .A2(n3825), .B1(n3827), .B2(n3664), .ZN(n3669)
         );
  INV_X1 U4448 ( .A(n3666), .ZN(n3667) );
  NAND2_X1 U4449 ( .A1(n3830), .A2(n3667), .ZN(n3668) );
  NAND4_X1 U4450 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(U3221)
         );
  INV_X1 U4451 ( .A(n3672), .ZN(n3674) );
  NAND2_X1 U4452 ( .A1(n3674), .A2(n3673), .ZN(n3675) );
  XNOR2_X1 U4453 ( .A(n3676), .B(n3675), .ZN(n3682) );
  AOI22_X1 U4454 ( .A1(n3827), .A2(n4104), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3678) );
  NAND2_X1 U4455 ( .A1(n4139), .A2(n3828), .ZN(n3677) );
  OAI211_X1 U4456 ( .C1(n3679), .C2(n3711), .A(n3678), .B(n3677), .ZN(n3680)
         );
  AOI21_X1 U4457 ( .B1(n4107), .B2(n3830), .A(n3680), .ZN(n3681) );
  OAI21_X1 U4458 ( .B1(n3682), .B2(n3818), .A(n3681), .ZN(U3222) );
  OAI21_X1 U4459 ( .B1(n3683), .B2(n3821), .A(n3820), .ZN(n3684) );
  XOR2_X1 U4460 ( .A(n3685), .B(n3684), .Z(n3686) );
  NAND2_X1 U4461 ( .A1(n3686), .A2(n3823), .ZN(n3691) );
  AND2_X1 U4462 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4412) );
  AOI21_X1 U4463 ( .B1(n4275), .B2(n3825), .A(n4412), .ZN(n3690) );
  AOI22_X1 U4464 ( .A1(n4000), .A2(n3828), .B1(n3827), .B2(n4272), .ZN(n3689)
         );
  NAND2_X1 U4465 ( .A1(n3830), .A2(n3687), .ZN(n3688) );
  NAND4_X1 U4466 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(U3223)
         );
  INV_X1 U4467 ( .A(n3693), .ZN(n3695) );
  NAND2_X1 U4468 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  XNOR2_X1 U4469 ( .A(n3692), .B(n3696), .ZN(n3697) );
  NAND2_X1 U4470 ( .A1(n3697), .A2(n3823), .ZN(n3703) );
  AND2_X1 U4471 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4423) );
  AOI21_X1 U4472 ( .B1(n3998), .B2(n3825), .A(n4423), .ZN(n3702) );
  AOI22_X1 U4473 ( .A1(n3999), .A2(n3828), .B1(n3827), .B2(n3698), .ZN(n3701)
         );
  NAND2_X1 U4474 ( .A1(n3830), .A2(n3699), .ZN(n3700) );
  NAND4_X1 U4475 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(U3225)
         );
  INV_X1 U4476 ( .A(n3705), .ZN(n3706) );
  NOR2_X1 U4477 ( .A1(n3704), .A2(n3706), .ZN(n3708) );
  XNOR2_X1 U4478 ( .A(n3708), .B(n3707), .ZN(n3714) );
  AOI22_X1 U4479 ( .A1(n4228), .A2(n3828), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3710) );
  NAND2_X1 U4480 ( .A1(n3827), .A2(n4227), .ZN(n3709) );
  OAI211_X1 U4481 ( .C1(n4231), .C2(n3711), .A(n3710), .B(n3709), .ZN(n3712)
         );
  AOI21_X1 U4482 ( .B1(n4121), .B2(n3830), .A(n3712), .ZN(n3713) );
  OAI21_X1 U4483 ( .B1(n3714), .B2(n3818), .A(n3713), .ZN(U3226) );
  AOI21_X1 U4484 ( .B1(n3715), .B2(n3716), .A(n3818), .ZN(n3718) );
  NAND2_X1 U4485 ( .A1(n3718), .A2(n3717), .ZN(n3727) );
  INV_X1 U4486 ( .A(n3719), .ZN(n3720) );
  AOI21_X1 U4487 ( .B1(n4006), .B2(n3828), .A(n3720), .ZN(n3726) );
  AOI22_X1 U4488 ( .A1(n3801), .A2(n3825), .B1(n3827), .B2(n3721), .ZN(n3725)
         );
  INV_X1 U4489 ( .A(n3722), .ZN(n3723) );
  NAND2_X1 U4490 ( .A1(n3830), .A2(n3723), .ZN(n3724) );
  NAND4_X1 U4491 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(U3227)
         );
  XNOR2_X1 U4492 ( .A(n3728), .B(n3729), .ZN(n3730) );
  NAND2_X1 U4493 ( .A1(n3730), .A2(n3823), .ZN(n3738) );
  NOR2_X1 U4494 ( .A1(STATE_REG_SCAN_IN), .A2(n3731), .ZN(n4351) );
  AOI21_X1 U4495 ( .B1(n4002), .B2(n3825), .A(n4351), .ZN(n3737) );
  AOI22_X1 U4496 ( .A1(n4003), .A2(n3828), .B1(n3827), .B2(n3732), .ZN(n3736)
         );
  INV_X1 U4497 ( .A(n3733), .ZN(n3734) );
  NAND2_X1 U4498 ( .A1(n3830), .A2(n3734), .ZN(n3735) );
  NAND4_X1 U4499 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(U3228)
         );
  NAND2_X1 U4500 ( .A1(n2175), .A2(n2035), .ZN(n3740) );
  AOI22_X1 U4501 ( .A1(n3742), .A2(n2035), .B1(n3741), .B2(n3740), .ZN(n3749)
         );
  NAND2_X1 U4502 ( .A1(n4257), .A2(n3825), .ZN(n3745) );
  AOI22_X1 U4503 ( .A1(n4179), .A2(n3828), .B1(n3743), .B2(n3827), .ZN(n3744)
         );
  OAI211_X1 U4504 ( .C1(STATE_REG_SCAN_IN), .C2(n3746), .A(n3745), .B(n3744), 
        .ZN(n3747) );
  AOI21_X1 U4505 ( .B1(n4183), .B2(n3830), .A(n3747), .ZN(n3748) );
  OAI21_X1 U4506 ( .B1(n3749), .B2(n3818), .A(n3748), .ZN(U3230) );
  XOR2_X1 U4507 ( .A(n3751), .B(n3750), .Z(n3752) );
  XNOR2_X1 U4508 ( .A(n3753), .B(n3752), .ZN(n3754) );
  NAND2_X1 U4509 ( .A1(n3754), .A2(n3823), .ZN(n3762) );
  AOI21_X1 U4510 ( .B1(n3776), .B2(n3828), .A(n3755), .ZN(n3761) );
  AOI22_X1 U4511 ( .A1(n4291), .A2(n3825), .B1(n3827), .B2(n3756), .ZN(n3760)
         );
  INV_X1 U4512 ( .A(n3757), .ZN(n3758) );
  NAND2_X1 U4513 ( .A1(n3830), .A2(n3758), .ZN(n3759) );
  NAND4_X1 U4514 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(U3231)
         );
  OAI21_X1 U4515 ( .B1(n3764), .B2(n3763), .A(n3586), .ZN(n3765) );
  NAND2_X1 U4516 ( .A1(n3765), .A2(n3823), .ZN(n3769) );
  AOI22_X1 U4517 ( .A1(n4257), .A2(n3828), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3768) );
  AOI22_X1 U4518 ( .A1(n4228), .A2(n3825), .B1(n4155), .B2(n3827), .ZN(n3767)
         );
  NAND2_X1 U4519 ( .A1(n4161), .A2(n3830), .ZN(n3766) );
  NAND4_X1 U4520 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(U3232)
         );
  XNOR2_X1 U4521 ( .A(n3772), .B(n3771), .ZN(n3773) );
  XNOR2_X1 U4522 ( .A(n3770), .B(n3773), .ZN(n3774) );
  NAND2_X1 U4523 ( .A1(n3774), .A2(n3823), .ZN(n3782) );
  NOR2_X1 U4524 ( .A1(STATE_REG_SCAN_IN), .A2(n3775), .ZN(n4370) );
  AOI21_X1 U4525 ( .B1(n3776), .B2(n3825), .A(n4370), .ZN(n3781) );
  AOI22_X1 U4526 ( .A1(n4002), .A2(n3828), .B1(n3827), .B2(n3777), .ZN(n3780)
         );
  NAND2_X1 U4527 ( .A1(n3830), .A2(n3778), .ZN(n3779) );
  NAND4_X1 U4528 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(U3233)
         );
  XNOR2_X1 U4529 ( .A(n3784), .B(n3783), .ZN(n3785) );
  XNOR2_X1 U4530 ( .A(n3615), .B(n3785), .ZN(n3786) );
  NAND2_X1 U4531 ( .A1(n3786), .A2(n3823), .ZN(n3794) );
  AOI21_X1 U4532 ( .B1(n4179), .B2(n3825), .A(n3787), .ZN(n3793) );
  AOI22_X1 U4533 ( .A1(n4275), .A2(n3828), .B1(n3827), .B2(n3788), .ZN(n3792)
         );
  INV_X1 U4534 ( .A(n3789), .ZN(n3790) );
  NAND2_X1 U4535 ( .A1(n3830), .A2(n3790), .ZN(n3791) );
  NAND4_X1 U4536 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(U3235)
         );
  XNOR2_X1 U4537 ( .A(n3796), .B(n3795), .ZN(n3797) );
  XNOR2_X1 U4538 ( .A(n3798), .B(n3797), .ZN(n3799) );
  NAND2_X1 U4539 ( .A1(n3799), .A2(n3823), .ZN(n3807) );
  AOI21_X1 U4540 ( .B1(n3801), .B2(n3828), .A(n3800), .ZN(n3806) );
  AOI22_X1 U4541 ( .A1(n4004), .A2(n3825), .B1(n3827), .B2(n3802), .ZN(n3805)
         );
  NAND2_X1 U4542 ( .A1(n3830), .A2(n3803), .ZN(n3804) );
  NAND4_X1 U4543 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(U3236)
         );
  INV_X1 U4544 ( .A(n3809), .ZN(n3810) );
  NOR2_X1 U4545 ( .A1(n3811), .A2(n3810), .ZN(n3812) );
  XNOR2_X1 U4546 ( .A(n3808), .B(n3812), .ZN(n3819) );
  NAND2_X1 U4547 ( .A1(n4120), .A2(n3828), .ZN(n3814) );
  AOI22_X1 U4548 ( .A1(n3827), .A2(n4085), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3813) );
  OAI211_X1 U4549 ( .C1(n4083), .C2(n3815), .A(n3814), .B(n3813), .ZN(n3816)
         );
  AOI21_X1 U4550 ( .B1(n4080), .B2(n3825), .A(n3816), .ZN(n3817) );
  OAI21_X1 U4551 ( .B1(n3819), .B2(n3818), .A(n3817), .ZN(U3237) );
  NAND2_X1 U4552 ( .A1(n2165), .A2(n3820), .ZN(n3822) );
  XNOR2_X1 U4553 ( .A(n3822), .B(n3821), .ZN(n3824) );
  NAND2_X1 U4554 ( .A1(n3824), .A2(n3823), .ZN(n3834) );
  AND2_X1 U4555 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4405) );
  AOI21_X1 U4556 ( .B1(n3999), .B2(n3825), .A(n4405), .ZN(n3833) );
  AOI22_X1 U4557 ( .A1(n4291), .A2(n3828), .B1(n3827), .B2(n3826), .ZN(n3832)
         );
  NAND2_X1 U4558 ( .A1(n3830), .A2(n3829), .ZN(n3831) );
  NAND4_X1 U4559 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(U3238)
         );
  INV_X1 U4560 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4561 ( .A1(n2418), .A2(REG2_REG_31__SCAN_IN), .ZN(n3836) );
  NAND2_X1 U4562 ( .A1(n3838), .A2(REG0_REG_31__SCAN_IN), .ZN(n3835) );
  OAI211_X1 U4563 ( .C1(n3842), .C2(n3837), .A(n3836), .B(n3835), .ZN(n4194)
         );
  NAND2_X1 U4564 ( .A1(n3906), .A2(DATAI_31_), .ZN(n4195) );
  AND2_X1 U4565 ( .A1(n4194), .A2(n4195), .ZN(n3917) );
  INV_X1 U4566 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4567 ( .A1(n2418), .A2(REG2_REG_30__SCAN_IN), .ZN(n3840) );
  NAND2_X1 U4568 ( .A1(n3838), .A2(REG0_REG_30__SCAN_IN), .ZN(n3839) );
  OAI211_X1 U4569 ( .C1(n3842), .C2(n3841), .A(n3840), .B(n3839), .ZN(n4042)
         );
  NAND2_X1 U4570 ( .A1(n3906), .A2(DATAI_30_), .ZN(n4199) );
  NAND2_X1 U4571 ( .A1(n4042), .A2(n4199), .ZN(n3976) );
  OR2_X1 U4572 ( .A1(n4194), .A2(n4195), .ZN(n3843) );
  AND2_X1 U4573 ( .A1(n3976), .A2(n3843), .ZN(n3938) );
  INV_X1 U4574 ( .A(n3844), .ZN(n3847) );
  OAI211_X1 U4575 ( .C1(n3847), .C2(n4334), .A(n3846), .B(n3845), .ZN(n3849)
         );
  NAND3_X1 U4576 ( .A1(n3849), .A2(n3848), .A3(n2661), .ZN(n3852) );
  NAND3_X1 U4577 ( .A1(n3852), .A2(n3851), .A3(n3850), .ZN(n3855) );
  NAND3_X1 U4578 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n3863) );
  INV_X1 U4579 ( .A(n3856), .ZN(n3858) );
  NOR3_X1 U4580 ( .A1(n3877), .A2(n3858), .A3(n3857), .ZN(n3862) );
  INV_X1 U4581 ( .A(n3859), .ZN(n3861) );
  AOI211_X1 U4582 ( .C1(n3863), .C2(n3862), .A(n3861), .B(n3860), .ZN(n3868)
         );
  NAND2_X1 U4583 ( .A1(n3865), .A2(n3864), .ZN(n3876) );
  OAI211_X1 U4584 ( .C1(n3868), .C2(n3876), .A(n3867), .B(n3866), .ZN(n3873)
         );
  NAND2_X1 U4585 ( .A1(n3870), .A2(n3869), .ZN(n3879) );
  INV_X1 U4586 ( .A(n3879), .ZN(n3872) );
  NAND3_X1 U4587 ( .A1(n3873), .A2(n3872), .A3(n3871), .ZN(n3887) );
  NOR4_X1 U4588 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3881)
         );
  INV_X1 U4589 ( .A(n3878), .ZN(n3880) );
  NAND2_X1 U4590 ( .A1(n3879), .A2(n3888), .ZN(n3953) );
  OAI21_X1 U4591 ( .B1(n3881), .B2(n3880), .A(n3953), .ZN(n3886) );
  INV_X1 U4592 ( .A(n3882), .ZN(n3885) );
  INV_X1 U4593 ( .A(n3883), .ZN(n3884) );
  AOI211_X1 U4594 ( .C1(n3887), .C2(n3886), .A(n3885), .B(n3884), .ZN(n3894)
         );
  NAND2_X1 U4595 ( .A1(n3889), .A2(n3888), .ZN(n3954) );
  INV_X1 U4596 ( .A(n3954), .ZN(n3891) );
  INV_X1 U4597 ( .A(n3953), .ZN(n3890) );
  AOI21_X1 U4598 ( .B1(n3892), .B2(n3891), .A(n3890), .ZN(n3893) );
  OAI21_X1 U4599 ( .B1(n3894), .B2(n3893), .A(n3956), .ZN(n3896) );
  AOI21_X1 U4600 ( .B1(n3896), .B2(n3958), .A(n3895), .ZN(n3900) );
  INV_X1 U4601 ( .A(n3897), .ZN(n3899) );
  OAI21_X1 U4602 ( .B1(n3900), .B2(n3899), .A(n3898), .ZN(n3902) );
  AOI21_X1 U4603 ( .B1(n3903), .B2(n3902), .A(n3901), .ZN(n3905) );
  INV_X1 U4604 ( .A(n3964), .ZN(n3904) );
  OAI21_X1 U4605 ( .B1(n3905), .B2(n3904), .A(n3971), .ZN(n3910) );
  NAND2_X1 U4606 ( .A1(n3906), .A2(DATAI_29_), .ZN(n4041) );
  NAND2_X1 U4607 ( .A1(n3996), .A2(n4041), .ZN(n3918) );
  NAND2_X1 U4608 ( .A1(n3918), .A2(n4037), .ZN(n3914) );
  NOR2_X1 U4609 ( .A1(n3907), .A2(n3914), .ZN(n3975) );
  INV_X1 U4610 ( .A(n3975), .ZN(n3908) );
  AOI211_X1 U4611 ( .C1(n3969), .C2(n3910), .A(n3909), .B(n3908), .ZN(n3915)
         );
  INV_X1 U4612 ( .A(n3911), .ZN(n3912) );
  NOR2_X1 U4613 ( .A1(n4036), .A2(n3912), .ZN(n3967) );
  INV_X1 U4614 ( .A(n4042), .ZN(n3913) );
  INV_X1 U4615 ( .A(n4199), .ZN(n4203) );
  AOI21_X1 U4616 ( .B1(n3913), .B2(n4203), .A(n3917), .ZN(n3968) );
  OR2_X1 U4617 ( .A1(n3996), .A2(n4041), .ZN(n3966) );
  OAI211_X1 U4618 ( .C1(n3967), .C2(n3914), .A(n3968), .B(n3966), .ZN(n3973)
         );
  OR2_X1 U4619 ( .A1(n3915), .A2(n3973), .ZN(n3916) );
  OAI21_X1 U4620 ( .B1(n3917), .B2(n3938), .A(n3916), .ZN(n3985) );
  NAND2_X1 U4621 ( .A1(n3966), .A2(n3918), .ZN(n4051) );
  INV_X1 U4622 ( .A(n4450), .ZN(n3919) );
  NAND4_X1 U4623 ( .A1(n4133), .A2(n2462), .A3(n3919), .A4(n3968), .ZN(n3923)
         );
  INV_X1 U4624 ( .A(n3920), .ZN(n3922) );
  OR4_X1 U4625 ( .A1(n3923), .A2(n4153), .A3(n3922), .A4(n3921), .ZN(n3952) );
  NOR4_X1 U4626 ( .A1(n3926), .A2(n2660), .A3(n3925), .A4(n3924), .ZN(n3951)
         );
  NOR4_X1 U4627 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3950)
         );
  NOR4_X1 U4628 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3949)
         );
  AND2_X1 U4629 ( .A1(n4074), .A2(n3937), .ZN(n4095) );
  AND4_X1 U4630 ( .A1(n3974), .A2(n4077), .A3(n4095), .A4(n3938), .ZN(n3945)
         );
  INV_X1 U4631 ( .A(n3939), .ZN(n3941) );
  AND2_X1 U4632 ( .A1(n3941), .A2(n3940), .ZN(n4175) );
  XNOR2_X1 U4633 ( .A(n4228), .B(n4143), .ZN(n4136) );
  NAND2_X1 U4634 ( .A1(n4093), .A2(n3942), .ZN(n4117) );
  NOR4_X1 U4635 ( .A1(n4175), .A2(n3943), .A3(n4136), .A4(n4117), .ZN(n3944)
         );
  OAI21_X1 U4636 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n3959) );
  INV_X1 U4637 ( .A(n3956), .ZN(n3957) );
  AOI21_X1 U4638 ( .B1(n3959), .B2(n3958), .A(n3957), .ZN(n3963) );
  INV_X1 U4639 ( .A(n3960), .ZN(n3962) );
  OAI21_X1 U4640 ( .B1(n3963), .B2(n3962), .A(n3961), .ZN(n3965) );
  NAND2_X1 U4641 ( .A1(n3965), .A2(n3964), .ZN(n3972) );
  NAND4_X1 U4642 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  AOI21_X1 U4643 ( .B1(n3972), .B2(n3971), .A(n3970), .ZN(n3979) );
  AOI21_X1 U4644 ( .B1(n3975), .B2(n3974), .A(n3973), .ZN(n3978) );
  AOI21_X1 U4645 ( .B1(n3976), .B2(n4194), .A(n4195), .ZN(n3977) );
  NOR3_X1 U4646 ( .A1(n3979), .A2(n3978), .A3(n3977), .ZN(n3980) );
  AOI21_X1 U4647 ( .B1(n4203), .B2(n4195), .A(n3980), .ZN(n3981) );
  MUX2_X1 U4648 ( .A(n3982), .B(n3981), .S(n4334), .Z(n3984) );
  MUX2_X1 U4649 ( .A(n3985), .B(n3984), .S(n3983), .Z(n3987) );
  XNOR2_X1 U4650 ( .A(n3987), .B(n3986), .ZN(n3995) );
  INV_X1 U4651 ( .A(n3988), .ZN(n3994) );
  NAND2_X1 U4652 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  OAI211_X1 U4653 ( .C1(n3992), .C2(n3994), .A(n3991), .B(B_REG_SCAN_IN), .ZN(
        n3993) );
  OAI21_X1 U4654 ( .B1(n3995), .B2(n3994), .A(n3993), .ZN(U3239) );
  MUX2_X1 U4655 ( .A(DATAO_REG_31__SCAN_IN), .B(n4194), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4656 ( .A(DATAO_REG_30__SCAN_IN), .B(n4042), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4657 ( .A(DATAO_REG_29__SCAN_IN), .B(n3996), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4658 ( .A(DATAO_REG_28__SCAN_IN), .B(n4212), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4659 ( .A(DATAO_REG_27__SCAN_IN), .B(n4080), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4660 ( .A(DATAO_REG_26__SCAN_IN), .B(n4211), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4661 ( .A(n4139), .B(DATAO_REG_24__SCAN_IN), .S(n4007), .Z(U3574)
         );
  MUX2_X1 U4662 ( .A(DATAO_REG_23__SCAN_IN), .B(n4228), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4663 ( .A(n3997), .B(DATAO_REG_22__SCAN_IN), .S(n4007), .Z(U3572)
         );
  MUX2_X1 U4664 ( .A(DATAO_REG_21__SCAN_IN), .B(n4257), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4665 ( .A(n4246), .B(DATAO_REG_20__SCAN_IN), .S(n4007), .Z(U3570)
         );
  MUX2_X1 U4666 ( .A(n4179), .B(DATAO_REG_19__SCAN_IN), .S(n4007), .Z(U3569)
         );
  MUX2_X1 U4667 ( .A(n3998), .B(DATAO_REG_18__SCAN_IN), .S(n4007), .Z(U3568)
         );
  MUX2_X1 U4668 ( .A(n4275), .B(DATAO_REG_17__SCAN_IN), .S(n4007), .Z(U3567)
         );
  MUX2_X1 U4669 ( .A(n3999), .B(DATAO_REG_16__SCAN_IN), .S(n4007), .Z(U3566)
         );
  MUX2_X1 U4670 ( .A(n4000), .B(DATAO_REG_15__SCAN_IN), .S(n4007), .Z(U3565)
         );
  MUX2_X1 U4671 ( .A(n4001), .B(DATAO_REG_11__SCAN_IN), .S(n4007), .Z(U3561)
         );
  MUX2_X1 U4672 ( .A(n4002), .B(DATAO_REG_10__SCAN_IN), .S(n4007), .Z(U3560)
         );
  MUX2_X1 U4673 ( .A(n4003), .B(DATAO_REG_8__SCAN_IN), .S(n4007), .Z(U3558) );
  MUX2_X1 U4674 ( .A(n4004), .B(DATAO_REG_7__SCAN_IN), .S(n4007), .Z(U3557) );
  MUX2_X1 U4675 ( .A(n4005), .B(DATAO_REG_4__SCAN_IN), .S(n4007), .Z(U3554) );
  MUX2_X1 U4676 ( .A(n4006), .B(DATAO_REG_3__SCAN_IN), .S(n4007), .Z(U3553) );
  MUX2_X1 U4677 ( .A(n2407), .B(DATAO_REG_1__SCAN_IN), .S(n4007), .Z(U3551) );
  MUX2_X1 U4678 ( .A(n4008), .B(DATAO_REG_0__SCAN_IN), .S(n4007), .Z(U3550) );
  AOI22_X1 U4679 ( .A1(n4424), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4022) );
  NAND2_X1 U4680 ( .A1(n4396), .A2(n4009), .ZN(n4021) );
  MUX2_X1 U4681 ( .A(REG1_REG_1__SCAN_IN), .B(n4512), .S(n4010), .Z(n4011) );
  OAI21_X1 U4682 ( .B1(n2045), .B2(n4012), .A(n4011), .ZN(n4013) );
  NAND3_X1 U4683 ( .A1(n4434), .A2(n4014), .A3(n4013), .ZN(n4020) );
  INV_X1 U4684 ( .A(n4015), .ZN(n4016) );
  OAI211_X1 U4685 ( .C1(n4018), .C2(n4017), .A(n4432), .B(n4016), .ZN(n4019)
         );
  NAND4_X1 U4686 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(U3241)
         );
  AOI22_X1 U4687 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4424), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4033) );
  AOI211_X1 U4688 ( .C1(n4025), .C2(n4024), .A(n4023), .B(n4389), .ZN(n4031)
         );
  XNOR2_X1 U4689 ( .A(n4027), .B(n4026), .ZN(n4029) );
  OAI22_X1 U4690 ( .A1(n4029), .A2(n4400), .B1(n4437), .B2(n4028), .ZN(n4030)
         );
  NOR2_X1 U4691 ( .A1(n4031), .A2(n4030), .ZN(n4032) );
  NAND3_X1 U4692 ( .A1(n4034), .A2(n4033), .A3(n4032), .ZN(U3242) );
  INV_X1 U4693 ( .A(n4035), .ZN(n4046) );
  AOI21_X1 U4694 ( .B1(n4038), .B2(n4037), .A(n4036), .ZN(n4039) );
  XOR2_X1 U4695 ( .A(n4051), .B(n4039), .Z(n4045) );
  AOI21_X1 U4696 ( .B1(n4040), .B2(B_REG_SCAN_IN), .A(n4286), .ZN(n4193) );
  INV_X1 U4697 ( .A(n4041), .ZN(n4054) );
  AOI22_X1 U4698 ( .A1(n4042), .A2(n4193), .B1(n4273), .B2(n4054), .ZN(n4044)
         );
  NAND2_X1 U4699 ( .A1(n4212), .A2(n4292), .ZN(n4043) );
  OAI211_X1 U4700 ( .C1(n4045), .C2(n4259), .A(n4044), .B(n4043), .ZN(n4206)
         );
  AOI21_X1 U4701 ( .B1(n4046), .B2(n4448), .A(n4206), .ZN(n4057) );
  XNOR2_X1 U4702 ( .A(n4052), .B(n4051), .ZN(n4205) );
  NAND2_X1 U4703 ( .A1(n4205), .A2(n4176), .ZN(n4056) );
  AOI21_X1 U4704 ( .B1(n4054), .B2(n4053), .A(n4200), .ZN(n4207) );
  AOI22_X1 U4705 ( .A1(n4207), .A2(n4439), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4182), .ZN(n4055) );
  OAI211_X1 U4706 ( .C1(n4182), .C2(n4057), .A(n4056), .B(n4055), .ZN(U3354)
         );
  XNOR2_X1 U4707 ( .A(n4058), .B(n4059), .ZN(n4218) );
  INV_X1 U4708 ( .A(n4218), .ZN(n4072) );
  XNOR2_X1 U4709 ( .A(n4060), .B(n4059), .ZN(n4061) );
  OR2_X1 U4710 ( .A1(n4084), .A2(n4062), .ZN(n4063) );
  NAND2_X1 U4711 ( .A1(n4064), .A2(n4063), .ZN(n4215) );
  NAND2_X1 U4712 ( .A1(n4211), .A2(n4180), .ZN(n4066) );
  AOI22_X1 U4713 ( .A1(n4119), .A2(n4210), .B1(n4182), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4065) );
  OAI211_X1 U4714 ( .C1(n4145), .C2(n4067), .A(n4066), .B(n4065), .ZN(n4068)
         );
  AOI21_X1 U4715 ( .B1(n4181), .B2(n4212), .A(n4068), .ZN(n4069) );
  OAI21_X1 U4716 ( .B1(n4215), .B2(n4164), .A(n4069), .ZN(n4070) );
  AOI21_X1 U4717 ( .B1(n4217), .B2(n2999), .A(n4070), .ZN(n4071) );
  OAI21_X1 U4718 ( .B1(n4072), .B2(n4169), .A(n4071), .ZN(U3263) );
  XNOR2_X1 U4719 ( .A(n4073), .B(n4077), .ZN(n4221) );
  INV_X1 U4720 ( .A(n4221), .ZN(n4091) );
  NAND2_X1 U4721 ( .A1(n4075), .A2(n4074), .ZN(n4076) );
  XOR2_X1 U4722 ( .A(n4077), .B(n4076), .Z(n4082) );
  OAI22_X1 U4723 ( .A1(n4231), .A2(n4277), .B1(n4078), .B2(n4285), .ZN(n4079)
         );
  AOI21_X1 U4724 ( .B1(n4080), .B2(n4274), .A(n4079), .ZN(n4081) );
  OAI21_X1 U4725 ( .B1(n4082), .B2(n4259), .A(n4081), .ZN(n4220) );
  OAI22_X1 U4726 ( .A1(n4083), .A2(n4145), .B1(n4620), .B2(n2999), .ZN(n4089)
         );
  INV_X1 U4727 ( .A(n4084), .ZN(n4087) );
  NAND2_X1 U4728 ( .A1(n4106), .A2(n4085), .ZN(n4086) );
  NAND2_X1 U4729 ( .A1(n4087), .A2(n4086), .ZN(n4307) );
  NOR2_X1 U4730 ( .A1(n4307), .A2(n4164), .ZN(n4088) );
  AOI211_X1 U4731 ( .C1(n2999), .C2(n4220), .A(n4089), .B(n4088), .ZN(n4090)
         );
  OAI21_X1 U4732 ( .B1(n4091), .B2(n4169), .A(n4090), .ZN(U3264) );
  XNOR2_X1 U4733 ( .A(n4092), .B(n4095), .ZN(n4224) );
  INV_X1 U4734 ( .A(n4224), .ZN(n4111) );
  NAND2_X1 U4735 ( .A1(n4094), .A2(n4093), .ZN(n4097) );
  INV_X1 U4736 ( .A(n4095), .ZN(n4096) );
  XNOR2_X1 U4737 ( .A(n4097), .B(n4096), .ZN(n4098) );
  NAND2_X1 U4738 ( .A1(n4098), .A2(n4159), .ZN(n4103) );
  OAI22_X1 U4739 ( .A1(n4100), .A2(n4277), .B1(n4099), .B2(n4285), .ZN(n4101)
         );
  AOI21_X1 U4740 ( .B1(n4211), .B2(n4274), .A(n4101), .ZN(n4102) );
  NAND2_X1 U4741 ( .A1(n4103), .A2(n4102), .ZN(n4223) );
  NAND2_X1 U4742 ( .A1(n2012), .A2(n4104), .ZN(n4105) );
  NAND2_X1 U4743 ( .A1(n4106), .A2(n4105), .ZN(n4311) );
  AOI22_X1 U4744 ( .A1(n4107), .A2(n4448), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4182), .ZN(n4108) );
  OAI21_X1 U4745 ( .B1(n4311), .B2(n4164), .A(n4108), .ZN(n4109) );
  AOI21_X1 U4746 ( .B1(n4223), .B2(n2999), .A(n4109), .ZN(n4110) );
  OAI21_X1 U4747 ( .B1(n4111), .B2(n4169), .A(n4110), .ZN(U3265) );
  NAND2_X1 U4748 ( .A1(n4113), .A2(n4112), .ZN(n4114) );
  XOR2_X1 U4749 ( .A(n4117), .B(n4114), .Z(n4115) );
  NAND2_X1 U4750 ( .A1(n4115), .A2(n4159), .ZN(n4230) );
  XNOR2_X1 U4751 ( .A(n4116), .B(n4117), .ZN(n4233) );
  NAND2_X1 U4752 ( .A1(n4233), .A2(n4176), .ZN(n4129) );
  NAND2_X1 U4753 ( .A1(n4142), .A2(n4227), .ZN(n4118) );
  NAND2_X1 U4754 ( .A1(n2012), .A2(n4118), .ZN(n4315) );
  INV_X1 U4755 ( .A(n4315), .ZN(n4127) );
  INV_X1 U4756 ( .A(n4180), .ZN(n4124) );
  AOI22_X1 U4757 ( .A1(n4120), .A2(n4181), .B1(n4119), .B2(n4227), .ZN(n4123)
         );
  AOI22_X1 U4758 ( .A1(n4121), .A2(n4448), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4182), .ZN(n4122) );
  OAI211_X1 U4759 ( .C1(n4125), .C2(n4124), .A(n4123), .B(n4122), .ZN(n4126)
         );
  AOI21_X1 U4760 ( .B1(n4127), .B2(n4439), .A(n4126), .ZN(n4128) );
  OAI211_X1 U4761 ( .C1(n4182), .C2(n4230), .A(n4129), .B(n4128), .ZN(U3266)
         );
  XOR2_X1 U4762 ( .A(n4136), .B(n4130), .Z(n4237) );
  INV_X1 U4763 ( .A(n4237), .ZN(n4150) );
  INV_X1 U4764 ( .A(n4131), .ZN(n4132) );
  AOI21_X1 U4765 ( .B1(n4134), .B2(n4133), .A(n4132), .ZN(n4154) );
  OAI21_X1 U4766 ( .B1(n4154), .B2(n4153), .A(n4135), .ZN(n4137) );
  XNOR2_X1 U4767 ( .A(n4137), .B(n4136), .ZN(n4141) );
  OAI22_X1 U4768 ( .A1(n4248), .A2(n4277), .B1(n4285), .B2(n4143), .ZN(n4138)
         );
  AOI21_X1 U4769 ( .B1(n4139), .B2(n4274), .A(n4138), .ZN(n4140) );
  OAI21_X1 U4770 ( .B1(n4141), .B2(n4259), .A(n4140), .ZN(n4236) );
  OAI21_X1 U4771 ( .B1(n4241), .B2(n4143), .A(n4142), .ZN(n4319) );
  NOR2_X1 U4772 ( .A1(n4319), .A2(n4164), .ZN(n4148) );
  INV_X1 U4773 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4144) );
  OAI22_X1 U4774 ( .A1(n4146), .A2(n4145), .B1(n4144), .B2(n2999), .ZN(n4147)
         );
  AOI211_X1 U4775 ( .C1(n4236), .C2(n2999), .A(n4148), .B(n4147), .ZN(n4149)
         );
  OAI21_X1 U4776 ( .B1(n4150), .B2(n4169), .A(n4149), .ZN(U3267) );
  OAI21_X1 U4777 ( .B1(n4152), .B2(n4153), .A(n4151), .ZN(n4244) );
  XNOR2_X1 U4778 ( .A(n4154), .B(n4153), .ZN(n4160) );
  NAND2_X1 U4779 ( .A1(n4228), .A2(n4274), .ZN(n4157) );
  AOI22_X1 U4780 ( .A1(n4257), .A2(n4292), .B1(n4155), .B2(n4273), .ZN(n4156)
         );
  NAND2_X1 U4781 ( .A1(n4157), .A2(n4156), .ZN(n4158) );
  AOI21_X1 U4782 ( .B1(n4160), .B2(n4159), .A(n4158), .ZN(n4243) );
  AOI22_X1 U4783 ( .A1(n4161), .A2(n4448), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4182), .ZN(n4166) );
  NOR2_X1 U4784 ( .A1(n4163), .A2(n4162), .ZN(n4240) );
  OR3_X1 U4785 ( .A1(n4241), .A2(n4240), .A3(n4164), .ZN(n4165) );
  OAI211_X1 U4786 ( .C1(n4243), .C2(n4182), .A(n4166), .B(n4165), .ZN(n4167)
         );
  INV_X1 U4787 ( .A(n4167), .ZN(n4168) );
  OAI21_X1 U4788 ( .B1(n4244), .B2(n4169), .A(n4168), .ZN(U3268) );
  INV_X1 U4789 ( .A(n4170), .ZN(n4171) );
  NAND2_X1 U4790 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  XNOR2_X1 U4791 ( .A(n4173), .B(n4175), .ZN(n4260) );
  XOR2_X1 U4792 ( .A(n4175), .B(n4174), .Z(n4262) );
  NAND2_X1 U4793 ( .A1(n4262), .A2(n4176), .ZN(n4190) );
  INV_X1 U4794 ( .A(n3332), .ZN(n4178) );
  OAI21_X1 U4795 ( .B1(n4178), .B2(n4254), .A(n4177), .ZN(n4325) );
  INV_X1 U4796 ( .A(n4325), .ZN(n4188) );
  AOI22_X1 U4797 ( .A1(n4257), .A2(n4181), .B1(n4180), .B2(n4179), .ZN(n4185)
         );
  AOI22_X1 U4798 ( .A1(n4183), .A2(n4448), .B1(REG2_REG_20__SCAN_IN), .B2(
        n4182), .ZN(n4184) );
  OAI211_X1 U4799 ( .C1(n4254), .C2(n4186), .A(n4185), .B(n4184), .ZN(n4187)
         );
  AOI21_X1 U4800 ( .B1(n4188), .B2(n4439), .A(n4187), .ZN(n4189) );
  OAI211_X1 U4801 ( .C1(n4260), .C2(n4191), .A(n4190), .B(n4189), .ZN(U3270)
         );
  NAND2_X1 U4802 ( .A1(n4200), .A2(n4199), .ZN(n4198) );
  XNOR2_X1 U4803 ( .A(n4198), .B(n4195), .ZN(n4343) );
  NAND2_X1 U4804 ( .A1(n4343), .A2(n4192), .ZN(n4197) );
  NAND2_X1 U4805 ( .A1(n4194), .A2(n4193), .ZN(n4201) );
  OAI21_X1 U4806 ( .B1(n4195), .B2(n4285), .A(n4201), .ZN(n4342) );
  NAND2_X1 U4807 ( .A1(n4342), .A2(n4518), .ZN(n4196) );
  OAI211_X1 U4808 ( .C1(n4518), .C2(n3837), .A(n4197), .B(n4196), .ZN(U3549)
         );
  OAI21_X1 U4809 ( .B1(n4200), .B2(n4199), .A(n4198), .ZN(n4345) );
  INV_X1 U4810 ( .A(n4201), .ZN(n4202) );
  AOI21_X1 U4811 ( .B1(n4203), .B2(n4273), .A(n4202), .ZN(n4348) );
  MUX2_X1 U4812 ( .A(n3841), .B(n4348), .S(n4518), .Z(n4204) );
  OAI21_X1 U4813 ( .B1(n4345), .B2(n4268), .A(n4204), .ZN(U3548) );
  NAND2_X1 U4814 ( .A1(n4205), .A2(n4502), .ZN(n4209) );
  NAND2_X1 U4815 ( .A1(n4209), .A2(n4208), .ZN(n4302) );
  MUX2_X1 U4816 ( .A(REG1_REG_29__SCAN_IN), .B(n4302), .S(n4518), .Z(U3547) );
  AOI22_X1 U4817 ( .A1(n4211), .A2(n4292), .B1(n4210), .B2(n4273), .ZN(n4214)
         );
  NAND2_X1 U4818 ( .A1(n4212), .A2(n4274), .ZN(n4213) );
  OAI211_X1 U4819 ( .C1(n4215), .C2(n4478), .A(n4214), .B(n4213), .ZN(n4216)
         );
  AOI211_X1 U4820 ( .C1(n4218), .C2(n4502), .A(n4217), .B(n4216), .ZN(n4219)
         );
  INV_X1 U4821 ( .A(n4219), .ZN(n4303) );
  MUX2_X1 U4822 ( .A(REG1_REG_27__SCAN_IN), .B(n4303), .S(n4518), .Z(U3545) );
  AOI21_X1 U4823 ( .B1(n4221), .B2(n4502), .A(n4220), .ZN(n4304) );
  MUX2_X1 U4824 ( .A(n4580), .B(n4304), .S(n4518), .Z(n4222) );
  OAI21_X1 U4825 ( .B1(n4268), .B2(n4307), .A(n4222), .ZN(U3544) );
  AOI21_X1 U4826 ( .B1(n4224), .B2(n4502), .A(n4223), .ZN(n4308) );
  MUX2_X1 U4827 ( .A(n4225), .B(n4308), .S(n4521), .Z(n4226) );
  OAI21_X1 U4828 ( .B1(n4268), .B2(n4311), .A(n4226), .ZN(U3543) );
  AOI22_X1 U4829 ( .A1(n4228), .A2(n4292), .B1(n4273), .B2(n4227), .ZN(n4229)
         );
  OAI211_X1 U4830 ( .C1(n4231), .C2(n4286), .A(n4230), .B(n4229), .ZN(n4232)
         );
  AOI21_X1 U4831 ( .B1(n4233), .B2(n4502), .A(n4232), .ZN(n4312) );
  MUX2_X1 U4832 ( .A(n4234), .B(n4312), .S(n4521), .Z(n4235) );
  OAI21_X1 U4833 ( .B1(n4268), .B2(n4315), .A(n4235), .ZN(U3542) );
  AOI21_X1 U4834 ( .B1(n4237), .B2(n4502), .A(n4236), .ZN(n4316) );
  MUX2_X1 U4835 ( .A(n4238), .B(n4316), .S(n4521), .Z(n4239) );
  OAI21_X1 U4836 ( .B1(n4268), .B2(n4319), .A(n4239), .ZN(U3541) );
  OR3_X1 U4837 ( .A1(n4241), .A2(n4240), .A3(n4478), .ZN(n4242) );
  OAI211_X1 U4838 ( .C1(n4244), .C2(n4490), .A(n4243), .B(n4242), .ZN(n4320)
         );
  MUX2_X1 U4839 ( .A(REG1_REG_22__SCAN_IN), .B(n4320), .S(n4521), .Z(U3540) );
  AOI22_X1 U4840 ( .A1(n4246), .A2(n4292), .B1(n4245), .B2(n4273), .ZN(n4247)
         );
  OAI21_X1 U4841 ( .B1(n4248), .B2(n4286), .A(n4247), .ZN(n4249) );
  AOI21_X1 U4842 ( .B1(n4250), .B2(n4504), .A(n4249), .ZN(n4252) );
  OAI211_X1 U4843 ( .C1(n4253), .C2(n4490), .A(n4252), .B(n4251), .ZN(n4321)
         );
  MUX2_X1 U4844 ( .A(REG1_REG_21__SCAN_IN), .B(n4321), .S(n4521), .Z(U3539) );
  OAI22_X1 U4845 ( .A1(n4255), .A2(n4277), .B1(n4254), .B2(n4285), .ZN(n4256)
         );
  AOI21_X1 U4846 ( .B1(n4274), .B2(n4257), .A(n4256), .ZN(n4258) );
  OAI21_X1 U4847 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(n4261) );
  AOI21_X1 U4848 ( .B1(n4262), .B2(n4502), .A(n4261), .ZN(n4322) );
  MUX2_X1 U4849 ( .A(n4578), .B(n4322), .S(n4521), .Z(n4263) );
  OAI21_X1 U4850 ( .B1(n4268), .B2(n4325), .A(n4263), .ZN(U3538) );
  AOI21_X1 U4851 ( .B1(n4265), .B2(n4502), .A(n4264), .ZN(n4326) );
  MUX2_X1 U4852 ( .A(n4266), .B(n4326), .S(n4521), .Z(n4267) );
  OAI21_X1 U4853 ( .B1(n4268), .B2(n4330), .A(n4267), .ZN(U3537) );
  OAI211_X1 U4854 ( .C1(n4271), .C2(n4490), .A(n4270), .B(n4269), .ZN(n4331)
         );
  MUX2_X1 U4855 ( .A(REG1_REG_18__SCAN_IN), .B(n4331), .S(n4521), .Z(U3536) );
  AOI22_X1 U4856 ( .A1(n4275), .A2(n4274), .B1(n4273), .B2(n4272), .ZN(n4276)
         );
  OAI21_X1 U4857 ( .B1(n4278), .B2(n4277), .A(n4276), .ZN(n4279) );
  AOI21_X1 U4858 ( .B1(n4280), .B2(n4504), .A(n4279), .ZN(n4282) );
  OAI211_X1 U4859 ( .C1(n4283), .C2(n4490), .A(n4282), .B(n4281), .ZN(n4332)
         );
  MUX2_X1 U4860 ( .A(REG1_REG_16__SCAN_IN), .B(n4332), .S(n4521), .Z(U3534) );
  OAI22_X1 U4861 ( .A1(n4287), .A2(n4286), .B1(n4285), .B2(n4284), .ZN(n4290)
         );
  NOR2_X1 U4862 ( .A1(n4288), .A2(n4478), .ZN(n4289) );
  AOI211_X1 U4863 ( .C1(n4292), .C2(n4291), .A(n4290), .B(n4289), .ZN(n4294)
         );
  OAI211_X1 U4864 ( .C1(n4295), .C2(n4490), .A(n4294), .B(n4293), .ZN(n4333)
         );
  MUX2_X1 U4865 ( .A(REG1_REG_15__SCAN_IN), .B(n4333), .S(n4521), .Z(U3533) );
  INV_X1 U4866 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4299) );
  NAND2_X1 U4867 ( .A1(n4343), .A2(n4296), .ZN(n4298) );
  NAND2_X1 U4868 ( .A1(n4342), .A2(n4511), .ZN(n4297) );
  OAI211_X1 U4869 ( .C1(n4511), .C2(n4299), .A(n4298), .B(n4297), .ZN(U3517)
         );
  INV_X1 U4870 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4300) );
  MUX2_X1 U4871 ( .A(n4300), .B(n4348), .S(n4511), .Z(n4301) );
  OAI21_X1 U4872 ( .B1(n4345), .B2(n4329), .A(n4301), .ZN(U3516) );
  MUX2_X1 U4873 ( .A(REG0_REG_29__SCAN_IN), .B(n4302), .S(n4511), .Z(U3515) );
  MUX2_X1 U4874 ( .A(REG0_REG_27__SCAN_IN), .B(n4303), .S(n4511), .Z(U3513) );
  INV_X1 U4875 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4305) );
  MUX2_X1 U4876 ( .A(n4305), .B(n4304), .S(n4511), .Z(n4306) );
  OAI21_X1 U4877 ( .B1(n4307), .B2(n4329), .A(n4306), .ZN(U3512) );
  INV_X1 U4878 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4309) );
  MUX2_X1 U4879 ( .A(n4309), .B(n4308), .S(n4511), .Z(n4310) );
  OAI21_X1 U4880 ( .B1(n4311), .B2(n4329), .A(n4310), .ZN(U3511) );
  INV_X1 U4881 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4313) );
  MUX2_X1 U4882 ( .A(n4313), .B(n4312), .S(n4511), .Z(n4314) );
  OAI21_X1 U4883 ( .B1(n4315), .B2(n4329), .A(n4314), .ZN(U3510) );
  INV_X1 U4884 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4317) );
  MUX2_X1 U4885 ( .A(n4317), .B(n4316), .S(n4511), .Z(n4318) );
  OAI21_X1 U4886 ( .B1(n4319), .B2(n4329), .A(n4318), .ZN(U3509) );
  MUX2_X1 U4887 ( .A(REG0_REG_22__SCAN_IN), .B(n4320), .S(n4511), .Z(U3508) );
  MUX2_X1 U4888 ( .A(REG0_REG_21__SCAN_IN), .B(n4321), .S(n4511), .Z(U3507) );
  INV_X1 U4889 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4323) );
  MUX2_X1 U4890 ( .A(n4323), .B(n4322), .S(n4511), .Z(n4324) );
  OAI21_X1 U4891 ( .B1(n4325), .B2(n4329), .A(n4324), .ZN(U3506) );
  INV_X1 U4892 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4327) );
  MUX2_X1 U4893 ( .A(n4327), .B(n4326), .S(n4511), .Z(n4328) );
  OAI21_X1 U4894 ( .B1(n4330), .B2(n4329), .A(n4328), .ZN(U3505) );
  MUX2_X1 U4895 ( .A(REG0_REG_18__SCAN_IN), .B(n4331), .S(n4511), .Z(U3503) );
  MUX2_X1 U4896 ( .A(REG0_REG_16__SCAN_IN), .B(n4332), .S(n4511), .Z(U3499) );
  MUX2_X1 U4897 ( .A(REG0_REG_15__SCAN_IN), .B(n4333), .S(n4511), .Z(U3497) );
  MUX2_X1 U4898 ( .A(n2392), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4899 ( .A(n4334), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  INV_X1 U4900 ( .A(n4335), .ZN(n4336) );
  MUX2_X1 U4901 ( .A(DATAI_7_), .B(n4336), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4902 ( .A(n4337), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4903 ( .A(DATAI_4_), .B(n4338), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4904 ( .A(n4339), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  INV_X1 U4905 ( .A(DATAI_28_), .ZN(n4340) );
  AOI22_X1 U4906 ( .A1(STATE_REG_SCAN_IN), .A2(n4341), .B1(n4340), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U4907 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U4908 ( .A1(n4343), .A2(n4439), .B1(n2999), .B2(n4342), .ZN(n4344)
         );
  OAI21_X1 U4909 ( .B1(n2999), .B2(n4637), .A(n4344), .ZN(U3260) );
  INV_X1 U4910 ( .A(n4345), .ZN(n4346) );
  AOI22_X1 U4911 ( .A1(n4346), .A2(n4439), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4182), .ZN(n4347) );
  OAI21_X1 U4912 ( .B1(n4182), .B2(n4348), .A(n4347), .ZN(U3261) );
  AOI211_X1 U4913 ( .C1(n2179), .C2(n4350), .A(n4349), .B(n4400), .ZN(n4352)
         );
  AOI211_X1 U4914 ( .C1(n4424), .C2(ADDR_REG_9__SCAN_IN), .A(n4352), .B(n4351), 
        .ZN(n4357) );
  OAI211_X1 U4915 ( .C1(n4355), .C2(n4354), .A(n4432), .B(n4353), .ZN(n4356)
         );
  OAI211_X1 U4916 ( .C1(n4437), .C2(n4469), .A(n4357), .B(n4356), .ZN(U3249)
         );
  AOI211_X1 U4917 ( .C1(n4360), .C2(n4359), .A(n4358), .B(n4400), .ZN(n4362)
         );
  AOI211_X1 U4918 ( .C1(n4424), .C2(ADDR_REG_10__SCAN_IN), .A(n4362), .B(n4361), .ZN(n4366) );
  OAI211_X1 U4919 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4364), .A(n4432), .B(n4363), .ZN(n4365) );
  OAI211_X1 U4920 ( .C1(n4437), .C2(n4467), .A(n4366), .B(n4365), .ZN(U3250)
         );
  AOI211_X1 U4921 ( .C1(n4369), .C2(n4368), .A(n4367), .B(n4400), .ZN(n4371)
         );
  AOI211_X1 U4922 ( .C1(n4424), .C2(ADDR_REG_11__SCAN_IN), .A(n4371), .B(n4370), .ZN(n4376) );
  OAI211_X1 U4923 ( .C1(n4374), .C2(n4373), .A(n4432), .B(n4372), .ZN(n4375)
         );
  OAI211_X1 U4924 ( .C1(n4437), .C2(n4377), .A(n4376), .B(n4375), .ZN(U3251)
         );
  AOI211_X1 U4925 ( .C1(n4380), .C2(n4379), .A(n4378), .B(n4400), .ZN(n4382)
         );
  AOI211_X1 U4926 ( .C1(n4424), .C2(ADDR_REG_12__SCAN_IN), .A(n4382), .B(n4381), .ZN(n4386) );
  OAI211_X1 U4927 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4384), .A(n4432), .B(n4383), .ZN(n4385) );
  OAI211_X1 U4928 ( .C1(n4437), .C2(n2343), .A(n4386), .B(n4385), .ZN(U3252)
         );
  NAND2_X1 U4929 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4424), .ZN(n4399) );
  AOI211_X1 U4930 ( .C1(n4392), .C2(n4391), .A(n4390), .B(n4389), .ZN(n4393)
         );
  AOI211_X1 U4931 ( .C1(n4396), .C2(n4395), .A(n4394), .B(n4393), .ZN(n4398)
         );
  NAND3_X1 U4932 ( .A1(n4399), .A2(n4398), .A3(n4397), .ZN(U3254) );
  AOI211_X1 U4933 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4404)
         );
  AOI211_X1 U4934 ( .C1(n4424), .C2(ADDR_REG_15__SCAN_IN), .A(n4405), .B(n4404), .ZN(n4411) );
  AOI21_X1 U4935 ( .B1(n4408), .B2(n4407), .A(n4406), .ZN(n4409) );
  NAND2_X1 U4936 ( .A1(n4432), .A2(n4409), .ZN(n4410) );
  OAI211_X1 U4937 ( .C1(n4437), .C2(n4461), .A(n4411), .B(n4410), .ZN(U3255)
         );
  AOI21_X1 U4938 ( .B1(n4424), .B2(ADDR_REG_16__SCAN_IN), .A(n4412), .ZN(n4422) );
  OAI21_X1 U4939 ( .B1(n4415), .B2(n4414), .A(n4413), .ZN(n4420) );
  OAI21_X1 U4940 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n4419) );
  AOI22_X1 U4941 ( .A1(n4434), .A2(n4420), .B1(n4432), .B2(n4419), .ZN(n4421)
         );
  OAI211_X1 U4942 ( .C1(n4459), .C2(n4437), .A(n4422), .B(n4421), .ZN(U3256)
         );
  AOI21_X1 U4943 ( .B1(n4424), .B2(ADDR_REG_17__SCAN_IN), .A(n4423), .ZN(n4436) );
  OAI21_X1 U4944 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n4433) );
  OAI21_X1 U4945 ( .B1(n4430), .B2(n4429), .A(n4428), .ZN(n4431) );
  AOI22_X1 U4946 ( .A1(n4434), .A2(n4433), .B1(n4432), .B2(n4431), .ZN(n4435)
         );
  OAI211_X1 U4947 ( .C1(n4458), .C2(n4437), .A(n4436), .B(n4435), .ZN(U3257)
         );
  AOI22_X1 U4948 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4182), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4448), .ZN(n4442) );
  AOI22_X1 U4949 ( .A1(n4440), .A2(n4449), .B1(n4439), .B2(n4438), .ZN(n4441)
         );
  OAI211_X1 U4950 ( .C1(n4182), .C2(n4443), .A(n4442), .B(n4441), .ZN(U3288)
         );
  NAND2_X1 U4951 ( .A1(n2722), .A2(n4444), .ZN(n4446) );
  AOI21_X1 U4952 ( .B1(n4447), .B2(n4446), .A(n4445), .ZN(n4453) );
  AOI22_X1 U4953 ( .A1(n4450), .A2(n4449), .B1(REG3_REG_0__SCAN_IN), .B2(n4448), .ZN(n4451) );
  OAI221_X1 U4954 ( .B1(n4182), .B2(n4453), .C1(n2999), .C2(n4452), .A(n4451), 
        .ZN(U3290) );
  AND2_X1 U4955 ( .A1(D_REG_31__SCAN_IN), .A2(n4634), .ZN(U3291) );
  AND2_X1 U4956 ( .A1(D_REG_30__SCAN_IN), .A2(n4634), .ZN(U3292) );
  AND2_X1 U4957 ( .A1(D_REG_29__SCAN_IN), .A2(n4634), .ZN(U3293) );
  AND2_X1 U4958 ( .A1(D_REG_28__SCAN_IN), .A2(n4634), .ZN(U3294) );
  AND2_X1 U4959 ( .A1(D_REG_27__SCAN_IN), .A2(n4634), .ZN(U3295) );
  AND2_X1 U4960 ( .A1(D_REG_26__SCAN_IN), .A2(n4634), .ZN(U3296) );
  INV_X1 U4961 ( .A(n4634), .ZN(n4454) );
  INV_X1 U4962 ( .A(D_REG_25__SCAN_IN), .ZN(n4549) );
  NOR2_X1 U4963 ( .A1(n4454), .A2(n4549), .ZN(U3297) );
  AND2_X1 U4964 ( .A1(D_REG_24__SCAN_IN), .A2(n4634), .ZN(U3298) );
  AND2_X1 U4965 ( .A1(D_REG_23__SCAN_IN), .A2(n4634), .ZN(U3299) );
  AND2_X1 U4966 ( .A1(D_REG_22__SCAN_IN), .A2(n4634), .ZN(U3300) );
  AND2_X1 U4967 ( .A1(D_REG_21__SCAN_IN), .A2(n4634), .ZN(U3301) );
  INV_X1 U4968 ( .A(D_REG_20__SCAN_IN), .ZN(n4548) );
  NOR2_X1 U4969 ( .A1(n4454), .A2(n4548), .ZN(U3302) );
  AND2_X1 U4970 ( .A1(D_REG_19__SCAN_IN), .A2(n4634), .ZN(U3303) );
  AND2_X1 U4971 ( .A1(D_REG_18__SCAN_IN), .A2(n4634), .ZN(U3304) );
  AND2_X1 U4972 ( .A1(D_REG_17__SCAN_IN), .A2(n4634), .ZN(U3305) );
  AND2_X1 U4973 ( .A1(D_REG_16__SCAN_IN), .A2(n4634), .ZN(U3306) );
  AND2_X1 U4974 ( .A1(D_REG_15__SCAN_IN), .A2(n4634), .ZN(U3307) );
  AND2_X1 U4975 ( .A1(D_REG_13__SCAN_IN), .A2(n4634), .ZN(U3309) );
  AND2_X1 U4976 ( .A1(D_REG_12__SCAN_IN), .A2(n4634), .ZN(U3310) );
  AND2_X1 U4977 ( .A1(D_REG_11__SCAN_IN), .A2(n4634), .ZN(U3311) );
  AND2_X1 U4978 ( .A1(D_REG_10__SCAN_IN), .A2(n4634), .ZN(U3312) );
  AND2_X1 U4979 ( .A1(D_REG_9__SCAN_IN), .A2(n4634), .ZN(U3313) );
  INV_X1 U4980 ( .A(D_REG_8__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U4981 ( .A1(n4454), .A2(n4551), .ZN(U3314) );
  AND2_X1 U4982 ( .A1(D_REG_7__SCAN_IN), .A2(n4634), .ZN(U3315) );
  AND2_X1 U4983 ( .A1(D_REG_6__SCAN_IN), .A2(n4634), .ZN(U3316) );
  AND2_X1 U4984 ( .A1(D_REG_5__SCAN_IN), .A2(n4634), .ZN(U3317) );
  AND2_X1 U4985 ( .A1(D_REG_4__SCAN_IN), .A2(n4634), .ZN(U3318) );
  INV_X1 U4986 ( .A(D_REG_3__SCAN_IN), .ZN(n4662) );
  NOR2_X1 U4987 ( .A1(n4454), .A2(n4662), .ZN(U3319) );
  AND2_X1 U4988 ( .A1(D_REG_2__SCAN_IN), .A2(n4634), .ZN(U3320) );
  INV_X1 U4989 ( .A(DATAI_23_), .ZN(n4456) );
  AOI21_X1 U4990 ( .B1(U3149), .B2(n4456), .A(n4455), .ZN(U3329) );
  INV_X1 U4991 ( .A(DATAI_18_), .ZN(n4523) );
  AOI22_X1 U4992 ( .A1(STATE_REG_SCAN_IN), .A2(n4457), .B1(n4523), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U4993 ( .A1(STATE_REG_SCAN_IN), .A2(n4458), .B1(n2555), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4994 ( .A(DATAI_16_), .ZN(n4656) );
  AOI22_X1 U4995 ( .A1(STATE_REG_SCAN_IN), .A2(n4459), .B1(n4656), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U4996 ( .A1(STATE_REG_SCAN_IN), .A2(n4461), .B1(n4460), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U4997 ( .A1(STATE_REG_SCAN_IN), .A2(n4462), .B1(n2527), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U4998 ( .A(DATAI_12_), .ZN(n4463) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n2343), .B1(n4463), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5000 ( .A1(U3149), .A2(n4464), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4465) );
  INV_X1 U5001 ( .A(n4465), .ZN(U3341) );
  INV_X1 U5002 ( .A(DATAI_10_), .ZN(n4466) );
  AOI22_X1 U5003 ( .A1(STATE_REG_SCAN_IN), .A2(n4467), .B1(n4466), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5004 ( .A(DATAI_9_), .ZN(n4468) );
  AOI22_X1 U5005 ( .A1(STATE_REG_SCAN_IN), .A2(n4469), .B1(n4468), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5006 ( .A1(STATE_REG_SCAN_IN), .A2(n2045), .B1(n2406), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5007 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5008 ( .A1(n4511), .A2(n4470), .B1(n4554), .B2(n4509), .ZN(U3467)
         );
  INV_X1 U5009 ( .A(n4471), .ZN(n4475) );
  OAI22_X1 U5010 ( .A1(n4473), .A2(n4479), .B1(n4478), .B2(n4472), .ZN(n4474)
         );
  NOR2_X1 U5011 ( .A1(n4475), .A2(n4474), .ZN(n4513) );
  INV_X1 U5012 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5013 ( .A1(n4511), .A2(n4513), .B1(n4476), .B2(n4509), .ZN(U3469)
         );
  OAI22_X1 U5014 ( .A1(n4480), .A2(n4479), .B1(n4478), .B2(n4477), .ZN(n4481)
         );
  NOR2_X1 U5015 ( .A1(n4482), .A2(n4481), .ZN(n4514) );
  INV_X1 U5016 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4553) );
  AOI22_X1 U5017 ( .A1(n4511), .A2(n4514), .B1(n4553), .B2(n4509), .ZN(U3473)
         );
  INV_X1 U5018 ( .A(n4483), .ZN(n4488) );
  INV_X1 U5019 ( .A(n4484), .ZN(n4486) );
  AOI211_X1 U5020 ( .C1(n4488), .C2(n4487), .A(n4486), .B(n4485), .ZN(n4515)
         );
  INV_X1 U5021 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U5022 ( .A1(n4511), .A2(n4515), .B1(n4489), .B2(n4509), .ZN(U3475)
         );
  NOR2_X1 U5023 ( .A1(n4491), .A2(n4490), .ZN(n4494) );
  INV_X1 U5024 ( .A(n4492), .ZN(n4493) );
  AOI211_X1 U5025 ( .C1(n4504), .C2(n4495), .A(n4494), .B(n4493), .ZN(n4516)
         );
  INV_X1 U5026 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5027 ( .A1(n4511), .A2(n4516), .B1(n4663), .B2(n4509), .ZN(U3477)
         );
  NAND3_X1 U5028 ( .A1(n2983), .A2(n4496), .A3(n4502), .ZN(n4498) );
  AND2_X1 U5029 ( .A1(n4498), .A2(n4497), .ZN(n4499) );
  AND2_X1 U5030 ( .A1(n4500), .A2(n4499), .ZN(n4517) );
  INV_X1 U5031 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5032 ( .A1(n4511), .A2(n4517), .B1(n4501), .B2(n4509), .ZN(U3481)
         );
  NAND2_X1 U5033 ( .A1(n4503), .A2(n4502), .ZN(n4508) );
  NAND2_X1 U5034 ( .A1(n4505), .A2(n4504), .ZN(n4506) );
  AND3_X1 U5035 ( .A1(n4508), .A2(n4507), .A3(n4506), .ZN(n4520) );
  INV_X1 U5036 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5037 ( .A1(n4511), .A2(n4520), .B1(n4510), .B2(n4509), .ZN(U3485)
         );
  AOI22_X1 U5038 ( .A1(n4518), .A2(n4513), .B1(n4512), .B2(n4519), .ZN(U3519)
         );
  AOI22_X1 U5039 ( .A1(n4518), .A2(n4514), .B1(n2421), .B2(n4519), .ZN(U3521)
         );
  AOI22_X1 U5040 ( .A1(n4521), .A2(n4515), .B1(n2428), .B2(n4519), .ZN(U3522)
         );
  AOI22_X1 U5041 ( .A1(n4521), .A2(n4516), .B1(n2436), .B2(n4519), .ZN(U3523)
         );
  AOI22_X1 U5042 ( .A1(n4518), .A2(n4517), .B1(n2457), .B2(n4519), .ZN(U3525)
         );
  AOI22_X1 U5043 ( .A1(n4521), .A2(n4520), .B1(n4644), .B2(n4519), .ZN(U3527)
         );
  INV_X1 U5044 ( .A(DATAI_21_), .ZN(n4524) );
  AOI22_X1 U5045 ( .A1(n4524), .A2(keyinput53), .B1(keyinput30), .B2(n4523), 
        .ZN(n4522) );
  OAI221_X1 U5046 ( .B1(n4524), .B2(keyinput53), .C1(n4523), .C2(keyinput30), 
        .A(n4522), .ZN(n4534) );
  AOI22_X1 U5047 ( .A1(n4526), .A2(keyinput26), .B1(n4656), .B2(keyinput5), 
        .ZN(n4525) );
  OAI221_X1 U5048 ( .B1(n4526), .B2(keyinput26), .C1(n4656), .C2(keyinput5), 
        .A(n4525), .ZN(n4533) );
  INV_X1 U5049 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5050 ( .A1(n4657), .A2(keyinput4), .B1(n4528), .B2(keyinput24), 
        .ZN(n4527) );
  OAI221_X1 U5051 ( .B1(n4657), .B2(keyinput4), .C1(n4528), .C2(keyinput24), 
        .A(n4527), .ZN(n4532) );
  XOR2_X1 U5052 ( .A(n2406), .B(keyinput55), .Z(n4530) );
  XNOR2_X1 U5053 ( .A(DATAI_3_), .B(keyinput6), .ZN(n4529) );
  NAND2_X1 U5054 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  NOR4_X1 U5055 ( .A1(n4534), .A2(n4533), .A3(n4532), .A4(n4531), .ZN(n4574)
         );
  XOR2_X1 U5056 ( .A(n2647), .B(keyinput42), .Z(n4540) );
  XOR2_X1 U5057 ( .A(n4535), .B(keyinput22), .Z(n4539) );
  INV_X1 U5058 ( .A(IR_REG_12__SCAN_IN), .ZN(n4536) );
  XOR2_X1 U5059 ( .A(n4536), .B(keyinput34), .Z(n4538) );
  XNOR2_X1 U5060 ( .A(IR_REG_24__SCAN_IN), .B(keyinput41), .ZN(n4537) );
  NAND4_X1 U5061 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4546)
         );
  XNOR2_X1 U5062 ( .A(IR_REG_6__SCAN_IN), .B(keyinput2), .ZN(n4544) );
  XNOR2_X1 U5063 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput63), .ZN(n4543) );
  XNOR2_X1 U5064 ( .A(IR_REG_18__SCAN_IN), .B(keyinput50), .ZN(n4542) );
  XNOR2_X1 U5065 ( .A(IR_REG_10__SCAN_IN), .B(keyinput9), .ZN(n4541) );
  NAND4_X1 U5066 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4545)
         );
  NOR2_X1 U5067 ( .A1(n4546), .A2(n4545), .ZN(n4573) );
  AOI22_X1 U5068 ( .A1(n4549), .A2(keyinput43), .B1(keyinput61), .B2(n4548), 
        .ZN(n4547) );
  OAI221_X1 U5069 ( .B1(n4549), .B2(keyinput43), .C1(n4548), .C2(keyinput61), 
        .A(n4547), .ZN(n4560) );
  AOI22_X1 U5070 ( .A1(n4551), .A2(keyinput7), .B1(keyinput1), .B2(n4662), 
        .ZN(n4550) );
  OAI221_X1 U5071 ( .B1(n4551), .B2(keyinput7), .C1(n4662), .C2(keyinput1), 
        .A(n4550), .ZN(n4559) );
  AOI22_X1 U5072 ( .A1(n4554), .A2(keyinput49), .B1(n4553), .B2(keyinput11), 
        .ZN(n4552) );
  OAI221_X1 U5073 ( .B1(n4554), .B2(keyinput49), .C1(n4553), .C2(keyinput11), 
        .A(n4552), .ZN(n4558) );
  XNOR2_X1 U5074 ( .A(D_REG_0__SCAN_IN), .B(keyinput38), .ZN(n4556) );
  XNOR2_X1 U5075 ( .A(IR_REG_31__SCAN_IN), .B(keyinput62), .ZN(n4555) );
  NAND2_X1 U5076 ( .A1(n4556), .A2(n4555), .ZN(n4557) );
  NOR4_X1 U5077 ( .A1(n4560), .A2(n4559), .A3(n4558), .A4(n4557), .ZN(n4572)
         );
  AOI22_X1 U5078 ( .A1(n4663), .A2(keyinput16), .B1(n4665), .B2(keyinput17), 
        .ZN(n4561) );
  OAI221_X1 U5079 ( .B1(n4663), .B2(keyinput16), .C1(n4665), .C2(keyinput17), 
        .A(n4561), .ZN(n4570) );
  INV_X1 U5080 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5081 ( .A1(n4563), .A2(keyinput0), .B1(n4664), .B2(keyinput56), 
        .ZN(n4562) );
  OAI221_X1 U5082 ( .B1(n4563), .B2(keyinput0), .C1(n4664), .C2(keyinput56), 
        .A(n4562), .ZN(n4569) );
  AOI22_X1 U5083 ( .A1(n2428), .A2(keyinput57), .B1(n4565), .B2(keyinput13), 
        .ZN(n4564) );
  OAI221_X1 U5084 ( .B1(n2428), .B2(keyinput57), .C1(n4565), .C2(keyinput13), 
        .A(n4564), .ZN(n4568) );
  AOI22_X1 U5085 ( .A1(n2448), .A2(keyinput40), .B1(n2457), .B2(keyinput15), 
        .ZN(n4566) );
  OAI221_X1 U5086 ( .B1(n2448), .B2(keyinput40), .C1(n2457), .C2(keyinput15), 
        .A(n4566), .ZN(n4567) );
  NOR4_X1 U5087 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(n4571)
         );
  NAND4_X1 U5088 ( .A1(n4574), .A2(n4573), .A3(n4572), .A4(n4571), .ZN(n4633)
         );
  AOI22_X1 U5089 ( .A1(n4576), .A2(keyinput23), .B1(keyinput60), .B2(n4644), 
        .ZN(n4575) );
  OAI221_X1 U5090 ( .B1(n4576), .B2(keyinput23), .C1(n4644), .C2(keyinput60), 
        .A(n4575), .ZN(n4587) );
  AOI22_X1 U5091 ( .A1(n4645), .A2(keyinput33), .B1(n4578), .B2(keyinput29), 
        .ZN(n4577) );
  OAI221_X1 U5092 ( .B1(n4645), .B2(keyinput33), .C1(n4578), .C2(keyinput29), 
        .A(n4577), .ZN(n4586) );
  AOI22_X1 U5093 ( .A1(n4581), .A2(keyinput51), .B1(n4580), .B2(keyinput28), 
        .ZN(n4579) );
  OAI221_X1 U5094 ( .B1(n4581), .B2(keyinput51), .C1(n4580), .C2(keyinput28), 
        .A(n4579), .ZN(n4585) );
  XNOR2_X1 U5095 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput35), .ZN(n4583) );
  XNOR2_X1 U5096 ( .A(keyinput32), .B(REG1_REG_30__SCAN_IN), .ZN(n4582) );
  NAND2_X1 U5097 ( .A1(n4583), .A2(n4582), .ZN(n4584) );
  NOR4_X1 U5098 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4631)
         );
  INV_X1 U5099 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4638) );
  INV_X1 U5100 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5101 ( .A1(n4638), .A2(keyinput58), .B1(n4589), .B2(keyinput37), 
        .ZN(n4588) );
  OAI221_X1 U5102 ( .B1(n4638), .B2(keyinput58), .C1(n4589), .C2(keyinput37), 
        .A(n4588), .ZN(n4599) );
  INV_X1 U5103 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5104 ( .A1(n4591), .A2(keyinput20), .B1(n3163), .B2(keyinput44), 
        .ZN(n4590) );
  OAI221_X1 U5105 ( .B1(n4591), .B2(keyinput20), .C1(n3163), .C2(keyinput44), 
        .A(n4590), .ZN(n4598) );
  AOI22_X1 U5106 ( .A1(n4637), .A2(keyinput46), .B1(n4144), .B2(keyinput47), 
        .ZN(n4592) );
  OAI221_X1 U5107 ( .B1(n4637), .B2(keyinput46), .C1(n4144), .C2(keyinput47), 
        .A(n4592), .ZN(n4597) );
  INV_X1 U5108 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4595) );
  INV_X1 U5109 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4594) );
  AOI22_X1 U5110 ( .A1(n4595), .A2(keyinput18), .B1(n4594), .B2(keyinput31), 
        .ZN(n4593) );
  OAI221_X1 U5111 ( .B1(n4595), .B2(keyinput18), .C1(n4594), .C2(keyinput31), 
        .A(n4593), .ZN(n4596) );
  NOR4_X1 U5112 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4630)
         );
  INV_X1 U5113 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4602) );
  INV_X1 U5114 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5115 ( .A1(n4602), .A2(keyinput10), .B1(n4601), .B2(keyinput59), 
        .ZN(n4600) );
  OAI221_X1 U5116 ( .B1(n4602), .B2(keyinput10), .C1(n4601), .C2(keyinput59), 
        .A(n4600), .ZN(n4611) );
  AOI22_X1 U5117 ( .A1(n4652), .A2(keyinput19), .B1(keyinput14), .B2(n4604), 
        .ZN(n4603) );
  OAI221_X1 U5118 ( .B1(n4652), .B2(keyinput19), .C1(n4604), .C2(keyinput14), 
        .A(n4603), .ZN(n4610) );
  AOI22_X1 U5119 ( .A1(n4654), .A2(keyinput21), .B1(n4655), .B2(keyinput3), 
        .ZN(n4605) );
  OAI221_X1 U5120 ( .B1(n4654), .B2(keyinput21), .C1(n4655), .C2(keyinput3), 
        .A(n4605), .ZN(n4609) );
  AOI22_X1 U5121 ( .A1(n4653), .A2(keyinput54), .B1(n4607), .B2(keyinput52), 
        .ZN(n4606) );
  OAI221_X1 U5122 ( .B1(n4653), .B2(keyinput54), .C1(n4607), .C2(keyinput52), 
        .A(n4606), .ZN(n4608) );
  NOR4_X1 U5123 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4629)
         );
  AOI22_X1 U5124 ( .A1(n4614), .A2(keyinput48), .B1(keyinput45), .B2(n4613), 
        .ZN(n4612) );
  OAI221_X1 U5125 ( .B1(n4614), .B2(keyinput48), .C1(n4613), .C2(keyinput45), 
        .A(n4612), .ZN(n4627) );
  AOI22_X1 U5126 ( .A1(n4617), .A2(keyinput36), .B1(keyinput8), .B2(n4616), 
        .ZN(n4615) );
  OAI221_X1 U5127 ( .B1(n4617), .B2(keyinput36), .C1(n4616), .C2(keyinput8), 
        .A(n4615), .ZN(n4626) );
  INV_X1 U5128 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5129 ( .A1(n4620), .A2(keyinput12), .B1(n4619), .B2(keyinput39), 
        .ZN(n4618) );
  OAI221_X1 U5130 ( .B1(n4620), .B2(keyinput12), .C1(n4619), .C2(keyinput39), 
        .A(n4618), .ZN(n4625) );
  INV_X1 U5131 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U5132 ( .A1(n4623), .A2(keyinput25), .B1(keyinput27), .B2(n4622), 
        .ZN(n4621) );
  OAI221_X1 U5133 ( .B1(n4623), .B2(keyinput25), .C1(n4622), .C2(keyinput27), 
        .A(n4621), .ZN(n4624) );
  NOR4_X1 U5134 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4628)
         );
  NAND4_X1 U5135 ( .A1(n4631), .A2(n4630), .A3(n4629), .A4(n4628), .ZN(n4632)
         );
  NOR2_X1 U5136 ( .A1(n4633), .A2(n4632), .ZN(n4636) );
  NAND2_X1 U5137 ( .A1(D_REG_14__SCAN_IN), .A2(n4634), .ZN(n4635) );
  XNOR2_X1 U5138 ( .A(n4636), .B(n4635), .ZN(n4677) );
  NOR3_X1 U5139 ( .A1(ADDR_REG_17__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        n4637), .ZN(n4675) );
  NAND4_X1 U5140 ( .A1(REG2_REG_8__SCAN_IN), .A2(REG2_REG_18__SCAN_IN), .A3(
        n3163), .A4(n4638), .ZN(n4643) );
  NAND3_X1 U5141 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .A3(
        IR_REG_31__SCAN_IN), .ZN(n4639) );
  OR4_X1 U5142 ( .A1(n4535), .A2(n4640), .A3(IR_REG_6__SCAN_IN), .A4(n4639), 
        .ZN(n4642) );
  INV_X1 U5143 ( .A(IR_REG_18__SCAN_IN), .ZN(n4641) );
  NOR4_X1 U5144 ( .A1(n4643), .A2(IR_REG_20__SCAN_IN), .A3(n4642), .A4(n4641), 
        .ZN(n4674) );
  NOR4_X1 U5145 ( .A1(REG1_REG_20__SCAN_IN), .A2(REG1_REG_11__SCAN_IN), .A3(
        n4645), .A4(n4644), .ZN(n4651) );
  NOR4_X1 U5146 ( .A1(REG3_REG_15__SCAN_IN), .A2(DATAO_REG_13__SCAN_IN), .A3(
        DATAO_REG_14__SCAN_IN), .A4(DATAO_REG_25__SCAN_IN), .ZN(n4650) );
  NOR4_X1 U5147 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .A3(
        REG2_REG_26__SCAN_IN), .A4(ADDR_REG_19__SCAN_IN), .ZN(n4646) );
  NAND3_X1 U5148 ( .A1(REG1_REG_26__SCAN_IN), .A2(n4646), .A3(
        REG1_REG_30__SCAN_IN), .ZN(n4648) );
  INV_X1 U5149 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4647) );
  NOR3_X1 U5150 ( .A1(n4648), .A2(n4647), .A3(REG1_REG_21__SCAN_IN), .ZN(n4649) );
  NAND3_X1 U5151 ( .A1(n4651), .A2(n4650), .A3(n4649), .ZN(n4672) );
  NOR4_X1 U5152 ( .A1(DATAO_REG_2__SCAN_IN), .A2(ADDR_REG_9__SCAN_IN), .A3(
        ADDR_REG_5__SCAN_IN), .A4(n4652), .ZN(n4661) );
  NOR4_X1 U5153 ( .A1(DATAO_REG_12__SCAN_IN), .A2(n4655), .A3(n4654), .A4(
        n4653), .ZN(n4660) );
  NOR4_X1 U5154 ( .A1(REG3_REG_17__SCAN_IN), .A2(DATAI_21_), .A3(DATAI_7_), 
        .A4(n4656), .ZN(n4659) );
  NOR4_X1 U5155 ( .A1(REG3_REG_21__SCAN_IN), .A2(DATAI_0_), .A3(DATAI_18_), 
        .A4(n4657), .ZN(n4658) );
  NAND4_X1 U5156 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4671)
         );
  NAND4_X1 U5157 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_0__SCAN_IN), .A3(
        REG0_REG_17__SCAN_IN), .A4(n4662), .ZN(n4670) );
  NOR4_X1 U5158 ( .A1(REG0_REG_10__SCAN_IN), .A2(DATAI_3_), .A3(n4664), .A4(
        n4663), .ZN(n4668) );
  NOR4_X1 U5159 ( .A1(REG1_REG_6__SCAN_IN), .A2(REG1_REG_7__SCAN_IN), .A3(
        n4665), .A4(n2428), .ZN(n4667) );
  NOR3_X1 U5160 ( .A1(D_REG_25__SCAN_IN), .A2(REG0_REG_3__SCAN_IN), .A3(
        REG0_REG_0__SCAN_IN), .ZN(n4666) );
  NAND4_X1 U5161 ( .A1(D_REG_20__SCAN_IN), .A2(n4668), .A3(n4667), .A4(n4666), 
        .ZN(n4669) );
  NOR4_X1 U5162 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4673)
         );
  NAND4_X1 U5163 ( .A1(REG2_REG_23__SCAN_IN), .A2(n4675), .A3(n4674), .A4(
        n4673), .ZN(n4676) );
  XNOR2_X1 U5164 ( .A(n4677), .B(n4676), .ZN(U3308) );
endmodule

