

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7418, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738;

  MUX2_X1 U7518 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n15561), .S(n16526), .Z(
        P2_U3528) );
  NAND2_X1 U7519 ( .A1(n14024), .A2(n14023), .ZN(n16025) );
  NOR2_X1 U7520 ( .A1(n8534), .A2(n13459), .ZN(n8533) );
  CLKBUF_X1 U7521 ( .A(n10837), .Z(n10915) );
  AND2_X1 U7522 ( .A1(n10024), .A2(n10023), .ZN(n12615) );
  INV_X2 U7523 ( .A(n10499), .ZN(n7420) );
  AND2_X4 U7524 ( .A1(n8994), .A2(n11277), .ZN(n8963) );
  INV_X2 U7525 ( .A(n13771), .ZN(n7421) );
  NAND2_X1 U7526 ( .A1(n11721), .A2(n10576), .ZN(n8284) );
  NAND2_X2 U7527 ( .A1(n14510), .A2(n10837), .ZN(n8994) );
  INV_X1 U7528 ( .A(n10208), .ZN(n10511) );
  NAND2_X1 U7529 ( .A1(n9797), .A2(n15612), .ZN(n9887) );
  NAND2_X1 U7530 ( .A1(n13712), .A2(n11277), .ZN(n11123) );
  AND2_X1 U7531 ( .A1(n10615), .A2(n10614), .ZN(n8033) );
  NAND2_X2 U7532 ( .A1(n8051), .A2(n8050), .ZN(n13599) );
  XNOR2_X2 U7533 ( .A(n8098), .B(n10664), .ZN(n10784) );
  NAND2_X2 U7534 ( .A1(n8911), .A2(n8910), .ZN(n9895) );
  OAI211_X1 U7535 ( .C1(n9078), .C2(n11271), .A(n8936), .B(n8935), .ZN(n12709)
         );
  INV_X1 U7536 ( .A(n8964), .ZN(n8616) );
  AND2_X1 U7537 ( .A1(n7673), .A2(n7672), .ZN(n14994) );
  NOR2_X1 U7538 ( .A1(n14994), .A2(n7468), .ZN(n14095) );
  INV_X1 U7539 ( .A(n9887), .ZN(n10514) );
  AOI21_X1 U7540 ( .B1(n15478), .B2(n15193), .A(n15259), .ZN(n15242) );
  INV_X1 U7541 ( .A(n9870), .ZN(n9909) );
  OAI21_X1 U7542 ( .B1(n10149), .B2(n9805), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9812) );
  INV_X1 U7543 ( .A(n11679), .ZN(n7695) );
  CLKBUF_X2 U7544 ( .A(n7460), .Z(n7418) );
  INV_X1 U7545 ( .A(n12917), .ZN(n12853) );
  AND2_X1 U7546 ( .A1(n10260), .A2(n10259), .ZN(n15595) );
  INV_X1 U7547 ( .A(n10569), .ZN(n13117) );
  INV_X2 U7548 ( .A(n10540), .ZN(n10220) );
  OAI22_X2 U7549 ( .A1(n13679), .A2(n8757), .B1(n13680), .B2(n8758), .ZN(
        n13683) );
  OAI21_X2 U7550 ( .B1(n9282), .B2(n8340), .A(n8337), .ZN(n14660) );
  NAND2_X2 U7551 ( .A1(n14701), .A2(n14705), .ZN(n9282) );
  XNOR2_X1 U7552 ( .A(n13582), .B(n15756), .ZN(n13855) );
  OR2_X1 U7553 ( .A1(n11250), .A2(n10569), .ZN(n7460) );
  AND2_X4 U7554 ( .A1(n14957), .A2(n14962), .ZN(n9277) );
  AOI21_X2 U7555 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n16366), .A(n16365), .ZN(
        n16374) );
  OAI21_X2 U7556 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n16404), .A(n16403), .ZN(
        n16412) );
  OR2_X4 U7557 ( .A1(n15604), .A2(n15605), .ZN(n9860) );
  NOR2_X2 U7558 ( .A1(n10516), .A2(n13431), .ZN(n11714) );
  NAND2_X1 U7559 ( .A1(n8386), .A2(n8385), .ZN(n15309) );
  NAND2_X1 U7560 ( .A1(n15199), .A2(n15198), .ZN(n15438) );
  AND2_X1 U7561 ( .A1(n10169), .A2(n10168), .ZN(n13348) );
  NAND4_X1 U7562 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        n15754) );
  INV_X2 U7563 ( .A(n13599), .ZN(n11762) );
  NAND4_X1 U7564 ( .A1(n8929), .A2(n8928), .A3(n8927), .A4(n8926), .ZN(n12279)
         );
  CLKBUF_X2 U7565 ( .A(n10677), .Z(n13810) );
  NOR2_X1 U7566 ( .A1(n8832), .A2(n8833), .ZN(n11226) );
  CLKBUF_X2 U7567 ( .A(n8937), .Z(n9326) );
  CLKBUF_X2 U7568 ( .A(n9890), .Z(n10463) );
  INV_X1 U7569 ( .A(n8862), .ZN(n14957) );
  AND2_X1 U7570 ( .A1(n10720), .A2(n10638), .ZN(n11106) );
  INV_X4 U7571 ( .A(n10674), .ZN(n11277) );
  NOR2_X1 U7572 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8628) );
  OAI21_X1 U7573 ( .B1(n13822), .B2(n13821), .A(n13820), .ZN(n13823) );
  NOR2_X1 U7574 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  AOI21_X1 U7575 ( .B1(n8124), .B2(n16529), .A(n7612), .ZN(n8315) );
  AND2_X1 U7576 ( .A1(n10409), .A2(n7434), .ZN(n7871) );
  NOR2_X1 U7577 ( .A1(n14832), .A2(n8106), .ZN(n14903) );
  NOR2_X1 U7578 ( .A1(n7426), .A2(n7618), .ZN(n7814) );
  OR2_X1 U7579 ( .A1(n15843), .A2(n7477), .ZN(n15831) );
  XNOR2_X1 U7580 ( .A(n14096), .B(n8204), .ZN(n14977) );
  NOR2_X1 U7581 ( .A1(n15869), .A2(n15873), .ZN(n15868) );
  NOR4_X1 U7582 ( .A1(n14496), .A2(n14495), .A3(n14494), .A4(n14634), .ZN(
        n14499) );
  NAND2_X1 U7583 ( .A1(n15051), .A2(n7595), .ZN(n15049) );
  NAND2_X1 U7584 ( .A1(n15309), .A2(n15217), .ZN(n15290) );
  XNOR2_X1 U7585 ( .A(n14095), .B(n14093), .ZN(n15051) );
  NAND2_X1 U7586 ( .A1(n15347), .A2(n8389), .ZN(n8386) );
  NAND2_X1 U7587 ( .A1(n15400), .A2(n15180), .ZN(n15383) );
  NAND2_X1 U7588 ( .A1(n14047), .A2(n14046), .ZN(n15971) );
  OAI21_X1 U7589 ( .B1(n14186), .B2(n14183), .A(n14182), .ZN(n13939) );
  OR2_X1 U7590 ( .A1(n14293), .A2(n14646), .ZN(n14326) );
  AND2_X1 U7591 ( .A1(n8305), .A2(n8304), .ZN(n8303) );
  NAND2_X1 U7592 ( .A1(n7647), .A2(n13350), .ZN(n15174) );
  NAND2_X1 U7593 ( .A1(n8403), .A2(n8404), .ZN(n15404) );
  AND2_X1 U7594 ( .A1(n15299), .A2(n15218), .ZN(n7646) );
  NAND2_X1 U7595 ( .A1(n10397), .A2(n10396), .ZN(n15299) );
  NAND2_X1 U7596 ( .A1(n16713), .A2(n16712), .ZN(n16711) );
  XNOR2_X1 U7597 ( .A(n8729), .B(n11122), .ZN(n16713) );
  NAND2_X1 U7598 ( .A1(n8083), .A2(n8730), .ZN(n8729) );
  NAND2_X1 U7599 ( .A1(n13231), .A2(n13230), .ZN(n13347) );
  NAND2_X1 U7600 ( .A1(n11180), .A2(n11179), .ZN(n16111) );
  NAND2_X1 U7601 ( .A1(n12881), .A2(n12880), .ZN(n16610) );
  OAI21_X1 U7602 ( .B1(n8053), .B2(n16570), .A(n8052), .ZN(n16612) );
  NAND2_X1 U7603 ( .A1(n12336), .A2(n10777), .ZN(n16575) );
  AOI21_X1 U7604 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n16397), .A(n16396), .ZN(
        n16402) );
  AND2_X1 U7605 ( .A1(n12495), .A2(n12615), .ZN(n12641) );
  NAND2_X1 U7606 ( .A1(n8841), .A2(n8840), .ZN(n9309) );
  NAND2_X1 U7607 ( .A1(n16493), .A2(n16494), .ZN(n16492) );
  INV_X2 U7608 ( .A(n14167), .ZN(n7422) );
  AND2_X1 U7609 ( .A1(n14379), .A2(n14378), .ZN(n14473) );
  INV_X2 U7610 ( .A(n13935), .ZN(n14163) );
  NAND2_X1 U7611 ( .A1(n10698), .A2(n10697), .ZN(n13607) );
  AND2_X1 U7612 ( .A1(n9913), .A2(n9912), .ZN(n12282) );
  NAND4_X1 U7613 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n15755) );
  INV_X2 U7614 ( .A(n13583), .ZN(n13836) );
  AND2_X1 U7615 ( .A1(n9934), .A2(n9933), .ZN(n12109) );
  INV_X2 U7616 ( .A(n9986), .ZN(n10540) );
  INV_X4 U7617 ( .A(n10875), .ZN(P3_U3897) );
  OAI211_X1 U7618 ( .C1(n11350), .C2(n10679), .A(n7528), .B(n10681), .ZN(
        n15756) );
  NAND2_X1 U7619 ( .A1(n11223), .A2(n13027), .ZN(n15443) );
  INV_X1 U7620 ( .A(n13579), .ZN(n13583) );
  AND3_X1 U7621 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(n14215) );
  NAND2_X1 U7622 ( .A1(n11714), .A2(n11248), .ZN(n9986) );
  INV_X2 U7623 ( .A(n11123), .ZN(n13838) );
  NAND4_X1 U7624 ( .A1(n8948), .A2(n8947), .A3(n8946), .A4(n8945), .ZN(n14366)
         );
  AND2_X2 U7625 ( .A1(n10637), .A2(n10814), .ZN(P1_U4016) );
  INV_X1 U7626 ( .A(n10679), .ZN(n13805) );
  NAND2_X1 U7627 ( .A1(n11199), .A2(n13850), .ZN(n16686) );
  NAND2_X2 U7628 ( .A1(n8862), .A2(n14962), .ZN(n12679) );
  NAND2_X2 U7629 ( .A1(n8994), .A2(n10674), .ZN(n9078) );
  AND2_X2 U7630 ( .A1(n13565), .A2(n10659), .ZN(n13829) );
  INV_X2 U7631 ( .A(n10650), .ZN(n16033) );
  OR2_X1 U7632 ( .A1(n13431), .A2(n11248), .ZN(n11250) );
  NAND2_X1 U7633 ( .A1(n10666), .A2(n10667), .ZN(n16170) );
  NAND2_X2 U7634 ( .A1(n15160), .A2(n10566), .ZN(n9870) );
  NAND2_X1 U7635 ( .A1(n10666), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8098) );
  XNOR2_X1 U7636 ( .A(n8749), .B(P1_IR_REG_22__SCAN_IN), .ZN(n16180) );
  XNOR2_X1 U7637 ( .A(n10643), .B(P1_IR_REG_21__SCAN_IN), .ZN(n13849) );
  OR2_X1 U7638 ( .A1(n10641), .A2(n10632), .ZN(n8088) );
  XNOR2_X1 U7639 ( .A(n7926), .B(P2_IR_REG_22__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U7640 ( .A1(n9829), .A2(n9830), .ZN(n15160) );
  XNOR2_X1 U7641 ( .A(n10630), .B(n10629), .ZN(n13516) );
  INV_X1 U7642 ( .A(n15612), .ZN(n9863) );
  NAND2_X1 U7643 ( .A1(n10548), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U7644 ( .A1(n8179), .A2(n10652), .ZN(n10666) );
  MUX2_X1 U7645 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10665), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n10667) );
  NAND2_X1 U7646 ( .A1(n9387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8232) );
  INV_X2 U7647 ( .A(n14952), .ZN(n14959) );
  XNOR2_X1 U7648 ( .A(n7885), .B(n7884), .ZN(n15612) );
  XNOR2_X1 U7649 ( .A(n10655), .B(n10654), .ZN(n13565) );
  MUX2_X1 U7650 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9828), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n9830) );
  INV_X1 U7651 ( .A(n10651), .ZN(n8179) );
  XNOR2_X1 U7652 ( .A(n9826), .B(n9825), .ZN(n10566) );
  NOR2_X1 U7653 ( .A1(n9165), .A2(n8857), .ZN(n8901) );
  NOR2_X1 U7654 ( .A1(n10149), .A2(n9809), .ZN(n9814) );
  AND3_X1 U7655 ( .A1(n7437), .A2(n7656), .A3(n7570), .ZN(n9793) );
  AND2_X1 U7656 ( .A1(n8852), .A2(n8905), .ZN(n8856) );
  AND2_X1 U7657 ( .A1(n9802), .A2(n7657), .ZN(n7656) );
  INV_X1 U7658 ( .A(n7459), .ZN(n8366) );
  AND2_X1 U7659 ( .A1(n8851), .A2(n9383), .ZN(n8905) );
  AND2_X1 U7660 ( .A1(n9792), .A2(n9791), .ZN(n7663) );
  NAND4_X1 U7661 ( .A1(n13391), .A2(n8906), .A3(n8907), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U7662 ( .A1(n8952), .A2(n8275), .ZN(n8964) );
  AND3_X1 U7663 ( .A1(n7658), .A2(n9806), .A3(n9790), .ZN(n7653) );
  AND3_X1 U7664 ( .A1(n8845), .A2(n7759), .A3(n7757), .ZN(n8617) );
  NAND4_X1 U7665 ( .A1(n8909), .A2(n8908), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n8910) );
  AND4_X1 U7666 ( .A1(n7655), .A2(n7654), .A3(n10255), .A4(n10549), .ZN(n7437)
         );
  AND2_X1 U7667 ( .A1(n7661), .A2(n7660), .ZN(n9802) );
  INV_X1 U7668 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7658) );
  NOR2_X1 U7669 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8221) );
  NOR2_X1 U7670 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n8222) );
  NOR2_X1 U7671 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n11102) );
  INV_X1 U7672 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7661) );
  NOR2_X2 U7673 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8952) );
  NOR2_X1 U7674 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8220) );
  NOR2_X1 U7675 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8849) );
  INV_X1 U7676 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9342) );
  NOR2_X2 U7677 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9831) );
  INV_X1 U7678 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9378) );
  INV_X1 U7679 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9379) );
  INV_X1 U7680 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10549) );
  NOR2_X2 U7681 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n10077) );
  XNOR2_X2 U7682 ( .A(n10646), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10650) );
  AOI22_X2 U7683 ( .A1(n15269), .A2(n15261), .B1(n15220), .B2(n15478), .ZN(
        n15252) );
  NOR2_X2 U7684 ( .A1(n9156), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9171) );
  INV_X2 U7685 ( .A(n9890), .ZN(n9840) );
  AOI211_X2 U7686 ( .C1(n15546), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15479) );
  AND2_X2 U7687 ( .A1(n8924), .A2(n8923), .ZN(n14661) );
  OAI21_X2 U7688 ( .B1(n12294), .B2(n7879), .A(n7876), .ZN(n12617) );
  INV_X1 U7689 ( .A(n10208), .ZN(n7423) );
  NAND2_X1 U7690 ( .A1(n9870), .A2(n10674), .ZN(n10208) );
  OR2_X1 U7691 ( .A1(n14293), .A2(n14674), .ZN(n9318) );
  NAND2_X1 U7692 ( .A1(n8777), .A2(n13646), .ZN(n8776) );
  OR2_X1 U7693 ( .A1(n14638), .A2(n14647), .ZN(n9371) );
  AND4_X1 U7694 ( .A1(n9342), .A2(n9378), .A3(n8850), .A4(n9379), .ZN(n9383)
         );
  INV_X1 U7695 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U7696 ( .A1(n16025), .A2(n8681), .ZN(n8025) );
  AND2_X1 U7697 ( .A1(n15991), .A2(n8682), .ZN(n8681) );
  NAND2_X1 U7698 ( .A1(n7703), .A2(n7708), .ZN(n12237) );
  INV_X1 U7699 ( .A(n7704), .ZN(n7701) );
  NOR2_X1 U7700 ( .A1(n9293), .A2(n8343), .ZN(n8342) );
  INV_X1 U7701 ( .A(n9281), .ZN(n8343) );
  NOR2_X1 U7702 ( .A1(n14645), .A2(n8363), .ZN(n8362) );
  INV_X1 U7703 ( .A(n8838), .ZN(n8363) );
  NAND2_X1 U7704 ( .A1(n9797), .A2(n9863), .ZN(n9890) );
  AND2_X1 U7705 ( .A1(n8293), .A2(n7551), .ZN(n8291) );
  INV_X1 U7706 ( .A(n9787), .ZN(n7651) );
  AND3_X1 U7707 ( .A1(n7650), .A2(n7531), .A3(n9831), .ZN(n7652) );
  AND4_X1 U7708 ( .A1(n7658), .A2(n9792), .A3(n9791), .A4(n9795), .ZN(n7650)
         );
  INV_X1 U7709 ( .A(n8668), .ZN(n8667) );
  AOI21_X1 U7710 ( .B1(n8668), .B2(n8666), .A(n8703), .ZN(n8665) );
  INV_X1 U7711 ( .A(n8670), .ZN(n8666) );
  OAI21_X1 U7712 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n10139) );
  NAND2_X1 U7713 ( .A1(n8351), .A2(n8349), .ZN(n13449) );
  NOR2_X1 U7714 ( .A1(n14483), .A2(n8350), .ZN(n8349) );
  INV_X1 U7715 ( .A(n8354), .ZN(n8350) );
  NAND2_X1 U7716 ( .A1(n15174), .A2(n8319), .ZN(n15442) );
  NOR2_X1 U7717 ( .A1(n15439), .A2(n8320), .ZN(n8319) );
  INV_X1 U7718 ( .A(n15173), .ZN(n8320) );
  NAND2_X1 U7719 ( .A1(n15688), .A2(n7988), .ZN(n7984) );
  NOR2_X1 U7720 ( .A1(n8737), .A2(n7989), .ZN(n7988) );
  INV_X1 U7721 ( .A(n7990), .ZN(n7989) );
  OR2_X1 U7722 ( .A1(n16697), .A2(n15643), .ZN(n13417) );
  INV_X1 U7723 ( .A(n8775), .ZN(n8773) );
  NAND2_X1 U7724 ( .A1(n7948), .A2(n7486), .ZN(n7944) );
  NOR2_X1 U7725 ( .A1(n8137), .A2(n8136), .ZN(n8135) );
  AND2_X1 U7726 ( .A1(n13676), .A2(n8138), .ZN(n8137) );
  NOR2_X1 U7727 ( .A1(n8770), .A2(n13673), .ZN(n8136) );
  INV_X1 U7728 ( .A(n13675), .ZN(n8138) );
  NAND2_X1 U7729 ( .A1(n8153), .A2(n13701), .ZN(n8151) );
  NOR2_X1 U7730 ( .A1(n8822), .A2(n10309), .ZN(n8821) );
  AOI21_X1 U7731 ( .B1(n8821), .B2(n8820), .A(n8819), .ZN(n8818) );
  NAND2_X1 U7732 ( .A1(n8822), .A2(n10309), .ZN(n8820) );
  AOI22_X1 U7733 ( .A1(n8814), .A2(n8817), .B1(n7469), .B2(n8821), .ZN(n8813)
         );
  INV_X1 U7734 ( .A(n8818), .ZN(n8817) );
  AND2_X1 U7735 ( .A1(n14323), .A2(n14689), .ZN(n8558) );
  NAND2_X1 U7736 ( .A1(n14664), .A2(n14682), .ZN(n7778) );
  INV_X1 U7737 ( .A(n12297), .ZN(n7880) );
  NOR2_X1 U7738 ( .A1(n8142), .A2(n7427), .ZN(n8140) );
  NOR2_X1 U7739 ( .A1(n8706), .A2(n8072), .ZN(n8071) );
  INV_X1 U7740 ( .A(n14040), .ZN(n8072) );
  INV_X1 U7741 ( .A(n8707), .ZN(n8706) );
  NAND2_X1 U7742 ( .A1(n8208), .A2(n10162), .ZN(n8207) );
  INV_X1 U7743 ( .A(n10182), .ZN(n8208) );
  OR2_X1 U7744 ( .A1(n13531), .A2(n8607), .ZN(n8606) );
  NAND2_X1 U7745 ( .A1(n11321), .A2(n10838), .ZN(n7919) );
  NAND2_X1 U7746 ( .A1(n7697), .A2(n10900), .ZN(n10901) );
  NAND2_X1 U7747 ( .A1(n8323), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U7748 ( .A1(n8322), .A2(n8326), .ZN(n7723) );
  OR2_X1 U7749 ( .A1(n14573), .A2(n7894), .ZN(n7893) );
  NOR2_X1 U7750 ( .A1(n7895), .A2(n14579), .ZN(n7894) );
  INV_X1 U7751 ( .A(n10920), .ZN(n7895) );
  AND2_X1 U7752 ( .A1(n8366), .A2(n8905), .ZN(n7902) );
  AND2_X1 U7753 ( .A1(n7774), .A2(n9023), .ZN(n7773) );
  NAND2_X1 U7754 ( .A1(n8874), .A2(n8875), .ZN(n7774) );
  NAND2_X1 U7755 ( .A1(n8528), .A2(n8530), .ZN(n8527) );
  INV_X1 U7756 ( .A(n8531), .ZN(n8528) );
  NOR2_X1 U7757 ( .A1(n15342), .A2(n8227), .ZN(n8226) );
  XNOR2_X1 U7758 ( .A(n12282), .B(n15096), .ZN(n11827) );
  NOR2_X1 U7759 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7655) );
  NOR2_X1 U7760 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7654) );
  OR2_X1 U7761 ( .A1(n10548), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n10556) );
  AND2_X1 U7762 ( .A1(n7662), .A2(n10255), .ZN(n9803) );
  INV_X1 U7763 ( .A(n13996), .ZN(n8721) );
  INV_X1 U7764 ( .A(n8738), .ZN(n8737) );
  INV_X1 U7765 ( .A(n8062), .ZN(n8061) );
  OAI21_X1 U7766 ( .B1(n8064), .B2(n8063), .A(n15927), .ZN(n8062) );
  INV_X1 U7767 ( .A(n8065), .ZN(n8063) );
  NAND2_X1 U7768 ( .A1(n8662), .A2(n13864), .ZN(n8661) );
  INV_X1 U7769 ( .A(n8663), .ZN(n8662) );
  AOI21_X1 U7770 ( .B1(n8715), .B2(n16574), .A(n7482), .ZN(n8052) );
  INV_X1 U7771 ( .A(n8715), .ZN(n8053) );
  NAND2_X1 U7772 ( .A1(n11762), .A2(n10675), .ZN(n13593) );
  NAND2_X1 U7773 ( .A1(n8669), .A2(n14027), .ZN(n8668) );
  INV_X1 U7774 ( .A(n8671), .ZN(n8669) );
  AOI21_X1 U7775 ( .B1(n16575), .B2(n10779), .A(n10778), .ZN(n12883) );
  NOR2_X1 U7776 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n11101) );
  NAND2_X1 U7777 ( .A1(n10460), .A2(n10459), .ZN(n10472) );
  INV_X1 U7778 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U7779 ( .A1(n8199), .A2(n10253), .ZN(n10275) );
  INV_X1 U7780 ( .A(n10254), .ZN(n10253) );
  INV_X1 U7781 ( .A(n10096), .ZN(n8638) );
  NAND2_X1 U7782 ( .A1(n10043), .A2(n10042), .ZN(n10075) );
  NOR2_X2 U7783 ( .A1(n10705), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n10720) );
  OR2_X1 U7784 ( .A1(n9823), .A2(n9903), .ZN(n9900) );
  NAND2_X1 U7785 ( .A1(n13532), .A2(n7465), .ZN(n8605) );
  AND4_X1 U7786 ( .A1(n8941), .A2(n8938), .A3(n8939), .A4(n8940), .ZN(n9355)
         );
  INV_X1 U7787 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U7788 ( .A1(n8013), .A2(n12189), .ZN(n8012) );
  NAND2_X1 U7789 ( .A1(n10850), .A2(n11259), .ZN(n12375) );
  NOR2_X1 U7790 ( .A1(n7705), .A2(n7710), .ZN(n7709) );
  OR2_X1 U7791 ( .A1(n10869), .A2(n10868), .ZN(n8100) );
  XNOR2_X1 U7792 ( .A(n7893), .B(n14590), .ZN(n10921) );
  AOI21_X1 U7793 ( .B1(n8261), .B2(n8263), .A(n8260), .ZN(n14316) );
  INV_X1 U7794 ( .A(n8262), .ZN(n8260) );
  AOI21_X1 U7795 ( .B1(n8263), .B2(n7777), .A(n14446), .ZN(n8262) );
  AOI21_X1 U7796 ( .B1(n8339), .B2(n8338), .A(n7541), .ZN(n8337) );
  INV_X1 U7797 ( .A(n8342), .ZN(n8338) );
  NAND2_X1 U7798 ( .A1(n9282), .A2(n8342), .ZN(n8341) );
  NAND2_X1 U7799 ( .A1(n7801), .A2(n7799), .ZN(n14734) );
  AOI21_X1 U7800 ( .B1(n7461), .B2(n14342), .A(n7800), .ZN(n7799) );
  INV_X1 U7801 ( .A(n14434), .ZN(n7800) );
  NAND2_X1 U7802 ( .A1(n9102), .A2(n8352), .ZN(n8351) );
  NOR2_X1 U7803 ( .A1(n8353), .A2(n9116), .ZN(n8352) );
  INV_X1 U7804 ( .A(n9101), .ZN(n8353) );
  INV_X1 U7805 ( .A(n16500), .ZN(n14817) );
  NAND2_X1 U7806 ( .A1(n9346), .A2(n14455), .ZN(n16495) );
  NAND2_X1 U7807 ( .A1(n14322), .A2(n9406), .ZN(n16500) );
  NAND2_X1 U7808 ( .A1(n9370), .A2(n14645), .ZN(n14650) );
  CLKBUF_X1 U7809 ( .A(n9078), .Z(n9323) );
  NAND2_X1 U7811 ( .A1(n9395), .A2(n9394), .ZN(n12266) );
  NAND2_X1 U7812 ( .A1(n9390), .A2(n7497), .ZN(n9395) );
  XNOR2_X1 U7813 ( .A(n8858), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U7814 ( .A1(n14950), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U7815 ( .A1(n8859), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8860) );
  OAI22_X1 U7816 ( .A1(n7776), .A2(n7775), .B1(P2_DATAO_REG_25__SCAN_IN), .B2(
        n15627), .ZN(n9306) );
  NAND2_X1 U7817 ( .A1(n9201), .A2(n7741), .ZN(n9337) );
  INV_X1 U7818 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7741) );
  AOI21_X1 U7819 ( .B1(n8561), .B2(n8563), .A(n7625), .ZN(n8560) );
  INV_X1 U7820 ( .A(n8889), .ZN(n8565) );
  OAI21_X1 U7821 ( .B1(n9056), .B2(n9055), .A(n8878), .ZN(n9077) );
  OR2_X1 U7822 ( .A1(n13177), .A2(n13178), .ZN(n13295) );
  NAND2_X1 U7823 ( .A1(n15049), .A2(n7510), .ZN(n14096) );
  INV_X1 U7824 ( .A(n15193), .ZN(n15220) );
  NOR2_X1 U7825 ( .A1(n14973), .A2(n8217), .ZN(n8216) );
  INV_X1 U7826 ( .A(n8548), .ZN(n8217) );
  OAI21_X1 U7827 ( .B1(n13177), .B2(n7677), .A(n7674), .ZN(n13468) );
  INV_X1 U7828 ( .A(n8533), .ZN(n7677) );
  AND2_X1 U7829 ( .A1(n7675), .A2(n13403), .ZN(n7674) );
  XNOR2_X1 U7830 ( .A(n12792), .B(n7695), .ZN(n12730) );
  OR3_X1 U7831 ( .A1(n10171), .A2(n13181), .A3(n10170), .ZN(n10191) );
  AND2_X1 U7832 ( .A1(n10325), .A2(n10324), .ZN(n15184) );
  NAND2_X1 U7833 ( .A1(n15246), .A2(n15470), .ZN(n15231) );
  AOI21_X1 U7834 ( .B1(n8291), .B2(n8289), .A(n7542), .ZN(n8288) );
  INV_X1 U7835 ( .A(n8294), .ZN(n8289) );
  INV_X1 U7836 ( .A(n8291), .ZN(n8290) );
  AND2_X1 U7837 ( .A1(n8387), .A2(n8392), .ZN(n8385) );
  INV_X1 U7838 ( .A(n15306), .ZN(n8392) );
  INV_X1 U7839 ( .A(n13344), .ZN(n7647) );
  NAND2_X1 U7840 ( .A1(n8297), .A2(n8296), .ZN(n12486) );
  NOR2_X1 U7841 ( .A1(n12298), .A2(n7648), .ZN(n8296) );
  INV_X1 U7842 ( .A(n8300), .ZN(n7648) );
  INV_X1 U7843 ( .A(n11226), .ZN(n15446) );
  NAND2_X1 U7844 ( .A1(n10490), .A2(n10489), .ZN(n15478) );
  AND2_X1 U7845 ( .A1(n15723), .A2(n8720), .ZN(n8719) );
  OR2_X1 U7846 ( .A1(n15673), .A2(n8721), .ZN(n8720) );
  NAND2_X1 U7847 ( .A1(n7984), .A2(n7983), .ZN(n15661) );
  NOR2_X1 U7848 ( .A1(n7986), .A2(n15664), .ZN(n7983) );
  AND2_X1 U7849 ( .A1(n8733), .A2(n7993), .ZN(n7992) );
  INV_X1 U7850 ( .A(n13015), .ZN(n8732) );
  AND2_X1 U7851 ( .A1(n8741), .A2(n8739), .ZN(n8738) );
  INV_X1 U7852 ( .A(n11203), .ZN(n8739) );
  OR2_X1 U7853 ( .A1(n11157), .A2(n11156), .ZN(n7990) );
  INV_X1 U7854 ( .A(n13810), .ZN(n13830) );
  NAND2_X1 U7855 ( .A1(n8645), .A2(n7641), .ZN(n13845) );
  NAND2_X1 U7856 ( .A1(n15603), .A2(n13838), .ZN(n8645) );
  INV_X1 U7857 ( .A(n16048), .ZN(n14031) );
  OR2_X1 U7858 ( .A1(n16082), .A2(n15737), .ZN(n8130) );
  NAND2_X1 U7859 ( .A1(n16088), .A2(n15917), .ZN(n8712) );
  NAND2_X1 U7860 ( .A1(n15921), .A2(n15665), .ZN(n8714) );
  NAND2_X1 U7861 ( .A1(n8191), .A2(n15665), .ZN(n8147) );
  OR2_X1 U7862 ( .A1(n15958), .A2(n15976), .ZN(n8689) );
  AND2_X1 U7863 ( .A1(n16111), .A2(n15996), .ZN(n8690) );
  NOR2_X1 U7864 ( .A1(n13420), .A2(n8145), .ZN(n8144) );
  INV_X1 U7865 ( .A(n13417), .ZN(n8145) );
  NAND2_X1 U7866 ( .A1(n12993), .A2(n8076), .ZN(n8075) );
  AND2_X1 U7867 ( .A1(n12992), .A2(n8660), .ZN(n8076) );
  INV_X2 U7868 ( .A(n10937), .ZN(n11178) );
  NAND2_X1 U7869 ( .A1(n16165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10653) );
  AND2_X1 U7870 ( .A1(n11102), .A2(n10612), .ZN(n10614) );
  AND2_X1 U7871 ( .A1(n10613), .A2(n11101), .ZN(n8032) );
  AND2_X1 U7872 ( .A1(n8756), .A2(n8755), .ZN(n10613) );
  NOR2_X1 U7873 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n8756) );
  NOR2_X1 U7874 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8755) );
  INV_X1 U7875 ( .A(n10430), .ZN(n7835) );
  INV_X1 U7876 ( .A(n7834), .ZN(n7833) );
  OAI21_X1 U7877 ( .B1(n7837), .B2(n7458), .A(n10436), .ZN(n7834) );
  OR2_X1 U7878 ( .A1(n10045), .A2(n10069), .ZN(n10068) );
  NAND2_X1 U7879 ( .A1(n8174), .A2(n16464), .ZN(n16352) );
  OAI21_X1 U7880 ( .B1(n16393), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7485), .ZN(
        n7867) );
  OAI21_X1 U7881 ( .B1(n16408), .B2(n16407), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n8175) );
  AOI21_X1 U7882 ( .B1(n14633), .B2(n9326), .A(n8865), .ZN(n14647) );
  NAND2_X1 U7883 ( .A1(n11996), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U7884 ( .A1(n8913), .A2(n8912), .ZN(n14638) );
  OR2_X1 U7885 ( .A1(n9078), .A2(n13916), .ZN(n8912) );
  INV_X1 U7886 ( .A(n14116), .ZN(n8212) );
  AOI21_X1 U7887 ( .B1(n15483), .B2(n15080), .A(n15079), .ZN(n7693) );
  INV_X1 U7888 ( .A(n8099), .ZN(n11764) );
  NAND3_X1 U7889 ( .A1(n7991), .A2(n13324), .A3(n8731), .ZN(n13323) );
  XNOR2_X1 U7890 ( .A(n7867), .B(n16398), .ZN(n7869) );
  OAI211_X1 U7891 ( .C1(n14306), .C2(n9604), .A(n8400), .B(n8399), .ZN(n8398)
         );
  AND2_X1 U7892 ( .A1(n8402), .A2(n8401), .ZN(n8400) );
  NAND2_X1 U7893 ( .A1(n14306), .A2(n9604), .ZN(n8399) );
  NAND2_X1 U7894 ( .A1(keyinput_0), .A2(P3_WR_REG_SCAN_IN), .ZN(n8402) );
  INV_X1 U7895 ( .A(n8397), .ZN(n8396) );
  OAI22_X1 U7896 ( .A1(n9605), .A2(n14960), .B1(SI_29_), .B2(keyinput_3), .ZN(
        n8397) );
  OAI22_X1 U7897 ( .A1(SI_25_), .A2(n9437), .B1(n13303), .B2(keyinput_135), 
        .ZN(n9438) );
  OAI21_X1 U7898 ( .B1(n8477), .B2(n9435), .A(n8475), .ZN(n9440) );
  INV_X1 U7899 ( .A(n8476), .ZN(n8475) );
  AOI21_X1 U7900 ( .B1(n9432), .B2(n9431), .A(n8478), .ZN(n8477) );
  OAI22_X1 U7901 ( .A1(n14969), .A2(keyinput_6), .B1(n9611), .B2(SI_26_), .ZN(
        n9612) );
  NAND2_X1 U7902 ( .A1(n12101), .A2(n10499), .ZN(n9835) );
  NOR2_X1 U7903 ( .A1(n13632), .A2(n13629), .ZN(n8156) );
  NAND2_X1 U7904 ( .A1(n13629), .A2(n13632), .ZN(n8155) );
  NAND2_X1 U7905 ( .A1(n8510), .A2(n8509), .ZN(n8508) );
  AOI22_X1 U7906 ( .A1(n12024), .A2(n9447), .B1(keyinput_141), .B2(SI_19_), 
        .ZN(n8509) );
  NAND2_X1 U7907 ( .A1(n8512), .A2(n8511), .ZN(n8510) );
  NOR3_X1 U7908 ( .A1(n9452), .A2(n9451), .A3(n9453), .ZN(n8507) );
  INV_X1 U7909 ( .A(n7923), .ZN(n7922) );
  AOI21_X1 U7910 ( .B1(n8440), .B2(n8439), .A(n9640), .ZN(n9643) );
  AND2_X1 U7911 ( .A1(n11263), .A2(keyinput_28), .ZN(n8453) );
  NAND2_X1 U7912 ( .A1(n9471), .A2(n9470), .ZN(n8506) );
  NOR2_X1 U7913 ( .A1(n9474), .A2(n7604), .ZN(n8505) );
  XNOR2_X1 U7914 ( .A(keyinput_165), .B(P3_REG3_REG_14__SCAN_IN), .ZN(n8504)
         );
  AND2_X1 U7915 ( .A1(n8776), .A2(n13653), .ZN(n8132) );
  NOR2_X1 U7916 ( .A1(n8777), .A2(n13646), .ZN(n8775) );
  INV_X1 U7917 ( .A(n13657), .ZN(n8786) );
  AOI21_X1 U7918 ( .B1(n9481), .B2(n8483), .A(n9488), .ZN(n8482) );
  AND2_X1 U7919 ( .A1(n9482), .A2(n8484), .ZN(n8483) );
  NAND2_X1 U7920 ( .A1(n9486), .A2(n9487), .ZN(n8481) );
  INV_X1 U7921 ( .A(n8480), .ZN(n8479) );
  OAI22_X1 U7922 ( .A1(n8984), .A2(keyinput_177), .B1(n9489), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n8480) );
  INV_X1 U7923 ( .A(n13660), .ZN(n8165) );
  NOR2_X1 U7924 ( .A1(n13663), .A2(n13660), .ZN(n8166) );
  NAND2_X1 U7925 ( .A1(n7947), .A2(n10094), .ZN(n7946) );
  INV_X1 U7926 ( .A(n10095), .ZN(n7947) );
  NAND2_X1 U7927 ( .A1(n10095), .A2(n7949), .ZN(n7948) );
  NOR2_X1 U7928 ( .A1(n8772), .A2(n13672), .ZN(n8771) );
  INV_X1 U7929 ( .A(n13678), .ZN(n8758) );
  NAND2_X1 U7930 ( .A1(n8519), .A2(n8518), .ZN(n8517) );
  AOI211_X1 U7931 ( .C1(n9503), .C2(n9504), .A(n9502), .B(n9501), .ZN(n8520)
         );
  NAND2_X1 U7932 ( .A1(keyinput_188), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8518)
         );
  INV_X1 U7933 ( .A(n9511), .ZN(n8514) );
  INV_X1 U7934 ( .A(n9510), .ZN(n8515) );
  AOI22_X1 U7935 ( .A1(n12380), .A2(n9506), .B1(keyinput_189), .B2(
        P3_REG3_REG_6__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U7936 ( .A1(n7951), .A2(n7950), .ZN(n10117) );
  AOI21_X1 U7937 ( .B1(n7431), .B2(n7931), .A(n7539), .ZN(n7930) );
  NOR2_X1 U7938 ( .A1(n10135), .A2(n10136), .ZN(n7931) );
  INV_X1 U7939 ( .A(n10159), .ZN(n8811) );
  NAND2_X1 U7940 ( .A1(n7431), .A2(n7933), .ZN(n7932) );
  NAND2_X1 U7941 ( .A1(n10135), .A2(n10136), .ZN(n7933) );
  OAI22_X1 U7942 ( .A1(n12263), .A2(keyinput_72), .B1(n9707), .B2(
        P3_DATAO_REG_24__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U7943 ( .A1(n8826), .A2(n10198), .ZN(n8825) );
  AND2_X1 U7944 ( .A1(n8781), .A2(n13690), .ZN(n8780) );
  INV_X1 U7945 ( .A(n13689), .ZN(n8781) );
  OAI21_X1 U7946 ( .B1(n9529), .B2(n8492), .A(n8491), .ZN(n8490) );
  AOI22_X1 U7947 ( .A1(n12056), .A2(n9531), .B1(keyinput_207), .B2(
        P3_DATAO_REG_17__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U7948 ( .A1(n8494), .A2(n8493), .ZN(n8492) );
  NAND2_X1 U7949 ( .A1(n9535), .A2(n9534), .ZN(n8488) );
  INV_X1 U7950 ( .A(n9536), .ZN(n8489) );
  AOI21_X1 U7951 ( .B1(n7602), .B2(n8425), .A(n8422), .ZN(n9719) );
  NAND2_X1 U7952 ( .A1(n8424), .A2(n8423), .ZN(n8422) );
  AOI22_X1 U7953 ( .A1(n12052), .A2(n9712), .B1(keyinput_78), .B2(
        P3_DATAO_REG_18__SCAN_IN), .ZN(n8425) );
  INV_X1 U7954 ( .A(n10310), .ZN(n8822) );
  OAI21_X1 U7955 ( .B1(n8472), .B2(n8469), .A(n9728), .ZN(n9730) );
  NAND2_X1 U7956 ( .A1(n8471), .A2(n8470), .ZN(n8469) );
  NOR2_X1 U7957 ( .A1(n9569), .A2(n9568), .ZN(n9576) );
  INV_X1 U7958 ( .A(n8813), .ZN(n8812) );
  AOI21_X1 U7959 ( .B1(n7941), .B2(n7439), .A(n7940), .ZN(n7939) );
  INV_X1 U7960 ( .A(n10368), .ZN(n7940) );
  OAI22_X1 U7961 ( .A1(n15576), .A2(n10540), .B1(n15188), .B2(n10499), .ZN(
        n10368) );
  NOR2_X1 U7962 ( .A1(n7439), .A2(n10367), .ZN(n7938) );
  INV_X1 U7963 ( .A(n7942), .ZN(n7941) );
  OAI21_X1 U7964 ( .B1(n7943), .B2(n7439), .A(n10367), .ZN(n7942) );
  INV_X1 U7965 ( .A(n7939), .ZN(n7936) );
  OR2_X1 U7966 ( .A1(n10340), .A2(n10341), .ZN(n7943) );
  INV_X1 U7967 ( .A(n7938), .ZN(n7935) );
  INV_X1 U7968 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n16308) );
  NOR3_X1 U7969 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(n9756) );
  NAND2_X1 U7970 ( .A1(n8557), .A2(n14333), .ZN(n8556) );
  NAND2_X1 U7971 ( .A1(n14492), .A2(n8558), .ZN(n8557) );
  OR2_X1 U7972 ( .A1(n14646), .A2(n14910), .ZN(n8838) );
  INV_X1 U7973 ( .A(n14393), .ZN(n7813) );
  AOI21_X1 U7974 ( .B1(n8251), .B2(n8252), .A(n8249), .ZN(n8248) );
  INV_X1 U7975 ( .A(n14404), .ZN(n8249) );
  NOR2_X1 U7976 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8848) );
  OR2_X1 U7977 ( .A1(n9112), .A2(n8582), .ZN(n8581) );
  INV_X1 U7978 ( .A(n8882), .ZN(n8582) );
  NOR2_X1 U7979 ( .A1(n10406), .A2(n10407), .ZN(n8794) );
  NAND2_X1 U7980 ( .A1(n8071), .A2(n8069), .ZN(n8068) );
  INV_X1 U7981 ( .A(n8709), .ZN(n8069) );
  INV_X1 U7982 ( .A(n8024), .ZN(n8023) );
  INV_X1 U7983 ( .A(n8651), .ZN(n8650) );
  OAI21_X1 U7984 ( .B1(n8653), .B2(n8652), .A(n13307), .ZN(n8651) );
  INV_X1 U7985 ( .A(n10369), .ZN(n8652) );
  AOI21_X1 U7986 ( .B1(n7828), .B2(n8205), .A(n7827), .ZN(n7826) );
  INV_X1 U7987 ( .A(n10201), .ZN(n7827) );
  INV_X1 U7988 ( .A(n7829), .ZN(n7828) );
  OR2_X1 U7989 ( .A1(n16320), .A2(n16321), .ZN(n7859) );
  INV_X1 U7990 ( .A(n13550), .ZN(n8607) );
  OR2_X1 U7991 ( .A1(n14357), .A2(n12468), .ZN(n12265) );
  NAND2_X1 U7992 ( .A1(n12009), .A2(n10881), .ZN(n10882) );
  NAND2_X1 U7993 ( .A1(n8009), .A2(n12259), .ZN(n8007) );
  INV_X1 U7994 ( .A(n10853), .ZN(n8009) );
  NAND2_X1 U7995 ( .A1(n8007), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U7996 ( .A1(n10856), .A2(n11289), .ZN(n10855) );
  INV_X1 U7997 ( .A(n12511), .ZN(n8017) );
  NAND2_X1 U7998 ( .A1(n7699), .A2(n7698), .ZN(n10894) );
  INV_X1 U7999 ( .A(n12506), .ZN(n7698) );
  NAND2_X1 U8000 ( .A1(n8079), .A2(n7615), .ZN(n10898) );
  NAND2_X1 U8001 ( .A1(n10861), .A2(n10862), .ZN(n10863) );
  NAND2_X1 U8002 ( .A1(n7696), .A2(n7904), .ZN(n8323) );
  NAND2_X1 U8003 ( .A1(n7721), .A2(n7720), .ZN(n8332) );
  NAND2_X1 U8004 ( .A1(n14553), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7720) );
  OR2_X1 U8005 ( .A1(n14854), .A2(n14737), .ZN(n14340) );
  NOR2_X1 U8006 ( .A1(n7790), .A2(n13542), .ZN(n7786) );
  INV_X1 U8007 ( .A(n8233), .ZN(n7790) );
  NOR2_X1 U8008 ( .A1(n8237), .A2(n8234), .ZN(n8233) );
  INV_X1 U8009 ( .A(n8235), .ZN(n7788) );
  AOI21_X1 U8010 ( .B1(n14797), .B2(n8236), .A(n7600), .ZN(n8235) );
  INV_X1 U8011 ( .A(n14343), .ZN(n8236) );
  INV_X1 U8012 ( .A(n14416), .ZN(n14816) );
  AND2_X1 U8013 ( .A1(n14411), .A2(n14410), .ZN(n14822) );
  AND4_X1 U8014 ( .A1(n8617), .A2(n8628), .A3(n8367), .A4(n8903), .ZN(n7797)
         );
  NAND2_X1 U8015 ( .A1(n8552), .A2(n8550), .ZN(n8895) );
  NAND2_X1 U8016 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n8551), .ZN(n8550) );
  NOR2_X1 U8017 ( .A1(n9200), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n9201) );
  NAND4_X1 U8018 ( .A1(n7438), .A2(n8366), .A3(n9151), .A4(n8616), .ZN(n9197)
         );
  AND2_X1 U8019 ( .A1(n7758), .A2(n8617), .ZN(n7438) );
  AND2_X1 U8020 ( .A1(n8628), .A2(n8367), .ZN(n7758) );
  INV_X1 U8021 ( .A(n8867), .ZN(n8570) );
  INV_X1 U8022 ( .A(n11975), .ZN(n8538) );
  INV_X1 U8023 ( .A(n13294), .ZN(n7676) );
  NOR2_X1 U8024 ( .A1(n8795), .A2(n10571), .ZN(n10532) );
  AOI21_X1 U8025 ( .B1(n7878), .B2(n7877), .A(n7517), .ZN(n7876) );
  NAND2_X1 U8026 ( .A1(n8750), .A2(n16686), .ZN(n13967) );
  NAND2_X1 U8027 ( .A1(n13800), .A2(n8767), .ZN(n8766) );
  INV_X1 U8028 ( .A(n13801), .ZN(n8767) );
  INV_X1 U8029 ( .A(n8677), .ZN(n8676) );
  OAI21_X1 U8030 ( .B1(n15856), .B2(n8678), .A(n15846), .ZN(n8677) );
  INV_X1 U8031 ( .A(n14028), .ZN(n8678) );
  AOI21_X1 U8032 ( .B1(n15873), .B2(n14049), .A(n15856), .ZN(n8702) );
  NOR2_X1 U8033 ( .A1(n13872), .A2(n8710), .ZN(n8709) );
  INV_X1 U8034 ( .A(n13499), .ZN(n8710) );
  NOR2_X1 U8035 ( .A1(n8658), .A2(n13607), .ZN(n8657) );
  INV_X1 U8036 ( .A(n10770), .ZN(n8658) );
  INV_X1 U8037 ( .A(n13587), .ZN(n10947) );
  AND2_X1 U8038 ( .A1(n14027), .A2(n15912), .ZN(n8670) );
  INV_X1 U8039 ( .A(n14044), .ZN(n8704) );
  NAND2_X1 U8040 ( .A1(n16022), .A2(n16026), .ZN(n8708) );
  INV_X1 U8041 ( .A(n8694), .ZN(n8693) );
  OAI21_X1 U8042 ( .B1(n10775), .B2(n8695), .A(n13860), .ZN(n8694) );
  INV_X1 U8043 ( .A(n10815), .ZN(n11199) );
  INV_X1 U8044 ( .A(n16180), .ZN(n13839) );
  INV_X1 U8045 ( .A(n7855), .ZN(n7854) );
  AOI21_X1 U8046 ( .B1(n7855), .B2(n7853), .A(n7852), .ZN(n7851) );
  INV_X1 U8047 ( .A(n10479), .ZN(n7852) );
  INV_X1 U8048 ( .A(n10471), .ZN(n7853) );
  NAND2_X1 U8049 ( .A1(n10472), .A2(n10471), .ZN(n7857) );
  NOR2_X1 U8050 ( .A1(n10507), .A2(n7856), .ZN(n7855) );
  INV_X1 U8051 ( .A(n10475), .ZN(n7856) );
  INV_X1 U8052 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U8053 ( .A1(n10370), .A2(n10369), .ZN(n10391) );
  AOI21_X1 U8054 ( .B1(n8632), .B2(n8633), .A(n7617), .ZN(n8630) );
  AOI21_X1 U8055 ( .B1(n10296), .B2(n8635), .A(n7619), .ZN(n8634) );
  NAND2_X1 U8056 ( .A1(n10720), .A2(n10635), .ZN(n10642) );
  NAND2_X1 U8057 ( .A1(n10275), .A2(n10274), .ZN(n10297) );
  NAND2_X1 U8058 ( .A1(n10206), .A2(SI_16_), .ZN(n8201) );
  NOR2_X1 U8059 ( .A1(n10206), .A2(SI_16_), .ZN(n8202) );
  INV_X1 U8060 ( .A(n10146), .ZN(n8209) );
  INV_X1 U8061 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10044) );
  AND2_X1 U8062 ( .A1(n9937), .A2(n7441), .ZN(n9924) );
  NAND2_X1 U8063 ( .A1(n9817), .A2(n8377), .ZN(n9819) );
  NAND2_X1 U8064 ( .A1(n9895), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U8065 ( .A1(n16339), .A2(n16338), .ZN(n16343) );
  INV_X1 U8066 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n16341) );
  AOI22_X1 U8067 ( .A1(n16351), .A2(n16350), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n12382), .ZN(n16357) );
  OR2_X1 U8068 ( .A1(n12382), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n16350) );
  NOR2_X1 U8069 ( .A1(n16436), .A2(n16435), .ZN(n16447) );
  AND2_X1 U8070 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n16434), .ZN(n16435) );
  INV_X1 U8071 ( .A(n14366), .ZN(n12544) );
  NAND2_X1 U8072 ( .A1(n7783), .A2(n12078), .ZN(n12711) );
  AOI21_X1 U8073 ( .B1(n7727), .B2(n7728), .A(n7726), .ZN(n7725) );
  INV_X1 U8074 ( .A(n13308), .ZN(n7726) );
  AOI21_X1 U8075 ( .B1(n7465), .B2(n8607), .A(n8604), .ZN(n8603) );
  INV_X1 U8076 ( .A(n13922), .ZN(n8604) );
  OAI211_X1 U8077 ( .C1(n14689), .C2(n14119), .A(n13944), .B(n14234), .ZN(
        n14236) );
  NAND2_X1 U8078 ( .A1(n13940), .A2(n8598), .ZN(n13944) );
  OAI21_X1 U8079 ( .B1(n13939), .B2(n8600), .A(n8599), .ZN(n8598) );
  NAND2_X1 U8080 ( .A1(n13942), .A2(n14267), .ZN(n8599) );
  INV_X1 U8081 ( .A(n9283), .ZN(n8841) );
  NAND2_X1 U8082 ( .A1(n14141), .A2(n8608), .ZN(n12796) );
  NOR2_X1 U8083 ( .A1(n12554), .A2(n8609), .ZN(n8608) );
  INV_X1 U8084 ( .A(n12548), .ZN(n8609) );
  NAND2_X1 U8085 ( .A1(n8623), .A2(n8621), .ZN(n14128) );
  NAND2_X1 U8086 ( .A1(n14274), .A2(n8625), .ZN(n14151) );
  NAND2_X1 U8087 ( .A1(n13087), .A2(n13086), .ZN(n8623) );
  NAND2_X1 U8088 ( .A1(n12273), .A2(n12274), .ZN(n14140) );
  NAND2_X1 U8089 ( .A1(n14210), .A2(n8619), .ZN(n12937) );
  NOR2_X1 U8090 ( .A1(n12940), .A2(n8620), .ZN(n8619) );
  INV_X1 U8091 ( .A(n12798), .ZN(n8620) );
  INV_X1 U8092 ( .A(n12722), .ZN(n14512) );
  INV_X1 U8093 ( .A(n14320), .ZN(n8245) );
  NAND2_X1 U8094 ( .A1(n8330), .A2(n12161), .ZN(n8329) );
  INV_X1 U8095 ( .A(n10882), .ZN(n8330) );
  NAND2_X1 U8096 ( .A1(n10882), .A2(n11262), .ZN(n12405) );
  INV_X1 U8097 ( .A(n8011), .ZN(n8010) );
  NAND2_X1 U8098 ( .A1(n8007), .A2(n12230), .ZN(n12254) );
  NAND2_X1 U8099 ( .A1(n10889), .A2(n12240), .ZN(n12241) );
  INV_X1 U8100 ( .A(n10855), .ZN(n8274) );
  OR2_X1 U8101 ( .A1(n12364), .A2(n8016), .ZN(n8014) );
  NAND2_X1 U8102 ( .A1(n8017), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U8103 ( .A1(n8274), .A2(n8017), .ZN(n8015) );
  NOR2_X1 U8104 ( .A1(n12364), .A2(n13226), .ZN(n12363) );
  OR2_X1 U8105 ( .A1(n12358), .A2(n10893), .ZN(n7699) );
  INV_X1 U8106 ( .A(n10891), .ZN(n10893) );
  INV_X1 U8107 ( .A(n10894), .ZN(n12504) );
  OR2_X1 U8108 ( .A1(n13056), .A2(n13057), .ZN(n10861) );
  OR2_X1 U8109 ( .A1(n12744), .A2(n12745), .ZN(n7918) );
  NAND2_X1 U8110 ( .A1(n7915), .A2(n7919), .ZN(n7914) );
  INV_X1 U8111 ( .A(n7917), .ZN(n7915) );
  INV_X1 U8112 ( .A(n7919), .ZN(n7916) );
  OR2_X1 U8113 ( .A1(n10898), .A2(n14531), .ZN(n7711) );
  NAND2_X1 U8114 ( .A1(n10898), .A2(n14531), .ZN(n10897) );
  AND3_X1 U8115 ( .A1(n7711), .A2(n10897), .A3(P3_REG2_REG_13__SCAN_IN), .ZN(
        n14521) );
  NOR2_X1 U8116 ( .A1(n14542), .A2(n7905), .ZN(n10916) );
  NOR2_X1 U8117 ( .A1(n7906), .A2(n14547), .ZN(n7905) );
  INV_X1 U8118 ( .A(n10841), .ZN(n7906) );
  XNOR2_X1 U8119 ( .A(n8332), .B(n11805), .ZN(n14581) );
  NOR2_X1 U8120 ( .A1(n7639), .A2(n8266), .ZN(n8001) );
  OR2_X1 U8121 ( .A1(n14561), .A2(n7898), .ZN(n7897) );
  NOR2_X1 U8122 ( .A1(n7900), .A2(n7899), .ZN(n7898) );
  INV_X1 U8123 ( .A(n10919), .ZN(n7900) );
  AND2_X1 U8124 ( .A1(n7897), .A2(n7896), .ZN(n14573) );
  INV_X1 U8125 ( .A(n14575), .ZN(n7896) );
  NOR2_X1 U8126 ( .A1(n14579), .A2(n10924), .ZN(n10925) );
  INV_X1 U8127 ( .A(n8332), .ZN(n10924) );
  NAND2_X1 U8128 ( .A1(n14963), .A2(n8963), .ZN(n8574) );
  NAND2_X1 U8129 ( .A1(n8341), .A2(n8345), .ZN(n14670) );
  INV_X1 U8130 ( .A(n14325), .ZN(n14690) );
  NOR2_X1 U8131 ( .A1(n14716), .A2(n8259), .ZN(n8258) );
  INV_X1 U8132 ( .A(n14438), .ZN(n8259) );
  NAND2_X1 U8133 ( .A1(n14734), .A2(n14733), .ZN(n14736) );
  AND2_X1 U8134 ( .A1(n14439), .A2(n14438), .ZN(n14733) );
  OAI21_X1 U8135 ( .B1(n9192), .B2(n8359), .A(n8358), .ZN(n14761) );
  INV_X1 U8136 ( .A(n8360), .ZN(n8359) );
  AOI21_X1 U8137 ( .B1(n8360), .B2(n14797), .A(n7614), .ZN(n8358) );
  NAND2_X1 U8138 ( .A1(n9364), .A2(n14346), .ZN(n14764) );
  NAND2_X1 U8139 ( .A1(n7791), .A2(n14426), .ZN(n14801) );
  NAND2_X1 U8140 ( .A1(n13539), .A2(n8370), .ZN(n7791) );
  NAND2_X1 U8141 ( .A1(n13541), .A2(n13542), .ZN(n13540) );
  INV_X1 U8142 ( .A(n14254), .ZN(n13526) );
  NAND2_X1 U8143 ( .A1(n13264), .A2(n9086), .ZN(n13365) );
  AND2_X1 U8144 ( .A1(n14353), .A2(n14406), .ZN(n14404) );
  INV_X1 U8145 ( .A(n13210), .ZN(n8257) );
  NAND2_X1 U8146 ( .A1(n12964), .A2(n14393), .ZN(n13210) );
  NAND2_X1 U8147 ( .A1(n12965), .A2(n14479), .ZN(n12964) );
  AND3_X1 U8148 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(n12815) );
  AND3_X1 U8149 ( .A1(n8981), .A2(n8980), .A3(n8979), .ZN(n12842) );
  AND2_X1 U8150 ( .A1(n14455), .A2(n12276), .ZN(n14779) );
  INV_X1 U8151 ( .A(n16495), .ZN(n14777) );
  XNOR2_X1 U8152 ( .A(n14366), .B(n16491), .ZN(n16494) );
  INV_X1 U8153 ( .A(n14330), .ZN(n8264) );
  AND2_X1 U8154 ( .A1(n8365), .A2(n8364), .ZN(n14629) );
  NAND2_X1 U8155 ( .A1(n14651), .A2(n8107), .ZN(n14832) );
  INV_X1 U8156 ( .A(n8108), .ZN(n8107) );
  OAI21_X1 U8157 ( .B1(n14653), .B2(n14817), .A(n14652), .ZN(n8108) );
  NAND2_X1 U8158 ( .A1(n12563), .A2(n12722), .ZN(n16663) );
  INV_X1 U8159 ( .A(n14779), .ZN(n16497) );
  INV_X1 U8160 ( .A(n8597), .ZN(n8596) );
  NAND2_X1 U8161 ( .A1(n8093), .A2(n8092), .ZN(n14299) );
  NAND2_X1 U8162 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n13802), .ZN(n8092) );
  NAND2_X1 U8163 ( .A1(n9320), .A2(n9321), .ZN(n8093) );
  INV_X1 U8164 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8903) );
  NOR2_X1 U8165 ( .A1(n9389), .A2(n9388), .ZN(n9411) );
  NAND2_X1 U8166 ( .A1(n7471), .A2(n8091), .ZN(n7776) );
  NAND2_X1 U8167 ( .A1(n7780), .A2(n8576), .ZN(n9271) );
  NAND2_X1 U8168 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n8577), .ZN(n8576) );
  NAND2_X1 U8169 ( .A1(n9258), .A2(n9256), .ZN(n7780) );
  OAI21_X1 U8170 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(n13256), .A(n8897), .ZN(
        n9258) );
  NAND2_X1 U8171 ( .A1(n9243), .A2(n9241), .ZN(n8897) );
  XNOR2_X1 U8172 ( .A(n7740), .B(P3_IR_REG_21__SCAN_IN), .ZN(n14357) );
  OAI21_X1 U8173 ( .B1(n9337), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7740) );
  XNOR2_X1 U8174 ( .A(n8895), .B(n13118), .ZN(n9229) );
  INV_X1 U8175 ( .A(n9201), .ZN(n9216) );
  NAND2_X1 U8176 ( .A1(n8893), .A2(n8892), .ZN(n9196) );
  INV_X1 U8177 ( .A(n7627), .ZN(n8562) );
  INV_X1 U8178 ( .A(n8094), .ZN(n8567) );
  NOR2_X1 U8179 ( .A1(n9094), .A2(n8584), .ZN(n8583) );
  INV_X1 U8180 ( .A(n8879), .ZN(n8584) );
  NAND2_X1 U8181 ( .A1(n9077), .A2(n9076), .ZN(n8880) );
  XNOR2_X1 U8182 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .ZN(n9076) );
  NAND2_X1 U8183 ( .A1(n7766), .A2(n7764), .ZN(n9056) );
  AOI21_X1 U8184 ( .B1(n7476), .B2(n7771), .A(n7765), .ZN(n7764) );
  INV_X1 U8185 ( .A(n8877), .ZN(n7765) );
  AOI21_X1 U8186 ( .B1(n7773), .B2(n7770), .A(n7536), .ZN(n7769) );
  INV_X1 U8187 ( .A(n8875), .ZN(n7770) );
  INV_X1 U8188 ( .A(n7773), .ZN(n7771) );
  XNOR2_X1 U8189 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .ZN(n9023) );
  NOR2_X1 U8190 ( .A1(n8952), .A2(n9386), .ZN(n8276) );
  NAND2_X1 U8191 ( .A1(n8930), .A2(n8866), .ZN(n8951) );
  NAND2_X1 U8192 ( .A1(n14104), .A2(n8549), .ZN(n8548) );
  INV_X1 U8193 ( .A(n14106), .ZN(n8549) );
  INV_X1 U8194 ( .A(n8530), .ZN(n8529) );
  INV_X1 U8195 ( .A(n14076), .ZN(n8540) );
  INV_X1 U8196 ( .A(n13475), .ZN(n8541) );
  NAND2_X1 U8197 ( .A1(n13468), .A2(n13467), .ZN(n13469) );
  NAND2_X1 U8198 ( .A1(n7688), .A2(n7687), .ZN(n15004) );
  NAND2_X1 U8199 ( .A1(n8084), .A2(n7690), .ZN(n7687) );
  OR2_X1 U8200 ( .A1(n10053), .A2(n10052), .ZN(n10088) );
  OR2_X1 U8201 ( .A1(n10301), .A2(n15044), .ZN(n10318) );
  NAND2_X1 U8202 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  INV_X1 U8203 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n13181) );
  NOR2_X1 U8204 ( .A1(n15059), .A2(n8219), .ZN(n8543) );
  INV_X1 U8205 ( .A(n14070), .ZN(n8219) );
  AOI21_X1 U8206 ( .B1(n13294), .B2(n13178), .A(n7496), .ZN(n8536) );
  AND2_X1 U8207 ( .A1(n10286), .A2(n10285), .ZN(n15181) );
  AND3_X1 U8208 ( .A1(n10265), .A2(n10264), .A3(n10263), .ZN(n15203) );
  AND4_X1 U8209 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n13352) );
  AND4_X1 U8210 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n12611) );
  AND3_X1 U8211 ( .A1(n7583), .A2(n9799), .A3(n7882), .ZN(n11723) );
  OR2_X1 U8212 ( .A1(n9887), .A2(n12096), .ZN(n7882) );
  AND2_X1 U8213 ( .A1(n16225), .A2(n16226), .ZN(n7739) );
  AND2_X1 U8214 ( .A1(n7745), .A2(n7744), .ZN(n11498) );
  NAND2_X1 U8215 ( .A1(n11520), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7744) );
  OR2_X1 U8216 ( .A1(n13435), .A2(n7636), .ZN(n7742) );
  NOR2_X1 U8217 ( .A1(n8286), .A2(n15261), .ZN(n8285) );
  INV_X1 U8218 ( .A(n8288), .ZN(n8286) );
  AOI21_X1 U8219 ( .B1(n8294), .B2(n7429), .A(n7540), .ZN(n8293) );
  NOR2_X1 U8220 ( .A1(n15289), .A2(n8295), .ZN(n8294) );
  NOR2_X1 U8221 ( .A1(n7429), .A2(n15306), .ZN(n8295) );
  AOI21_X1 U8222 ( .B1(n8389), .B2(n8388), .A(n7521), .ZN(n8387) );
  INV_X1 U8223 ( .A(n7463), .ZN(n8388) );
  NAND2_X1 U8224 ( .A1(n8390), .A2(n8393), .ZN(n15322) );
  NAND2_X1 U8225 ( .A1(n8391), .A2(n7463), .ZN(n8390) );
  INV_X1 U8226 ( .A(n15347), .ZN(n8391) );
  NAND2_X1 U8227 ( .A1(n8308), .A2(n7424), .ZN(n8305) );
  AOI21_X1 U8228 ( .B1(n8412), .B2(n8411), .A(n7519), .ZN(n8410) );
  INV_X1 U8229 ( .A(n15209), .ZN(n8411) );
  AND2_X1 U8230 ( .A1(n7442), .A2(n15182), .ZN(n8311) );
  AOI21_X1 U8231 ( .B1(n8406), .B2(n8405), .A(n7518), .ZN(n8404) );
  NAND2_X1 U8232 ( .A1(n12635), .A2(n12618), .ZN(n12620) );
  NAND2_X1 U8233 ( .A1(n12620), .A2(n12619), .ZN(n12919) );
  NAND2_X1 U8234 ( .A1(n12294), .A2(n12293), .ZN(n7881) );
  INV_X1 U8235 ( .A(n11829), .ZN(n8280) );
  XNOR2_X1 U8236 ( .A(n16521), .B(n11723), .ZN(n12091) );
  INV_X1 U8237 ( .A(n12091), .ZN(n12102) );
  NAND2_X1 U8238 ( .A1(n9829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9826) );
  XNOR2_X1 U8239 ( .A(n11662), .B(n13431), .ZN(n11223) );
  AND2_X1 U8240 ( .A1(n9949), .A2(n9948), .ZN(n11968) );
  AND2_X1 U8241 ( .A1(n9788), .A2(n9789), .ZN(n7649) );
  INV_X1 U8242 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U8243 ( .A1(n10557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U8244 ( .A1(n10561), .A2(n10560), .ZN(n10563) );
  OR2_X1 U8245 ( .A1(n9946), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9997) );
  AOI21_X1 U8246 ( .B1(n8719), .B2(n8721), .A(n7512), .ZN(n8717) );
  NAND2_X1 U8247 ( .A1(n13481), .A2(n7509), .ZN(n8083) );
  INV_X1 U8248 ( .A(n15739), .ZN(n15976) );
  AOI21_X1 U8249 ( .B1(n8717), .B2(n7979), .A(n7978), .ZN(n7977) );
  INV_X1 U8250 ( .A(n8719), .ZN(n7979) );
  INV_X1 U8251 ( .A(n15631), .ZN(n7978) );
  NAND2_X1 U8252 ( .A1(n15687), .A2(n7990), .ZN(n7987) );
  AOI21_X1 U8253 ( .B1(n8738), .B2(n8736), .A(n7490), .ZN(n8735) );
  INV_X1 U8254 ( .A(n8725), .ZN(n8724) );
  OAI21_X1 U8255 ( .B1(n15705), .B2(n8726), .A(n15649), .ZN(n8725) );
  INV_X1 U8256 ( .A(n13975), .ZN(n8726) );
  OAI21_X1 U8257 ( .B1(n11032), .B2(n11031), .A(n11866), .ZN(n11039) );
  NAND2_X1 U8258 ( .A1(n15661), .A2(n13966), .ZN(n15704) );
  XNOR2_X1 U8259 ( .A(n11012), .B(n11072), .ZN(n11020) );
  NAND2_X1 U8260 ( .A1(n7962), .A2(n12068), .ZN(n7961) );
  INV_X1 U8261 ( .A(n7964), .ZN(n7962) );
  OR2_X1 U8262 ( .A1(n7965), .A2(n11986), .ZN(n7964) );
  INV_X1 U8263 ( .A(n7968), .ZN(n7965) );
  INV_X1 U8264 ( .A(n13829), .ZN(n13807) );
  OR2_X1 U8265 ( .A1(n10679), .A2(n10669), .ZN(n8159) );
  OR2_X1 U8266 ( .A1(n11079), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10953) );
  AND2_X1 U8267 ( .A1(n11305), .A2(n13712), .ZN(n11330) );
  NAND2_X1 U8268 ( .A1(n15887), .A2(n8193), .ZN(n15834) );
  NOR2_X1 U8269 ( .A1(n16054), .A2(n8195), .ZN(n8193) );
  AND2_X1 U8270 ( .A1(n14026), .A2(n7484), .ZN(n8671) );
  NAND2_X1 U8271 ( .A1(n15901), .A2(n15912), .ZN(n8672) );
  AOI21_X1 U8272 ( .B1(n8061), .B2(n8063), .A(n7538), .ZN(n8058) );
  NOR2_X1 U8273 ( .A1(n15934), .A2(n8110), .ZN(n8064) );
  NAND2_X1 U8274 ( .A1(n8066), .A2(n8149), .ZN(n8065) );
  OAI21_X1 U8275 ( .B1(n15966), .B2(n8063), .A(n8061), .ZN(n15926) );
  NOR2_X1 U8276 ( .A1(n15927), .A2(n8043), .ZN(n8042) );
  INV_X1 U8277 ( .A(n8045), .ZN(n8043) );
  NAND2_X1 U8278 ( .A1(n10939), .A2(n10938), .ZN(n15958) );
  NAND2_X1 U8279 ( .A1(n15951), .A2(n15963), .ZN(n15950) );
  NAND2_X1 U8280 ( .A1(n15990), .A2(n14045), .ZN(n14047) );
  NOR2_X1 U8281 ( .A1(n16129), .A2(n8187), .ZN(n8185) );
  OR2_X1 U8282 ( .A1(n16718), .A2(n16030), .ZN(n14023) );
  NAND2_X1 U8283 ( .A1(n14041), .A2(n14040), .ZN(n16022) );
  NAND2_X1 U8284 ( .A1(n13500), .A2(n8709), .ZN(n14041) );
  AND2_X1 U8285 ( .A1(n11072), .A2(n10649), .ZN(n12431) );
  INV_X1 U8286 ( .A(n13870), .ZN(n13420) );
  OR2_X1 U8287 ( .A1(n13659), .A2(n13221), .ZN(n13139) );
  NOR2_X1 U8288 ( .A1(n13869), .A2(n8074), .ZN(n8073) );
  INV_X1 U8289 ( .A(n13150), .ZN(n8074) );
  OR2_X1 U8290 ( .A1(n7589), .A2(n8661), .ZN(n12996) );
  AOI21_X1 U8291 ( .B1(n8661), .B2(n12995), .A(n8660), .ZN(n8659) );
  AND2_X1 U8292 ( .A1(n10808), .A2(n15761), .ZN(n15955) );
  NAND2_X1 U8293 ( .A1(n11061), .A2(n11060), .ZN(n13649) );
  NAND2_X1 U8294 ( .A1(n8041), .A2(n15750), .ZN(n8040) );
  AND2_X1 U8295 ( .A1(n13863), .A2(n10753), .ZN(n8715) );
  NAND2_X1 U8296 ( .A1(n16570), .A2(n16569), .ZN(n10754) );
  NAND2_X1 U8297 ( .A1(n10742), .A2(n10741), .ZN(n13633) );
  INV_X1 U8298 ( .A(n13858), .ZN(n10775) );
  INV_X1 U8299 ( .A(n10937), .ZN(n8048) );
  NAND2_X1 U8300 ( .A1(n11763), .A2(n13854), .ZN(n11778) );
  INV_X1 U8301 ( .A(n11576), .ZN(n11763) );
  OR2_X1 U8302 ( .A1(n15761), .A2(n13840), .ZN(n16029) );
  NOR2_X1 U8303 ( .A1(n11760), .A2(n8018), .ZN(n11768) );
  AND2_X1 U8304 ( .A1(n13854), .A2(n11761), .ZN(n8018) );
  NAND2_X1 U8305 ( .A1(n11764), .A2(n13584), .ZN(n11576) );
  NAND2_X1 U8306 ( .A1(n12431), .A2(n16033), .ZN(n16619) );
  NAND2_X1 U8307 ( .A1(n10971), .A2(n10970), .ZN(n16697) );
  OR2_X1 U8308 ( .A1(n13828), .A2(n10782), .ZN(n16623) );
  NAND2_X1 U8309 ( .A1(n16619), .A2(n16602), .ZN(n16705) );
  NAND2_X1 U8310 ( .A1(n11200), .A2(n11199), .ZN(n16684) );
  NAND2_X1 U8311 ( .A1(n7832), .A2(n7831), .ZN(n10460) );
  AOI21_X1 U8312 ( .B1(n7833), .B2(n7458), .A(n7634), .ZN(n7831) );
  NAND2_X1 U8313 ( .A1(n8031), .A2(n8030), .ZN(n10651) );
  NAND2_X1 U8314 ( .A1(n10625), .A2(n10621), .ZN(n7959) );
  INV_X1 U8315 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8748) );
  OAI21_X1 U8316 ( .B1(n10645), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10641) );
  INV_X1 U8317 ( .A(n10642), .ZN(n8087) );
  AND2_X1 U8318 ( .A1(n10275), .A2(n8198), .ZN(n12847) );
  NAND2_X1 U8319 ( .A1(n7825), .A2(n8205), .ZN(n10202) );
  NAND2_X1 U8320 ( .A1(n10139), .A2(n7829), .ZN(n7825) );
  NAND2_X1 U8321 ( .A1(n10139), .A2(n10138), .ZN(n10142) );
  NAND2_X1 U8322 ( .A1(n10142), .A2(n7466), .ZN(n10163) );
  OR2_X1 U8323 ( .A1(n10074), .A2(n8643), .ZN(n8642) );
  NAND2_X1 U8324 ( .A1(n10066), .A2(n8111), .ZN(n10045) );
  NAND2_X1 U8325 ( .A1(n8113), .A2(n8112), .ZN(n8111) );
  INV_X1 U8326 ( .A(n10075), .ZN(n8113) );
  NAND2_X1 U8327 ( .A1(n10013), .A2(n10012), .ZN(n10018) );
  OAI21_X1 U8328 ( .B1(n9995), .B2(n7686), .A(n7684), .ZN(n10043) );
  INV_X1 U8329 ( .A(n7685), .ZN(n7684) );
  INV_X1 U8330 ( .A(n10012), .ZN(n7686) );
  NAND2_X1 U8331 ( .A1(n9995), .A2(n9994), .ZN(n10013) );
  INV_X1 U8332 ( .A(n10674), .ZN(n8230) );
  AND2_X1 U8333 ( .A1(n9900), .A2(n9824), .ZN(n11290) );
  INV_X1 U8334 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n16310) );
  OAI21_X1 U8335 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(P1_ADDR_REG_1__SCAN_IN), 
        .A(n8173), .ZN(n8172) );
  NAND2_X1 U8336 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n8173) );
  NAND2_X1 U8337 ( .A1(n16333), .A2(n16334), .ZN(n16348) );
  NAND2_X1 U8338 ( .A1(n16355), .A2(n16356), .ZN(n16368) );
  AOI21_X1 U8339 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16376), .A(n16375), .ZN(
        n16388) );
  AND2_X1 U8340 ( .A1(n16423), .A2(n7849), .ZN(n7846) );
  INV_X1 U8341 ( .A(n7848), .ZN(n7845) );
  NAND2_X1 U8342 ( .A1(n7850), .A2(n13113), .ZN(n7849) );
  NAND2_X1 U8343 ( .A1(n16417), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U8344 ( .A1(n8589), .A2(n16446), .ZN(n16454) );
  NAND2_X1 U8345 ( .A1(n16444), .A2(n16445), .ZN(n8589) );
  NOR2_X1 U8346 ( .A1(n14284), .A2(n7522), .ZN(n8611) );
  AND3_X1 U8347 ( .A1(n8968), .A2(n8967), .A3(n8966), .ZN(n14145) );
  OR2_X1 U8348 ( .A1(n9078), .A2(SI_3_), .ZN(n8967) );
  NAND2_X1 U8349 ( .A1(n9220), .A2(n9219), .ZN(n14160) );
  NAND2_X1 U8350 ( .A1(n8615), .A2(n13953), .ZN(n8612) );
  NAND2_X1 U8351 ( .A1(n8615), .A2(n8614), .ZN(n8613) );
  INV_X1 U8352 ( .A(n14285), .ZN(n8614) );
  OR2_X1 U8353 ( .A1(n12350), .A2(n12351), .ZN(n12348) );
  OR2_X1 U8354 ( .A1(n12354), .A2(n7782), .ZN(n7781) );
  AND2_X1 U8355 ( .A1(n7422), .A2(n7783), .ZN(n7782) );
  NAND2_X1 U8356 ( .A1(n7736), .A2(n7735), .ZN(n14186) );
  AOI21_X1 U8357 ( .B1(n7737), .B2(n8626), .A(n7603), .ZN(n7735) );
  NAND2_X1 U8358 ( .A1(n9245), .A2(n9244), .ZN(n14191) );
  AOI21_X1 U8359 ( .B1(n7732), .B2(n7734), .A(n7731), .ZN(n7730) );
  INV_X1 U8360 ( .A(n14225), .ZN(n7731) );
  NAND2_X1 U8361 ( .A1(n8610), .A2(n14140), .ZN(n14141) );
  AND2_X1 U8362 ( .A1(n14142), .A2(n14139), .ZN(n8610) );
  OAI21_X1 U8363 ( .B1(n14276), .B2(n8626), .A(n7737), .ZN(n14245) );
  NAND2_X2 U8364 ( .A1(n12126), .A2(n12125), .ZN(n14287) );
  NAND2_X1 U8365 ( .A1(n12137), .A2(n14792), .ZN(n14292) );
  NAND4_X1 U8366 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n12556)
         );
  INV_X1 U8367 ( .A(n9355), .ZN(n7783) );
  OAI21_X1 U8368 ( .B1(n12164), .B2(n12165), .A(n7491), .ZN(n12017) );
  NOR2_X1 U8369 ( .A1(n8964), .A2(n8618), .ZN(n8995) );
  NAND2_X1 U8370 ( .A1(n8845), .A2(n7759), .ZN(n8618) );
  NOR2_X1 U8371 ( .A1(n12359), .A2(n9050), .ZN(n12358) );
  INV_X1 U8372 ( .A(n8100), .ZN(n10929) );
  XNOR2_X1 U8373 ( .A(n10916), .B(n7904), .ZN(n10843) );
  NOR2_X1 U8374 ( .A1(n10843), .A2(n10842), .ZN(n10917) );
  INV_X1 U8375 ( .A(n14604), .ZN(n14574) );
  NAND2_X1 U8376 ( .A1(n8100), .A2(n10928), .ZN(n8267) );
  INV_X1 U8377 ( .A(n7721), .ZN(n14557) );
  NOR2_X1 U8378 ( .A1(n14569), .A2(n14570), .ZN(n14568) );
  INV_X1 U8379 ( .A(n14610), .ZN(n8077) );
  XNOR2_X1 U8380 ( .A(n7892), .B(n14596), .ZN(n7891) );
  NOR2_X1 U8381 ( .A1(n14591), .A2(n8102), .ZN(n7892) );
  NOR2_X1 U8382 ( .A1(n10875), .A2(n10874), .ZN(n14604) );
  AOI21_X1 U8383 ( .B1(n9354), .B2(n16500), .A(n9353), .ZN(n14621) );
  NAND2_X1 U8384 ( .A1(n8574), .A2(n8917), .ZN(n14655) );
  NAND2_X1 U8385 ( .A1(n9297), .A2(n9296), .ZN(n14681) );
  OR2_X1 U8386 ( .A1(n9078), .A2(n13303), .ZN(n9296) );
  NAND2_X1 U8387 ( .A1(n9155), .A2(n9154), .ZN(n14886) );
  AND2_X1 U8388 ( .A1(n9115), .A2(n9114), .ZN(n16673) );
  AND2_X1 U8389 ( .A1(n14650), .A2(n8263), .ZN(n14637) );
  NAND2_X1 U8390 ( .A1(n16666), .A2(n16724), .ZN(n7818) );
  NAND2_X1 U8391 ( .A1(n7821), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7820) );
  INV_X1 U8392 ( .A(n14636), .ZN(n7819) );
  NOR2_X1 U8393 ( .A1(n10606), .A2(n14938), .ZN(n9418) );
  OAI21_X1 U8394 ( .B1(n9167), .B2(n9166), .A(n9181), .ZN(n14553) );
  INV_X1 U8395 ( .A(SI_12_), .ZN(n11319) );
  AND2_X1 U8396 ( .A1(n15078), .A2(n8548), .ZN(n8547) );
  AND2_X1 U8397 ( .A1(n14977), .A2(n8203), .ZN(n14983) );
  NOR2_X1 U8398 ( .A1(n14117), .A2(n7499), .ZN(n8213) );
  INV_X1 U8399 ( .A(n8218), .ZN(n8214) );
  INV_X1 U8400 ( .A(n8216), .ZN(n8215) );
  AND2_X1 U8401 ( .A1(n15078), .A2(n8216), .ZN(n14972) );
  NAND2_X1 U8402 ( .A1(n13469), .A2(n13475), .ZN(n14071) );
  NAND2_X1 U8403 ( .A1(n10332), .A2(n10331), .ZN(n15342) );
  NAND2_X1 U8404 ( .A1(n11689), .A2(n15427), .ZN(n15080) );
  NAND2_X1 U8405 ( .A1(n9837), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U8406 ( .A1(n9866), .A2(n9865), .ZN(n15099) );
  INV_X1 U8407 ( .A(n7745), .ZN(n11509) );
  INV_X1 U8408 ( .A(n7750), .ZN(n12653) );
  NOR2_X1 U8409 ( .A1(n13101), .A2(n13100), .ZN(n13435) );
  XNOR2_X1 U8410 ( .A(n7742), .B(n15117), .ZN(n13437) );
  INV_X1 U8411 ( .A(n7747), .ZN(n16250) );
  NAND2_X1 U8412 ( .A1(n15254), .A2(n15253), .ZN(n15472) );
  NAND2_X1 U8413 ( .A1(n8408), .A2(n8406), .ZN(n15421) );
  NAND2_X1 U8414 ( .A1(n15442), .A2(n15176), .ZN(n15417) );
  NAND2_X1 U8415 ( .A1(n8297), .A2(n8300), .ZN(n12291) );
  NAND2_X1 U8416 ( .A1(n15463), .A2(n15464), .ZN(n15553) );
  AND2_X1 U8417 ( .A1(n8103), .A2(n7594), .ZN(n7873) );
  AND2_X1 U8418 ( .A1(n15469), .A2(n8104), .ZN(n8103) );
  NAND2_X1 U8419 ( .A1(n15236), .A2(n15546), .ZN(n8104) );
  OAI21_X1 U8420 ( .B1(n11450), .B2(n10208), .A(n10051), .ZN(n12792) );
  NAND2_X1 U8421 ( .A1(n7822), .A2(n10482), .ZN(n15552) );
  NAND2_X1 U8422 ( .A1(n15603), .A2(n7423), .ZN(n7822) );
  OR2_X1 U8423 ( .A1(n15553), .A2(n16527), .ZN(n7671) );
  INV_X1 U8424 ( .A(n15471), .ZN(n8124) );
  NAND2_X1 U8425 ( .A1(n15222), .A2(n7425), .ZN(n8314) );
  NOR2_X1 U8426 ( .A1(n15222), .A2(n7425), .ZN(n8313) );
  NAND2_X1 U8427 ( .A1(n15586), .A2(n15546), .ZN(n15594) );
  OAI21_X1 U8428 ( .B1(n11234), .B2(P2_D_REG_0__SCAN_IN), .A(n11233), .ZN(
        n16222) );
  INV_X1 U8429 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U8430 ( .A1(n10810), .A2(n10631), .ZN(n11015) );
  NOR2_X1 U8431 ( .A1(n16176), .A2(n13516), .ZN(n10631) );
  NAND2_X1 U8432 ( .A1(n10960), .A2(n10959), .ZN(n16137) );
  NAND2_X1 U8433 ( .A1(n13732), .A2(n13731), .ZN(n16088) );
  NAND2_X1 U8434 ( .A1(n12894), .A2(n7993), .ZN(n13016) );
  INV_X1 U8435 ( .A(n15756), .ZN(n13581) );
  NAND2_X1 U8436 ( .A1(n13989), .A2(n13988), .ZN(n15672) );
  NAND2_X1 U8437 ( .A1(n15696), .A2(n15697), .ZN(n13989) );
  OR2_X1 U8438 ( .A1(n11039), .A2(n11038), .ZN(n11901) );
  NAND2_X1 U8439 ( .A1(n8740), .A2(n8741), .ZN(n11202) );
  NAND2_X1 U8440 ( .A1(n15713), .A2(n8743), .ZN(n8740) );
  NAND2_X1 U8441 ( .A1(n8118), .A2(n8117), .ZN(n8116) );
  INV_X1 U8442 ( .A(n11095), .ZN(n8117) );
  INV_X1 U8443 ( .A(n11094), .ZN(n8118) );
  NAND2_X1 U8444 ( .A1(n13776), .A2(n13775), .ZN(n16069) );
  OR2_X1 U8445 ( .A1(n11537), .A2(P1_U3086), .ZN(n16723) );
  INV_X1 U8446 ( .A(n13914), .ZN(n8164) );
  INV_X1 U8447 ( .A(n13913), .ZN(n8163) );
  NAND2_X1 U8448 ( .A1(n11189), .A2(n11188), .ZN(n15954) );
  OR2_X1 U8449 ( .A1(n10677), .A2(n10656), .ZN(n8691) );
  AND2_X1 U8450 ( .A1(n13569), .A2(n13568), .ZN(n16048) );
  INV_X1 U8451 ( .A(n14052), .ZN(n8027) );
  INV_X1 U8452 ( .A(n14030), .ZN(n8028) );
  XNOR2_X1 U8453 ( .A(n16348), .B(n16347), .ZN(n16349) );
  XNOR2_X1 U8454 ( .A(n16368), .B(n8587), .ZN(n16370) );
  INV_X1 U8455 ( .A(n16369), .ZN(n8587) );
  AOI21_X1 U8456 ( .B1(n16381), .B2(n16380), .A(n16379), .ZN(n16384) );
  AND2_X1 U8457 ( .A1(n8585), .A2(n7547), .ZN(n16408) );
  NAND2_X1 U8458 ( .A1(n7869), .A2(n7868), .ZN(n8585) );
  INV_X1 U8459 ( .A(n7867), .ZN(n16399) );
  NAND2_X1 U8460 ( .A1(n16408), .A2(n16407), .ZN(n16409) );
  NOR2_X1 U8461 ( .A1(n16424), .A2(n16423), .ZN(n16431) );
  NAND2_X1 U8462 ( .A1(n7843), .A2(n7848), .ZN(n16424) );
  NAND2_X1 U8463 ( .A1(n16416), .A2(n7849), .ZN(n7843) );
  AOI21_X1 U8464 ( .B1(n8178), .B2(n8177), .A(n16431), .ZN(n16439) );
  INV_X1 U8465 ( .A(n16430), .ZN(n8178) );
  XNOR2_X1 U8466 ( .A(n16454), .B(n8588), .ZN(n16453) );
  INV_X1 U8467 ( .A(n16455), .ZN(n8588) );
  NAND2_X1 U8468 ( .A1(n16453), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U8469 ( .A1(keyinput_2), .A2(SI_30_), .ZN(n8401) );
  INV_X1 U8470 ( .A(n9430), .ZN(n9431) );
  OAI22_X1 U8471 ( .A1(n9433), .A2(n13916), .B1(SI_28_), .B2(keyinput_132), 
        .ZN(n8478) );
  OAI22_X1 U8472 ( .A1(n14969), .A2(keyinput_134), .B1(n9436), .B2(SI_26_), 
        .ZN(n8476) );
  NAND2_X1 U8473 ( .A1(n8395), .A2(n9608), .ZN(n9609) );
  OAI21_X1 U8474 ( .B1(n9603), .B2(n8398), .A(n8396), .ZN(n8395) );
  OAI22_X1 U8475 ( .A1(SI_28_), .A2(n9606), .B1(n13916), .B2(keyinput_4), .ZN(
        n9607) );
  NAND2_X1 U8476 ( .A1(n9445), .A2(n9446), .ZN(n8512) );
  NOR2_X1 U8477 ( .A1(n9444), .A2(n9443), .ZN(n8511) );
  NAND2_X1 U8478 ( .A1(n9622), .A2(n9623), .ZN(n8446) );
  NOR2_X1 U8479 ( .A1(n9621), .A2(n9620), .ZN(n8445) );
  NAND2_X1 U8480 ( .A1(n12024), .A2(keyinput_13), .ZN(n8443) );
  NAND2_X1 U8481 ( .A1(n8444), .A2(n8441), .ZN(n8440) );
  AND2_X1 U8482 ( .A1(n8443), .A2(n8442), .ZN(n8441) );
  NAND2_X1 U8483 ( .A1(n8446), .A2(n8445), .ZN(n8444) );
  NAND2_X1 U8484 ( .A1(n9624), .A2(SI_19_), .ZN(n8442) );
  NOR3_X1 U8485 ( .A1(n9628), .A2(n9630), .A3(n9629), .ZN(n8439) );
  INV_X1 U8486 ( .A(n13634), .ZN(n8779) );
  AOI21_X1 U8487 ( .B1(n8508), .B2(n8507), .A(n9462), .ZN(n9465) );
  NAND2_X1 U8488 ( .A1(n9886), .A2(n7925), .ZN(n8806) );
  NAND2_X1 U8489 ( .A1(n8452), .A2(n9650), .ZN(n8451) );
  OAI21_X1 U8490 ( .B1(n9646), .B2(n8453), .A(n9645), .ZN(n8452) );
  NOR2_X1 U8491 ( .A1(n9648), .A2(n9649), .ZN(n8450) );
  AOI22_X1 U8492 ( .A1(n9477), .A2(n9476), .B1(keyinput_167), .B2(
        P3_REG3_REG_10__SCAN_IN), .ZN(n9478) );
  AOI21_X1 U8493 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n9477) );
  XNOR2_X1 U8494 ( .A(n8485), .B(P3_REG3_REG_19__SCAN_IN), .ZN(n8484) );
  INV_X1 U8495 ( .A(keyinput_169), .ZN(n8485) );
  NAND2_X1 U8496 ( .A1(n8449), .A2(n8447), .ZN(n9653) );
  NOR2_X1 U8497 ( .A1(n9652), .A2(n8448), .ZN(n8447) );
  NAND2_X1 U8498 ( .A1(n8451), .A2(n8450), .ZN(n8449) );
  XNOR2_X1 U8499 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n8448) );
  INV_X1 U8500 ( .A(n10010), .ZN(n8803) );
  NAND2_X1 U8501 ( .A1(n8786), .A2(n13658), .ZN(n8785) );
  NAND2_X1 U8502 ( .A1(n8784), .A2(n13657), .ZN(n8783) );
  INV_X1 U8503 ( .A(n13658), .ZN(n8784) );
  AND2_X1 U8504 ( .A1(n9660), .A2(n8420), .ZN(n8419) );
  XNOR2_X1 U8505 ( .A(n8421), .B(P3_REG3_REG_8__SCAN_IN), .ZN(n8420) );
  INV_X1 U8506 ( .A(keyinput_43), .ZN(n8421) );
  OAI22_X1 U8507 ( .A1(n8984), .A2(n9668), .B1(P3_REG3_REG_5__SCAN_IN), .B2(
        keyinput_49), .ZN(n8416) );
  INV_X1 U8508 ( .A(n13672), .ZN(n8770) );
  OAI21_X1 U8509 ( .B1(n8482), .B2(n8481), .A(n8479), .ZN(n9490) );
  OAI21_X1 U8510 ( .B1(n8418), .B2(n8417), .A(n8415), .ZN(n9673) );
  INV_X1 U8511 ( .A(n8416), .ZN(n8415) );
  NAND2_X1 U8512 ( .A1(n9666), .A2(n9665), .ZN(n8417) );
  AOI21_X1 U8513 ( .B1(n9659), .B2(n8419), .A(n9667), .ZN(n8418) );
  INV_X1 U8514 ( .A(n13673), .ZN(n8772) );
  NAND2_X1 U8515 ( .A1(n9689), .A2(n9505), .ZN(n8519) );
  INV_X1 U8516 ( .A(n7948), .ZN(n7945) );
  NAND2_X1 U8517 ( .A1(n8438), .A2(n9688), .ZN(n8437) );
  NAND2_X1 U8518 ( .A1(n9681), .A2(n9680), .ZN(n8438) );
  NOR2_X1 U8519 ( .A1(n9687), .A2(n9686), .ZN(n8436) );
  NAND2_X1 U8520 ( .A1(n12380), .A2(n9691), .ZN(n8431) );
  NAND2_X1 U8521 ( .A1(keyinput_61), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8430)
         );
  NAND2_X1 U8522 ( .A1(n9689), .A2(keyinput_60), .ZN(n8434) );
  NAND2_X1 U8523 ( .A1(n9690), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U8524 ( .A1(n10200), .A2(n10199), .ZN(n8827) );
  AND2_X1 U8525 ( .A1(n13680), .A2(n8758), .ZN(n8757) );
  AOI21_X1 U8526 ( .B1(n7513), .B2(n8516), .A(n8513), .ZN(n9516) );
  AOI21_X1 U8527 ( .B1(n8435), .B2(n8432), .A(n8429), .ZN(n9700) );
  AND2_X1 U8528 ( .A1(n8434), .A2(n8433), .ZN(n8432) );
  NAND2_X1 U8529 ( .A1(n8431), .A2(n8430), .ZN(n8429) );
  NAND2_X1 U8530 ( .A1(n8437), .A2(n8436), .ZN(n8435) );
  AOI21_X1 U8531 ( .B1(n7930), .B2(n7932), .A(n7928), .ZN(n7927) );
  INV_X1 U8532 ( .A(n10200), .ZN(n8826) );
  NAND2_X1 U8533 ( .A1(n12052), .A2(n9530), .ZN(n8494) );
  NAND2_X1 U8534 ( .A1(keyinput_206), .A2(P3_DATAO_REG_18__SCAN_IN), .ZN(n8493) );
  AOI21_X1 U8535 ( .B1(n9706), .B2(n8427), .A(n7640), .ZN(n8426) );
  INV_X1 U8536 ( .A(n8428), .ZN(n8427) );
  NAND2_X1 U8537 ( .A1(n12056), .A2(keyinput_79), .ZN(n8424) );
  NAND2_X1 U8538 ( .A1(n9713), .A2(P3_DATAO_REG_17__SCAN_IN), .ZN(n8423) );
  OAI22_X1 U8539 ( .A1(n12036), .A2(keyinput_213), .B1(n9537), .B2(
        P3_DATAO_REG_11__SCAN_IN), .ZN(n8486) );
  AOI21_X1 U8540 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8487) );
  NAND2_X1 U8541 ( .A1(keyinput_87), .A2(P3_DATAO_REG_9__SCAN_IN), .ZN(n8474)
         );
  OAI22_X1 U8542 ( .A1(n15595), .A2(n10540), .B1(n15203), .B2(n10499), .ZN(
        n10269) );
  NAND2_X1 U8543 ( .A1(n13707), .A2(n13709), .ZN(n8759) );
  NAND2_X1 U8544 ( .A1(n11661), .A2(n9729), .ZN(n8471) );
  NAND2_X1 U8545 ( .A1(keyinput_90), .A2(P3_DATAO_REG_6__SCAN_IN), .ZN(n8470)
         );
  AOI21_X1 U8546 ( .B1(n9723), .B2(n9722), .A(n8473), .ZN(n8472) );
  INV_X1 U8547 ( .A(n13741), .ZN(n8764) );
  AOI21_X1 U8548 ( .B1(n8818), .B2(n8816), .A(n8815), .ZN(n8814) );
  INV_X1 U8549 ( .A(n10327), .ZN(n8815) );
  INV_X1 U8550 ( .A(n8820), .ZN(n8816) );
  NOR2_X1 U8551 ( .A1(n9740), .A2(n9739), .ZN(n9745) );
  AND2_X1 U8552 ( .A1(n13788), .A2(n8143), .ZN(n8142) );
  INV_X1 U8553 ( .A(n13787), .ZN(n8143) );
  OAI21_X1 U8554 ( .B1(n9576), .B2(n9575), .A(n8834), .ZN(n9579) );
  NAND2_X1 U8555 ( .A1(n9768), .A2(keyinput_246), .ZN(n8501) );
  NAND2_X1 U8556 ( .A1(n9586), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U8557 ( .A1(n9765), .A2(keyinput_114), .ZN(n8468) );
  INV_X1 U8558 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8851) );
  NOR2_X1 U8559 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8855) );
  NOR2_X1 U8560 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8854) );
  NOR2_X1 U8561 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n8853) );
  AOI21_X1 U8562 ( .B1(n7937), .B2(n7489), .A(n7934), .ZN(n10385) );
  OAI22_X1 U8563 ( .A1(n7936), .A2(n7941), .B1(n7943), .B2(n7935), .ZN(n7934)
         );
  INV_X1 U8564 ( .A(n10342), .ZN(n7937) );
  INV_X1 U8565 ( .A(n8795), .ZN(n8790) );
  NAND2_X1 U8566 ( .A1(n8797), .A2(n8796), .ZN(n8795) );
  NAND2_X1 U8567 ( .A1(n10525), .A2(n10526), .ZN(n8796) );
  INV_X1 U8568 ( .A(n10527), .ZN(n8797) );
  NAND2_X1 U8569 ( .A1(n8800), .A2(n8799), .ZN(n8798) );
  INV_X1 U8570 ( .A(n10503), .ZN(n8799) );
  INV_X1 U8571 ( .A(n10504), .ZN(n8800) );
  INV_X1 U8572 ( .A(n12293), .ZN(n7877) );
  NAND2_X1 U8573 ( .A1(n13787), .A2(n13789), .ZN(n8141) );
  NOR2_X1 U8574 ( .A1(n8686), .A2(n8683), .ZN(n8682) );
  INV_X1 U8575 ( .A(n8688), .ZN(n8683) );
  NAND2_X1 U8576 ( .A1(n8685), .A2(n8688), .ZN(n8684) );
  OAI21_X1 U8577 ( .B1(n8687), .B2(n8686), .A(n16015), .ZN(n8685) );
  NOR2_X1 U8578 ( .A1(n16633), .A2(n13637), .ZN(n8183) );
  AOI21_X1 U8579 ( .B1(n8634), .B2(n8636), .A(n10328), .ZN(n8632) );
  INV_X1 U8580 ( .A(n8634), .ZN(n8633) );
  INV_X1 U8581 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10638) );
  INV_X1 U8582 ( .A(n10312), .ZN(n10313) );
  OAI21_X1 U8583 ( .B1(n10674), .B2(n8115), .A(n8114), .ZN(n9923) );
  NAND2_X1 U8584 ( .A1(n10674), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8114) );
  OAI21_X1 U8585 ( .B1(n9895), .B2(n8868), .A(n8082), .ZN(n9896) );
  NAND2_X1 U8586 ( .A1(n9895), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8082) );
  INV_X1 U8587 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8906) );
  INV_X1 U8588 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8907) );
  INV_X1 U8589 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8909) );
  INV_X1 U8590 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8908) );
  AND2_X1 U8591 ( .A1(n8170), .A2(n7550), .ZN(n16318) );
  NAND2_X1 U8592 ( .A1(n8172), .A2(n8171), .ZN(n8170) );
  NOR2_X1 U8593 ( .A1(n16310), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n8171) );
  INV_X1 U8594 ( .A(n7858), .ZN(n16336) );
  OAI21_X1 U8595 ( .B1(n16324), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7534), .ZN(
        n7858) );
  INV_X1 U8596 ( .A(n7859), .ZN(n16323) );
  AOI21_X1 U8597 ( .B1(n8503), .B2(n8502), .A(n8499), .ZN(n8498) );
  NAND2_X1 U8598 ( .A1(n8501), .A2(n8500), .ZN(n8499) );
  NOR2_X1 U8599 ( .A1(n9583), .A2(n9582), .ZN(n8502) );
  NAND2_X1 U8600 ( .A1(n9585), .A2(n9584), .ZN(n8503) );
  OR2_X1 U8601 ( .A1(n9764), .A2(n8466), .ZN(n8465) );
  NAND2_X1 U8602 ( .A1(n8468), .A2(n8467), .ZN(n8466) );
  NAND2_X1 U8603 ( .A1(n9766), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8467) );
  INV_X1 U8604 ( .A(n9767), .ZN(n8464) );
  INV_X1 U8605 ( .A(keyinput_117), .ZN(n8462) );
  NAND2_X1 U8606 ( .A1(n9768), .A2(keyinput_118), .ZN(n8460) );
  NAND2_X1 U8607 ( .A1(n9769), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8459) );
  OR2_X1 U8608 ( .A1(n13941), .A2(n14720), .ZN(n13942) );
  NAND2_X1 U8609 ( .A1(n13942), .A2(n8601), .ZN(n8600) );
  INV_X1 U8610 ( .A(n13938), .ZN(n8601) );
  OAI211_X1 U8611 ( .C1(n14339), .C2(n14455), .A(n14444), .B(n8555), .ZN(
        n14450) );
  OR2_X1 U8612 ( .A1(n12154), .A2(n16534), .ZN(n12153) );
  NAND2_X1 U8613 ( .A1(n8012), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8011) );
  OR2_X1 U8614 ( .A1(n8336), .A2(n11309), .ZN(n7719) );
  AND2_X1 U8615 ( .A1(n14553), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U8616 ( .A1(n8574), .A2(n8572), .ZN(n14329) );
  NOR2_X1 U8617 ( .A1(n14661), .A2(n8573), .ZN(n8572) );
  INV_X1 U8618 ( .A(n8917), .ZN(n8573) );
  NAND2_X1 U8619 ( .A1(n14918), .A2(n14702), .ZN(n8345) );
  NOR2_X1 U8620 ( .A1(n7591), .A2(n7794), .ZN(n7793) );
  INV_X1 U8621 ( .A(n14340), .ZN(n7794) );
  OR2_X1 U8622 ( .A1(n14700), .A2(n7591), .ZN(n7796) );
  AND2_X1 U8623 ( .A1(n7806), .A2(n14353), .ZN(n7805) );
  OAI21_X1 U8624 ( .B1(n7813), .B2(n8250), .A(n8248), .ZN(n7806) );
  INV_X1 U8625 ( .A(n14822), .ZN(n7809) );
  NAND2_X1 U8626 ( .A1(n12807), .A2(n12806), .ZN(n8357) );
  NAND2_X1 U8627 ( .A1(n8348), .A2(n8346), .ZN(n12594) );
  AND2_X1 U8628 ( .A1(n8347), .A2(n8982), .ZN(n8346) );
  INV_X1 U8629 ( .A(n14473), .ZN(n8347) );
  NAND2_X1 U8630 ( .A1(n12556), .A2(n16530), .ZN(n14368) );
  NAND2_X1 U8631 ( .A1(n16498), .A2(n14145), .ZN(n14373) );
  AOI21_X1 U8632 ( .B1(n14663), .B2(n14664), .A(n7784), .ZN(n9370) );
  INV_X1 U8633 ( .A(n14326), .ZN(n7784) );
  NAND2_X1 U8634 ( .A1(n14655), .A2(n14661), .ZN(n14330) );
  NAND2_X1 U8635 ( .A1(n8365), .A2(n8361), .ZN(n14628) );
  AND2_X1 U8636 ( .A1(n14634), .A2(n8364), .ZN(n8361) );
  NAND2_X1 U8637 ( .A1(n14906), .A2(n14661), .ZN(n8364) );
  NAND2_X1 U8638 ( .A1(n9319), .A2(n8838), .ZN(n14644) );
  NAND2_X1 U8639 ( .A1(n8251), .A2(n7804), .ZN(n7803) );
  NOR2_X1 U8640 ( .A1(n7811), .A2(n7813), .ZN(n7804) );
  INV_X1 U8641 ( .A(n8248), .ZN(n7812) );
  NAND2_X1 U8642 ( .A1(n14777), .A2(n7783), .ZN(n12714) );
  INV_X1 U8643 ( .A(n8857), .ZN(n7798) );
  INV_X1 U8644 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U8645 ( .A1(n9415), .A2(n8592), .ZN(n12116) );
  AND2_X1 U8646 ( .A1(n8886), .A2(n8561), .ZN(n7762) );
  INV_X1 U8647 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8847) );
  INV_X1 U8648 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8846) );
  OAI21_X1 U8649 ( .B1(n8880), .B2(n8581), .A(n8579), .ZN(n8885) );
  INV_X1 U8650 ( .A(n8580), .ZN(n8579) );
  OAI21_X1 U8651 ( .B1(n8583), .B2(n8581), .A(n8883), .ZN(n8580) );
  INV_X1 U8652 ( .A(n9039), .ZN(n7767) );
  NOR2_X1 U8653 ( .A1(n15027), .A2(n8532), .ZN(n7689) );
  NAND2_X1 U8654 ( .A1(n9837), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9800) );
  INV_X1 U8655 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9857) );
  INV_X1 U8656 ( .A(n15348), .ZN(n8304) );
  NAND2_X1 U8657 ( .A1(n15207), .A2(n15209), .ZN(n8414) );
  INV_X1 U8658 ( .A(n7464), .ZN(n8405) );
  INV_X1 U8659 ( .A(n12978), .ZN(n8384) );
  INV_X1 U8660 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9789) );
  INV_X1 U8661 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9788) );
  XNOR2_X1 U8662 ( .A(n10550), .B(n10549), .ZN(n11456) );
  INV_X1 U8663 ( .A(n8743), .ZN(n8736) );
  NAND2_X1 U8664 ( .A1(n13587), .A2(n11015), .ZN(n13968) );
  NOR2_X1 U8665 ( .A1(n16069), .A2(n16074), .ZN(n8197) );
  NOR2_X1 U8666 ( .A1(n8701), .A2(n15846), .ZN(n8698) );
  AND2_X1 U8667 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n13743), .ZN(n13742) );
  INV_X1 U8668 ( .A(n15912), .ZN(n8711) );
  NOR2_X1 U8669 ( .A1(n16111), .A2(n15958), .ZN(n8190) );
  NOR2_X1 U8670 ( .A1(n11147), .A2(n11146), .ZN(n11145) );
  INV_X1 U8671 ( .A(n8071), .ZN(n8070) );
  AND2_X1 U8672 ( .A1(n8068), .A2(n8705), .ZN(n8067) );
  AOI21_X1 U8673 ( .B1(n8707), .B2(n8687), .A(n7478), .ZN(n8705) );
  NOR2_X1 U8674 ( .A1(n10974), .A2(n10962), .ZN(n10961) );
  NOR2_X1 U8675 ( .A1(n8131), .A2(n8038), .ZN(n8037) );
  INV_X1 U8676 ( .A(n8040), .ZN(n8038) );
  NOR2_X1 U8677 ( .A1(n16633), .A2(n13019), .ZN(n8131) );
  AND2_X1 U8678 ( .A1(n10940), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11062) );
  NOR2_X1 U8679 ( .A1(n8182), .A2(n13649), .ZN(n8181) );
  INV_X1 U8680 ( .A(n8183), .ZN(n8182) );
  INV_X1 U8681 ( .A(n16612), .ZN(n12881) );
  XNOR2_X1 U8682 ( .A(n15754), .B(n13611), .ZN(n13616) );
  XNOR2_X1 U8683 ( .A(n15755), .B(n13607), .ZN(n13856) );
  NAND2_X1 U8684 ( .A1(n15887), .A2(n15871), .ZN(n15870) );
  NAND2_X1 U8685 ( .A1(n8680), .A2(n15991), .ZN(n8024) );
  INV_X1 U8686 ( .A(n8684), .ZN(n8680) );
  NAND2_X1 U8687 ( .A1(n8679), .A2(n8684), .ZN(n15992) );
  NAND2_X1 U8688 ( .A1(n16025), .A2(n8682), .ZN(n8679) );
  NAND2_X1 U8689 ( .A1(n8146), .A2(n7480), .ZN(n14024) );
  NAND2_X1 U8690 ( .A1(n16571), .A2(n8183), .ZN(n16614) );
  NAND2_X1 U8691 ( .A1(n13580), .A2(n8180), .ZN(n11793) );
  INV_X1 U8692 ( .A(n11784), .ZN(n8180) );
  NAND3_X1 U8693 ( .A1(n10611), .A2(n10610), .A3(n10609), .ZN(n11103) );
  OAI21_X1 U8694 ( .B1(n10391), .B2(n13307), .A(n10392), .ZN(n10410) );
  NOR2_X1 U8695 ( .A1(n10353), .A2(n8654), .ZN(n8653) );
  INV_X1 U8696 ( .A(n10348), .ZN(n8654) );
  OR2_X1 U8697 ( .A1(n10251), .A2(SI_18_), .ZN(n10252) );
  AOI21_X1 U8698 ( .B1(n7826), .B2(n8206), .A(n7532), .ZN(n7824) );
  NAND2_X1 U8699 ( .A1(n10204), .A2(n11753), .ZN(n10205) );
  NOR2_X1 U8700 ( .A1(n8207), .A2(n7830), .ZN(n7829) );
  INV_X1 U8701 ( .A(n10138), .ZN(n7830) );
  NAND2_X1 U8702 ( .A1(n8090), .A2(n8089), .ZN(n10705) );
  INV_X1 U8703 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8089) );
  XNOR2_X1 U8704 ( .A(n16318), .B(n16317), .ZN(n16319) );
  XNOR2_X1 U8705 ( .A(n7859), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n16324) );
  XNOR2_X1 U8706 ( .A(n16336), .B(n16335), .ZN(n16337) );
  OAI21_X1 U8707 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n16390), .A(n16389), .ZN(
        n16394) );
  OAI21_X1 U8708 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n16429), .A(n16428), .ZN(
        n16433) );
  AOI21_X1 U8709 ( .B1(n8497), .B2(n8496), .A(n8495), .ZN(n9595) );
  XNOR2_X1 U8710 ( .A(n11100), .B(keyinput_249), .ZN(n8495) );
  INV_X1 U8711 ( .A(n9587), .ZN(n8496) );
  INV_X1 U8712 ( .A(n8498), .ZN(n8497) );
  AOI21_X1 U8713 ( .B1(n8463), .B2(n8461), .A(n8458), .ZN(n9774) );
  NAND2_X1 U8714 ( .A1(n8460), .A2(n8459), .ZN(n8458) );
  XNOR2_X1 U8715 ( .A(n10610), .B(n8462), .ZN(n8461) );
  NAND2_X1 U8716 ( .A1(n8465), .A2(n8464), .ZN(n8463) );
  NAND3_X1 U8717 ( .A1(n9412), .A2(n9411), .A3(n9410), .ZN(n12117) );
  NAND2_X1 U8718 ( .A1(n14264), .A2(n13940), .ZN(n14120) );
  INV_X1 U8719 ( .A(n13954), .ZN(n8615) );
  INV_X1 U8720 ( .A(n7733), .ZN(n7732) );
  OAI21_X1 U8721 ( .B1(n8603), .B2(n7734), .A(n13925), .ZN(n7733) );
  INV_X1 U8722 ( .A(n14203), .ZN(n7734) );
  NAND2_X1 U8723 ( .A1(n14120), .A2(n14119), .ZN(n14232) );
  NAND2_X1 U8724 ( .A1(n7783), .A2(n12674), .ZN(n14355) );
  AOI21_X1 U8725 ( .B1(n8625), .B2(n7738), .A(n7516), .ZN(n7737) );
  INV_X1 U8726 ( .A(n14275), .ZN(n7738) );
  INV_X1 U8727 ( .A(n13933), .ZN(n8624) );
  INV_X1 U8728 ( .A(n14154), .ZN(n8627) );
  NOR2_X1 U8729 ( .A1(n9221), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9233) );
  AND2_X1 U8730 ( .A1(n9233), .A2(n9232), .ZN(n9246) );
  OR2_X1 U8731 ( .A1(n13939), .A2(n13938), .ZN(n8602) );
  AOI21_X1 U8732 ( .B1(n13247), .B2(n8622), .A(n7440), .ZN(n7727) );
  INV_X1 U8733 ( .A(n13247), .ZN(n7728) );
  NAND2_X1 U8734 ( .A1(n12348), .A2(n12272), .ZN(n12273) );
  OR2_X1 U8735 ( .A1(n9206), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U8736 ( .A1(n14211), .A2(n14212), .ZN(n14210) );
  OR2_X1 U8737 ( .A1(n9001), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9016) );
  AND2_X1 U8738 ( .A1(n8242), .A2(n9785), .ZN(n8240) );
  NOR2_X1 U8739 ( .A1(n14322), .A2(n14605), .ZN(n8242) );
  NOR2_X1 U8740 ( .A1(n10844), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11998) );
  OR2_X1 U8741 ( .A1(n12172), .A2(n8925), .ZN(n12174) );
  NAND2_X1 U8742 ( .A1(n7909), .A2(n7908), .ZN(n11996) );
  NAND2_X1 U8743 ( .A1(n10915), .A2(n10844), .ZN(n7908) );
  OR2_X1 U8744 ( .A1(n10915), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7909) );
  INV_X1 U8745 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n16317) );
  OAI21_X1 U8746 ( .B1(n10878), .B2(P3_REG1_REG_2__SCAN_IN), .A(n8101), .ZN(
        n12008) );
  NAND2_X1 U8747 ( .A1(n10878), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U8748 ( .A1(n8329), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8328) );
  INV_X1 U8749 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n16335) );
  NAND2_X1 U8750 ( .A1(n8008), .A2(n12229), .ZN(n12233) );
  NAND2_X1 U8751 ( .A1(n8005), .A2(n12230), .ZN(n12252) );
  INV_X1 U8752 ( .A(n8006), .ZN(n8005) );
  NAND2_X1 U8753 ( .A1(n7707), .A2(n7705), .ZN(n12238) );
  NAND2_X1 U8754 ( .A1(n12241), .A2(n10890), .ZN(n10892) );
  NAND2_X1 U8755 ( .A1(n10892), .A2(n11289), .ZN(n10891) );
  NAND2_X1 U8756 ( .A1(n7717), .A2(n7719), .ZN(n12746) );
  AND2_X1 U8757 ( .A1(n7717), .A2(n7718), .ZN(n13060) );
  NOR2_X1 U8758 ( .A1(n13067), .A2(n7921), .ZN(n7917) );
  NAND2_X1 U8759 ( .A1(n7997), .A2(n10839), .ZN(n8270) );
  NAND2_X1 U8760 ( .A1(n8270), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8269) );
  NOR2_X1 U8761 ( .A1(n14521), .A2(n10899), .ZN(n14536) );
  INV_X1 U8762 ( .A(n10897), .ZN(n10899) );
  INV_X1 U8763 ( .A(n8323), .ZN(n8325) );
  NAND2_X1 U8764 ( .A1(n7723), .A2(n7722), .ZN(n7721) );
  INV_X1 U8765 ( .A(n14555), .ZN(n7722) );
  INV_X1 U8766 ( .A(n7723), .ZN(n14554) );
  NOR2_X1 U8767 ( .A1(n14579), .A2(n14551), .ZN(n8003) );
  NOR2_X1 U8768 ( .A1(n14579), .A2(n8004), .ZN(n8002) );
  INV_X1 U8769 ( .A(n8265), .ZN(n8004) );
  OR2_X1 U8770 ( .A1(n10926), .A2(n14794), .ZN(n8335) );
  INV_X1 U8771 ( .A(n7893), .ZN(n14593) );
  OR2_X1 U8772 ( .A1(n8919), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n14615) );
  OR2_X1 U8773 ( .A1(n9078), .A2(n14964), .ZN(n8917) );
  OR3_X1 U8774 ( .A1(n9309), .A2(P3_REG3_REG_26__SCAN_IN), .A3(
        P3_REG3_REG_25__SCAN_IN), .ZN(n9310) );
  AND2_X1 U8775 ( .A1(n14326), .A2(n14324), .ZN(n14664) );
  NAND2_X1 U8776 ( .A1(n9282), .A2(n9281), .ZN(n14688) );
  INV_X1 U8777 ( .A(n7795), .ZN(n14686) );
  AOI21_X1 U8778 ( .B1(n14706), .B2(n14700), .A(n7591), .ZN(n7795) );
  NAND2_X1 U8779 ( .A1(n14713), .A2(n14340), .ZN(n14706) );
  OR2_X1 U8780 ( .A1(n9261), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9275) );
  OR2_X1 U8781 ( .A1(n9275), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9283) );
  AND2_X1 U8782 ( .A1(n14776), .A2(n9193), .ZN(n8360) );
  AOI21_X1 U8783 ( .B1(n8233), .B2(n7789), .A(n7788), .ZN(n7787) );
  INV_X1 U8784 ( .A(n14426), .ZN(n7789) );
  AOI21_X1 U8785 ( .B1(n8371), .B2(n8370), .A(n7613), .ZN(n8369) );
  NAND2_X1 U8786 ( .A1(n9192), .A2(n8237), .ZN(n14789) );
  INV_X1 U8787 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9662) );
  OR2_X1 U8788 ( .A1(n9140), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9156) );
  OR2_X1 U8789 ( .A1(n9087), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9103) );
  NOR2_X1 U8790 ( .A1(n9103), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9127) );
  OR2_X1 U8791 ( .A1(n9069), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U8792 ( .A1(n8357), .A2(n9030), .ZN(n12962) );
  AND2_X1 U8793 ( .A1(n14383), .A2(n14382), .ZN(n14474) );
  NAND2_X1 U8794 ( .A1(n8348), .A2(n8982), .ZN(n12596) );
  OAI21_X1 U8795 ( .B1(n16490), .B2(n16494), .A(n9357), .ZN(n14360) );
  NAND2_X1 U8796 ( .A1(n14360), .A2(n14468), .ZN(n12774) );
  NAND2_X1 U8797 ( .A1(n9102), .A2(n9101), .ZN(n14814) );
  INV_X1 U8798 ( .A(n16503), .ZN(n16678) );
  NAND2_X1 U8799 ( .A1(n9390), .A2(n9411), .ZN(n8597) );
  AND2_X1 U8800 ( .A1(n12116), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11545) );
  OAI21_X1 U8801 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n15620), .A(n8899), .ZN(
        n9320) );
  NAND2_X1 U8802 ( .A1(n8127), .A2(n8125), .ZN(n8916) );
  NAND2_X1 U8803 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n8126), .ZN(n8125) );
  NAND2_X1 U8804 ( .A1(n9306), .A2(n9304), .ZN(n8127) );
  NOR2_X1 U8805 ( .A1(n9413), .A2(P3_IR_REG_23__SCAN_IN), .ZN(n8593) );
  INV_X1 U8806 ( .A(n7779), .ZN(n9290) );
  OAI21_X1 U8807 ( .B1(n9271), .B2(n9272), .A(n8575), .ZN(n7779) );
  NAND2_X1 U8808 ( .A1(n13339), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8575) );
  NOR2_X1 U8809 ( .A1(n7901), .A2(n8368), .ZN(n9343) );
  NAND2_X1 U8810 ( .A1(n7435), .A2(n8366), .ZN(n7901) );
  NAND2_X1 U8811 ( .A1(n7763), .A2(n8896), .ZN(n9243) );
  NAND2_X1 U8812 ( .A1(n9229), .A2(n13167), .ZN(n7763) );
  NAND2_X1 U8813 ( .A1(n8894), .A2(n8553), .ZN(n9214) );
  NAND2_X1 U8814 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n8554), .ZN(n8553) );
  NAND2_X1 U8815 ( .A1(n8081), .A2(n9198), .ZN(n9200) );
  INV_X1 U8816 ( .A(n9197), .ZN(n8081) );
  NOR2_X1 U8817 ( .A1(n8368), .A2(n7459), .ZN(n9118) );
  INV_X1 U8818 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9119) );
  OR2_X1 U8819 ( .A1(n9080), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9109) );
  INV_X1 U8820 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7757) );
  XNOR2_X1 U8821 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .ZN(n8991) );
  XNOR2_X1 U8822 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .ZN(n8975) );
  NAND2_X1 U8823 ( .A1(n7760), .A2(n8569), .ZN(n8977) );
  AOI21_X1 U8824 ( .B1(n8570), .B2(n8960), .A(n7537), .ZN(n8569) );
  AND2_X1 U8825 ( .A1(n9868), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8931) );
  NOR2_X1 U8826 ( .A1(n12207), .A2(n8538), .ZN(n8537) );
  XNOR2_X1 U8827 ( .A(n14066), .B(n11672), .ZN(n11664) );
  AND2_X1 U8828 ( .A1(n15443), .A2(n11662), .ZN(n11672) );
  INV_X1 U8829 ( .A(n14993), .ZN(n7672) );
  OR2_X1 U8830 ( .A1(n10359), .A2(n10358), .ZN(n10375) );
  AND2_X1 U8831 ( .A1(n14096), .A2(n7596), .ZN(n8084) );
  NAND2_X1 U8832 ( .A1(n8523), .A2(n8522), .ZN(n8521) );
  INV_X1 U8833 ( .A(n11809), .ZN(n8522) );
  OR2_X1 U8834 ( .A1(n12581), .A2(n12580), .ZN(n8531) );
  NAND2_X1 U8835 ( .A1(n12581), .A2(n12580), .ZN(n8530) );
  OR2_X1 U8836 ( .A1(n10106), .A2(n10105), .ZN(n10128) );
  NAND3_X1 U8837 ( .A1(n8525), .A2(n8524), .A3(n7502), .ZN(n7680) );
  NAND2_X1 U8838 ( .A1(n7679), .A2(n7467), .ZN(n7678) );
  INV_X1 U8839 ( .A(n13035), .ZN(n7679) );
  OR2_X1 U8840 ( .A1(n10261), .A2(n15127), .ZN(n10280) );
  NAND2_X1 U8841 ( .A1(n10190), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10233) );
  INV_X1 U8842 ( .A(n8536), .ZN(n8534) );
  NAND2_X1 U8843 ( .A1(n13177), .A2(n13294), .ZN(n8535) );
  NAND2_X1 U8844 ( .A1(n13117), .A2(n11248), .ZN(n11662) );
  NAND2_X1 U8845 ( .A1(n10506), .A2(n7447), .ZN(n8791) );
  NOR2_X1 U8846 ( .A1(n8793), .A2(n10533), .ZN(n8792) );
  NAND2_X1 U8847 ( .A1(n10506), .A2(n7871), .ZN(n7870) );
  NAND2_X1 U8848 ( .A1(n9812), .A2(n9806), .ZN(n9807) );
  XNOR2_X1 U8849 ( .A(n15552), .B(n10524), .ZN(n10571) );
  AND2_X1 U8850 ( .A1(n10308), .A2(n10307), .ZN(n15183) );
  AND4_X1 U8851 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        n12921) );
  AND4_X1 U8852 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n12621) );
  AND4_X1 U8853 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n11969)
         );
  NOR2_X1 U8854 ( .A1(n7739), .A2(n7472), .ZN(n11466) );
  NOR2_X1 U8855 ( .A1(n11494), .A2(n7505), .ZN(n11511) );
  OR2_X1 U8856 ( .A1(n11511), .A2(n11510), .ZN(n7745) );
  NOR2_X1 U8857 ( .A1(n11498), .A2(n11497), .ZN(n11546) );
  OR2_X1 U8858 ( .A1(n11739), .A2(n11738), .ZN(n7753) );
  NOR2_X1 U8859 ( .A1(n16263), .A2(n7751), .ZN(n12539) );
  AND2_X1 U8860 ( .A1(n16269), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7751) );
  OR2_X1 U8861 ( .A1(n12539), .A2(n12538), .ZN(n7750) );
  AND2_X1 U8862 ( .A1(n7750), .A2(n7749), .ZN(n12655) );
  NAND2_X1 U8863 ( .A1(n12654), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U8864 ( .A1(n12655), .A2(n12656), .ZN(n12945) );
  NOR2_X1 U8865 ( .A1(n16238), .A2(n7748), .ZN(n16252) );
  AND2_X1 U8866 ( .A1(n16243), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7748) );
  OR2_X1 U8867 ( .A1(n16252), .A2(n16251), .ZN(n7747) );
  AND2_X1 U8868 ( .A1(n7747), .A2(n7746), .ZN(n15136) );
  NAND2_X1 U8869 ( .A1(n16255), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7746) );
  NOR2_X1 U8870 ( .A1(n15136), .A2(n15135), .ZN(n15141) );
  AND2_X1 U8871 ( .A1(n11682), .A2(n11463), .ZN(n15225) );
  NAND2_X1 U8872 ( .A1(n15372), .A2(n7444), .ZN(n15312) );
  NAND2_X1 U8873 ( .A1(n15372), .A2(n8226), .ZN(n15340) );
  NAND2_X1 U8874 ( .A1(n15372), .A2(n15360), .ZN(n15355) );
  NAND2_X1 U8875 ( .A1(n7883), .A2(n15206), .ZN(n15392) );
  NAND2_X1 U8876 ( .A1(n8408), .A2(n15201), .ZN(n15419) );
  INV_X1 U8877 ( .A(n15201), .ZN(n8407) );
  NAND2_X1 U8878 ( .A1(n8409), .A2(n7464), .ZN(n8408) );
  INV_X1 U8879 ( .A(n15438), .ZN(n8409) );
  NAND2_X1 U8880 ( .A1(n15448), .A2(n15457), .ZN(n15449) );
  NAND2_X1 U8881 ( .A1(n7872), .A2(n13349), .ZN(n15195) );
  NAND2_X1 U8882 ( .A1(n13343), .A2(n13342), .ZN(n13344) );
  AND2_X1 U8883 ( .A1(n13234), .A2(n13348), .ZN(n13358) );
  INV_X1 U8884 ( .A(n13232), .ZN(n13340) );
  NAND2_X1 U8885 ( .A1(n12635), .A2(n7886), .ZN(n7888) );
  NOR2_X1 U8886 ( .A1(n8383), .A2(n7887), .ZN(n7886) );
  INV_X1 U8887 ( .A(n12618), .ZN(n7887) );
  NAND2_X1 U8888 ( .A1(n12643), .A2(n12917), .ZN(n12926) );
  AND2_X1 U8889 ( .A1(n12789), .A2(n12641), .ZN(n12643) );
  NAND2_X1 U8890 ( .A1(n12613), .A2(n12612), .ZN(n12634) );
  XNOR2_X1 U8891 ( .A(n12792), .B(n12621), .ZN(n12638) );
  NAND2_X1 U8892 ( .A1(n8301), .A2(n12295), .ZN(n8300) );
  NOR2_X1 U8893 ( .A1(n12293), .A2(n8299), .ZN(n8298) );
  INV_X1 U8894 ( .A(n11952), .ZN(n8299) );
  NAND2_X1 U8895 ( .A1(n7666), .A2(n8301), .ZN(n12303) );
  INV_X1 U8896 ( .A(n11961), .ZN(n7666) );
  NAND2_X1 U8897 ( .A1(n11937), .A2(n11968), .ZN(n11961) );
  NAND2_X1 U8898 ( .A1(n11716), .A2(n11225), .ZN(n11722) );
  NAND2_X1 U8899 ( .A1(n13117), .A2(n10515), .ZN(n10516) );
  INV_X1 U8900 ( .A(n11250), .ZN(n11918) );
  NAND2_X1 U8901 ( .A1(n15381), .A2(n15182), .ZN(n15376) );
  NAND2_X1 U8902 ( .A1(n10214), .A2(n10213), .ZN(n15539) );
  AND2_X1 U8903 ( .A1(n11224), .A2(n11735), .ZN(n12204) );
  AND2_X1 U8904 ( .A1(n10608), .A2(n11456), .ZN(n11692) );
  INV_X1 U8905 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10560) );
  OAI21_X1 U8906 ( .B1(n10556), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10565) );
  INV_X1 U8907 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10564) );
  INV_X1 U8908 ( .A(n11456), .ZN(n10607) );
  NAND2_X1 U8909 ( .A1(n9814), .A2(n9813), .ZN(n10548) );
  OR3_X1 U8910 ( .A1(n10079), .A2(P2_IR_REG_9__SCAN_IN), .A3(n10078), .ZN(
        n10081) );
  OR2_X1 U8911 ( .A1(n9927), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9929) );
  INV_X1 U8912 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U8913 ( .A1(n8121), .A2(n8120), .ZN(n8119) );
  INV_X1 U8914 ( .A(n11097), .ZN(n8120) );
  INV_X1 U8915 ( .A(n11096), .ZN(n8121) );
  NAND2_X1 U8916 ( .A1(n7995), .A2(n7994), .ZN(n7993) );
  INV_X1 U8917 ( .A(n11057), .ZN(n7994) );
  NAND2_X1 U8918 ( .A1(n8123), .A2(n8122), .ZN(n11866) );
  INV_X1 U8919 ( .A(n11869), .ZN(n8122) );
  AOI21_X1 U8920 ( .B1(n7977), .B2(n7980), .A(n7514), .ZN(n7975) );
  INV_X1 U8921 ( .A(n8717), .ZN(n7980) );
  NOR2_X1 U8922 ( .A1(n15655), .A2(n8744), .ZN(n8743) );
  INV_X1 U8923 ( .A(n15714), .ZN(n8744) );
  INV_X1 U8924 ( .A(n8742), .ZN(n8741) );
  OAI21_X1 U8925 ( .B1(n15655), .B2(n8747), .A(n8746), .ZN(n8742) );
  NAND2_X1 U8926 ( .A1(n15704), .A2(n15705), .ZN(n15703) );
  INV_X1 U8927 ( .A(n13217), .ZN(n8734) );
  NAND2_X1 U8928 ( .A1(n11098), .A2(n11099), .ZN(n8730) );
  INV_X1 U8929 ( .A(n13967), .ZN(n14012) );
  OR2_X1 U8930 ( .A1(n7432), .A2(n7477), .ZN(n8055) );
  NAND2_X1 U8931 ( .A1(n16054), .A2(n15733), .ZN(n8056) );
  NOR2_X1 U8932 ( .A1(n16062), .A2(n15734), .ZN(n8128) );
  AND4_X1 U8933 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n15827) );
  AOI21_X1 U8934 ( .B1(n8676), .B2(n8678), .A(n7504), .ZN(n8674) );
  NAND2_X1 U8935 ( .A1(n15887), .A2(n8197), .ZN(n15858) );
  INV_X1 U8936 ( .A(n13733), .ZN(n13743) );
  AND2_X1 U8937 ( .A1(n15904), .A2(n15889), .ZN(n15887) );
  NOR2_X1 U8938 ( .A1(n15919), .A2(n16088), .ZN(n15904) );
  NAND2_X1 U8939 ( .A1(n15998), .A2(n8189), .ZN(n15919) );
  AND2_X1 U8940 ( .A1(n15921), .A2(n7473), .ZN(n8189) );
  AOI21_X1 U8941 ( .B1(n15934), .B2(n8046), .A(n8148), .ZN(n8045) );
  INV_X1 U8942 ( .A(n8689), .ZN(n8046) );
  NOR2_X1 U8943 ( .A1(n15937), .A2(n8149), .ZN(n8148) );
  NAND2_X1 U8944 ( .A1(n15998), .A2(n8190), .ZN(n15952) );
  NAND2_X1 U8945 ( .A1(n15998), .A2(n15985), .ZN(n15983) );
  NAND2_X1 U8946 ( .A1(n13422), .A2(n7445), .ZN(n16007) );
  OR2_X1 U8947 ( .A1(n11129), .A2(n11128), .ZN(n11147) );
  OR2_X1 U8948 ( .A1(n10988), .A2(n10972), .ZN(n10974) );
  INV_X1 U8949 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U8950 ( .A1(n13422), .A2(n13425), .ZN(n13508) );
  NOR2_X1 U8951 ( .A1(n13203), .A2(n16697), .ZN(n13422) );
  INV_X1 U8952 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10986) );
  OR2_X1 U8953 ( .A1(n11085), .A2(n10986), .ZN(n10988) );
  NAND2_X1 U8954 ( .A1(n13138), .A2(n13137), .ZN(n13198) );
  INV_X1 U8955 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U8956 ( .A1(n16571), .A2(n8041), .ZN(n16613) );
  NOR2_X1 U8957 ( .A1(n12342), .A2(n13633), .ZN(n16571) );
  INV_X1 U8958 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10760) );
  OR2_X1 U8959 ( .A1(n10761), .A2(n10760), .ZN(n10788) );
  NAND2_X1 U8960 ( .A1(n8656), .A2(n11775), .ZN(n8655) );
  NOR2_X1 U8961 ( .A1(n11793), .A2(n13607), .ZN(n12448) );
  INV_X1 U8962 ( .A(n13616), .ZN(n13857) );
  INV_X1 U8963 ( .A(n13856), .ZN(n11797) );
  NAND2_X1 U8964 ( .A1(n11762), .A2(n16474), .ZN(n11784) );
  NAND2_X1 U8965 ( .A1(n8664), .A2(n8668), .ZN(n15874) );
  NAND2_X1 U8966 ( .A1(n15901), .A2(n8670), .ZN(n8664) );
  NAND2_X1 U8967 ( .A1(n7616), .A2(n8021), .ZN(n15973) );
  NAND2_X1 U8968 ( .A1(n8708), .A2(n8707), .ZN(n16016) );
  NAND2_X1 U8969 ( .A1(n12481), .A2(n10776), .ZN(n12337) );
  XNOR2_X1 U8970 ( .A(n8646), .B(n10481), .ZN(n15603) );
  OAI21_X1 U8971 ( .B1(n10472), .B2(n7854), .A(n7851), .ZN(n8646) );
  AND2_X1 U8972 ( .A1(n10510), .A2(n10509), .ZN(n13919) );
  NAND2_X1 U8973 ( .A1(n7857), .A2(n7855), .ZN(n10510) );
  NAND2_X1 U8974 ( .A1(n7857), .A2(n10475), .ZN(n10508) );
  NOR2_X1 U8975 ( .A1(n10431), .A2(n7838), .ZN(n7837) );
  INV_X1 U8976 ( .A(n10414), .ZN(n7838) );
  AND2_X1 U8977 ( .A1(n10624), .A2(n10651), .ZN(n10810) );
  MUX2_X1 U8978 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10622), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10624) );
  NAND2_X1 U8979 ( .A1(n7959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10622) );
  INV_X1 U8980 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10629) );
  NAND2_X1 U8981 ( .A1(n8033), .A2(n8032), .ZN(n10639) );
  XNOR2_X1 U8982 ( .A(n10636), .B(P1_IR_REG_23__SCAN_IN), .ZN(n11304) );
  NAND2_X1 U8983 ( .A1(n8631), .A2(n8634), .ZN(n10329) );
  NAND2_X1 U8984 ( .A1(n10297), .A2(n8635), .ZN(n8631) );
  OAI21_X1 U8985 ( .B1(n10297), .B2(n10296), .A(n7428), .ZN(n10314) );
  OR2_X1 U8986 ( .A1(n11139), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n11158) );
  OR2_X1 U8987 ( .A1(n10204), .A2(n11753), .ZN(n10226) );
  NAND2_X1 U8988 ( .A1(n10163), .A2(n10162), .ZN(n10183) );
  NAND2_X1 U8989 ( .A1(n9990), .A2(n9989), .ZN(n9995) );
  AND2_X1 U8990 ( .A1(n10012), .A2(n9993), .ZN(n9994) );
  AND2_X1 U8991 ( .A1(n9989), .A2(n9970), .ZN(n9971) );
  AND2_X1 U8992 ( .A1(n9966), .A2(n7443), .ZN(n9941) );
  AND2_X1 U8993 ( .A1(n9938), .A2(n9926), .ZN(n11312) );
  NAND2_X1 U8994 ( .A1(n9818), .A2(n11271), .ZN(n9820) );
  AND3_X1 U8995 ( .A1(n8376), .A2(SI_0_), .A3(n8374), .ZN(n9845) );
  NAND2_X1 U8996 ( .A1(n9895), .A2(n8375), .ZN(n8374) );
  OR2_X1 U8997 ( .A1(n9895), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8376) );
  XNOR2_X1 U8998 ( .A(n16337), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n16330) );
  NOR2_X1 U8999 ( .A1(n16345), .A2(n16344), .ZN(n16351) );
  NAND2_X1 U9000 ( .A1(n8167), .A2(n8168), .ZN(n16391) );
  NAND2_X1 U9001 ( .A1(n16383), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8168) );
  OR2_X1 U9002 ( .A1(n16383), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8169) );
  OR2_X1 U9003 ( .A1(n16451), .A2(n16450), .ZN(n16457) );
  NAND2_X1 U9004 ( .A1(n14251), .A2(n13530), .ZN(n13532) );
  NAND2_X1 U9005 ( .A1(n13532), .A2(n13531), .ZN(n13551) );
  NAND2_X1 U9006 ( .A1(n9274), .A2(n9273), .ZN(n14323) );
  NAND2_X1 U9007 ( .A1(n14128), .A2(n13247), .ZN(n14129) );
  NAND2_X1 U9008 ( .A1(n14274), .A2(n13931), .ZN(n14153) );
  NAND2_X1 U9009 ( .A1(n12906), .A2(n12905), .ZN(n13087) );
  INV_X1 U9010 ( .A(n14674), .ZN(n14646) );
  AOI21_X1 U9011 ( .B1(n14236), .B2(n14195), .A(n14194), .ZN(n14197) );
  NAND2_X1 U9012 ( .A1(n8605), .A2(n8603), .ZN(n14204) );
  NAND2_X1 U9013 ( .A1(n14204), .A2(n14203), .ZN(n14202) );
  OAI21_X1 U9014 ( .B1(n8605), .B2(n7734), .A(n7732), .ZN(n14226) );
  NAND2_X1 U9015 ( .A1(n8623), .A2(n13089), .ZN(n13092) );
  NAND2_X1 U9016 ( .A1(n14151), .A2(n13933), .ZN(n14244) );
  NAND2_X1 U9017 ( .A1(n8602), .A2(n13940), .ZN(n14266) );
  OAI21_X1 U9018 ( .B1(n8623), .B2(n7728), .A(n7727), .ZN(n13309) );
  INV_X1 U9019 ( .A(n12556), .ZN(n16498) );
  NAND2_X1 U9020 ( .A1(n14224), .A2(n13928), .ZN(n14276) );
  NAND2_X1 U9021 ( .A1(n14276), .A2(n14275), .ZN(n14274) );
  NAND2_X1 U9022 ( .A1(n14210), .A2(n12798), .ZN(n12939) );
  NAND2_X1 U9023 ( .A1(n9308), .A2(n9307), .ZN(n14293) );
  OR2_X1 U9024 ( .A1(n9078), .A2(n14969), .ZN(n9307) );
  NAND2_X1 U9025 ( .A1(n13551), .A2(n13550), .ZN(n13921) );
  NAND2_X1 U9026 ( .A1(n8239), .A2(n8246), .ZN(n8096) );
  OR2_X1 U9027 ( .A1(n14514), .A2(n14513), .ZN(n8246) );
  NAND2_X1 U9028 ( .A1(n8245), .A2(n14500), .ZN(n8244) );
  NAND2_X1 U9029 ( .A1(n9303), .A2(n9302), .ZN(n14325) );
  NOR2_X1 U9030 ( .A1(n10879), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n12002) );
  AOI21_X1 U9031 ( .B1(n12017), .B2(n12016), .A(n7907), .ZN(n12151) );
  AND2_X1 U9032 ( .A1(n10823), .A2(n10878), .ZN(n7907) );
  NAND2_X1 U9033 ( .A1(n8327), .A2(n12405), .ZN(n12407) );
  INV_X1 U9034 ( .A(n8328), .ZN(n8327) );
  NAND2_X1 U9035 ( .A1(n8329), .A2(n12405), .ZN(n12157) );
  NAND2_X1 U9036 ( .A1(n8964), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8965) );
  OR2_X1 U9037 ( .A1(n12185), .A2(n8986), .ZN(n12386) );
  NAND2_X1 U9038 ( .A1(n8012), .A2(n12375), .ZN(n12182) );
  NAND2_X1 U9039 ( .A1(n7706), .A2(n7708), .ZN(n12251) );
  OAI22_X1 U9040 ( .A1(n12247), .A2(n12248), .B1(n10830), .B2(n7705), .ZN(
        n12226) );
  NAND2_X1 U9041 ( .A1(n8014), .A2(n8015), .ZN(n12510) );
  INV_X1 U9042 ( .A(n7699), .ZN(n12505) );
  INV_X1 U9043 ( .A(n10861), .ZN(n13055) );
  NAND2_X1 U9044 ( .A1(n7918), .A2(n7920), .ZN(n13066) );
  AOI21_X1 U9045 ( .B1(n7914), .B2(n7593), .A(n7913), .ZN(n7912) );
  INV_X1 U9046 ( .A(n14517), .ZN(n7913) );
  NAND2_X1 U9047 ( .A1(n7911), .A2(n7914), .ZN(n14518) );
  OR2_X1 U9048 ( .A1(n12744), .A2(n7593), .ZN(n7911) );
  NAND2_X1 U9049 ( .A1(n7711), .A2(n10897), .ZN(n14523) );
  AND2_X1 U9050 ( .A1(n8268), .A2(n8269), .ZN(n14534) );
  NOR2_X1 U9051 ( .A1(n14543), .A2(n14544), .ZN(n14542) );
  NAND3_X1 U9052 ( .A1(n7999), .A2(n7998), .A3(n8000), .ZN(n14569) );
  NOR2_X1 U9053 ( .A1(n8002), .A2(n8001), .ZN(n8000) );
  INV_X1 U9054 ( .A(n7897), .ZN(n14576) );
  OR2_X1 U9055 ( .A1(n10933), .A2(n10932), .ZN(n14588) );
  OAI21_X1 U9056 ( .B1(n7715), .B2(n14599), .A(n14603), .ZN(n7714) );
  NOR2_X1 U9057 ( .A1(n8331), .A2(n7716), .ZN(n7715) );
  OR2_X1 U9058 ( .A1(n10925), .A2(n8334), .ZN(n7716) );
  INV_X1 U9059 ( .A(n7713), .ZN(n7712) );
  OAI21_X1 U9060 ( .B1(n10927), .B2(n14574), .A(n7635), .ZN(n7713) );
  AND2_X1 U9061 ( .A1(n14308), .A2(n14307), .ZN(n14617) );
  NAND2_X1 U9062 ( .A1(n8341), .A2(n8339), .ZN(n14672) );
  NAND2_X1 U9063 ( .A1(n14736), .A2(n14438), .ZN(n14711) );
  NAND2_X1 U9064 ( .A1(n9260), .A2(n9259), .ZN(n14854) );
  NAND2_X1 U9065 ( .A1(n7802), .A2(n7461), .ZN(n14748) );
  AND2_X1 U9066 ( .A1(n7802), .A2(n14466), .ZN(n14749) );
  OR2_X1 U9067 ( .A1(n14764), .A2(n14342), .ZN(n7802) );
  NAND2_X1 U9068 ( .A1(n9205), .A2(n9204), .ZN(n14873) );
  NAND2_X1 U9069 ( .A1(n8238), .A2(n14343), .ZN(n14798) );
  NAND2_X1 U9070 ( .A1(n14801), .A2(n14803), .ZN(n8238) );
  NAND2_X1 U9071 ( .A1(n9185), .A2(n9184), .ZN(n14796) );
  NAND2_X1 U9072 ( .A1(n13540), .A2(n9163), .ZN(n14802) );
  NAND2_X1 U9073 ( .A1(n8351), .A2(n8354), .ZN(n13447) );
  NAND2_X1 U9074 ( .A1(n8247), .A2(n8251), .ZN(n13370) );
  NAND2_X1 U9075 ( .A1(n13210), .A2(n8253), .ZN(n8247) );
  NOR2_X2 U9076 ( .A1(n12673), .A2(n12672), .ZN(n14821) );
  NAND2_X1 U9077 ( .A1(n8255), .A2(n13208), .ZN(n13260) );
  NAND2_X1 U9078 ( .A1(n8257), .A2(n8256), .ZN(n8255) );
  INV_X2 U9079 ( .A(n14819), .ZN(n16517) );
  NAND2_X1 U9080 ( .A1(n12136), .A2(n12135), .ZN(n14792) );
  INV_X1 U9081 ( .A(n14821), .ZN(n14809) );
  INV_X1 U9082 ( .A(n14617), .ZN(n16735) );
  OAI21_X1 U9083 ( .B1(n14956), .B2(n14312), .A(n14311), .ZN(n16726) );
  INV_X1 U9084 ( .A(n14638), .ZN(n14902) );
  AOI21_X1 U9085 ( .B1(n7819), .B2(n7816), .A(n14829), .ZN(n14899) );
  NOR2_X1 U9086 ( .A1(n14637), .A2(n14894), .ZN(n7816) );
  AND2_X1 U9087 ( .A1(n14833), .A2(n16643), .ZN(n8106) );
  INV_X1 U9088 ( .A(n14655), .ZN(n14906) );
  INV_X1 U9089 ( .A(n14293), .ZN(n14910) );
  INV_X1 U9090 ( .A(n14681), .ZN(n14914) );
  INV_X1 U9091 ( .A(n14323), .ZN(n14922) );
  INV_X1 U9092 ( .A(n14191), .ZN(n14930) );
  AND2_X1 U9093 ( .A1(n9231), .A2(n9230), .ZN(n14934) );
  OR2_X1 U9094 ( .A1(n9078), .A2(n12466), .ZN(n9230) );
  INV_X1 U9095 ( .A(n14160), .ZN(n14939) );
  AND3_X1 U9096 ( .A1(n9065), .A2(n9064), .A3(n9063), .ZN(n13213) );
  INV_X1 U9097 ( .A(n12078), .ZN(n12674) );
  NAND2_X1 U9098 ( .A1(n16727), .A2(n16672), .ZN(n14938) );
  AND2_X2 U9099 ( .A1(n9416), .A2(n12135), .ZN(n16727) );
  AND2_X1 U9100 ( .A1(n9392), .A2(n9391), .ZN(n14946) );
  INV_X1 U9101 ( .A(n11545), .ZN(n14947) );
  INV_X1 U9102 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8373) );
  INV_X1 U9103 ( .A(SI_29_), .ZN(n14960) );
  INV_X1 U9104 ( .A(n8861), .ZN(n14962) );
  INV_X1 U9105 ( .A(SI_28_), .ZN(n13916) );
  INV_X1 U9106 ( .A(SI_27_), .ZN(n14964) );
  INV_X1 U9107 ( .A(SI_25_), .ZN(n13303) );
  XNOR2_X1 U9108 ( .A(n9380), .B(n9379), .ZN(n13304) );
  OAI21_X1 U9109 ( .B1(n8592), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9380) );
  INV_X1 U9110 ( .A(n7776), .ZN(n9295) );
  INV_X1 U9111 ( .A(n14357), .ZN(n12563) );
  XNOR2_X1 U9112 ( .A(n9339), .B(n9338), .ZN(n12468) );
  INV_X1 U9113 ( .A(SI_18_), .ZN(n11896) );
  NAND2_X1 U9114 ( .A1(n8559), .A2(n8561), .ZN(n9164) );
  NAND2_X1 U9115 ( .A1(n8094), .A2(n8564), .ZN(n8559) );
  INV_X1 U9116 ( .A(SI_15_), .ZN(n11603) );
  NAND2_X1 U9117 ( .A1(n8566), .A2(n8889), .ZN(n9150) );
  NAND2_X1 U9118 ( .A1(n8567), .A2(n7627), .ZN(n8566) );
  INV_X1 U9119 ( .A(SI_14_), .ZN(n11532) );
  INV_X1 U9120 ( .A(SI_13_), .ZN(n11452) );
  NAND2_X1 U9121 ( .A1(n8578), .A2(n8882), .ZN(n9113) );
  NAND2_X1 U9122 ( .A1(n8880), .A2(n8583), .ZN(n8578) );
  INV_X1 U9123 ( .A(SI_11_), .ZN(n11307) );
  NAND2_X1 U9124 ( .A1(n8880), .A2(n8879), .ZN(n9096) );
  INV_X1 U9125 ( .A(SI_10_), .ZN(n11296) );
  NAND2_X1 U9126 ( .A1(n7768), .A2(n7769), .ZN(n9040) );
  OR2_X1 U9127 ( .A1(n9009), .A2(n7771), .ZN(n7768) );
  NAND2_X1 U9128 ( .A1(n7772), .A2(n8875), .ZN(n9024) );
  OR2_X1 U9129 ( .A1(n9009), .A2(n8874), .ZN(n7772) );
  INV_X1 U9130 ( .A(SI_6_), .ZN(n11267) );
  XNOR2_X1 U9131 ( .A(n8978), .B(P3_IR_REG_4__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U9132 ( .A1(n8571), .A2(n8867), .ZN(n8962) );
  XNOR2_X1 U9133 ( .A(n8933), .B(n8934), .ZN(n12166) );
  NAND2_X1 U9134 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8933) );
  NOR2_X1 U9135 ( .A1(n10608), .A2(n10607), .ZN(n11459) );
  AND4_X1 U9136 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n13284) );
  INV_X1 U9137 ( .A(n13348), .ZN(n15545) );
  NAND2_X1 U9138 ( .A1(n13295), .A2(n13294), .ZN(n13395) );
  INV_X1 U9139 ( .A(n7596), .ZN(n8204) );
  NAND2_X1 U9140 ( .A1(n7681), .A2(n8525), .ZN(n13036) );
  NOR2_X1 U9141 ( .A1(n7683), .A2(n7682), .ZN(n7681) );
  INV_X1 U9142 ( .A(n12731), .ZN(n7682) );
  INV_X1 U9143 ( .A(n8524), .ZN(n7683) );
  AOI21_X1 U9144 ( .B1(n8543), .B2(n8541), .A(n8540), .ZN(n8539) );
  AND2_X1 U9145 ( .A1(n8521), .A2(n7475), .ZN(n11820) );
  XNOR2_X1 U9146 ( .A(n12730), .B(n12728), .ZN(n12726) );
  NAND2_X1 U9147 ( .A1(n8526), .A2(n8530), .ZN(n12727) );
  NAND2_X1 U9148 ( .A1(n12582), .A2(n8531), .ZN(n8526) );
  NAND2_X1 U9149 ( .A1(n13041), .A2(n13040), .ZN(n13043) );
  NAND2_X1 U9150 ( .A1(n13036), .A2(n13035), .ZN(n13041) );
  AND2_X2 U9151 ( .A1(n9834), .A2(n7665), .ZN(n16521) );
  NAND2_X1 U9152 ( .A1(n11290), .A2(n7423), .ZN(n7665) );
  NAND2_X1 U9153 ( .A1(n14071), .A2(n8543), .ZN(n15061) );
  NAND2_X1 U9154 ( .A1(n14071), .A2(n14070), .ZN(n15060) );
  NAND2_X1 U9155 ( .A1(n15015), .A2(n11975), .ZN(n12206) );
  INV_X1 U9156 ( .A(n15076), .ZN(n15033) );
  NAND2_X1 U9157 ( .A1(n8535), .A2(n8536), .ZN(n13460) );
  INV_X1 U9158 ( .A(n10470), .ZN(n15083) );
  NAND2_X1 U9159 ( .A1(n10498), .A2(n10497), .ZN(n15193) );
  INV_X1 U9160 ( .A(n15184), .ZN(n15212) );
  INV_X1 U9161 ( .A(n13284), .ZN(n15086) );
  XNOR2_X1 U9162 ( .A(n15100), .B(n11460), .ZN(n15108) );
  NOR2_X1 U9163 ( .A1(n7739), .A2(n16227), .ZN(n16229) );
  AOI21_X1 U9164 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n11547), .A(n11546), .ZN(
        n11550) );
  NOR2_X1 U9165 ( .A1(n11736), .A2(n7754), .ZN(n11739) );
  AND2_X1 U9166 ( .A1(n11740), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7754) );
  INV_X1 U9167 ( .A(n7753), .ZN(n11847) );
  NAND2_X1 U9168 ( .A1(n11850), .A2(n11849), .ZN(n12533) );
  AND2_X1 U9169 ( .A1(n7753), .A2(n7752), .ZN(n11850) );
  NAND2_X1 U9170 ( .A1(n11853), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7752) );
  NOR2_X1 U9171 ( .A1(n13099), .A2(n7743), .ZN(n13101) );
  AND2_X1 U9172 ( .A1(n13105), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7743) );
  NOR2_X1 U9173 ( .A1(n15134), .A2(n15133), .ZN(n16240) );
  INV_X1 U9174 ( .A(n7742), .ZN(n15132) );
  NAND2_X1 U9175 ( .A1(n11478), .A2(n11464), .ZN(n16264) );
  NAND2_X1 U9176 ( .A1(n15157), .A2(n15232), .ZN(n15463) );
  NAND2_X1 U9177 ( .A1(n7875), .A2(n15446), .ZN(n7874) );
  NAND2_X1 U9178 ( .A1(n8287), .A2(n8288), .ZN(n15260) );
  AND2_X1 U9179 ( .A1(n10491), .A2(n10420), .ZN(n15281) );
  NAND2_X1 U9180 ( .A1(n8292), .A2(n8293), .ZN(n15274) );
  NAND2_X1 U9181 ( .A1(n15305), .A2(n8294), .ZN(n8292) );
  AOI21_X1 U9182 ( .B1(n15305), .B2(n15306), .A(n7429), .ZN(n15288) );
  NAND2_X1 U9183 ( .A1(n8386), .A2(n8387), .ZN(n15307) );
  AND2_X1 U9184 ( .A1(n15326), .A2(n15325), .ZN(n15501) );
  NAND2_X1 U9185 ( .A1(n8390), .A2(n8389), .ZN(n15324) );
  NAND2_X1 U9186 ( .A1(n8306), .A2(n8305), .ZN(n15339) );
  NAND2_X1 U9187 ( .A1(n8307), .A2(n8310), .ZN(n15354) );
  NAND2_X1 U9188 ( .A1(n15381), .A2(n8311), .ZN(n8307) );
  NAND2_X1 U9189 ( .A1(n15174), .A2(n15173), .ZN(n15440) );
  NAND2_X1 U9190 ( .A1(n12919), .A2(n12918), .ZN(n12920) );
  NAND2_X1 U9191 ( .A1(n7881), .A2(n12297), .ZN(n12490) );
  NAND2_X1 U9192 ( .A1(n11953), .A2(n11952), .ZN(n12290) );
  NAND2_X1 U9193 ( .A1(n8282), .A2(n11829), .ZN(n11936) );
  AND2_X1 U9194 ( .A1(n15429), .A2(n11686), .ZN(n15316) );
  INV_X1 U9195 ( .A(n15316), .ZN(n15456) );
  INV_X1 U9196 ( .A(n12615), .ZN(n12521) );
  NAND2_X1 U9197 ( .A1(n10001), .A2(n10000), .ZN(n12488) );
  NAND2_X1 U9198 ( .A1(n8229), .A2(n9870), .ZN(n8228) );
  AND2_X1 U9199 ( .A1(n16526), .A2(n15546), .ZN(n15536) );
  AND2_X2 U9200 ( .A1(n11908), .A2(n11713), .ZN(n16526) );
  INV_X1 U9201 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8317) );
  OAI211_X1 U9202 ( .C1(n15475), .C2(n15550), .A(n8457), .B(n8456), .ZN(n15562) );
  NOR2_X1 U9203 ( .A1(n15473), .A2(n7605), .ZN(n8456) );
  INV_X1 U9204 ( .A(n15472), .ZN(n8457) );
  INV_X1 U9205 ( .A(n15299), .ZN(n15568) );
  AND2_X1 U9206 ( .A1(n10277), .A2(n10276), .ZN(n15590) );
  OR3_X1 U9207 ( .A1(n15534), .A2(n15533), .A3(n15532), .ZN(n15596) );
  NAND2_X1 U9208 ( .A1(n10231), .A2(n10230), .ZN(n15598) );
  AND2_X1 U9209 ( .A1(n10189), .A2(n10188), .ZN(n15197) );
  NAND2_X1 U9210 ( .A1(n10104), .A2(n10103), .ZN(n13052) );
  INV_X1 U9211 ( .A(n12792), .ZN(n12789) );
  AND2_X1 U9212 ( .A1(n11692), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16223) );
  NAND2_X1 U9213 ( .A1(n9796), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7885) );
  INV_X1 U9214 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n15620) );
  XNOR2_X1 U9215 ( .A(n10559), .B(n10558), .ZN(n15622) );
  NAND2_X1 U9216 ( .A1(n10563), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10559) );
  INV_X1 U9217 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15627) );
  NAND2_X1 U9218 ( .A1(n10563), .A2(n10562), .ZN(n15625) );
  OR2_X1 U9219 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  XNOR2_X1 U9220 ( .A(n10565), .B(n10564), .ZN(n13513) );
  INV_X1 U9221 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13339) );
  INV_X1 U9222 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13256) );
  INV_X1 U9223 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13118) );
  INV_X1 U9224 ( .A(n10515), .ZN(n13027) );
  INV_X1 U9225 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11843) );
  INV_X1 U9226 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11634) );
  INV_X1 U9227 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n11542) );
  INV_X1 U9228 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n11316) );
  INV_X1 U9229 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n11310) );
  AND2_X1 U9230 ( .A1(n9947), .A2(n9997), .ZN(n11520) );
  INV_X1 U9231 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n11313) );
  AND2_X1 U9232 ( .A1(n11277), .A2(P2_U3088), .ZN(n15608) );
  XNOR2_X1 U9233 ( .A(n7756), .B(n7755), .ZN(n15100) );
  INV_X1 U9234 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7755) );
  NOR2_X1 U9235 ( .A1(n15103), .A2(n15605), .ZN(n7756) );
  NOR2_X1 U9236 ( .A1(n11304), .A2(P1_U3086), .ZN(n10814) );
  NAND2_X1 U9237 ( .A1(n7963), .A2(n7507), .ZN(n12417) );
  NAND2_X1 U9238 ( .A1(n11046), .A2(n7967), .ZN(n7966) );
  NAND2_X1 U9239 ( .A1(n7976), .A2(n8717), .ZN(n15630) );
  INV_X1 U9240 ( .A(n8083), .ZN(n15638) );
  NAND2_X1 U9241 ( .A1(n13481), .A2(n8119), .ZN(n15639) );
  NAND2_X1 U9242 ( .A1(n15703), .A2(n13975), .ZN(n15648) );
  NAND2_X1 U9243 ( .A1(n13016), .A2(n13015), .ZN(n13014) );
  AOI21_X1 U9244 ( .B1(n15713), .B2(n15714), .A(n8745), .ZN(n15654) );
  OAI21_X1 U9245 ( .B1(n7975), .B2(n7981), .A(n7971), .ZN(n7970) );
  NAND2_X1 U9246 ( .A1(n7975), .A2(n7972), .ZN(n7971) );
  NAND2_X1 U9247 ( .A1(n7973), .A2(n14017), .ZN(n7972) );
  INV_X1 U9248 ( .A(n7977), .ZN(n7973) );
  NAND2_X1 U9249 ( .A1(n7975), .A2(n14017), .ZN(n7974) );
  NAND2_X1 U9250 ( .A1(n7984), .A2(n7985), .ZN(n15663) );
  AND2_X1 U9251 ( .A1(n8731), .A2(n7991), .ZN(n13325) );
  NAND2_X1 U9252 ( .A1(n16711), .A2(n8727), .ZN(n15680) );
  NAND2_X1 U9253 ( .A1(n8729), .A2(n8728), .ZN(n8727) );
  INV_X1 U9254 ( .A(n11122), .ZN(n8728) );
  NAND2_X1 U9255 ( .A1(n11901), .A2(n11897), .ZN(n11987) );
  NAND2_X1 U9256 ( .A1(n8723), .A2(n8722), .ZN(n15696) );
  AOI21_X1 U9257 ( .B1(n8724), .B2(n8726), .A(n7511), .ZN(n8722) );
  NAND2_X1 U9258 ( .A1(n13752), .A2(n13751), .ZN(n16082) );
  AND2_X1 U9259 ( .A1(n12895), .A2(n7452), .ZN(n8751) );
  NAND2_X1 U9260 ( .A1(n13014), .A2(n11078), .ZN(n13216) );
  NAND2_X1 U9261 ( .A1(n11605), .A2(n11606), .ZN(n11604) );
  OAI21_X1 U9262 ( .B1(n15688), .B2(n15687), .A(n7990), .ZN(n15713) );
  NAND2_X1 U9263 ( .A1(n11161), .A2(n11160), .ZN(n16118) );
  AND2_X1 U9264 ( .A1(n7963), .A2(n7961), .ZN(n12067) );
  NAND2_X1 U9265 ( .A1(n7960), .A2(n7964), .ZN(n12069) );
  NAND2_X1 U9266 ( .A1(n8718), .A2(n13996), .ZN(n15722) );
  NAND2_X1 U9267 ( .A1(n15672), .A2(n15673), .ZN(n8718) );
  NAND2_X1 U9268 ( .A1(n11206), .A2(n16036), .ZN(n16719) );
  OAI21_X1 U9269 ( .B1(n15959), .B2(n10700), .A(n10946), .ZN(n15739) );
  NAND2_X1 U9270 ( .A1(n11170), .A2(n11169), .ZN(n15740) );
  INV_X1 U9271 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n11333) );
  INV_X1 U9272 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13391) );
  INV_X1 U9273 ( .A(n13845), .ZN(n16042) );
  INV_X1 U9274 ( .A(n13852), .ZN(n16045) );
  NAND2_X1 U9275 ( .A1(n8675), .A2(n14028), .ZN(n15845) );
  NAND2_X1 U9276 ( .A1(n15857), .A2(n15856), .ZN(n8675) );
  AND2_X1 U9277 ( .A1(n8713), .A2(n8712), .ZN(n15896) );
  NAND2_X1 U9278 ( .A1(n8672), .A2(n8671), .ZN(n15885) );
  NAND2_X1 U9279 ( .A1(n15926), .A2(n8714), .ZN(n15911) );
  NAND2_X1 U9280 ( .A1(n8060), .A2(n8065), .ZN(n15928) );
  NAND2_X1 U9281 ( .A1(n15966), .A2(n8064), .ZN(n8060) );
  AND2_X1 U9282 ( .A1(n15933), .A2(n15934), .ZN(n15935) );
  NAND2_X1 U9283 ( .A1(n15950), .A2(n8689), .ZN(n15933) );
  NAND2_X1 U9284 ( .A1(n15966), .A2(n8109), .ZN(n15932) );
  NAND2_X1 U9285 ( .A1(n16023), .A2(n8837), .ZN(n16010) );
  NAND2_X1 U9286 ( .A1(n13500), .A2(n13499), .ZN(n13503) );
  NAND2_X1 U9287 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  NAND2_X1 U9288 ( .A1(n8075), .A2(n13150), .ZN(n13196) );
  NAND2_X1 U9289 ( .A1(n10984), .A2(n10983), .ZN(n13659) );
  NAND2_X1 U9290 ( .A1(n12993), .A2(n12992), .ZN(n13149) );
  NAND2_X1 U9291 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  NAND2_X1 U9292 ( .A1(n8039), .A2(n8040), .ZN(n16617) );
  NAND2_X1 U9293 ( .A1(n10754), .A2(n8715), .ZN(n12879) );
  NAND2_X1 U9294 ( .A1(n10754), .A2(n10753), .ZN(n10767) );
  INV_X1 U9295 ( .A(n15825), .ZN(n16636) );
  NAND2_X1 U9296 ( .A1(n8696), .A2(n10775), .ZN(n12481) );
  INV_X1 U9297 ( .A(n11931), .ZN(n8696) );
  INV_X2 U9298 ( .A(n16631), .ZN(n16036) );
  NAND2_X1 U9299 ( .A1(n8048), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8050) );
  OAI21_X1 U9300 ( .B1(n13854), .B2(n11763), .A(n11778), .ZN(n11766) );
  AND2_X1 U9301 ( .A1(n11207), .A2(n11303), .ZN(n16631) );
  INV_X2 U9302 ( .A(n16707), .ZN(n16708) );
  OAI211_X1 U9303 ( .C1(n16053), .C2(n16702), .A(n16052), .B(n8129), .ZN(
        n16146) );
  AND2_X1 U9304 ( .A1(n7587), .A2(n10654), .ZN(n8154) );
  NAND2_X1 U9305 ( .A1(n8034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U9306 ( .A1(n10460), .A2(n10442), .ZN(n15613) );
  OAI21_X1 U9307 ( .B1(n10415), .B2(n7458), .A(n7833), .ZN(n10440) );
  XNOR2_X1 U9308 ( .A(n10488), .B(n10487), .ZN(n16169) );
  NAND2_X1 U9309 ( .A1(n7836), .A2(n10430), .ZN(n10488) );
  NAND2_X1 U9310 ( .A1(n10415), .A2(n7837), .ZN(n7836) );
  INV_X1 U9311 ( .A(n10810), .ZN(n16175) );
  MUX2_X1 U9312 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10627), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n10628) );
  OR2_X1 U9313 ( .A1(n13710), .A2(n10674), .ZN(n13711) );
  NAND2_X1 U9314 ( .A1(n10644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8749) );
  NOR2_X1 U9315 ( .A1(n8087), .A2(n8086), .ZN(n8085) );
  NOR2_X1 U9316 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8086) );
  NAND2_X1 U9317 ( .A1(n10142), .A2(n10141), .ZN(n10147) );
  INV_X1 U9318 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n11455) );
  OAI21_X1 U9319 ( .B1(n10018), .B2(n8642), .A(n8640), .ZN(n10097) );
  AND2_X1 U9320 ( .A1(n11058), .A2(n10998), .ZN(n11587) );
  NAND2_X1 U9321 ( .A1(n10068), .A2(n10046), .ZN(n11450) );
  INV_X1 U9322 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n11325) );
  INV_X1 U9323 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n11300) );
  INV_X1 U9324 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n11280) );
  INV_X1 U9325 ( .A(n8172), .ZN(n16309) );
  XNOR2_X1 U9326 ( .A(n16330), .B(n8590), .ZN(n16332) );
  INV_X1 U9327 ( .A(n7839), .ZN(n16465) );
  OAI21_X1 U9328 ( .B1(n16349), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7488), .ZN(
        n7839) );
  XNOR2_X1 U9329 ( .A(n16352), .B(n8591), .ZN(n16354) );
  INV_X1 U9330 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U9331 ( .A1(n8586), .A2(n16371), .ZN(n16377) );
  NAND2_X1 U9332 ( .A1(n16370), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n8586) );
  XNOR2_X1 U9333 ( .A(n16391), .B(n16392), .ZN(n16393) );
  OAI211_X1 U9334 ( .C1(n8175), .C2(n7842), .A(n7844), .B(n7841), .ZN(n16430)
         );
  NAND2_X1 U9335 ( .A1(n7845), .A2(n16423), .ZN(n7844) );
  INV_X1 U9336 ( .A(n7846), .ZN(n7842) );
  OAI21_X1 U9337 ( .B1(n16442), .B2(n16441), .A(n16440), .ZN(n16444) );
  XNOR2_X1 U9338 ( .A(n8378), .B(n9786), .ZN(P3_U3150) );
  AOI21_X1 U9339 ( .B1(n8379), .B2(n7644), .A(n9782), .ZN(n8378) );
  NOR2_X1 U9340 ( .A1(n8611), .A2(n14175), .ZN(n13959) );
  OR2_X1 U9341 ( .A1(n14175), .A2(n14165), .ZN(n14181) );
  NOR2_X1 U9342 ( .A1(n12355), .A2(n7781), .ZN(n12356) );
  OR2_X1 U9343 ( .A1(n14918), .A2(n14282), .ZN(n8080) );
  NAND2_X1 U9344 ( .A1(n14141), .A2(n12548), .ZN(n12555) );
  NAND2_X1 U9345 ( .A1(n8241), .A2(n8095), .ZN(P3_U3296) );
  AOI21_X1 U9346 ( .B1(n7450), .B2(n8097), .A(n8096), .ZN(n8095) );
  NAND2_X1 U9347 ( .A1(n14508), .A2(n9785), .ZN(n8241) );
  INV_X1 U9348 ( .A(n14321), .ZN(n8097) );
  NAND2_X1 U9349 ( .A1(P3_U3897), .A2(n7783), .ZN(n12063) );
  OR4_X1 U9350 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(
        P3_U3197) );
  INV_X1 U9351 ( .A(n8267), .ZN(n14552) );
  NAND2_X1 U9352 ( .A1(n8272), .A2(n8271), .ZN(P3_U3200) );
  NAND2_X1 U9353 ( .A1(n8273), .A2(n14528), .ZN(n8272) );
  AND2_X1 U9354 ( .A1(n7714), .A2(n7712), .ZN(n8271) );
  NAND2_X1 U9355 ( .A1(n10934), .A2(n14588), .ZN(n8273) );
  NAND2_X1 U9356 ( .A1(n7891), .A2(n14604), .ZN(n7890) );
  NAND2_X1 U9357 ( .A1(n14602), .A2(n14603), .ZN(n8078) );
  NOR2_X1 U9358 ( .A1(n7501), .A2(n8077), .ZN(n7889) );
  NAND2_X1 U9359 ( .A1(n8356), .A2(n8355), .ZN(P3_U3488) );
  NOR2_X1 U9360 ( .A1(n7626), .A2(n7456), .ZN(n8355) );
  NAND2_X1 U9361 ( .A1(n10605), .A2(n16724), .ZN(n8356) );
  NAND2_X1 U9362 ( .A1(n7815), .A2(n7814), .ZN(P3_U3487) );
  NAND2_X1 U9363 ( .A1(n7819), .A2(n7817), .ZN(n7815) );
  NOR2_X1 U9364 ( .A1(n14637), .A2(n7818), .ZN(n7817) );
  NOR2_X1 U9365 ( .A1(n9419), .A2(n9418), .ZN(n9420) );
  OAI21_X1 U9366 ( .B1(n8545), .B2(n14972), .A(n8544), .ZN(P2_U3186) );
  INV_X1 U9367 ( .A(n14976), .ZN(n8544) );
  OAI21_X1 U9368 ( .B1(n8547), .B2(n8546), .A(n15070), .ZN(n8545) );
  AOI21_X1 U9369 ( .B1(n8213), .B2(n8215), .A(n8212), .ZN(n8211) );
  OAI21_X1 U9370 ( .B1(n15078), .B2(n15077), .A(n7693), .ZN(n7692) );
  NAND2_X1 U9371 ( .A1(n8225), .A2(n8223), .ZN(P2_U3530) );
  AOI21_X1 U9372 ( .B1(n15552), .B2(n15536), .A(n8224), .ZN(n8223) );
  NAND2_X1 U9373 ( .A1(n15553), .A2(n16526), .ZN(n8225) );
  NOR2_X1 U9374 ( .A1(n16526), .A2(n10483), .ZN(n8224) );
  NAND2_X1 U9375 ( .A1(n8455), .A2(n8454), .ZN(P2_U3527) );
  OR2_X1 U9376 ( .A1(n16526), .A2(n10452), .ZN(n8454) );
  NAND2_X1 U9377 ( .A1(n15562), .A2(n16526), .ZN(n8455) );
  NAND2_X1 U9378 ( .A1(n7671), .A2(n7670), .ZN(n15555) );
  NAND2_X1 U9379 ( .A1(n16527), .A2(n15554), .ZN(n7670) );
  OAI21_X1 U9380 ( .B1(n8839), .B2(n8316), .A(n8315), .ZN(P2_U3496) );
  NAND2_X1 U9381 ( .A1(n16529), .A2(n16523), .ZN(n8316) );
  OR4_X1 U9382 ( .A1(n11222), .A2(n11221), .A3(n11220), .A4(n11219), .ZN(
        P1_U3233) );
  AOI21_X1 U9383 ( .B1(n8648), .B2(n8647), .A(n13911), .ZN(n8161) );
  NAND2_X1 U9384 ( .A1(n16384), .A2(n16383), .ZN(n16385) );
  INV_X1 U9385 ( .A(n7869), .ZN(n16400) );
  INV_X1 U9386 ( .A(n16416), .ZN(n7847) );
  XNOR2_X1 U9387 ( .A(n16463), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8176) );
  NAND2_X1 U9388 ( .A1(n7866), .A2(n16456), .ZN(n7865) );
  AND2_X2 U9389 ( .A1(n14957), .A2(n8861), .ZN(n9031) );
  INV_X2 U9390 ( .A(n9977), .ZN(n10499) );
  OR2_X1 U9391 ( .A1(n15360), .A2(n15184), .ZN(n7424) );
  AND2_X1 U9392 ( .A1(n15248), .A2(n10572), .ZN(n7425) );
  AND2_X1 U9393 ( .A1(n14829), .A2(n16724), .ZN(n7426) );
  AND2_X1 U9394 ( .A1(n13772), .A2(n13774), .ZN(n7427) );
  INV_X1 U9395 ( .A(n14797), .ZN(n8237) );
  INV_X1 U9396 ( .A(n16417), .ZN(n7850) );
  OR2_X1 U9397 ( .A1(n10295), .A2(SI_19_), .ZN(n7428) );
  INV_X1 U9398 ( .A(n14579), .ZN(n11805) );
  XNOR2_X1 U9399 ( .A(n8276), .B(n8275), .ZN(n10878) );
  INV_X1 U9400 ( .A(n16026), .ZN(n8687) );
  NAND2_X1 U9401 ( .A1(n9811), .A2(n9810), .ZN(n10569) );
  AND2_X1 U9402 ( .A1(n15496), .A2(n15191), .ZN(n7429) );
  XOR2_X1 U9403 ( .A(n14110), .B(n7695), .Z(n7430) );
  INV_X1 U9404 ( .A(n12296), .ZN(n8301) );
  NOR2_X1 U9405 ( .A1(n8394), .A2(n15333), .ZN(n8389) );
  INV_X1 U9406 ( .A(n8626), .ZN(n8625) );
  NAND2_X1 U9407 ( .A1(n8627), .A2(n13931), .ZN(n8626) );
  OR2_X1 U9408 ( .A1(n10159), .A2(n10161), .ZN(n7431) );
  AND2_X1 U9409 ( .A1(n8698), .A2(n8697), .ZN(n7432) );
  OR2_X1 U9410 ( .A1(n15675), .A2(n15865), .ZN(n7433) );
  AOI21_X1 U9411 ( .B1(n8732), .B2(n8733), .A(n7543), .ZN(n8731) );
  XNOR2_X1 U9412 ( .A(n8860), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U9413 ( .A1(n8798), .A2(n8794), .ZN(n7434) );
  AND2_X1 U9414 ( .A1(n8628), .A2(n7474), .ZN(n7435) );
  AND2_X1 U9415 ( .A1(n8226), .A2(n15576), .ZN(n7436) );
  AND2_X1 U9416 ( .A1(n10340), .A2(n10341), .ZN(n7439) );
  XNOR2_X1 U9417 ( .A(n7481), .B(n9378), .ZN(n9393) );
  NAND2_X1 U9418 ( .A1(n10444), .A2(n10443), .ZN(n15474) );
  AND2_X1 U9419 ( .A1(n13249), .A2(n14403), .ZN(n7440) );
  NAND2_X1 U9420 ( .A1(n14789), .A2(n8360), .ZN(n14775) );
  OR2_X1 U9421 ( .A1(n9923), .A2(SI_4_), .ZN(n7441) );
  NAND2_X1 U9422 ( .A1(n15585), .A2(n15183), .ZN(n7442) );
  OR2_X1 U9423 ( .A1(n9939), .A2(SI_5_), .ZN(n7443) );
  AND2_X1 U9424 ( .A1(n10153), .A2(n10152), .ZN(n13240) );
  INV_X1 U9425 ( .A(n13240), .ZN(n13274) );
  INV_X1 U9426 ( .A(n15027), .ZN(n7690) );
  NAND2_X1 U9427 ( .A1(n11127), .A2(n11126), .ZN(n16129) );
  INV_X1 U9428 ( .A(n14048), .ZN(n15974) );
  AND2_X1 U9429 ( .A1(n15572), .A2(n7436), .ZN(n7444) );
  INV_X1 U9430 ( .A(n8206), .ZN(n8205) );
  OAI21_X1 U9431 ( .B1(n7466), .B2(n8207), .A(n10186), .ZN(n8206) );
  INV_X1 U9432 ( .A(n14702), .ZN(n14673) );
  AND2_X1 U9433 ( .A1(n9289), .A2(n9288), .ZN(n14702) );
  AND2_X1 U9434 ( .A1(n8185), .A2(n8184), .ZN(n7445) );
  AND2_X1 U9435 ( .A1(n8159), .A2(n10670), .ZN(n7446) );
  AND2_X1 U9436 ( .A1(n7434), .A2(n7524), .ZN(n7447) );
  NAND2_X1 U9437 ( .A1(n7874), .A2(n7594), .ZN(n7448) );
  AND3_X1 U9438 ( .A1(n8244), .A2(n8243), .A3(n14509), .ZN(n7449) );
  INV_X1 U9439 ( .A(n16054), .ZN(n15839) );
  NAND2_X1 U9440 ( .A1(n13804), .A2(n13803), .ZN(n16054) );
  AND2_X1 U9441 ( .A1(n7449), .A2(n9785), .ZN(n7450) );
  AND2_X1 U9442 ( .A1(n9884), .A2(n9883), .ZN(n7451) );
  NAND2_X1 U9443 ( .A1(n9371), .A2(n14445), .ZN(n14634) );
  AND2_X1 U9444 ( .A1(n10462), .A2(n10461), .ZN(n15470) );
  INV_X1 U9445 ( .A(n15470), .ZN(n15236) );
  INV_X1 U9446 ( .A(n13968), .ZN(n14005) );
  NAND2_X1 U9447 ( .A1(n11055), .A2(n11054), .ZN(n7452) );
  NAND2_X1 U9448 ( .A1(n16137), .A2(n13505), .ZN(n7453) );
  INV_X1 U9449 ( .A(n13209), .ZN(n8256) );
  INV_X1 U9450 ( .A(n15192), .ZN(n15219) );
  AND2_X1 U9451 ( .A1(n10426), .A2(n10425), .ZN(n15192) );
  NAND2_X1 U9452 ( .A1(n13708), .A2(n8761), .ZN(n7454) );
  INV_X1 U9453 ( .A(n13542), .ZN(n8370) );
  INV_X1 U9454 ( .A(n15937), .ZN(n8066) );
  INV_X1 U9455 ( .A(n16062), .ZN(n8196) );
  NAND2_X1 U9456 ( .A1(n13712), .A2(n16181), .ZN(n15921) );
  INV_X1 U9457 ( .A(n15921), .ZN(n8191) );
  NAND2_X1 U9458 ( .A1(n9118), .A2(n9119), .ZN(n9121) );
  OR2_X1 U9459 ( .A1(n8269), .A2(n10864), .ZN(n7455) );
  INV_X1 U9460 ( .A(n8636), .ZN(n8635) );
  NAND2_X1 U9461 ( .A1(n7620), .A2(n7428), .ZN(n8636) );
  NOR2_X1 U9462 ( .A1(n10606), .A2(n14872), .ZN(n7456) );
  NAND2_X1 U9463 ( .A1(n8887), .A2(n8886), .ZN(n8094) );
  AND2_X1 U9464 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n8568), .ZN(n7457) );
  INV_X1 U9465 ( .A(n15077), .ZN(n15070) );
  OR2_X1 U9466 ( .A1(n10487), .A2(n7835), .ZN(n7458) );
  INV_X1 U9467 ( .A(n14551), .ZN(n8266) );
  OR2_X1 U9468 ( .A1(n13587), .A2(n10647), .ZN(n11072) );
  INV_X1 U9469 ( .A(n15222), .ZN(n15223) );
  INV_X1 U9470 ( .A(n8963), .ZN(n14312) );
  NAND4_X1 U9471 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), .ZN(n7459)
         );
  INV_X1 U9472 ( .A(n13866), .ZN(n8660) );
  NAND2_X1 U9473 ( .A1(n14057), .A2(n13565), .ZN(n10677) );
  AND2_X1 U9474 ( .A1(n9365), .A2(n14466), .ZN(n7461) );
  INV_X1 U9475 ( .A(n15832), .ZN(n8057) );
  XNOR2_X1 U9476 ( .A(n9812), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10515) );
  NAND2_X1 U9477 ( .A1(n8059), .A2(n8058), .ZN(n8713) );
  INV_X1 U9478 ( .A(n10326), .ZN(n8819) );
  NOR2_X1 U9479 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n10672) );
  INV_X1 U9480 ( .A(n14017), .ZN(n7981) );
  AND2_X1 U9481 ( .A1(n12594), .A2(n9000), .ZN(n7462) );
  INV_X1 U9482 ( .A(n15576), .ZN(n15503) );
  OR2_X1 U9483 ( .A1(n15342), .A2(n15214), .ZN(n7463) );
  OR2_X1 U9484 ( .A1(n15539), .A2(n15200), .ZN(n7464) );
  INV_X1 U9485 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9386) );
  AND2_X1 U9486 ( .A1(n8606), .A2(n13920), .ZN(n7465) );
  AND2_X1 U9487 ( .A1(n8209), .A2(n10141), .ZN(n7466) );
  INV_X1 U9488 ( .A(n10178), .ZN(n7928) );
  AND2_X1 U9489 ( .A1(n13040), .A2(n13042), .ZN(n7467) );
  INV_X1 U9490 ( .A(n8284), .ZN(n11716) );
  AND2_X1 U9491 ( .A1(n14091), .A2(n14092), .ZN(n7468) );
  INV_X1 U9492 ( .A(n14803), .ZN(n8234) );
  AND2_X1 U9493 ( .A1(n8820), .A2(n8819), .ZN(n7469) );
  AND2_X1 U9494 ( .A1(n15887), .A2(n8194), .ZN(n7470) );
  OR2_X1 U9495 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n9290), .ZN(n7471) );
  INV_X1 U9496 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8845) );
  INV_X1 U9497 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15103) );
  AND2_X1 U9498 ( .A1(n16228), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7472) );
  AND2_X1 U9499 ( .A1(n8190), .A2(n8066), .ZN(n7473) );
  AND4_X1 U9500 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n9151), .ZN(n7474)
         );
  NAND2_X1 U9501 ( .A1(n11813), .A2(n11812), .ZN(n7475) );
  AND2_X1 U9502 ( .A1(n7769), .A2(n7767), .ZN(n7476) );
  INV_X1 U9503 ( .A(n8383), .ZN(n8382) );
  NAND2_X1 U9504 ( .A1(n12918), .A2(n8384), .ZN(n8383) );
  OR2_X1 U9505 ( .A1(n8057), .A2(n8128), .ZN(n7477) );
  AND2_X1 U9506 ( .A1(n10316), .A2(n10315), .ZN(n15360) );
  INV_X1 U9507 ( .A(n15360), .ZN(n8227) );
  AND2_X1 U9508 ( .A1(n16123), .A2(n15741), .ZN(n7478) );
  AND2_X1 U9509 ( .A1(n14687), .A2(n7796), .ZN(n7479) );
  INV_X1 U9510 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n16322) );
  AND2_X1 U9511 ( .A1(n13872), .A2(n7453), .ZN(n7480) );
  OR2_X1 U9512 ( .A1(n8593), .A2(n9386), .ZN(n7481) );
  AND2_X1 U9513 ( .A1(n13637), .A2(n15750), .ZN(n7482) );
  AND2_X1 U9514 ( .A1(n8960), .A2(n8949), .ZN(n7483) );
  INV_X1 U9515 ( .A(n8837), .ZN(n8686) );
  INV_X1 U9516 ( .A(n10094), .ZN(n7949) );
  OR2_X1 U9517 ( .A1(n15905), .A2(n15917), .ZN(n7484) );
  OR2_X1 U9518 ( .A1(n16392), .A2(n16391), .ZN(n7485) );
  AND2_X1 U9519 ( .A1(n10061), .A2(n10062), .ZN(n7486) );
  OR2_X1 U9520 ( .A1(n13712), .A2(n11341), .ZN(n7487) );
  NAND2_X1 U9521 ( .A1(n11000), .A2(n10999), .ZN(n16633) );
  NAND2_X1 U9522 ( .A1(n13706), .A2(n13705), .ZN(n15937) );
  INV_X1 U9523 ( .A(n9876), .ZN(n14066) );
  NAND2_X1 U9524 ( .A1(n8228), .A2(n8231), .ZN(n9876) );
  OR2_X1 U9525 ( .A1(n16348), .A2(n16347), .ZN(n7488) );
  OR2_X1 U9526 ( .A1(n7939), .A2(n7938), .ZN(n7489) );
  AND2_X1 U9527 ( .A1(n13962), .A2(n13961), .ZN(n7490) );
  OR2_X1 U9528 ( .A1(n10821), .A2(n12166), .ZN(n7491) );
  NOR2_X1 U9529 ( .A1(n14634), .A2(n8264), .ZN(n8263) );
  AND2_X1 U9530 ( .A1(n8527), .A2(n12726), .ZN(n7492) );
  AND3_X1 U9531 ( .A1(n8366), .A2(n8616), .A3(n7797), .ZN(n7493) );
  NAND2_X1 U9532 ( .A1(n13799), .A2(n13798), .ZN(n16062) );
  NAND2_X1 U9533 ( .A1(n8616), .A2(n8617), .ZN(n9010) );
  NOR2_X1 U9534 ( .A1(n14983), .A2(n8084), .ZN(n7494) );
  NOR2_X1 U9535 ( .A1(n15843), .A2(n8128), .ZN(n7495) );
  NAND2_X1 U9536 ( .A1(n13770), .A2(n13769), .ZN(n16074) );
  INV_X1 U9537 ( .A(n10406), .ZN(n8801) );
  AND2_X1 U9538 ( .A1(n13394), .A2(n13393), .ZN(n7496) );
  AND2_X1 U9539 ( .A1(n9411), .A2(n8594), .ZN(n7497) );
  INV_X1 U9540 ( .A(n14973), .ZN(n8546) );
  AND2_X1 U9541 ( .A1(n8210), .A2(n8211), .ZN(n7498) );
  AND2_X1 U9542 ( .A1(n8216), .A2(n8214), .ZN(n7499) );
  NOR2_X1 U9543 ( .A1(n14550), .A2(n8265), .ZN(n7500) );
  NOR2_X1 U9544 ( .A1(n14612), .A2(n14611), .ZN(n7501) );
  AND2_X1 U9545 ( .A1(n7467), .A2(n12731), .ZN(n7502) );
  INV_X1 U9546 ( .A(n7777), .ZN(n14645) );
  NAND2_X1 U9547 ( .A1(n14330), .A2(n14329), .ZN(n7777) );
  INV_X1 U9548 ( .A(n7664), .ZN(n15263) );
  NOR2_X1 U9549 ( .A1(n15280), .A2(n15478), .ZN(n7664) );
  INV_X1 U9550 ( .A(n13648), .ZN(n8777) );
  AND2_X1 U9551 ( .A1(n13754), .A2(n13753), .ZN(n7503) );
  AND2_X1 U9552 ( .A1(n16062), .A2(n15828), .ZN(n7504) );
  INV_X1 U9553 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9790) );
  AND2_X1 U9554 ( .A1(n11495), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7505) );
  AND2_X1 U9555 ( .A1(n8740), .A2(n8738), .ZN(n7506) );
  INV_X1 U9556 ( .A(n8622), .ZN(n8621) );
  NAND2_X1 U9557 ( .A1(n13090), .A2(n13089), .ZN(n8622) );
  INV_X1 U9558 ( .A(n7986), .ZN(n7985) );
  OAI21_X1 U9559 ( .B1(n8737), .B2(n7987), .A(n8735), .ZN(n7986) );
  NOR2_X1 U9560 ( .A1(n14581), .A2(n14794), .ZN(n8331) );
  AND2_X1 U9561 ( .A1(n7961), .A2(n7966), .ZN(n7507) );
  NAND2_X1 U9562 ( .A1(n8672), .A2(n7484), .ZN(n7508) );
  INV_X1 U9563 ( .A(n8394), .ZN(n8393) );
  NOR2_X1 U9564 ( .A1(n15580), .A2(n15215), .ZN(n8394) );
  AND2_X1 U9565 ( .A1(n10513), .A2(n10512), .ZN(n15560) );
  INV_X1 U9566 ( .A(n15560), .ZN(n15467) );
  AND2_X1 U9567 ( .A1(n7982), .A2(n8119), .ZN(n7509) );
  OR2_X1 U9568 ( .A1(n14095), .A2(n14094), .ZN(n7510) );
  AND2_X1 U9569 ( .A1(n14340), .A2(n14341), .ZN(n14493) );
  AND2_X1 U9570 ( .A1(n13981), .A2(n13980), .ZN(n7511) );
  AND2_X1 U9571 ( .A1(n14004), .A2(n14003), .ZN(n7512) );
  OR2_X1 U9572 ( .A1(n16025), .A2(n16026), .ZN(n16023) );
  OR2_X1 U9573 ( .A1(n8520), .A2(n8517), .ZN(n7513) );
  INV_X1 U9574 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8275) );
  INV_X1 U9575 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10664) );
  AND2_X1 U9576 ( .A1(n14011), .A2(n14010), .ZN(n7514) );
  OR2_X1 U9577 ( .A1(n8801), .A2(n10408), .ZN(n7515) );
  INV_X1 U9578 ( .A(n8251), .ZN(n8250) );
  AOI21_X1 U9579 ( .B1(n8253), .B2(n13209), .A(n7598), .ZN(n8251) );
  OR2_X1 U9580 ( .A1(n14243), .A2(n8624), .ZN(n7516) );
  NOR2_X1 U9581 ( .A1(n12488), .A2(n12487), .ZN(n7517) );
  NOR2_X1 U9582 ( .A1(n15598), .A2(n15202), .ZN(n7518) );
  NOR2_X1 U9583 ( .A1(n15585), .A2(n15210), .ZN(n7519) );
  AND2_X1 U9584 ( .A1(n11942), .A2(n12109), .ZN(n7520) );
  AND2_X1 U9585 ( .A1(n15576), .A2(n15216), .ZN(n7521) );
  OR2_X1 U9586 ( .A1(n8615), .A2(n13953), .ZN(n7522) );
  INV_X1 U9587 ( .A(n8110), .ZN(n8109) );
  NOR2_X1 U9588 ( .A1(n16104), .A2(n15976), .ZN(n8110) );
  OAI22_X1 U9589 ( .A1(SI_27_), .A2(n9434), .B1(n14964), .B2(keyinput_133), 
        .ZN(n9435) );
  INV_X1 U9590 ( .A(n7433), .ZN(n8701) );
  INV_X1 U9591 ( .A(n8026), .ZN(n8022) );
  OR2_X1 U9592 ( .A1(n16118), .A2(n15977), .ZN(n8026) );
  OR2_X1 U9593 ( .A1(n10639), .A2(n8035), .ZN(n7523) );
  NAND2_X1 U9594 ( .A1(n8798), .A2(n7515), .ZN(n7524) );
  NAND2_X1 U9595 ( .A1(n10672), .A2(n10620), .ZN(n10695) );
  INV_X1 U9596 ( .A(n10695), .ZN(n8090) );
  AND2_X1 U9597 ( .A1(n8044), .A2(n8045), .ZN(n7525) );
  NOR2_X1 U9598 ( .A1(n15585), .A2(n15183), .ZN(n7526) );
  NAND2_X1 U9599 ( .A1(n10226), .A2(n10205), .ZN(n7527) );
  INV_X1 U9600 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n15605) );
  AND2_X1 U9601 ( .A1(n10680), .A2(n10682), .ZN(n7528) );
  INV_X1 U9602 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9151) );
  INV_X1 U9603 ( .A(n15284), .ZN(n15483) );
  AND2_X1 U9604 ( .A1(n10417), .A2(n10416), .ZN(n15284) );
  OR2_X1 U9605 ( .A1(n10010), .A2(n10011), .ZN(n7529) );
  NAND2_X1 U9606 ( .A1(n9820), .A2(n9821), .ZN(n7530) );
  INV_X1 U9607 ( .A(n8187), .ZN(n8186) );
  NAND2_X1 U9608 ( .A1(n13425), .A2(n8188), .ZN(n8187) );
  INV_X1 U9609 ( .A(n8195), .ZN(n8194) );
  NAND2_X1 U9610 ( .A1(n8196), .A2(n8197), .ZN(n8195) );
  AND4_X1 U9611 ( .A1(n9788), .A2(n9789), .A3(n9806), .A4(n9790), .ZN(n7531)
         );
  AND2_X1 U9612 ( .A1(n10203), .A2(n11603), .ZN(n7532) );
  AND4_X1 U9613 ( .A1(n7661), .A2(n7660), .A3(n7662), .A4(n10255), .ZN(n7533)
         );
  OR2_X1 U9614 ( .A1(n16323), .A2(n16322), .ZN(n7534) );
  INV_X1 U9615 ( .A(n8413), .ZN(n8412) );
  INV_X1 U9616 ( .A(n8340), .ZN(n8339) );
  NAND2_X1 U9617 ( .A1(n8344), .A2(n8345), .ZN(n8340) );
  NAND2_X1 U9618 ( .A1(n9292), .A2(n9345), .ZN(n14918) );
  INV_X1 U9619 ( .A(n8747), .ZN(n8745) );
  NAND2_X1 U9620 ( .A1(n11176), .A2(n11175), .ZN(n8747) );
  BUF_X1 U9621 ( .A(n13582), .Z(n8105) );
  AND2_X1 U9622 ( .A1(n12211), .A2(n12210), .ZN(n7535) );
  AND2_X1 U9623 ( .A1(n11300), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7536) );
  AND2_X1 U9624 ( .A1(n8868), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U9625 ( .A1(n8711), .A2(n8714), .ZN(n7538) );
  NOR2_X1 U9626 ( .A1(n8811), .A2(n10160), .ZN(n7539) );
  NOR2_X1 U9627 ( .A1(n15568), .A2(n15218), .ZN(n7540) );
  NOR2_X1 U9628 ( .A1(n14914), .A2(n14690), .ZN(n7541) );
  AND2_X1 U9629 ( .A1(n15284), .A2(n15192), .ZN(n7542) );
  AND2_X1 U9630 ( .A1(n11093), .A2(n11092), .ZN(n7543) );
  OAI21_X1 U9631 ( .B1(n8311), .B2(n8309), .A(n15185), .ZN(n8308) );
  AND2_X1 U9632 ( .A1(n8160), .A2(n8158), .ZN(n7544) );
  INV_X1 U9633 ( .A(n8310), .ZN(n8309) );
  NAND2_X1 U9634 ( .A1(n7526), .A2(n7442), .ZN(n8310) );
  NAND2_X1 U9635 ( .A1(n8769), .A2(n13801), .ZN(n7545) );
  INV_X1 U9636 ( .A(n15496), .ZN(n15572) );
  NAND2_X1 U9637 ( .A1(n10373), .A2(n10372), .ZN(n15496) );
  INV_X1 U9638 ( .A(n13700), .ZN(n8153) );
  INV_X1 U9639 ( .A(n13863), .ZN(n10780) );
  OR2_X1 U9640 ( .A1(n10061), .A2(n10062), .ZN(n7546) );
  OR2_X1 U9641 ( .A1(n16399), .A2(n16398), .ZN(n7547) );
  NOR2_X1 U9642 ( .A1(n15868), .A2(n14050), .ZN(n7548) );
  AND2_X1 U9643 ( .A1(n7977), .A2(n7981), .ZN(n7549) );
  OR2_X1 U9644 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n16308), .ZN(n7550) );
  OR2_X1 U9645 ( .A1(n15284), .A2(n15192), .ZN(n7551) );
  AND2_X1 U9646 ( .A1(n7968), .A2(n12068), .ZN(n7552) );
  AND3_X1 U9647 ( .A1(n9795), .A2(n9825), .A3(n7884), .ZN(n7553) );
  AND2_X1 U9648 ( .A1(n7958), .A2(n9964), .ZN(n7554) );
  AND2_X1 U9649 ( .A1(n15895), .A2(n8712), .ZN(n7555) );
  INV_X1 U9650 ( .A(n9987), .ZN(n7958) );
  AND2_X1 U9651 ( .A1(n9085), .A2(n9067), .ZN(n7556) );
  INV_X1 U9652 ( .A(n14353), .ZN(n7811) );
  AND2_X1 U9653 ( .A1(n8827), .A2(n10180), .ZN(n7557) );
  OR2_X1 U9654 ( .A1(n8814), .A2(n7469), .ZN(n7558) );
  NOR2_X1 U9655 ( .A1(n15418), .A2(n8407), .ZN(n8406) );
  AND2_X1 U9656 ( .A1(n8037), .A2(n12995), .ZN(n7559) );
  OR2_X1 U9657 ( .A1(n8487), .A2(n8486), .ZN(n7560) );
  AND2_X1 U9658 ( .A1(n9836), .A2(n9835), .ZN(n7561) );
  AND2_X1 U9659 ( .A1(n8321), .A2(n8326), .ZN(n7562) );
  INV_X1 U9660 ( .A(n10776), .ZN(n8695) );
  AND2_X1 U9661 ( .A1(n8697), .A2(n7433), .ZN(n7563) );
  INV_X1 U9662 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10632) );
  AND2_X1 U9663 ( .A1(n9045), .A2(n9030), .ZN(n7564) );
  AND2_X1 U9664 ( .A1(n8021), .A2(n8024), .ZN(n7565) );
  AND2_X1 U9665 ( .A1(n14789), .A2(n9193), .ZN(n7566) );
  AND2_X1 U9666 ( .A1(n11819), .A2(n7475), .ZN(n7567) );
  OR2_X1 U9667 ( .A1(n13741), .A2(n8765), .ZN(n7568) );
  AND2_X1 U9668 ( .A1(n8827), .A2(n7928), .ZN(n7569) );
  AND2_X1 U9669 ( .A1(n7653), .A2(n7663), .ZN(n7570) );
  OR2_X1 U9670 ( .A1(n13636), .A2(n13634), .ZN(n7571) );
  AND2_X1 U9671 ( .A1(n13677), .A2(n13675), .ZN(n7572) );
  AND2_X1 U9672 ( .A1(n7847), .A2(n7850), .ZN(n7573) );
  OR2_X1 U9673 ( .A1(n8964), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n7574) );
  AND2_X1 U9674 ( .A1(n7944), .A2(n7946), .ZN(n7575) );
  AND2_X1 U9675 ( .A1(n11078), .A2(n8734), .ZN(n8733) );
  AND2_X1 U9676 ( .A1(n7454), .A2(n8152), .ZN(n7576) );
  AND2_X1 U9677 ( .A1(n8903), .A2(n8373), .ZN(n7577) );
  NAND2_X1 U9678 ( .A1(n13773), .A2(n8762), .ZN(n7578) );
  INV_X1 U9679 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10654) );
  AND2_X1 U9680 ( .A1(n8055), .A2(n8056), .ZN(n7579) );
  AND2_X1 U9681 ( .A1(n8310), .A2(n7424), .ZN(n7580) );
  AND2_X1 U9682 ( .A1(n7545), .A2(n8141), .ZN(n7581) );
  AND2_X1 U9683 ( .A1(n10205), .A2(n10206), .ZN(n7582) );
  AND2_X1 U9684 ( .A1(n9800), .A2(n9801), .ZN(n7583) );
  OR2_X1 U9685 ( .A1(n8803), .A2(n8804), .ZN(n7584) );
  INV_X1 U9686 ( .A(n12259), .ZN(n7705) );
  INV_X1 U9687 ( .A(n8372), .ZN(n8371) );
  NAND2_X1 U9688 ( .A1(n8234), .A2(n9163), .ZN(n8372) );
  INV_X1 U9689 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7884) );
  OR2_X1 U9690 ( .A1(n13740), .A2(n8764), .ZN(n7585) );
  NAND2_X1 U9691 ( .A1(n10530), .A2(n10531), .ZN(n7586) );
  INV_X1 U9692 ( .A(n7879), .ZN(n7878) );
  OR2_X1 U9693 ( .A1(n12489), .A2(n7880), .ZN(n7879) );
  AND2_X1 U9694 ( .A1(n10652), .A2(n10664), .ZN(n7587) );
  NAND2_X1 U9695 ( .A1(n10947), .A2(n11015), .ZN(n13969) );
  INV_X1 U9696 ( .A(n15934), .ZN(n8047) );
  OR2_X1 U9697 ( .A1(n12883), .A2(n13863), .ZN(n8039) );
  INV_X1 U9698 ( .A(n14682), .ZN(n8344) );
  INV_X1 U9699 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10611) );
  AND2_X1 U9700 ( .A1(n13422), .A2(n8186), .ZN(n7588) );
  AND2_X1 U9701 ( .A1(n8039), .A2(n8037), .ZN(n7589) );
  INV_X1 U9702 ( .A(n13208), .ZN(n8254) );
  NOR2_X1 U9703 ( .A1(n16015), .A2(n8704), .ZN(n8707) );
  AND2_X1 U9704 ( .A1(n8535), .A2(n8533), .ZN(n7590) );
  INV_X1 U9705 ( .A(SI_16_), .ZN(n11753) );
  AND2_X1 U9706 ( .A1(n14922), .A2(n14720), .ZN(n7591) );
  AND2_X1 U9707 ( .A1(n15372), .A2(n7436), .ZN(n7592) );
  OR2_X1 U9708 ( .A1(n12745), .A2(n7916), .ZN(n7593) );
  INV_X1 U9709 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8568) );
  AND2_X1 U9710 ( .A1(n15230), .A2(n15229), .ZN(n7594) );
  AND2_X1 U9711 ( .A1(n15215), .A2(n7418), .ZN(n7595) );
  AND3_X1 U9712 ( .A1(n9265), .A2(n9264), .A3(n9263), .ZN(n14737) );
  INV_X1 U9713 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8367) );
  INV_X1 U9714 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8375) );
  INV_X1 U9715 ( .A(n10206), .ZN(n8644) );
  XOR2_X1 U9716 ( .A(n15576), .B(n11679), .Z(n7596) );
  OR2_X1 U9717 ( .A1(n14902), .A2(n14872), .ZN(n7597) );
  AND2_X1 U9718 ( .A1(n9358), .A2(n14402), .ZN(n7598) );
  NAND2_X1 U9719 ( .A1(n10455), .A2(n10454), .ZN(n15226) );
  AND2_X1 U9720 ( .A1(n13422), .A2(n8185), .ZN(n7599) );
  AND2_X1 U9721 ( .A1(n14796), .A2(n14806), .ZN(n7600) );
  OR2_X1 U9722 ( .A1(n14906), .A2(n14872), .ZN(n7601) );
  OR3_X1 U9723 ( .A1(n8426), .A2(n9711), .A3(n9710), .ZN(n7602) );
  AND2_X1 U9724 ( .A1(n13934), .A2(n14187), .ZN(n7603) );
  XOR2_X1 U9725 ( .A(n12249), .B(n9472), .Z(n7604) );
  AND2_X1 U9726 ( .A1(n15474), .A2(n15546), .ZN(n7605) );
  AND2_X1 U9727 ( .A1(n8708), .A2(n14044), .ZN(n7606) );
  INV_X1 U9728 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9729 ( .A1(n15998), .A2(n7473), .ZN(n8192) );
  OR2_X1 U9730 ( .A1(n7718), .A2(n10896), .ZN(n7607) );
  AND2_X1 U9731 ( .A1(n8268), .A2(n8270), .ZN(n7608) );
  NAND2_X1 U9732 ( .A1(n8146), .A2(n7453), .ZN(n7609) );
  AND2_X1 U9733 ( .A1(n13540), .A2(n8371), .ZN(n7610) );
  AND2_X1 U9734 ( .A1(n12919), .A2(n8382), .ZN(n7611) );
  NOR2_X1 U9735 ( .A1(n16529), .A2(n8317), .ZN(n7612) );
  NOR2_X1 U9736 ( .A1(n14882), .A2(n14227), .ZN(n7613) );
  NOR2_X1 U9737 ( .A1(n14873), .A2(n14156), .ZN(n7614) );
  OR2_X1 U9738 ( .A1(n13070), .A2(n10877), .ZN(n7615) );
  INV_X1 U9739 ( .A(n7921), .ZN(n7920) );
  NOR2_X1 U9740 ( .A1(n11309), .A2(n10836), .ZN(n7921) );
  NOR2_X1 U9741 ( .A1(n8023), .A2(n8022), .ZN(n7616) );
  AND2_X1 U9742 ( .A1(n10330), .A2(SI_21_), .ZN(n7617) );
  INV_X1 U9743 ( .A(n8532), .ZN(n8203) );
  OR2_X1 U9744 ( .A1(n15188), .A2(n15232), .ZN(n8532) );
  NAND2_X1 U9745 ( .A1(n7597), .A2(n7820), .ZN(n7618) );
  AND2_X1 U9746 ( .A1(n10313), .A2(SI_20_), .ZN(n7619) );
  AND2_X1 U9747 ( .A1(n10863), .A2(n14531), .ZN(n10864) );
  OR2_X1 U9748 ( .A1(n10313), .A2(SI_20_), .ZN(n7620) );
  OR2_X1 U9749 ( .A1(n14902), .A2(n14938), .ZN(n7621) );
  OR2_X1 U9750 ( .A1(n14906), .A2(n14938), .ZN(n7622) );
  AOI21_X1 U9751 ( .B1(n8562), .B2(n8564), .A(n7457), .ZN(n8561) );
  NAND2_X1 U9752 ( .A1(n11297), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7623) );
  INV_X1 U9753 ( .A(n13656), .ZN(n13136) );
  NAND2_X1 U9754 ( .A1(n11081), .A2(n11080), .ZN(n13656) );
  INV_X1 U9755 ( .A(n16724), .ZN(n7821) );
  NAND2_X1 U9756 ( .A1(n11217), .A2(n11216), .ZN(n15957) );
  INV_X1 U9757 ( .A(n15957), .ZN(n8149) );
  NAND2_X1 U9758 ( .A1(n7680), .A2(n7678), .ZN(n7624) );
  INV_X1 U9759 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8577) );
  INV_X1 U9760 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8551) );
  XOR2_X1 U9761 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .Z(n7625) );
  AND2_X1 U9762 ( .A1(n7821), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7626) );
  AND2_X1 U9763 ( .A1(n8889), .A2(n8888), .ZN(n7627) );
  NAND2_X1 U9764 ( .A1(n11109), .A2(n11108), .ZN(n16718) );
  INV_X1 U9765 ( .A(n16718), .ZN(n8188) );
  NAND2_X1 U9766 ( .A1(n11144), .A2(n11143), .ZN(n16123) );
  INV_X1 U9767 ( .A(n16123), .ZN(n8184) );
  AND2_X1 U9768 ( .A1(n8181), .A2(n16571), .ZN(n7628) );
  OAI21_X1 U9769 ( .B1(n8248), .B2(n7811), .A(n7803), .ZN(n7810) );
  NAND2_X1 U9770 ( .A1(n9068), .A2(n9067), .ZN(n13261) );
  NOR2_X1 U9771 ( .A1(n12363), .A2(n8274), .ZN(n7629) );
  INV_X1 U9772 ( .A(n7669), .ZN(n12983) );
  NOR2_X1 U9773 ( .A1(n12926), .A2(n13052), .ZN(n7669) );
  INV_X1 U9774 ( .A(n8564), .ZN(n8563) );
  NOR2_X1 U9775 ( .A1(n9148), .A2(n8565), .ZN(n8564) );
  INV_X1 U9776 ( .A(n7667), .ZN(n13129) );
  NAND2_X1 U9777 ( .A1(n7669), .A2(n7668), .ZN(n7667) );
  INV_X1 U9778 ( .A(n8253), .ZN(n8252) );
  NOR2_X1 U9779 ( .A1(n9085), .A2(n8254), .ZN(n8253) );
  AND2_X1 U9780 ( .A1(n7918), .A2(n7917), .ZN(n7630) );
  INV_X1 U9781 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7662) );
  XNOR2_X1 U9782 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n7631)
         );
  AND2_X1 U9783 ( .A1(n13014), .A2(n8733), .ZN(n7632) );
  AND2_X1 U9784 ( .A1(n7888), .A2(n8380), .ZN(n7633) );
  NAND2_X1 U9785 ( .A1(n10459), .A2(n10439), .ZN(n7634) );
  NOR2_X1 U9786 ( .A1(n10936), .A2(n10935), .ZN(n7635) );
  AND2_X1 U9787 ( .A1(n8336), .A2(n11309), .ZN(n10896) );
  INV_X1 U9788 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12878) );
  INV_X1 U9789 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13434) );
  AND2_X1 U9790 ( .A1(n13436), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7636) );
  INV_X1 U9791 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8554) );
  AND2_X1 U9792 ( .A1(n8752), .A2(n7452), .ZN(n7637) );
  INV_X1 U9793 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U9794 ( .A1(n14357), .A2(n14512), .ZN(n14451) );
  INV_X1 U9795 ( .A(n14451), .ZN(n14455) );
  AND2_X1 U9796 ( .A1(n10906), .A2(n10905), .ZN(n14603) );
  AND2_X1 U9797 ( .A1(n8010), .A2(n12375), .ZN(n7638) );
  OR2_X1 U9798 ( .A1(n16180), .A2(n13849), .ZN(n10815) );
  INV_X1 U9799 ( .A(n10926), .ZN(n8334) );
  INV_X1 U9800 ( .A(n9294), .ZN(n7775) );
  NAND2_X1 U9801 ( .A1(n10125), .A2(n10124), .ZN(n13191) );
  INV_X1 U9802 ( .A(n13191), .ZN(n7668) );
  INV_X1 U9803 ( .A(n11715), .ZN(n8283) );
  INV_X1 U9804 ( .A(n16520), .ZN(n15546) );
  OR2_X1 U9805 ( .A1(n11805), .A2(n8265), .ZN(n7639) );
  XNOR2_X1 U9806 ( .A(n12026), .B(keyinput_73), .ZN(n7640) );
  OR2_X1 U9807 ( .A1(n10937), .A2(n16163), .ZN(n7641) );
  INV_X1 U9808 ( .A(SI_24_), .ZN(n13307) );
  INV_X1 U9809 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15623) );
  NAND2_X2 U9810 ( .A1(n10659), .A2(n10658), .ZN(n10700) );
  OR2_X1 U9811 ( .A1(n9405), .A2(n9404), .ZN(n7642) );
  INV_X1 U9812 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10610) );
  INV_X1 U9813 ( .A(n14553), .ZN(n7899) );
  NAND2_X1 U9814 ( .A1(n9217), .A2(n9337), .ZN(n14605) );
  INV_X1 U9815 ( .A(n14605), .ZN(n14500) );
  AND3_X1 U9816 ( .A1(n9794), .A2(n7553), .A3(n9793), .ZN(n15604) );
  INV_X1 U9817 ( .A(n9797), .ZN(n13918) );
  OR2_X1 U9818 ( .A1(keyinput_87), .A2(P3_DATAO_REG_9__SCAN_IN), .ZN(n7643) );
  AND3_X1 U9819 ( .A1(n9781), .A2(n9779), .A3(n9780), .ZN(n7644) );
  INV_X1 U9820 ( .A(SI_9_), .ZN(n8112) );
  INV_X1 U9821 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8115) );
  INV_X1 U9822 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8590) );
  INV_X1 U9823 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U9824 ( .A1(n10901), .A2(n11601), .ZN(n8326) );
  AOI21_X1 U9825 ( .B1(n11601), .B2(n10918), .A(n10917), .ZN(n14563) );
  INV_X1 U9826 ( .A(n11601), .ZN(n7904) );
  NAND2_X1 U9827 ( .A1(n10349), .A2(n10348), .ZN(n10354) );
  OAI21_X1 U9828 ( .B1(n10017), .B2(n8642), .A(n8829), .ZN(n8641) );
  AOI21_X1 U9829 ( .B1(n8640), .B2(n8642), .A(n8638), .ZN(n8637) );
  OAI22_X2 U9830 ( .A1(n13661), .A2(n8166), .B1(n13662), .B2(n8165), .ZN(
        n13666) );
  OAI21_X1 U9831 ( .B1(n7503), .B2(n7645), .A(n8140), .ZN(n8139) );
  NAND2_X1 U9832 ( .A1(n13759), .A2(n7578), .ZN(n7645) );
  BUF_X4 U9833 ( .A(n13583), .Z(n13771) );
  NAND2_X1 U9834 ( .A1(n8157), .A2(n8778), .ZN(n13640) );
  NAND2_X1 U9835 ( .A1(n8760), .A2(n8759), .ZN(n13724) );
  NAND2_X1 U9836 ( .A1(n8763), .A2(n7568), .ZN(n13755) );
  NAND2_X1 U9837 ( .A1(n13688), .A2(n13687), .ZN(n13691) );
  NAND2_X1 U9838 ( .A1(n8134), .A2(n8133), .ZN(n13679) );
  NAND2_X1 U9839 ( .A1(n8768), .A2(n8766), .ZN(n13816) );
  NAND2_X1 U9840 ( .A1(n8164), .A2(n8163), .ZN(n8162) );
  OAI21_X1 U9841 ( .B1(n13825), .B2(n13824), .A(n13823), .ZN(n13914) );
  OAI21_X4 U9842 ( .B1(n15363), .B2(n15211), .A(n15213), .ZN(n15347) );
  AOI21_X2 U9843 ( .B1(n15290), .B2(n15289), .A(n7646), .ZN(n15275) );
  NAND2_X1 U9844 ( .A1(n13125), .A2(n13237), .ZN(n13231) );
  NAND2_X1 U9845 ( .A1(n15404), .A2(n15204), .ZN(n7883) );
  NAND2_X1 U9846 ( .A1(n13347), .A2(n13346), .ZN(n7872) );
  OAI22_X1 U9847 ( .A1(n12617), .A2(n12616), .B1(n12615), .B2(n15091), .ZN(
        n12637) );
  NAND2_X2 U9848 ( .A1(n15190), .A2(n15189), .ZN(n15305) );
  NAND2_X2 U9849 ( .A1(n15383), .A2(n15382), .ZN(n15381) );
  NAND2_X1 U9850 ( .A1(n12981), .A2(n12980), .ZN(n13120) );
  NAND2_X1 U9851 ( .A1(n8278), .A2(n13121), .ZN(n13239) );
  NAND2_X1 U9852 ( .A1(n8277), .A2(n12614), .ZN(n12914) );
  NAND2_X1 U9853 ( .A1(n7649), .A2(n9831), .ZN(n7659) );
  NOR2_X2 U9854 ( .A1(n9787), .A2(n7659), .ZN(n9794) );
  NAND4_X1 U9855 ( .A1(n7652), .A2(n7656), .A3(n7437), .A4(n7651), .ZN(n9829)
         );
  NAND3_X1 U9856 ( .A1(n7653), .A2(n7663), .A3(n7533), .ZN(n9809) );
  AND2_X1 U9857 ( .A1(n7662), .A2(n9813), .ZN(n7657) );
  INV_X1 U9858 ( .A(n9794), .ZN(n10149) );
  NOR2_X2 U9859 ( .A1(n15231), .A2(n15467), .ZN(n15166) );
  NOR2_X2 U9860 ( .A1(n15263), .A2(n15474), .ZN(n15246) );
  NOR2_X2 U9861 ( .A1(n12303), .A2(n12488), .ZN(n12495) );
  NOR2_X2 U9862 ( .A1(n7667), .A2(n13274), .ZN(n13234) );
  NOR2_X2 U9863 ( .A1(n15312), .A2(n15299), .ZN(n15295) );
  AND2_X2 U9864 ( .A1(n15384), .A2(n15585), .ZN(n15372) );
  AND2_X2 U9865 ( .A1(n15407), .A2(n15590), .ZN(n15384) );
  NAND2_X1 U9866 ( .A1(n15040), .A2(n14090), .ZN(n7673) );
  NAND2_X1 U9867 ( .A1(n8533), .A2(n7676), .ZN(n7675) );
  NAND3_X1 U9868 ( .A1(n7680), .A2(n7678), .A3(n13080), .ZN(n13176) );
  OAI21_X1 U9869 ( .B1(n9994), .B2(n7686), .A(n10017), .ZN(n7685) );
  NAND2_X1 U9870 ( .A1(n14977), .A2(n7689), .ZN(n7688) );
  NAND2_X1 U9871 ( .A1(n7694), .A2(n7691), .ZN(P2_U3212) );
  INV_X1 U9872 ( .A(n7692), .ZN(n7691) );
  NAND2_X1 U9873 ( .A1(n15006), .A2(n8218), .ZN(n15078) );
  OR2_X1 U9874 ( .A1(n15082), .A2(n15081), .ZN(n7694) );
  INV_X1 U9875 ( .A(n10901), .ZN(n7696) );
  INV_X1 U9876 ( .A(n14535), .ZN(n7697) );
  AOI21_X1 U9877 ( .B1(n7700), .B2(n7705), .A(n7701), .ZN(n7703) );
  INV_X1 U9878 ( .A(n12388), .ZN(n7700) );
  NAND2_X1 U9879 ( .A1(n7702), .A2(n7705), .ZN(n7706) );
  NAND2_X1 U9880 ( .A1(n12388), .A2(n10888), .ZN(n7702) );
  NAND2_X1 U9881 ( .A1(n12388), .A2(n7709), .ZN(n7708) );
  AOI21_X1 U9882 ( .B1(n7705), .B2(n7710), .A(n9018), .ZN(n7704) );
  NAND2_X1 U9883 ( .A1(n12388), .A2(n10888), .ZN(n7707) );
  INV_X1 U9884 ( .A(n10888), .ZN(n7710) );
  OAI21_X1 U9885 ( .B1(n14581), .B2(n8335), .A(n8333), .ZN(n14599) );
  NAND2_X1 U9886 ( .A1(n7719), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7718) );
  INV_X1 U9887 ( .A(n10896), .ZN(n7717) );
  NAND2_X1 U9888 ( .A1(n8623), .A2(n7727), .ZN(n7724) );
  NAND2_X1 U9889 ( .A1(n7724), .A2(n7725), .ZN(n13313) );
  NAND2_X1 U9890 ( .A1(n8605), .A2(n7732), .ZN(n7729) );
  NAND2_X1 U9891 ( .A1(n7729), .A2(n7730), .ZN(n14224) );
  NAND2_X1 U9892 ( .A1(n14276), .A2(n7737), .ZN(n7736) );
  NAND3_X1 U9893 ( .A1(n7438), .A2(n8366), .A3(n8616), .ZN(n9165) );
  NAND2_X1 U9894 ( .A1(n8977), .A2(n8975), .ZN(n8870) );
  NAND2_X1 U9895 ( .A1(n7483), .A2(n8951), .ZN(n7760) );
  NAND2_X1 U9896 ( .A1(n8887), .A2(n7762), .ZN(n7761) );
  NAND2_X1 U9897 ( .A1(n7761), .A2(n8560), .ZN(n8891) );
  NAND2_X1 U9898 ( .A1(n9009), .A2(n7476), .ZN(n7766) );
  AND2_X2 U9899 ( .A1(n14336), .A2(n14687), .ZN(n14492) );
  NOR2_X2 U9900 ( .A1(n7778), .A2(n7777), .ZN(n14336) );
  NAND2_X1 U9901 ( .A1(n14650), .A2(n14330), .ZN(n14635) );
  NAND2_X1 U9902 ( .A1(n13539), .A2(n7786), .ZN(n7785) );
  NAND2_X1 U9903 ( .A1(n7785), .A2(n7787), .ZN(n14771) );
  NAND2_X1 U9904 ( .A1(n7792), .A2(n7479), .ZN(n9367) );
  NAND2_X1 U9905 ( .A1(n14713), .A2(n7793), .ZN(n7792) );
  NAND2_X1 U9906 ( .A1(n7798), .A2(n7493), .ZN(n8859) );
  NAND2_X1 U9907 ( .A1(n14764), .A2(n7461), .ZN(n7801) );
  NAND2_X1 U9908 ( .A1(n12964), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U9909 ( .A1(n7808), .A2(n7807), .ZN(n9360) );
  AOI21_X1 U9910 ( .B1(n7810), .B2(n7812), .A(n7809), .ZN(n7808) );
  OAI21_X1 U9911 ( .B1(n12964), .B2(n7812), .A(n7810), .ZN(n14823) );
  NOR2_X1 U9912 ( .A1(n14636), .A2(n14637), .ZN(n14830) );
  NAND2_X1 U9913 ( .A1(n10139), .A2(n7826), .ZN(n7823) );
  NAND2_X1 U9914 ( .A1(n7823), .A2(n7824), .ZN(n10204) );
  NAND2_X1 U9915 ( .A1(n10415), .A2(n7833), .ZN(n7832) );
  NAND2_X1 U9916 ( .A1(n10415), .A2(n10414), .ZN(n10432) );
  INV_X1 U9917 ( .A(n16409), .ZN(n7840) );
  NAND2_X1 U9918 ( .A1(n8175), .A2(n16409), .ZN(n16416) );
  NAND2_X1 U9919 ( .A1(n7840), .A2(n7846), .ZN(n7841) );
  NAND3_X1 U9920 ( .A1(n7861), .A2(n7860), .A3(n10592), .ZN(P2_U3328) );
  OAI21_X1 U9921 ( .B1(n7864), .B2(n10569), .A(n10591), .ZN(n7860) );
  OAI211_X1 U9922 ( .C1(n7864), .C2(n7863), .A(n7862), .B(n10555), .ZN(n7861)
         );
  NAND2_X1 U9923 ( .A1(n7864), .A2(n10554), .ZN(n7862) );
  INV_X1 U9924 ( .A(n10547), .ZN(n7863) );
  NAND2_X1 U9925 ( .A1(n10545), .A2(n10544), .ZN(n7864) );
  XNOR2_X1 U9926 ( .A(n7865), .B(n8176), .ZN(SUB_1596_U4) );
  INV_X1 U9927 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7868) );
  NAND3_X1 U9928 ( .A1(n8792), .A2(n8791), .A3(n7870), .ZN(n10539) );
  OAI21_X1 U9929 ( .B1(n8839), .B2(n15550), .A(n15471), .ZN(n15561) );
  AND2_X2 U9930 ( .A1(n7874), .A2(n7873), .ZN(n15471) );
  XNOR2_X1 U9931 ( .A(n15224), .B(n15223), .ZN(n7875) );
  OAI21_X2 U9932 ( .B1(n15392), .B2(n8413), .A(n8410), .ZN(n15363) );
  NAND3_X1 U9933 ( .A1(n7888), .A2(n8380), .A3(n12982), .ZN(n13124) );
  NAND3_X1 U9934 ( .A1(n7890), .A2(n8078), .A3(n7889), .ZN(P3_U3201) );
  INV_X1 U9935 ( .A(n8368), .ZN(n7903) );
  NAND3_X1 U9936 ( .A1(n7903), .A2(n7435), .A3(n7902), .ZN(n9387) );
  NAND2_X1 U9937 ( .A1(n7910), .A2(n7912), .ZN(n14516) );
  NAND2_X1 U9938 ( .A1(n12744), .A2(n7914), .ZN(n7910) );
  OAI21_X1 U9939 ( .B1(n8806), .B2(n7924), .A(n7922), .ZN(n8808) );
  OAI21_X1 U9940 ( .B1(n8805), .B2(n7924), .A(n9936), .ZN(n7923) );
  INV_X1 U9941 ( .A(n9935), .ZN(n7924) );
  OR2_X1 U9942 ( .A1(n9914), .A2(n8809), .ZN(n8805) );
  AOI22_X1 U9943 ( .A1(n9914), .A2(n8809), .B1(n7451), .B2(n7561), .ZN(n7925)
         );
  OAI21_X1 U9944 ( .B1(n10137), .B2(n7932), .A(n7930), .ZN(n10177) );
  NAND2_X1 U9945 ( .A1(n7929), .A2(n7927), .ZN(n10181) );
  NAND2_X1 U9946 ( .A1(n10137), .A2(n7930), .ZN(n7929) );
  OAI21_X1 U9947 ( .B1(n8810), .B2(n7945), .A(n7575), .ZN(n10114) );
  INV_X1 U9948 ( .A(n10113), .ZN(n7950) );
  INV_X1 U9949 ( .A(n10114), .ZN(n7951) );
  NAND2_X1 U9950 ( .A1(n9965), .A2(n7554), .ZN(n7953) );
  NAND2_X1 U9951 ( .A1(n9963), .A2(n7958), .ZN(n7954) );
  NAND3_X1 U9952 ( .A1(n7955), .A2(n7529), .A3(n7952), .ZN(n8802) );
  NAND3_X1 U9953 ( .A1(n7954), .A2(n7953), .A3(n9988), .ZN(n7952) );
  NAND3_X1 U9954 ( .A1(n7956), .A2(n7957), .A3(n9987), .ZN(n7955) );
  NAND2_X1 U9955 ( .A1(n9965), .A2(n9964), .ZN(n7956) );
  INV_X1 U9956 ( .A(n9963), .ZN(n7957) );
  NAND2_X1 U9957 ( .A1(n10628), .A2(n7959), .ZN(n16176) );
  NAND3_X1 U9958 ( .A1(n11901), .A2(n11897), .A3(n7968), .ZN(n7960) );
  NAND3_X1 U9959 ( .A1(n11901), .A2(n11897), .A3(n7552), .ZN(n7963) );
  INV_X1 U9960 ( .A(n11047), .ZN(n7967) );
  NAND2_X1 U9961 ( .A1(n11045), .A2(n11044), .ZN(n7968) );
  NAND2_X1 U9962 ( .A1(n15672), .A2(n7549), .ZN(n7969) );
  OAI211_X1 U9963 ( .C1(n15672), .C2(n7974), .A(n7970), .B(n7969), .ZN(n14022)
         );
  NAND2_X1 U9964 ( .A1(n15672), .A2(n8719), .ZN(n7976) );
  INV_X1 U9965 ( .A(n15640), .ZN(n7982) );
  NAND2_X1 U9966 ( .A1(n12894), .A2(n7992), .ZN(n7991) );
  INV_X1 U9967 ( .A(n11056), .ZN(n7995) );
  NAND2_X1 U9968 ( .A1(n8090), .A2(n8836), .ZN(n8035) );
  AND2_X1 U9969 ( .A1(n8836), .A2(n10629), .ZN(n7996) );
  NAND4_X1 U9970 ( .A1(n7996), .A2(n8090), .A3(n8032), .A4(n8033), .ZN(n10626)
         );
  INV_X1 U9971 ( .A(n10863), .ZN(n7997) );
  NOR2_X1 U9972 ( .A1(n12751), .A2(n10860), .ZN(n13056) );
  AND2_X1 U9973 ( .A1(n8267), .A2(n8266), .ZN(n14550) );
  NAND2_X1 U9974 ( .A1(n8267), .A2(n8003), .ZN(n7998) );
  OR2_X1 U9975 ( .A1(n8267), .A2(n7639), .ZN(n7999) );
  NAND2_X1 U9976 ( .A1(n8006), .A2(n12230), .ZN(n8008) );
  NAND2_X1 U9977 ( .A1(n8011), .A2(n12375), .ZN(n10851) );
  INV_X1 U9978 ( .A(n10850), .ZN(n8013) );
  NAND3_X1 U9979 ( .A1(n8014), .A2(n8015), .A3(n7623), .ZN(n10859) );
  NAND4_X1 U9980 ( .A1(n13856), .A2(n13855), .A3(n16473), .A4(n13854), .ZN(
        n13859) );
  NOR2_X2 U9981 ( .A1(n15972), .A2(n8690), .ZN(n15951) );
  AND2_X2 U9982 ( .A1(n8019), .A2(n8025), .ZN(n15972) );
  NOR2_X1 U9983 ( .A1(n8023), .A2(n8020), .ZN(n8019) );
  NAND2_X1 U9984 ( .A1(n14048), .A2(n8026), .ZN(n8020) );
  CLKBUF_X1 U9985 ( .A(n8025), .Z(n8021) );
  XNOR2_X2 U9986 ( .A(n8028), .B(n8027), .ZN(n16053) );
  AND3_X1 U9987 ( .A1(n8033), .A2(n8032), .A3(n10623), .ZN(n8031) );
  AND2_X1 U9988 ( .A1(n8090), .A2(n8836), .ZN(n8030) );
  AND2_X1 U9989 ( .A1(n10623), .A2(n7587), .ZN(n8029) );
  NAND4_X1 U9990 ( .A1(n8030), .A2(n8032), .A3(n8029), .A4(n8033), .ZN(n8034)
         );
  NAND2_X1 U9991 ( .A1(n7559), .A2(n8039), .ZN(n8036) );
  NAND2_X1 U9992 ( .A1(n8659), .A2(n8036), .ZN(n13138) );
  INV_X1 U9993 ( .A(n13637), .ZN(n8041) );
  NAND2_X1 U9994 ( .A1(n8044), .A2(n8042), .ZN(n15915) );
  OR2_X2 U9995 ( .A1(n15950), .A2(n8047), .ZN(n8044) );
  OAI21_X1 U9996 ( .B1(n11123), .B2(n11318), .A(n7487), .ZN(n8049) );
  INV_X1 U9997 ( .A(n8049), .ZN(n8051) );
  INV_X1 U9998 ( .A(n15757), .ZN(n10675) );
  NAND2_X2 U9999 ( .A1(n7544), .A2(n7446), .ZN(n15757) );
  NAND2_X1 U10000 ( .A1(n15757), .A2(n13599), .ZN(n13596) );
  NAND2_X1 U10001 ( .A1(n13596), .A2(n13593), .ZN(n13854) );
  OR2_X1 U10002 ( .A1(n8699), .A2(n7477), .ZN(n8054) );
  NAND2_X1 U10003 ( .A1(n8054), .A2(n7579), .ZN(n14053) );
  AND2_X1 U10004 ( .A1(n8699), .A2(n7432), .ZN(n15843) );
  NAND2_X1 U10005 ( .A1(n15966), .A2(n8061), .ZN(n8059) );
  OAI21_X1 U10006 ( .B1(n13500), .B2(n8070), .A(n8067), .ZN(n15990) );
  NAND2_X1 U10007 ( .A1(n8075), .A2(n8073), .ZN(n13194) );
  NAND2_X1 U10008 ( .A1(n13415), .A2(n13420), .ZN(n13500) );
  NAND2_X1 U10009 ( .A1(n15894), .A2(n8130), .ZN(n15869) );
  OAI22_X1 U10010 ( .A1(n15971), .A2(n14048), .B1(n16111), .B2(n15954), .ZN(
        n15964) );
  NAND2_X1 U10011 ( .A1(n10739), .A2(n10738), .ZN(n16570) );
  AOI21_X2 U10012 ( .B1(n13414), .B2(n13868), .A(n13413), .ZN(n13415) );
  NAND2_X1 U10013 ( .A1(n12454), .A2(n13857), .ZN(n12453) );
  NAND2_X1 U10014 ( .A1(n10676), .A2(n8716), .ZN(n11759) );
  NAND2_X1 U10015 ( .A1(n13194), .A2(n13151), .ZN(n13414) );
  NAND2_X1 U10016 ( .A1(n16610), .A2(n12882), .ZN(n12991) );
  NAND2_X1 U10017 ( .A1(n11773), .A2(n10688), .ZN(n11798) );
  NAND2_X1 U10018 ( .A1(n12453), .A2(n10709), .ZN(n11927) );
  NAND2_X1 U10019 ( .A1(n11927), .A2(n13858), .ZN(n11926) );
  OR2_X2 U10020 ( .A1(n10659), .A2(n13565), .ZN(n10679) );
  NAND2_X1 U10021 ( .A1(n10687), .A2(n10686), .ZN(n13582) );
  NAND2_X2 U10022 ( .A1(n13712), .A2(n10674), .ZN(n10937) );
  NAND2_X1 U10023 ( .A1(n11926), .A2(n10725), .ZN(n12335) );
  NAND2_X1 U10024 ( .A1(n11796), .A2(n10699), .ZN(n12454) );
  NAND2_X1 U10025 ( .A1(n9876), .A2(n10575), .ZN(n11721) );
  OAI22_X1 U10026 ( .A1(n15275), .A2(n15276), .B1(n15284), .B2(n15219), .ZN(
        n15269) );
  NAND2_X1 U10027 ( .A1(n11759), .A2(n13593), .ZN(n11774) );
  NAND2_X1 U10028 ( .A1(n12991), .A2(n12990), .ZN(n12993) );
  NAND2_X1 U10029 ( .A1(n10894), .A2(n10895), .ZN(n8336) );
  NAND2_X1 U10030 ( .A1(n10883), .A2(n12404), .ZN(n12409) );
  NAND2_X1 U10031 ( .A1(n12011), .A2(n12010), .ZN(n12009) );
  INV_X1 U10032 ( .A(n13059), .ZN(n8079) );
  NOR2_X1 U10033 ( .A1(n14536), .A2(n14537), .ZN(n14535) );
  INV_X1 U10034 ( .A(n13855), .ZN(n11777) );
  NAND3_X1 U10035 ( .A1(n14242), .A2(n14241), .A3(n8080), .ZN(P3_U3169) );
  NAND3_X1 U10036 ( .A1(n8602), .A2(n14737), .A3(n13940), .ZN(n14264) );
  NAND2_X1 U10037 ( .A1(n14081), .A2(n14984), .ZN(n15037) );
  OAI21_X1 U10038 ( .B1(n15004), .B2(n14103), .A(n15005), .ZN(n15006) );
  OAI21_X1 U10039 ( .B1(n10204), .B2(n8202), .A(n8201), .ZN(n10245) );
  NAND2_X1 U10040 ( .A1(n9967), .A2(n9966), .ZN(n9972) );
  NAND2_X1 U10041 ( .A1(n12417), .A2(n12416), .ZN(n12415) );
  NAND2_X1 U10042 ( .A1(n12415), .A2(n8753), .ZN(n8752) );
  NAND2_X1 U10043 ( .A1(n11613), .A2(n11612), .ZN(n11611) );
  AOI22_X2 U10044 ( .A1(n15680), .A2(n15681), .B1(n11138), .B2(n11137), .ZN(
        n15688) );
  NAND2_X2 U10045 ( .A1(n10784), .A2(n16170), .ZN(n13712) );
  NAND2_X1 U10046 ( .A1(n14087), .A2(n15036), .ZN(n15040) );
  NAND2_X1 U10047 ( .A1(n13483), .A2(n13482), .ZN(n13481) );
  INV_X1 U10048 ( .A(n8543), .ZN(n8542) );
  NAND2_X1 U10049 ( .A1(n14075), .A2(n14076), .ZN(n15059) );
  INV_X1 U10050 ( .A(n10245), .ZN(n10250) );
  NAND2_X1 U10051 ( .A1(n9925), .A2(n9924), .ZN(n9938) );
  NAND2_X2 U10052 ( .A1(n8088), .A2(n8085), .ZN(n13850) );
  NAND2_X1 U10053 ( .A1(n13323), .A2(n8116), .ZN(n13483) );
  NAND2_X1 U10054 ( .A1(n8898), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U10055 ( .A1(n8916), .A2(n8914), .ZN(n8899) );
  NAND2_X1 U10056 ( .A1(n8873), .A2(n8872), .ZN(n9009) );
  NAND2_X1 U10057 ( .A1(n8870), .A2(n8869), .ZN(n8993) );
  NAND2_X1 U10058 ( .A1(n11798), .A2(n11797), .ZN(n11796) );
  NAND4_X1 U10059 ( .A1(n10661), .A2(n8691), .A3(n10660), .A4(n10662), .ZN(
        n8099) );
  INV_X1 U10060 ( .A(n8716), .ZN(n11761) );
  NAND2_X1 U10061 ( .A1(n14901), .A2(n7621), .ZN(P3_U3455) );
  NAND2_X1 U10062 ( .A1(n14588), .A2(n14587), .ZN(n14589) );
  NAND2_X1 U10063 ( .A1(n12374), .A2(n10852), .ZN(n10853) );
  NAND2_X1 U10064 ( .A1(n12006), .A2(n10846), .ZN(n10847) );
  OR2_X1 U10065 ( .A1(n14532), .A2(n10866), .ZN(n10867) );
  NAND2_X1 U10066 ( .A1(n10867), .A2(n11601), .ZN(n10928) );
  AND2_X1 U10067 ( .A1(n14593), .A2(n14592), .ZN(n8102) );
  NAND2_X1 U10068 ( .A1(n8521), .A2(n7567), .ZN(n11967) );
  AOI21_X1 U10069 ( .B1(n15015), .B2(n8537), .A(n7535), .ZN(n12218) );
  NAND2_X1 U10070 ( .A1(n12325), .A2(n12324), .ZN(n12582) );
  INV_X1 U10071 ( .A(n8641), .ZN(n8640) );
  AOI21_X1 U10072 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(n10251) );
  INV_X1 U10073 ( .A(n10042), .ZN(n8643) );
  NAND2_X1 U10074 ( .A1(n8639), .A2(n8637), .ZN(n10122) );
  NAND2_X1 U10075 ( .A1(n15375), .A2(n8414), .ZN(n8413) );
  INV_X1 U10076 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10609) );
  INV_X1 U10077 ( .A(n11103), .ZN(n10615) );
  NAND2_X1 U10078 ( .A1(n12007), .A2(n12008), .ZN(n12006) );
  NOR2_X1 U10079 ( .A1(n12752), .A2(n16668), .ZN(n12751) );
  NOR2_X1 U10080 ( .A1(n14568), .A2(n10931), .ZN(n10933) );
  NAND2_X1 U10081 ( .A1(n14835), .A2(n7601), .ZN(P3_U3486) );
  NAND2_X1 U10082 ( .A1(n14905), .A2(n7622), .ZN(P3_U3454) );
  AND2_X1 U10083 ( .A1(n8808), .A2(n8807), .ZN(n9962) );
  AOI21_X1 U10084 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(n10242) );
  NAND3_X1 U10085 ( .A1(n8824), .A2(n8823), .A3(n8825), .ZN(n10222) );
  AOI21_X1 U10086 ( .B1(n10311), .B2(n7558), .A(n8812), .ZN(n10342) );
  AOI21_X1 U10087 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(n10137) );
  NAND2_X1 U10088 ( .A1(n8802), .A2(n7584), .ZN(n10036) );
  NAND2_X1 U10089 ( .A1(n12092), .A2(n12091), .ZN(n12090) );
  INV_X1 U10090 ( .A(n10626), .ZN(n10625) );
  NAND2_X1 U10091 ( .A1(n11604), .A2(n11030), .ZN(n11868) );
  NAND2_X1 U10092 ( .A1(n7492), .A2(n8529), .ZN(n8524) );
  INV_X1 U10093 ( .A(n13565), .ZN(n10658) );
  INV_X1 U10094 ( .A(n11868), .ZN(n8123) );
  OR2_X1 U10095 ( .A1(n10700), .A2(n12423), .ZN(n8158) );
  NAND2_X1 U10096 ( .A1(n8752), .A2(n8751), .ZN(n12894) );
  NAND2_X1 U10097 ( .A1(n16051), .A2(n16705), .ZN(n8129) );
  NAND2_X1 U10098 ( .A1(n13584), .A2(n8099), .ZN(n8716) );
  NAND2_X1 U10099 ( .A1(n8713), .A2(n7555), .ZN(n15894) );
  NAND2_X1 U10100 ( .A1(n9196), .A2(n9194), .ZN(n8894) );
  NAND2_X1 U10101 ( .A1(n9214), .A2(n9212), .ZN(n8552) );
  NAND2_X1 U10102 ( .A1(n10036), .A2(n10037), .ZN(n10035) );
  OAI21_X1 U10103 ( .B1(n13647), .B2(n8775), .A(n8132), .ZN(n13654) );
  NAND2_X1 U10104 ( .A1(n13645), .A2(n13644), .ZN(n13647) );
  AOI21_X1 U10105 ( .B1(n8135), .B2(n8771), .A(n7572), .ZN(n8133) );
  NAND2_X1 U10106 ( .A1(n13674), .A2(n8135), .ZN(n8134) );
  NAND2_X1 U10107 ( .A1(n8139), .A2(n7581), .ZN(n8768) );
  NAND2_X1 U10108 ( .A1(n13418), .A2(n8144), .ZN(n8146) );
  INV_X1 U10109 ( .A(n8146), .ZN(n13504) );
  OAI21_X2 U10110 ( .B1(n15901), .B2(n8667), .A(n8665), .ZN(n15872) );
  NAND2_X2 U10111 ( .A1(n15915), .A2(n8147), .ZN(n15901) );
  NAND3_X1 U10112 ( .A1(n13699), .A2(n13698), .A3(n8151), .ZN(n8150) );
  NAND2_X1 U10113 ( .A1(n8150), .A2(n7576), .ZN(n8760) );
  NAND2_X1 U10114 ( .A1(n13700), .A2(n13702), .ZN(n8152) );
  NAND2_X1 U10115 ( .A1(n8179), .A2(n8154), .ZN(n16165) );
  OAI211_X1 U10116 ( .C1(n8156), .C2(n13630), .A(n7571), .B(n8155), .ZN(n8157)
         );
  OR2_X1 U10117 ( .A1(n10677), .A2(n10668), .ZN(n8160) );
  NAND3_X1 U10118 ( .A1(n8649), .A2(n8162), .A3(n8161), .ZN(P1_U3242) );
  NAND2_X1 U10119 ( .A1(n13666), .A2(n13667), .ZN(n13665) );
  NAND2_X1 U10120 ( .A1(n16384), .A2(n8169), .ZN(n8167) );
  NAND2_X1 U10121 ( .A1(n16465), .A2(n16466), .ZN(n16464) );
  OAI21_X1 U10122 ( .B1(n16465), .B2(n16466), .A(P2_ADDR_REG_6__SCAN_IN), .ZN(
        n8174) );
  NAND3_X1 U10123 ( .A1(n8181), .A2(n13136), .A3(n16571), .ZN(n13201) );
  INV_X1 U10124 ( .A(n8192), .ZN(n15940) );
  NAND2_X1 U10125 ( .A1(n8200), .A2(n10254), .ZN(n8198) );
  INV_X1 U10126 ( .A(n8200), .ZN(n8199) );
  NAND2_X1 U10127 ( .A1(n10252), .A2(n10274), .ZN(n8200) );
  NAND2_X1 U10128 ( .A1(n15006), .A2(n8213), .ZN(n8210) );
  AND2_X1 U10129 ( .A1(n15081), .A2(n14105), .ZN(n8218) );
  MUX2_X1 U10130 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10674), .Z(n9939) );
  NAND4_X1 U10131 ( .A1(n10077), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n9787) );
  NOR2_X2 U10132 ( .A1(n11839), .A2(n11938), .ZN(n11937) );
  NOR2_X2 U10133 ( .A1(n15449), .A2(n15598), .ZN(n15426) );
  AND2_X2 U10134 ( .A1(n13358), .A2(n15197), .ZN(n15448) );
  NAND2_X1 U10135 ( .A1(n9793), .A2(n9794), .ZN(n9827) );
  NAND2_X1 U10136 ( .A1(n9870), .A2(n11277), .ZN(n10101) );
  OAI22_X1 U10137 ( .A1(n11318), .A2(n11277), .B1(n10674), .B2(n11257), .ZN(
        n8229) );
  NAND3_X1 U10138 ( .A1(n15160), .A2(n10566), .A3(n15100), .ZN(n8231) );
  XNOR2_X2 U10139 ( .A(n8232), .B(n8852), .ZN(n10837) );
  NAND3_X1 U10140 ( .A1(n14321), .A2(n8240), .A3(n8243), .ZN(n8239) );
  NAND2_X1 U10141 ( .A1(n14320), .A2(n14605), .ZN(n8243) );
  NAND2_X1 U10142 ( .A1(n14736), .A2(n8258), .ZN(n14713) );
  NAND2_X1 U10143 ( .A1(n12774), .A2(n14373), .ZN(n12836) );
  INV_X1 U10144 ( .A(n9370), .ZN(n8261) );
  NAND3_X1 U10145 ( .A1(n8616), .A2(n8617), .A3(n8367), .ZN(n8368) );
  INV_X1 U10146 ( .A(n10864), .ZN(n8268) );
  NAND2_X1 U10147 ( .A1(n12914), .A2(n12913), .ZN(n12916) );
  NAND2_X1 U10148 ( .A1(n12634), .A2(n12638), .ZN(n8277) );
  NAND2_X1 U10149 ( .A1(n13239), .A2(n13238), .ZN(n13242) );
  NAND2_X1 U10150 ( .A1(n13120), .A2(n13119), .ZN(n8278) );
  NAND2_X1 U10151 ( .A1(n11828), .A2(n11827), .ZN(n8282) );
  OAI21_X1 U10152 ( .B1(n8282), .B2(n8281), .A(n8279), .ZN(n11951) );
  AOI21_X1 U10153 ( .B1(n11935), .B2(n8280), .A(n7520), .ZN(n8279) );
  INV_X1 U10154 ( .A(n11935), .ZN(n8281) );
  NAND2_X1 U10155 ( .A1(n8284), .A2(n8283), .ZN(n11718) );
  AND2_X2 U10156 ( .A1(n8287), .A2(n8285), .ZN(n15259) );
  OR2_X2 U10157 ( .A1(n15305), .A2(n8290), .ZN(n8287) );
  NAND2_X1 U10158 ( .A1(n12486), .A2(n12485), .ZN(n12610) );
  NAND2_X1 U10159 ( .A1(n11953), .A2(n8298), .ZN(n8297) );
  INV_X1 U10160 ( .A(n15381), .ZN(n8302) );
  NAND2_X1 U10161 ( .A1(n8302), .A2(n7580), .ZN(n8306) );
  NAND2_X1 U10162 ( .A1(n8306), .A2(n8303), .ZN(n15187) );
  NAND2_X1 U10163 ( .A1(n15240), .A2(n8313), .ZN(n8312) );
  OAI211_X2 U10164 ( .C1(n15240), .C2(n15223), .A(n8314), .B(n8312), .ZN(n8839) );
  NAND2_X1 U10165 ( .A1(n15442), .A2(n8318), .ZN(n15179) );
  AND2_X1 U10166 ( .A1(n15418), .A2(n15176), .ZN(n8318) );
  INV_X1 U10167 ( .A(n8322), .ZN(n8321) );
  OR2_X1 U10168 ( .A1(n8325), .A2(n8324), .ZN(n10903) );
  INV_X1 U10169 ( .A(n8326), .ZN(n8324) );
  NAND2_X1 U10170 ( .A1(n8328), .A2(n12405), .ZN(n10883) );
  NAND2_X1 U10171 ( .A1(n10925), .A2(n8334), .ZN(n8333) );
  MUX2_X1 U10172 ( .A(n14971), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U10173 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14971), .S(n8994), .Z(n12078)
         );
  MUX2_X1 U10174 ( .A(n11997), .B(n14606), .S(P3_IR_REG_0__SCAN_IN), .Z(n12004) );
  NAND2_X1 U10175 ( .A1(n12834), .A2(n12833), .ZN(n8348) );
  OR2_X1 U10176 ( .A1(n16673), .A2(n14254), .ZN(n8354) );
  NAND2_X1 U10177 ( .A1(n9068), .A2(n7556), .ZN(n13264) );
  NAND2_X1 U10178 ( .A1(n8357), .A2(n7564), .ZN(n12960) );
  NAND2_X1 U10179 ( .A1(n9319), .A2(n8362), .ZN(n8365) );
  INV_X1 U10180 ( .A(n8365), .ZN(n14643) );
  OAI21_X1 U10181 ( .B1(n13541), .B2(n8372), .A(n8369), .ZN(n14785) );
  NAND2_X1 U10182 ( .A1(n8901), .A2(n7577), .ZN(n14950) );
  NAND2_X1 U10183 ( .A1(n15195), .A2(n15194), .ZN(n15199) );
  NAND2_X1 U10184 ( .A1(n9819), .A2(SI_1_), .ZN(n9821) );
  NAND3_X1 U10185 ( .A1(n9820), .A2(n9845), .A3(n9821), .ZN(n9848) );
  NAND3_X1 U10186 ( .A1(n8911), .A2(n8910), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n8377) );
  NAND3_X1 U10187 ( .A1(n9777), .A2(n9775), .A3(n9776), .ZN(n8379) );
  INV_X1 U10188 ( .A(n8381), .ZN(n8380) );
  OAI21_X1 U10189 ( .B1(n12619), .B2(n8383), .A(n12975), .ZN(n8381) );
  NAND2_X1 U10190 ( .A1(n15438), .A2(n8406), .ZN(n8403) );
  OAI21_X1 U10191 ( .B1(n15392), .B2(n15207), .A(n15209), .ZN(n15368) );
  NAND3_X1 U10192 ( .A1(n9725), .A2(n7643), .A3(n8474), .ZN(n8473) );
  INV_X1 U10193 ( .A(n9674), .ZN(n9675) );
  NOR2_X2 U10194 ( .A1(n16118), .A2(n16007), .ZN(n15998) );
  NOR2_X2 U10195 ( .A1(n14031), .A2(n15834), .ZN(n15820) );
  NAND3_X1 U10196 ( .A1(n8515), .A2(n7631), .A3(n8514), .ZN(n8513) );
  INV_X1 U10197 ( .A(n11808), .ZN(n8523) );
  NAND2_X1 U10198 ( .A1(n12582), .A2(n7492), .ZN(n8525) );
  INV_X2 U10199 ( .A(n11672), .ZN(n11679) );
  NAND2_X1 U10200 ( .A1(n15016), .A2(n15017), .ZN(n15015) );
  OAI21_X1 U10201 ( .B1(n13469), .B2(n8542), .A(n8539), .ZN(n14081) );
  AOI21_X1 U10202 ( .B1(n8556), .B2(n14455), .A(n14634), .ZN(n8555) );
  NAND2_X1 U10203 ( .A1(n8951), .A2(n8949), .ZN(n8571) );
  INV_X1 U10204 ( .A(n8593), .ZN(n8592) );
  INV_X1 U10205 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10206 ( .A1(n8596), .A2(n8595), .ZN(n9392) );
  INV_X1 U10207 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10208 ( .A1(n8596), .A2(n7642), .ZN(n10593) );
  NAND2_X1 U10209 ( .A1(n8597), .A2(n11545), .ZN(n11750) );
  NOR2_X1 U10210 ( .A1(n14286), .A2(n14285), .ZN(n14284) );
  OAI21_X1 U10211 ( .B1(n14286), .B2(n8613), .A(n8612), .ZN(n14175) );
  NAND2_X1 U10212 ( .A1(n10297), .A2(n8632), .ZN(n8629) );
  NAND2_X1 U10213 ( .A1(n8629), .A2(n8630), .ZN(n10346) );
  NAND2_X1 U10214 ( .A1(n10018), .A2(n8640), .ZN(n8639) );
  NAND2_X1 U10215 ( .A1(n7582), .A2(n10226), .ZN(n10227) );
  AOI21_X1 U10216 ( .B1(n13909), .B2(n13910), .A(n13908), .ZN(n8647) );
  INV_X1 U10217 ( .A(n13907), .ZN(n8648) );
  NAND2_X1 U10218 ( .A1(n13887), .A2(n13888), .ZN(n13907) );
  NAND2_X1 U10219 ( .A1(n13912), .A2(n13914), .ZN(n8649) );
  OAI21_X1 U10220 ( .B1(n10349), .B2(n8652), .A(n8650), .ZN(n10390) );
  NAND2_X1 U10221 ( .A1(n10349), .A2(n8653), .ZN(n10370) );
  NAND2_X1 U10222 ( .A1(n10771), .A2(n8655), .ZN(n12446) );
  NAND2_X1 U10223 ( .A1(n11780), .A2(n8657), .ZN(n8656) );
  NAND2_X1 U10224 ( .A1(n11780), .A2(n10770), .ZN(n11790) );
  NAND2_X1 U10225 ( .A1(n12446), .A2(n13616), .ZN(n10774) );
  NOR2_X1 U10226 ( .A1(n7589), .A2(n8663), .ZN(n12884) );
  AND2_X1 U10227 ( .A1(n16633), .A2(n13019), .ZN(n8663) );
  NAND2_X1 U10228 ( .A1(n15857), .A2(n8676), .ZN(n8673) );
  NAND2_X1 U10229 ( .A1(n8673), .A2(n8674), .ZN(n15826) );
  NAND2_X1 U10230 ( .A1(n16123), .A2(n16028), .ZN(n8688) );
  NAND2_X1 U10231 ( .A1(n11931), .A2(n10776), .ZN(n8692) );
  NAND2_X1 U10232 ( .A1(n8692), .A2(n8693), .ZN(n12336) );
  INV_X1 U10233 ( .A(n15869), .ZN(n8700) );
  NAND2_X1 U10234 ( .A1(n8699), .A2(n7563), .ZN(n15844) );
  NAND2_X1 U10235 ( .A1(n8702), .A2(n14050), .ZN(n8697) );
  NAND2_X1 U10236 ( .A1(n8700), .A2(n8702), .ZN(n8699) );
  INV_X1 U10237 ( .A(n15873), .ZN(n8703) );
  INV_X1 U10238 ( .A(n8713), .ZN(n15910) );
  NAND2_X1 U10239 ( .A1(n15704), .A2(n8724), .ZN(n8723) );
  OR2_X1 U10240 ( .A1(n11195), .A2(n11194), .ZN(n8746) );
  NAND3_X1 U10241 ( .A1(n10720), .A2(n10635), .A3(n8748), .ZN(n10644) );
  INV_X2 U10242 ( .A(n13969), .ZN(n8750) );
  NAND2_X1 U10243 ( .A1(n12415), .A2(n11052), .ZN(n12571) );
  INV_X1 U10244 ( .A(n8752), .ZN(n12570) );
  NOR2_X1 U10245 ( .A1(n12572), .A2(n8754), .ZN(n8753) );
  INV_X1 U10246 ( .A(n11052), .ZN(n8754) );
  INV_X1 U10247 ( .A(n13683), .ZN(n13686) );
  INV_X1 U10248 ( .A(n13707), .ZN(n8761) );
  INV_X1 U10249 ( .A(n13772), .ZN(n8762) );
  NAND3_X1 U10250 ( .A1(n13728), .A2(n13727), .A3(n7585), .ZN(n8763) );
  INV_X1 U10251 ( .A(n13740), .ZN(n8765) );
  INV_X1 U10252 ( .A(n13800), .ZN(n8769) );
  NAND2_X1 U10253 ( .A1(n13647), .A2(n8776), .ZN(n8774) );
  NAND3_X1 U10254 ( .A1(n8774), .A2(n8773), .A3(n13652), .ZN(n13651) );
  OR2_X1 U10255 ( .A1(n8779), .A2(n13635), .ZN(n8778) );
  OAI22_X2 U10256 ( .A1(n13691), .A2(n8780), .B1(n13690), .B2(n8781), .ZN(
        n13694) );
  INV_X1 U10257 ( .A(n13694), .ZN(n13697) );
  NAND3_X1 U10258 ( .A1(n13655), .A2(n13654), .A3(n8785), .ZN(n8782) );
  NAND2_X1 U10259 ( .A1(n8782), .A2(n8783), .ZN(n13661) );
  NAND2_X1 U10260 ( .A1(n8789), .A2(n8787), .ZN(n8793) );
  NAND2_X1 U10261 ( .A1(n8790), .A2(n8788), .ZN(n8787) );
  NOR2_X1 U10262 ( .A1(n10571), .A2(n7586), .ZN(n8788) );
  NAND2_X1 U10263 ( .A1(n10534), .A2(n10535), .ZN(n8789) );
  INV_X1 U10264 ( .A(n10011), .ZN(n8804) );
  NAND3_X1 U10265 ( .A1(n8806), .A2(n7924), .A3(n8805), .ZN(n8807) );
  INV_X1 U10266 ( .A(n9915), .ZN(n8809) );
  NAND3_X1 U10267 ( .A1(n10041), .A2(n10040), .A3(n7546), .ZN(n8810) );
  NAND2_X1 U10268 ( .A1(n10179), .A2(n7569), .ZN(n8823) );
  NAND2_X1 U10269 ( .A1(n10181), .A2(n7557), .ZN(n8824) );
  NAND4_X1 U10270 ( .A1(n9793), .A2(n9794), .A3(n9795), .A4(n9825), .ZN(n9796)
         );
  NAND2_X1 U10271 ( .A1(n14061), .A2(n14062), .ZN(n14060) );
  AND2_X1 U10272 ( .A1(n11667), .A2(n11671), .ZN(n14061) );
  NAND2_X1 U10273 ( .A1(n9376), .A2(n16666), .ZN(n9377) );
  NAND2_X1 U10274 ( .A1(n9369), .A2(n9368), .ZN(n14663) );
  INV_X1 U10275 ( .A(n9387), .ZN(n9388) );
  XNOR2_X1 U10276 ( .A(n12109), .B(n15095), .ZN(n11935) );
  NAND2_X1 U10277 ( .A1(n10605), .A2(n16727), .ZN(n9421) );
  OAI211_X1 U10278 ( .C1(n12679), .C2(n9280), .A(n9279), .B(n9278), .ZN(n14720) );
  OR2_X1 U10279 ( .A1(n12679), .A2(n8955), .ZN(n8956) );
  OR2_X1 U10280 ( .A1(n12679), .A2(n8944), .ZN(n8945) );
  AOI21_X1 U10281 ( .B1(n13528), .B2(n8830), .A(n8831), .ZN(n14253) );
  NAND2_X1 U10282 ( .A1(n9344), .A2(n9413), .ZN(n12722) );
  OR2_X1 U10283 ( .A1(n12269), .A2(n16496), .ZN(n12270) );
  NAND2_X1 U10284 ( .A1(n13939), .A2(n13938), .ZN(n13940) );
  OAI21_X1 U10285 ( .B1(n10644), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10636) );
  NAND2_X1 U10286 ( .A1(n13671), .A2(n13670), .ZN(n13674) );
  INV_X1 U10287 ( .A(n16686), .ZN(n16698) );
  OR2_X1 U10288 ( .A1(n12320), .A2(n11123), .ZN(n11127) );
  INV_X1 U10289 ( .A(n10659), .ZN(n14057) );
  NAND2_X1 U10290 ( .A1(n10539), .A2(n10538), .ZN(n10545) );
  OR2_X1 U10291 ( .A1(n9888), .A2(n9798), .ZN(n9799) );
  NAND2_X1 U10292 ( .A1(n10385), .A2(n10384), .ZN(n10386) );
  AND2_X1 U10293 ( .A1(n8862), .A2(n8861), .ZN(n8937) );
  OAI22_X2 U10294 ( .A1(n14761), .A2(n9228), .B1(n14750), .B2(n14939), .ZN(
        n14747) );
  AND2_X1 U10295 ( .A1(n10114), .A2(n10113), .ZN(n10115) );
  NAND2_X1 U10296 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  NAND2_X2 U10297 ( .A1(n12673), .A2(n14792), .ZN(n14819) );
  NAND2_X2 U10298 ( .A1(n15427), .A2(n11246), .ZN(n15429) );
  INV_X1 U10299 ( .A(n14746), .ZN(n9365) );
  NOR2_X1 U10300 ( .A1(n14112), .A2(n15077), .ZN(n8828) );
  AND2_X1 U10301 ( .A1(n10073), .A2(n10072), .ZN(n8829) );
  OR2_X1 U10302 ( .A1(n13527), .A2(n13526), .ZN(n8830) );
  AND2_X1 U10303 ( .A1(n13527), .A2(n13526), .ZN(n8831) );
  AND2_X1 U10304 ( .A1(n13431), .A2(n10515), .ZN(n8832) );
  AND2_X1 U10305 ( .A1(n10569), .A2(n11248), .ZN(n8833) );
  AND3_X1 U10306 ( .A1(n9574), .A2(n9573), .A3(n9572), .ZN(n8834) );
  AND2_X1 U10307 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8835) );
  INV_X2 U10308 ( .A(n9895), .ZN(n10674) );
  AND4_X1 U10309 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n8836) );
  NAND2_X2 U10310 ( .A1(n14035), .A2(n16036), .ZN(n16014) );
  INV_X2 U10311 ( .A(n16014), .ZN(n16642) );
  OR2_X1 U10312 ( .A1(n14043), .A2(n15742), .ZN(n8837) );
  INV_X1 U10313 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11568) );
  INV_X1 U10314 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n16366) );
  INV_X1 U10315 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16376) );
  INV_X1 U10316 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9126) );
  INV_X1 U10317 ( .A(n16523), .ZN(n15550) );
  INV_X1 U10318 ( .A(n14483), .ZN(n9133) );
  AND2_X1 U10319 ( .A1(n16503), .A2(n16676), .ZN(n14894) );
  INV_X4 U10320 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U10321 ( .A(n9343), .ZN(n9382) );
  INV_X1 U10322 ( .A(n13649), .ZN(n12994) );
  INV_X1 U10323 ( .A(n11072), .ZN(n10648) );
  INV_X1 U10324 ( .A(n13596), .ZN(n13597) );
  INV_X1 U10325 ( .A(n13593), .ZN(n13594) );
  NAND2_X1 U10326 ( .A1(n13627), .A2(n13626), .ZN(n13630) );
  OAI22_X1 U10327 ( .A1(SI_30_), .A2(keyinput_130), .B1(SI_31_), .B2(
        keyinput_129), .ZN(n9425) );
  OAI22_X1 U10328 ( .A1(SI_29_), .A2(n9429), .B1(n14960), .B2(keyinput_131), 
        .ZN(n9430) );
  INV_X1 U10329 ( .A(n9607), .ZN(n9608) );
  INV_X1 U10330 ( .A(n9612), .ZN(n9613) );
  NAND2_X1 U10331 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  INV_X1 U10332 ( .A(n9438), .ZN(n9439) );
  NAND2_X1 U10333 ( .A1(n9440), .A2(n9439), .ZN(n9445) );
  OAI22_X1 U10334 ( .A1(n12615), .A2(n7420), .B1(n12611), .B2(n10220), .ZN(
        n10037) );
  INV_X1 U10335 ( .A(keyinput_163), .ZN(n9472) );
  OAI22_X1 U10336 ( .A1(n14146), .A2(keyinput_40), .B1(n9655), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n9656) );
  INV_X1 U10337 ( .A(n9656), .ZN(n9657) );
  NAND2_X1 U10338 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  XNOR2_X1 U10339 ( .A(keyinput_52), .B(P3_REG3_REG_4__SCAN_IN), .ZN(n9671) );
  AOI21_X1 U10340 ( .B1(n9673), .B2(n9672), .A(n9671), .ZN(n9674) );
  OAI22_X1 U10341 ( .A1(n9678), .A2(n9677), .B1(P3_REG3_REG_0__SCAN_IN), .B2(
        keyinput_54), .ZN(n9679) );
  INV_X1 U10342 ( .A(n9679), .ZN(n9680) );
  INV_X1 U10343 ( .A(n9496), .ZN(n9497) );
  NAND2_X1 U10344 ( .A1(n9498), .A2(n9497), .ZN(n9503) );
  XNOR2_X1 U10345 ( .A(keyinput_71), .B(P3_DATAO_REG_25__SCAN_IN), .ZN(n9702)
         );
  AND2_X1 U10346 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  AOI21_X1 U10347 ( .B1(n9704), .B2(n9703), .A(n9702), .ZN(n9705) );
  INV_X1 U10348 ( .A(n9705), .ZN(n9706) );
  OAI22_X1 U10349 ( .A1(n12263), .A2(keyinput_200), .B1(n9519), .B2(
        P3_DATAO_REG_24__SCAN_IN), .ZN(n9520) );
  INV_X1 U10350 ( .A(n9520), .ZN(n9521) );
  NAND2_X1 U10351 ( .A1(n9522), .A2(n9521), .ZN(n9527) );
  OAI21_X1 U10352 ( .B1(keyinput_101), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n9742), 
        .ZN(n9743) );
  OAI22_X1 U10353 ( .A1(n15576), .A2(n10499), .B1(n10540), .B2(n15188), .ZN(
        n10367) );
  AND2_X1 U10354 ( .A1(n11685), .A2(n11248), .ZN(n10517) );
  INV_X1 U10355 ( .A(n12679), .ZN(n9328) );
  INV_X1 U10356 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9485) );
  AND2_X1 U10357 ( .A1(n10532), .A2(n10505), .ZN(n10506) );
  INV_X1 U10358 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10358) );
  INV_X1 U10359 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9795) );
  AND2_X1 U10360 ( .A1(n14318), .A2(n16735), .ZN(n14319) );
  NAND2_X1 U10361 ( .A1(n9246), .A2(n9485), .ZN(n9261) );
  NAND2_X1 U10362 ( .A1(n16496), .A2(n12709), .ZN(n14363) );
  INV_X1 U10363 ( .A(n14396), .ZN(n9085) );
  INV_X1 U10364 ( .A(n14474), .ZN(n9014) );
  NAND2_X1 U10365 ( .A1(n8856), .A2(n7474), .ZN(n8857) );
  INV_X1 U10366 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U10367 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  AND2_X1 U10368 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n10234) );
  INV_X1 U10369 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10105) );
  INV_X1 U10370 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9813) );
  AND2_X1 U10371 ( .A1(n13742), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n13760) );
  INV_X1 U10372 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11146) );
  NOR3_X1 U10373 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n10623) );
  OR2_X1 U10374 ( .A1(n10071), .A2(SI_9_), .ZN(n10072) );
  OAI21_X1 U10375 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9777) );
  INV_X1 U10376 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9670) );
  INV_X1 U10377 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9047) );
  OR2_X1 U10378 ( .A1(n14319), .A2(n14464), .ZN(n14320) );
  INV_X1 U10379 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12228) );
  OR2_X1 U10380 ( .A1(n14160), .A2(n14750), .ZN(n14466) );
  INV_X1 U10381 ( .A(SI_22_), .ZN(n10343) );
  NAND2_X1 U10382 ( .A1(n12468), .A2(n14500), .ZN(n16509) );
  AND3_X1 U10383 ( .A1(n14948), .A2(n14946), .A3(n10593), .ZN(n12134) );
  NAND2_X1 U10384 ( .A1(n9343), .A2(n9342), .ZN(n9413) );
  INV_X1 U10385 ( .A(n13044), .ZN(n13042) );
  OR2_X1 U10386 ( .A1(n10333), .A2(n15053), .ZN(n10359) );
  OR2_X1 U10387 ( .A1(n10419), .A2(n10418), .ZN(n10491) );
  AND2_X1 U10388 ( .A1(n13431), .A2(n11248), .ZN(n11682) );
  INV_X1 U10389 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10255) );
  INV_X1 U10390 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13750) );
  INV_X1 U10391 ( .A(n11075), .ZN(n11076) );
  INV_X1 U10392 ( .A(n10648), .ZN(n13999) );
  AND2_X1 U10393 ( .A1(n13760), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n13792) );
  INV_X1 U10394 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11128) );
  INV_X1 U10395 ( .A(n13713), .ZN(n13734) );
  OR2_X1 U10396 ( .A1(n11182), .A2(n11181), .ZN(n11184) );
  INV_X1 U10397 ( .A(n13872), .ZN(n13501) );
  INV_X1 U10398 ( .A(n16618), .ZN(n12880) );
  OR2_X1 U10399 ( .A1(n11124), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n11139) );
  AND2_X1 U10400 ( .A1(n9032), .A2(n12228), .ZN(n9048) );
  AND2_X1 U10401 ( .A1(n9171), .A2(n9662), .ZN(n9186) );
  NAND2_X1 U10402 ( .A1(n9186), .A2(n9670), .ZN(n9206) );
  INV_X1 U10403 ( .A(n14719), .ZN(n14751) );
  INV_X1 U10404 ( .A(n14780), .ZN(n14750) );
  NAND2_X1 U10405 ( .A1(n12132), .A2(n12276), .ZN(n14290) );
  OR2_X1 U10406 ( .A1(n12679), .A2(n8925), .ZN(n8926) );
  OR2_X1 U10407 ( .A1(n12135), .A2(n9785), .ZN(n10871) );
  AND2_X1 U10408 ( .A1(n10872), .A2(n10871), .ZN(n10906) );
  AND2_X1 U10409 ( .A1(n12683), .A2(n9334), .ZN(n14632) );
  INV_X1 U10410 ( .A(n14493), .ZN(n14716) );
  INV_X1 U10411 ( .A(n14156), .ZN(n14786) );
  INV_X1 U10412 ( .A(n14205), .ZN(n14805) );
  OR2_X1 U10413 ( .A1(n16663), .A2(n14504), .ZN(n12672) );
  NAND2_X1 U10414 ( .A1(n12670), .A2(n12669), .ZN(n12673) );
  NOR2_X1 U10415 ( .A1(n16663), .A2(n16509), .ZN(n12136) );
  INV_X1 U10416 ( .A(n13213), .ZN(n14397) );
  INV_X1 U10417 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9417) );
  INV_X1 U10418 ( .A(n12806), .ZN(n14475) );
  AND2_X1 U10419 ( .A1(n9375), .A2(n10596), .ZN(n16503) );
  NAND2_X1 U10420 ( .A1(n13117), .A2(n13027), .ZN(n11685) );
  AOI21_X1 U10421 ( .B1(n15474), .B2(n15080), .A(n14115), .ZN(n14116) );
  INV_X1 U10422 ( .A(n9875), .ZN(n10575) );
  INV_X1 U10423 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n15127) );
  INV_X1 U10424 ( .A(n15268), .ZN(n15261) );
  INV_X1 U10425 ( .A(n15162), .ZN(n15073) );
  INV_X1 U10426 ( .A(n10516), .ZN(n11922) );
  NAND2_X1 U10427 ( .A1(n11918), .A2(n11685), .ZN(n16520) );
  OR2_X1 U10428 ( .A1(n10166), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n10209) );
  OR2_X1 U10429 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  NAND2_X1 U10430 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NOR2_X1 U10431 ( .A1(n11184), .A2(n11209), .ZN(n11210) );
  INV_X1 U10432 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n16421) );
  NOR2_X1 U10433 ( .A1(n11208), .A2(P1_U3086), .ZN(n11218) );
  INV_X1 U10434 ( .A(n10784), .ZN(n15761) );
  INV_X1 U10435 ( .A(n15745), .ZN(n15643) );
  AND2_X1 U10436 ( .A1(n10781), .A2(n13849), .ZN(n13828) );
  INV_X1 U10437 ( .A(n15750), .ZN(n12896) );
  INV_X1 U10438 ( .A(n15955), .ZN(n16031) );
  NOR2_X1 U10439 ( .A1(n16686), .A2(n16033), .ZN(n11207) );
  INV_X1 U10440 ( .A(n16684), .ZN(n16696) );
  INV_X1 U10441 ( .A(n13611), .ZN(n16546) );
  INV_X1 U10442 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10621) );
  AND2_X1 U10443 ( .A1(n10042), .A2(n10016), .ZN(n10017) );
  INV_X1 U10444 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10620) );
  NAND2_X1 U10445 ( .A1(n12937), .A2(n12800), .ZN(n12902) );
  AND3_X1 U10446 ( .A1(n9084), .A2(n9083), .A3(n9082), .ZN(n14402) );
  INV_X1 U10447 ( .A(n14295), .ZN(n14273) );
  NAND2_X1 U10448 ( .A1(n9317), .A2(n9316), .ZN(n14674) );
  INV_X1 U10449 ( .A(n14737), .ZN(n14267) );
  OR2_X1 U10450 ( .A1(n12117), .A2(n14947), .ZN(n10875) );
  INV_X1 U10451 ( .A(n14606), .ZN(n14580) );
  NAND2_X1 U10452 ( .A1(n10870), .A2(n10871), .ZN(n14572) );
  INV_X1 U10453 ( .A(n10906), .ZN(n10876) );
  AND2_X1 U10454 ( .A1(n14350), .A2(n14343), .ZN(n14803) );
  INV_X1 U10455 ( .A(n14792), .ZN(n16508) );
  INV_X1 U10456 ( .A(n14813), .ZN(n14824) );
  AND2_X1 U10457 ( .A1(n14819), .A2(n12773), .ZN(n14758) );
  AND2_X1 U10458 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  INV_X1 U10459 ( .A(n14894), .ZN(n16666) );
  INV_X1 U10460 ( .A(n16676), .ZN(n16643) );
  AND2_X1 U10461 ( .A1(n12117), .A2(n11545), .ZN(n12135) );
  INV_X1 U10462 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9338) );
  INV_X1 U10463 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9166) );
  AND2_X1 U10464 ( .A1(n11277), .A2(P3_U3151), .ZN(n12874) );
  OR3_X1 U10465 ( .A1(n15622), .A2(n15625), .A3(n13513), .ZN(n10608) );
  AND2_X1 U10466 ( .A1(n11694), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15074) );
  AND2_X1 U10467 ( .A1(n10366), .A2(n10365), .ZN(n15188) );
  AND3_X1 U10468 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n15172) );
  INV_X1 U10469 ( .A(n12535), .ZN(n16269) );
  AND2_X1 U10470 ( .A1(n11478), .A2(n11477), .ZN(n16270) );
  AND2_X1 U10471 ( .A1(n11478), .A2(n11468), .ZN(n16257) );
  INV_X1 U10472 ( .A(n15197), .ZN(n13463) );
  INV_X1 U10473 ( .A(n15318), .ZN(n15461) );
  NAND2_X1 U10474 ( .A1(n16223), .A2(n11230), .ZN(n15427) );
  NOR2_X1 U10475 ( .A1(n16215), .A2(n11712), .ZN(n11908) );
  NAND2_X1 U10476 ( .A1(n15543), .A2(n15443), .ZN(n16523) );
  INV_X1 U10477 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10558) );
  AND2_X1 U10478 ( .A1(n10228), .A2(n10212), .ZN(n16243) );
  INV_X1 U10479 ( .A(n15626), .ZN(n15617) );
  OR2_X1 U10480 ( .A1(n15691), .A2(n16029), .ZN(n15717) );
  INV_X1 U10481 ( .A(n15729), .ZN(n16714) );
  OR2_X1 U10482 ( .A1(n10700), .A2(n15860), .ZN(n13784) );
  AND4_X1 U10483 ( .A1(n13719), .A2(n13718), .A3(n13717), .A4(n13716), .ZN(
        n15665) );
  INV_X1 U10484 ( .A(n16297), .ZN(n15807) );
  AND2_X1 U10485 ( .A1(n13387), .A2(n15761), .ZN(n15797) );
  NOR2_X1 U10486 ( .A1(n16285), .A2(n15761), .ZN(n16294) );
  INV_X1 U10487 ( .A(n16029), .ZN(n15956) );
  INV_X1 U10488 ( .A(n14025), .ZN(n15963) );
  INV_X1 U10489 ( .A(n15970), .ZN(n15948) );
  INV_X1 U10490 ( .A(n16040), .ZN(n15929) );
  INV_X1 U10491 ( .A(n16587), .ZN(n16632) );
  OAI21_X1 U10492 ( .B1(n11281), .B2(P1_D_REG_0__SCAN_IN), .A(n10813), .ZN(
        n11770) );
  INV_X1 U10493 ( .A(n16623), .ZN(n16702) );
  INV_X1 U10494 ( .A(n16705), .ZN(n16142) );
  AND2_X1 U10495 ( .A1(n10814), .A2(n11015), .ZN(n11303) );
  INV_X1 U10496 ( .A(n16174), .ZN(n12848) );
  INV_X1 U10497 ( .A(n13259), .ZN(n13335) );
  INV_X1 U10498 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n16358) );
  INV_X1 U10499 ( .A(n14292), .ZN(n14282) );
  NAND2_X1 U10500 ( .A1(n12130), .A2(n12135), .ZN(n14295) );
  INV_X1 U10501 ( .A(n14603), .ZN(n14541) );
  OR2_X1 U10502 ( .A1(n10876), .A2(n14594), .ZN(n14611) );
  AND2_X1 U10503 ( .A1(n14676), .A2(n14675), .ZN(n14842) );
  NAND2_X1 U10504 ( .A1(n16724), .A2(n16672), .ZN(n14872) );
  AND2_X2 U10505 ( .A1(n12670), .A2(n10604), .ZN(n16724) );
  INV_X1 U10506 ( .A(n16727), .ZN(n16733) );
  OR2_X1 U10507 ( .A1(n11688), .A2(n11684), .ZN(n15077) );
  INV_X1 U10508 ( .A(n10524), .ZN(n15163) );
  INV_X1 U10509 ( .A(n15188), .ZN(n15216) );
  INV_X1 U10510 ( .A(n13352), .ZN(n15085) );
  INV_X1 U10511 ( .A(n12611), .ZN(n15091) );
  INV_X2 U10512 ( .A(P2_U3947), .ZN(n15098) );
  INV_X1 U10513 ( .A(n16224), .ZN(n16278) );
  NAND2_X1 U10514 ( .A1(n15429), .A2(n13027), .ZN(n15318) );
  NAND2_X1 U10515 ( .A1(n15429), .A2(n12081), .ZN(n15435) );
  INV_X1 U10516 ( .A(n15429), .ZN(n15454) );
  INV_X1 U10517 ( .A(n15536), .ZN(n15530) );
  INV_X1 U10518 ( .A(n16526), .ZN(n16525) );
  AND2_X1 U10519 ( .A1(n11908), .A2(n16222), .ZN(n15586) );
  INV_X1 U10520 ( .A(n15342), .ZN(n15580) );
  INV_X1 U10521 ( .A(n15586), .ZN(n16527) );
  INV_X1 U10522 ( .A(n16527), .ZN(n16529) );
  OR2_X1 U10523 ( .A1(n16220), .A2(n16218), .ZN(n16219) );
  INV_X1 U10524 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n15616) );
  INV_X1 U10525 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11995) );
  INV_X1 U10526 ( .A(n16633), .ZN(n16616) );
  NAND2_X1 U10527 ( .A1(n11205), .A2(n11201), .ZN(n15729) );
  INV_X1 U10528 ( .A(n15827), .ZN(n15732) );
  INV_X1 U10529 ( .A(n15665), .ZN(n15738) );
  INV_X1 U10530 ( .A(n15797), .ZN(n16291) );
  INV_X1 U10531 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n16429) );
  OR2_X1 U10532 ( .A1(n14035), .A2(n10650), .ZN(n15825) );
  OR2_X1 U10533 ( .A1(n16642), .A2(n12432), .ZN(n16040) );
  OR2_X1 U10534 ( .A1(n16642), .A2(n13843), .ZN(n16006) );
  OR2_X1 U10535 ( .A1(n16642), .A2(n16702), .ZN(n15970) );
  OR2_X1 U10536 ( .A1(n11771), .A2(n11770), .ZN(n16707) );
  OR2_X1 U10537 ( .A1(n11771), .A2(n11574), .ZN(n16709) );
  AND2_X2 U10538 ( .A1(n11281), .A2(n11303), .ZN(n16214) );
  INV_X1 U10539 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13730) );
  INV_X1 U10540 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n12567) );
  INV_X1 U10541 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n11636) );
  NAND2_X1 U10542 ( .A1(n8230), .A2(P1_U3086), .ZN(n13259) );
  NAND2_X1 U10543 ( .A1(n9421), .A2(n9420), .ZN(P3_U3456) );
  AND2_X1 U10544 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11459), .ZN(P2_U3947) );
  OR4_X1 U10545 ( .A1(n10820), .A2(n10819), .A3(n10818), .A4(n10817), .ZN(
        P1_U3285) );
  NOR2_X1 U10546 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8983) );
  INV_X1 U10547 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U10548 ( .A1(n8983), .A2(n8984), .ZN(n9001) );
  NOR2_X1 U10549 ( .A1(n9016), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U10550 ( .A1(n9048), .A2(n9047), .ZN(n9069) );
  NAND2_X1 U10551 ( .A1(n9127), .A2(n9126), .ZN(n9140) );
  INV_X1 U10552 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9232) );
  INV_X1 U10553 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8840) );
  INV_X1 U10554 ( .A(n9310), .ZN(n8843) );
  INV_X1 U10555 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U10556 ( .A1(n8843), .A2(n8842), .ZN(n8919) );
  NAND2_X1 U10557 ( .A1(n8919), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U10558 ( .A1(n14615), .A2(n8844), .ZN(n14633) );
  INV_X1 U10559 ( .A(n9031), .ZN(n9332) );
  INV_X1 U10560 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U10561 ( .A1(n9328), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U10562 ( .A1(n9277), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8863) );
  OAI211_X1 U10563 ( .C1(n9332), .C2(n14831), .A(n8864), .B(n8863), .ZN(n8865)
         );
  INV_X1 U10564 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16172) );
  AOI22_X1 U10565 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n15620), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16172), .ZN(n8914) );
  AOI22_X1 U10566 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n15623), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8126), .ZN(n9304) );
  AOI22_X1 U10567 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n13339), .B2(n13730), .ZN(n9272) );
  AOI22_X1 U10568 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n13434), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8577), .ZN(n9256) );
  INV_X1 U10569 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U10570 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n13256), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n13704), .ZN(n9241) );
  AOI22_X1 U10571 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11568), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n8551), .ZN(n9212) );
  XNOR2_X1 U10572 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .ZN(n9194) );
  XNOR2_X1 U10573 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8932) );
  NAND2_X1 U10574 ( .A1(n8932), .A2(n8931), .ZN(n8930) );
  INV_X1 U10575 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n11257) );
  NAND2_X1 U10576 ( .A1(n11257), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U10577 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .ZN(n8949) );
  INV_X1 U10578 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U10579 ( .A1(n9822), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8867) );
  XNOR2_X1 U10580 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .ZN(n8960) );
  INV_X1 U10581 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U10582 ( .A1(n11313), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U10583 ( .A1(n8993), .A2(n8991), .ZN(n8873) );
  INV_X1 U10584 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10585 ( .A1(n8871), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8872) );
  AND2_X1 U10586 ( .A1(n11310), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U10587 ( .A1(n11280), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U10588 ( .A1(n11316), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U10589 ( .A1(n11325), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U10590 ( .A1(n8877), .A2(n8876), .ZN(n9039) );
  XNOR2_X1 U10591 ( .A(n10044), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U10592 ( .A1(n10044), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U10593 ( .A1(n11455), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U10594 ( .A1(n11542), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8882) );
  INV_X1 U10595 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n11544) );
  NAND2_X1 U10596 ( .A1(n11544), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U10597 ( .A1(n8882), .A2(n8881), .ZN(n9094) );
  XNOR2_X1 U10598 ( .A(n11636), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10599 ( .A1(n11636), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U10600 ( .A(n8885), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U10601 ( .A1(n9117), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8887) );
  INV_X1 U10602 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U10603 ( .A1(n8885), .A2(n8884), .ZN(n8886) );
  NAND2_X1 U10604 ( .A1(n11843), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8889) );
  INV_X1 U10605 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11846) );
  NAND2_X1 U10606 ( .A1(n11846), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8888) );
  XNOR2_X1 U10607 ( .A(n8568), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n9148) );
  INV_X1 U10608 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U10609 ( .A1(n12318), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U10610 ( .A1(n8891), .A2(n8890), .ZN(n9180) );
  XNOR2_X1 U10611 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .ZN(n9178) );
  NAND2_X1 U10612 ( .A1(n9180), .A2(n9178), .ZN(n8893) );
  NAND2_X1 U10613 ( .A1(n12567), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U10614 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8895), .ZN(n8896) );
  INV_X1 U10615 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U10616 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n9290), .ZN(n8898) );
  INV_X1 U10617 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16179) );
  AOI22_X1 U10618 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n15627), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16179), .ZN(n9294) );
  INV_X1 U10619 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U10620 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n15616), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n13802), .ZN(n9321) );
  INV_X1 U10621 ( .A(n9321), .ZN(n8900) );
  XNOR2_X1 U10622 ( .A(n9320), .B(n8900), .ZN(n13915) );
  INV_X1 U10623 ( .A(n8901), .ZN(n8902) );
  NAND2_X1 U10624 ( .A1(n8902), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8904) );
  XNOR2_X2 U10625 ( .A(n8904), .B(n8903), .ZN(n14510) );
  NAND2_X1 U10626 ( .A1(n13915), .A2(n8963), .ZN(n8913) );
  INV_X1 U10627 ( .A(n8914), .ZN(n8915) );
  XNOR2_X1 U10628 ( .A(n8916), .B(n8915), .ZN(n14963) );
  NAND2_X1 U10629 ( .A1(n9310), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U10630 ( .A1(n8919), .A2(n8918), .ZN(n14654) );
  NAND2_X1 U10631 ( .A1(n14654), .A2(n9326), .ZN(n8924) );
  INV_X1 U10632 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n14834) );
  NAND2_X1 U10633 ( .A1(n9328), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U10634 ( .A1(n9277), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8920) );
  OAI211_X1 U10635 ( .C1(n9332), .C2(n14834), .A(n8921), .B(n8920), .ZN(n8922)
         );
  INV_X1 U10636 ( .A(n8922), .ZN(n8923) );
  NAND2_X1 U10637 ( .A1(n8937), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U10638 ( .A1(n9277), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U10639 ( .A1(n9031), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8927) );
  INV_X1 U10640 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8925) );
  INV_X1 U10641 ( .A(SI_1_), .ZN(n11271) );
  OAI21_X1 U10642 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n11270) );
  NAND2_X1 U10643 ( .A1(n8963), .A2(n11270), .ZN(n8936) );
  INV_X1 U10644 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8934) );
  OR2_X1 U10645 ( .A1(n8994), .A2(n12166), .ZN(n8935) );
  INV_X1 U10646 ( .A(n12709), .ZN(n12352) );
  NAND2_X1 U10647 ( .A1(n12279), .A2(n12352), .ZN(n14356) );
  NAND2_X1 U10648 ( .A1(n14363), .A2(n14356), .ZN(n12707) );
  NAND2_X1 U10649 ( .A1(n8937), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U10650 ( .A1(n9277), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U10651 ( .A1(n9031), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8939) );
  INV_X1 U10652 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10879) );
  OR2_X1 U10653 ( .A1(n12679), .A2(n10879), .ZN(n8938) );
  XNOR2_X1 U10654 ( .A(n9868), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n8942) );
  MUX2_X1 U10655 ( .A(SI_0_), .B(n8942), .S(n11277), .Z(n14971) );
  NAND2_X1 U10656 ( .A1(n12707), .A2(n12711), .ZN(n12710) );
  INV_X2 U10657 ( .A(n12279), .ZN(n16496) );
  NAND2_X1 U10658 ( .A1(n16496), .A2(n12352), .ZN(n8943) );
  NAND2_X1 U10659 ( .A1(n12710), .A2(n8943), .ZN(n16493) );
  NAND2_X1 U10660 ( .A1(n8937), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U10661 ( .A1(n9277), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U10662 ( .A1(n9031), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8946) );
  INV_X1 U10663 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n8944) );
  INV_X1 U10664 ( .A(n8949), .ZN(n8950) );
  XNOR2_X1 U10665 ( .A(n8951), .B(n8950), .ZN(n11302) );
  NAND2_X1 U10666 ( .A1(n8963), .A2(n11302), .ZN(n8954) );
  OR2_X1 U10667 ( .A1(n8994), .A2(n10878), .ZN(n8953) );
  OAI211_X1 U10668 ( .C1(n9078), .C2(SI_2_), .A(n8954), .B(n8953), .ZN(n16491)
         );
  INV_X1 U10669 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U10670 ( .A1(n8937), .A2(n14146), .ZN(n8959) );
  NAND2_X1 U10671 ( .A1(n9277), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U10672 ( .A1(n9031), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8957) );
  INV_X1 U10673 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8955) );
  INV_X1 U10674 ( .A(n8960), .ZN(n8961) );
  XNOR2_X1 U10675 ( .A(n8962), .B(n8961), .ZN(n11261) );
  NAND2_X1 U10676 ( .A1(n8963), .A2(n11261), .ZN(n8968) );
  XNOR2_X1 U10677 ( .A(n8965), .B(P3_IR_REG_3__SCAN_IN), .ZN(n12161) );
  OR2_X1 U10678 ( .A1(n8994), .A2(n12161), .ZN(n8966) );
  INV_X1 U10679 ( .A(n14145), .ZN(n16530) );
  NAND2_X1 U10680 ( .A1(n14373), .A2(n14368), .ZN(n12776) );
  NAND2_X1 U10681 ( .A1(n12544), .A2(n16491), .ZN(n12777) );
  AND2_X1 U10682 ( .A1(n12776), .A2(n12777), .ZN(n8969) );
  NAND2_X1 U10683 ( .A1(n16492), .A2(n8969), .ZN(n12775) );
  NAND2_X1 U10684 ( .A1(n12556), .A2(n14145), .ZN(n8970) );
  NAND2_X1 U10685 ( .A1(n12775), .A2(n8970), .ZN(n12834) );
  NAND2_X1 U10686 ( .A1(n9031), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U10687 ( .A1(n9277), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8973) );
  OR2_X1 U10688 ( .A1(n8835), .A2(n8983), .ZN(n12841) );
  NAND2_X1 U10689 ( .A1(n8937), .A2(n12841), .ZN(n8972) );
  INV_X1 U10690 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10884) );
  OR2_X1 U10691 ( .A1(n12679), .A2(n10884), .ZN(n8971) );
  NAND4_X1 U10692 ( .A1(n8974), .A2(n8973), .A3(n8972), .A4(n8971), .ZN(n14216) );
  INV_X1 U10693 ( .A(n14216), .ZN(n12549) );
  INV_X1 U10694 ( .A(n8975), .ZN(n8976) );
  XNOR2_X1 U10695 ( .A(n8977), .B(n8976), .ZN(n11264) );
  NAND2_X1 U10696 ( .A1(n8963), .A2(n11264), .ZN(n8981) );
  OR2_X1 U10697 ( .A1(n9323), .A2(SI_4_), .ZN(n8980) );
  NAND2_X1 U10698 ( .A1(n7574), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8978) );
  OR2_X1 U10699 ( .A1(n8994), .A2(n12412), .ZN(n8979) );
  NAND2_X1 U10700 ( .A1(n12549), .A2(n12842), .ZN(n14375) );
  INV_X1 U10701 ( .A(n12842), .ZN(n16537) );
  NAND2_X1 U10702 ( .A1(n14216), .A2(n16537), .ZN(n14374) );
  NAND2_X1 U10703 ( .A1(n14375), .A2(n14374), .ZN(n12833) );
  NAND2_X1 U10704 ( .A1(n14216), .A2(n12842), .ZN(n8982) );
  NAND2_X1 U10705 ( .A1(n9031), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U10706 ( .A1(n9277), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8989) );
  OR2_X1 U10707 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  NAND2_X1 U10708 ( .A1(n9001), .A2(n8985), .ZN(n14219) );
  NAND2_X1 U10709 ( .A1(n8937), .A2(n14219), .ZN(n8988) );
  INV_X1 U10710 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8986) );
  OR2_X1 U10711 ( .A1(n12679), .A2(n8986), .ZN(n8987) );
  NAND4_X1 U10712 ( .A1(n8990), .A2(n8989), .A3(n8988), .A4(n8987), .ZN(n12933) );
  INV_X1 U10713 ( .A(n12933), .ZN(n12837) );
  INV_X1 U10714 ( .A(n8991), .ZN(n8992) );
  XNOR2_X1 U10715 ( .A(n8993), .B(n8992), .ZN(n11258) );
  NAND2_X1 U10716 ( .A1(n8963), .A2(n11258), .ZN(n8999) );
  OR2_X1 U10717 ( .A1(n9078), .A2(SI_5_), .ZN(n8998) );
  OR2_X1 U10718 ( .A1(n8995), .A2(n9386), .ZN(n8996) );
  XNOR2_X1 U10719 ( .A(n8996), .B(P3_IR_REG_5__SCAN_IN), .ZN(n12189) );
  OR2_X1 U10720 ( .A1(n9345), .A2(n12189), .ZN(n8997) );
  NAND2_X1 U10721 ( .A1(n12837), .A2(n14215), .ZN(n14379) );
  INV_X1 U10722 ( .A(n14215), .ZN(n12604) );
  NAND2_X1 U10723 ( .A1(n12933), .A2(n12604), .ZN(n14378) );
  NAND2_X1 U10724 ( .A1(n12837), .A2(n12604), .ZN(n9000) );
  NAND2_X1 U10725 ( .A1(n9031), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U10726 ( .A1(n9277), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U10727 ( .A1(n9001), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U10728 ( .A1(n9016), .A2(n9002), .ZN(n12943) );
  NAND2_X1 U10729 ( .A1(n9326), .A2(n12943), .ZN(n9005) );
  INV_X1 U10730 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9003) );
  OR2_X1 U10731 ( .A1(n12679), .A2(n9003), .ZN(n9004) );
  NAND4_X1 U10732 ( .A1(n9007), .A2(n9006), .A3(n9005), .A4(n9004), .ZN(n14217) );
  INV_X1 U10733 ( .A(n14217), .ZN(n12810) );
  XNOR2_X1 U10734 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n9008) );
  XNOR2_X1 U10735 ( .A(n9009), .B(n9008), .ZN(n11266) );
  NAND2_X1 U10736 ( .A1(n8963), .A2(n11266), .ZN(n9013) );
  NAND2_X1 U10737 ( .A1(n9010), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9011) );
  XNOR2_X1 U10738 ( .A(n9011), .B(n8367), .ZN(n11269) );
  OR2_X1 U10739 ( .A1(n9345), .A2(n11269), .ZN(n9012) );
  OAI211_X1 U10740 ( .C1(n9323), .C2(n11267), .A(n9013), .B(n9012), .ZN(n12827) );
  NAND2_X1 U10741 ( .A1(n12810), .A2(n12827), .ZN(n14383) );
  INV_X1 U10742 ( .A(n12827), .ZN(n12936) );
  NAND2_X1 U10743 ( .A1(n14217), .A2(n12936), .ZN(n14382) );
  NAND2_X1 U10744 ( .A1(n7462), .A2(n9014), .ZN(n12761) );
  NAND2_X1 U10745 ( .A1(n14217), .A2(n12827), .ZN(n9015) );
  NAND2_X1 U10746 ( .A1(n12761), .A2(n9015), .ZN(n12807) );
  NAND2_X1 U10747 ( .A1(n9031), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U10748 ( .A1(n9277), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9021) );
  AND2_X1 U10749 ( .A1(n9016), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9017) );
  OR2_X1 U10750 ( .A1(n9017), .A2(n9032), .ZN(n12814) );
  NAND2_X1 U10751 ( .A1(n9326), .A2(n12814), .ZN(n9020) );
  INV_X1 U10752 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9018) );
  OR2_X1 U10753 ( .A1(n12679), .A2(n9018), .ZN(n9019) );
  NAND4_X1 U10754 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n12963) );
  INV_X1 U10755 ( .A(n12963), .ZN(n9029) );
  XNOR2_X1 U10756 ( .A(n9024), .B(n9023), .ZN(n11299) );
  NAND2_X1 U10757 ( .A1(n8963), .A2(n11299), .ZN(n9028) );
  OR2_X1 U10758 ( .A1(n9323), .A2(SI_7_), .ZN(n9027) );
  NAND2_X1 U10759 ( .A1(n8368), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9025) );
  XNOR2_X1 U10760 ( .A(n9025), .B(P3_IR_REG_7__SCAN_IN), .ZN(n12259) );
  OR2_X1 U10761 ( .A1(n9345), .A2(n12259), .ZN(n9026) );
  NAND2_X1 U10762 ( .A1(n9029), .A2(n12815), .ZN(n14387) );
  INV_X1 U10763 ( .A(n12815), .ZN(n16562) );
  NAND2_X1 U10764 ( .A1(n12963), .A2(n16562), .ZN(n14386) );
  NAND2_X1 U10765 ( .A1(n14387), .A2(n14386), .ZN(n12806) );
  NAND2_X1 U10766 ( .A1(n12963), .A2(n12815), .ZN(n9030) );
  NAND2_X1 U10767 ( .A1(n9031), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U10768 ( .A1(n9277), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9037) );
  NOR2_X1 U10769 ( .A1(n9032), .A2(n12228), .ZN(n9033) );
  OR2_X1 U10770 ( .A1(n9048), .A2(n9033), .ZN(n12969) );
  NAND2_X1 U10771 ( .A1(n9326), .A2(n12969), .ZN(n9036) );
  INV_X1 U10772 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n9034) );
  OR2_X1 U10773 ( .A1(n12679), .A2(n9034), .ZN(n9035) );
  NAND4_X1 U10774 ( .A1(n9038), .A2(n9037), .A3(n9036), .A4(n9035), .ZN(n14391) );
  INV_X1 U10775 ( .A(SI_8_), .ZN(n11274) );
  XNOR2_X1 U10776 ( .A(n9040), .B(n9039), .ZN(n11273) );
  NAND2_X1 U10777 ( .A1(n8963), .A2(n11273), .ZN(n9044) );
  OR2_X1 U10778 ( .A1(n8368), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10779 ( .A1(n9057), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9042) );
  INV_X1 U10780 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9041) );
  XNOR2_X1 U10781 ( .A(n9042), .B(n9041), .ZN(n11276) );
  OR2_X1 U10782 ( .A1(n9345), .A2(n11276), .ZN(n9043) );
  OAI211_X1 U10783 ( .C1(n9323), .C2(n11274), .A(n9044), .B(n9043), .ZN(n12970) );
  XNOR2_X1 U10784 ( .A(n14391), .B(n12970), .ZN(n14479) );
  INV_X1 U10785 ( .A(n14479), .ZN(n9045) );
  INV_X1 U10786 ( .A(n14391), .ZN(n12907) );
  INV_X1 U10787 ( .A(n12970), .ZN(n16595) );
  NAND2_X1 U10788 ( .A1(n12907), .A2(n16595), .ZN(n9046) );
  NAND2_X1 U10789 ( .A1(n12960), .A2(n9046), .ZN(n13211) );
  NAND2_X1 U10790 ( .A1(n9277), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9054) );
  OR2_X1 U10791 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  NAND2_X1 U10792 ( .A1(n9069), .A2(n9049), .ZN(n13277) );
  NAND2_X1 U10793 ( .A1(n9326), .A2(n13277), .ZN(n9053) );
  NAND2_X1 U10794 ( .A1(n9031), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9052) );
  INV_X1 U10795 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9050) );
  OR2_X1 U10796 ( .A1(n12679), .A2(n9050), .ZN(n9051) );
  NAND4_X1 U10797 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n14398) );
  XNOR2_X1 U10798 ( .A(n9056), .B(n9055), .ZN(n11288) );
  NAND2_X1 U10799 ( .A1(n8963), .A2(n11288), .ZN(n9065) );
  OR2_X1 U10800 ( .A1(n9323), .A2(SI_9_), .ZN(n9064) );
  NOR2_X1 U10801 ( .A1(n9057), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9060) );
  NOR2_X1 U10802 ( .A1(n9060), .A2(n9386), .ZN(n9058) );
  MUX2_X1 U10803 ( .A(n9386), .B(n9058), .S(P3_IR_REG_9__SCAN_IN), .Z(n9062)
         );
  INV_X1 U10804 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U10805 ( .A1(n9060), .A2(n9059), .ZN(n9080) );
  INV_X1 U10806 ( .A(n9080), .ZN(n9061) );
  NOR2_X1 U10807 ( .A1(n9062), .A2(n9061), .ZN(n12368) );
  OR2_X1 U10808 ( .A1(n9345), .A2(n12368), .ZN(n9063) );
  NAND2_X1 U10809 ( .A1(n14398), .A2(n13213), .ZN(n9066) );
  NAND2_X1 U10810 ( .A1(n13211), .A2(n9066), .ZN(n9068) );
  INV_X1 U10811 ( .A(n14398), .ZN(n13262) );
  NAND2_X1 U10812 ( .A1(n13262), .A2(n14397), .ZN(n9067) );
  NAND2_X1 U10813 ( .A1(n9277), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U10814 ( .A1(n9031), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U10815 ( .A1(n9069), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U10816 ( .A1(n9087), .A2(n9070), .ZN(n14134) );
  NAND2_X1 U10817 ( .A1(n9326), .A2(n14134), .ZN(n9073) );
  INV_X1 U10818 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9071) );
  OR2_X1 U10819 ( .A1(n12679), .A2(n9071), .ZN(n9072) );
  NAND4_X1 U10820 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n14403) );
  XNOR2_X1 U10821 ( .A(n9077), .B(n9076), .ZN(n11295) );
  NAND2_X1 U10822 ( .A1(n8963), .A2(n11295), .ZN(n9084) );
  OR2_X1 U10823 ( .A1(n9323), .A2(SI_10_), .ZN(n9083) );
  NAND2_X1 U10824 ( .A1(n9080), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9079) );
  MUX2_X1 U10825 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9079), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n9081) );
  NAND2_X1 U10826 ( .A1(n9081), .A2(n9109), .ZN(n11297) );
  INV_X1 U10827 ( .A(n11297), .ZN(n12515) );
  OR2_X1 U10828 ( .A1(n8994), .A2(n12515), .ZN(n9082) );
  XNOR2_X1 U10829 ( .A(n14403), .B(n14402), .ZN(n14396) );
  NAND2_X1 U10830 ( .A1(n14403), .A2(n14402), .ZN(n9086) );
  NAND2_X1 U10831 ( .A1(n9277), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U10832 ( .A1(n9087), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U10833 ( .A1(n9103), .A2(n9088), .ZN(n13367) );
  NAND2_X1 U10834 ( .A1(n9326), .A2(n13367), .ZN(n9092) );
  NAND2_X1 U10835 ( .A1(n9031), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9091) );
  INV_X1 U10836 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9089) );
  OR2_X1 U10837 ( .A1(n12679), .A2(n9089), .ZN(n9090) );
  NAND4_X1 U10838 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(n14133) );
  INV_X1 U10839 ( .A(n14133), .ZN(n14815) );
  INV_X1 U10840 ( .A(n9094), .ZN(n9095) );
  XNOR2_X1 U10841 ( .A(n9096), .B(n9095), .ZN(n11308) );
  NAND2_X1 U10842 ( .A1(n8963), .A2(n11308), .ZN(n9099) );
  NAND2_X1 U10843 ( .A1(n9109), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U10844 ( .A(n9097), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12756) );
  OR2_X1 U10845 ( .A1(n9345), .A2(n12756), .ZN(n9098) );
  OAI211_X1 U10846 ( .C1(n9323), .C2(SI_11_), .A(n9099), .B(n9098), .ZN(n16664) );
  NAND2_X1 U10847 ( .A1(n14815), .A2(n16664), .ZN(n9100) );
  NAND2_X1 U10848 ( .A1(n13365), .A2(n9100), .ZN(n9102) );
  INV_X1 U10849 ( .A(n16664), .ZN(n13250) );
  NAND2_X1 U10850 ( .A1(n14133), .A2(n13250), .ZN(n9101) );
  NAND2_X1 U10851 ( .A1(n9031), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U10852 ( .A1(n9277), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9107) );
  AND2_X1 U10853 ( .A1(n9103), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9104) );
  OR2_X1 U10854 ( .A1(n9104), .A2(n9127), .ZN(n14820) );
  NAND2_X1 U10855 ( .A1(n9326), .A2(n14820), .ZN(n9106) );
  INV_X1 U10856 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10877) );
  OR2_X1 U10857 ( .A1(n12679), .A2(n10877), .ZN(n9105) );
  NAND4_X1 U10858 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n14254) );
  OAI21_X1 U10859 ( .B1(n9109), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9110) );
  XNOR2_X1 U10860 ( .A(n9110), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13070) );
  OAI22_X1 U10861 ( .A1(n9323), .A2(SI_12_), .B1(n13070), .B2(n9345), .ZN(
        n9111) );
  INV_X1 U10862 ( .A(n9111), .ZN(n9115) );
  XNOR2_X1 U10863 ( .A(n9113), .B(n9112), .ZN(n11320) );
  NAND2_X1 U10864 ( .A1(n11320), .A2(n8963), .ZN(n9114) );
  AND2_X1 U10865 ( .A1(n14254), .A2(n16673), .ZN(n9116) );
  XNOR2_X1 U10866 ( .A(n9117), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n11451) );
  NAND2_X1 U10867 ( .A1(n11451), .A2(n8963), .ZN(n9125) );
  OR2_X1 U10868 ( .A1(n9118), .A2(n9386), .ZN(n9120) );
  MUX2_X1 U10869 ( .A(n9120), .B(P3_IR_REG_31__SCAN_IN), .S(n9119), .Z(n9122)
         );
  NAND2_X1 U10870 ( .A1(n9122), .A2(n9121), .ZN(n14531) );
  INV_X1 U10871 ( .A(n14531), .ZN(n10839) );
  OAI22_X1 U10872 ( .A1(n9323), .A2(SI_13_), .B1(n10839), .B2(n9345), .ZN(
        n9123) );
  INV_X1 U10873 ( .A(n9123), .ZN(n9124) );
  NAND2_X1 U10874 ( .A1(n9125), .A2(n9124), .ZN(n14898) );
  NAND2_X1 U10875 ( .A1(n9031), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U10876 ( .A1(n9277), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9131) );
  OR2_X1 U10877 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U10878 ( .A1(n9140), .A2(n9128), .ZN(n14259) );
  NAND2_X1 U10879 ( .A1(n9326), .A2(n14259), .ZN(n9130) );
  INV_X1 U10880 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14522) );
  OR2_X1 U10881 ( .A1(n12679), .A2(n14522), .ZN(n9129) );
  NAND4_X1 U10882 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n14416) );
  XNOR2_X1 U10883 ( .A(n14898), .B(n14816), .ZN(n14483) );
  OR2_X1 U10884 ( .A1(n14816), .A2(n14898), .ZN(n9134) );
  NAND2_X1 U10885 ( .A1(n13449), .A2(n9134), .ZN(n13519) );
  XNOR2_X1 U10886 ( .A(n8094), .B(n7627), .ZN(n11533) );
  NAND2_X1 U10887 ( .A1(n11533), .A2(n8963), .ZN(n9139) );
  NAND2_X1 U10888 ( .A1(n9121), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9135) );
  MUX2_X1 U10889 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9135), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n9136) );
  NAND2_X1 U10890 ( .A1(n9136), .A2(n9165), .ZN(n11534) );
  INV_X1 U10891 ( .A(n11534), .ZN(n14547) );
  OAI22_X1 U10892 ( .A1(n9323), .A2(SI_14_), .B1(n14547), .B2(n9345), .ZN(
        n9137) );
  INV_X1 U10893 ( .A(n9137), .ZN(n9138) );
  NAND2_X1 U10894 ( .A1(n9139), .A2(n9138), .ZN(n14889) );
  NAND2_X1 U10895 ( .A1(n9277), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U10896 ( .A1(n9140), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U10897 ( .A1(n9156), .A2(n9141), .ZN(n13536) );
  NAND2_X1 U10898 ( .A1(n9326), .A2(n13536), .ZN(n9145) );
  NAND2_X1 U10899 ( .A1(n9031), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9144) );
  INV_X1 U10900 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n9142) );
  OR2_X1 U10901 ( .A1(n12679), .A2(n9142), .ZN(n9143) );
  NAND4_X1 U10902 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(n13557) );
  OR2_X1 U10903 ( .A1(n14889), .A2(n13557), .ZN(n14423) );
  NAND2_X1 U10904 ( .A1(n14889), .A2(n13557), .ZN(n14422) );
  NAND2_X1 U10905 ( .A1(n14423), .A2(n14422), .ZN(n14484) );
  NAND2_X1 U10906 ( .A1(n13519), .A2(n14484), .ZN(n13518) );
  INV_X1 U10907 ( .A(n13557), .ZN(n14256) );
  OR2_X1 U10908 ( .A1(n14889), .A2(n14256), .ZN(n9147) );
  NAND2_X1 U10909 ( .A1(n13518), .A2(n9147), .ZN(n13541) );
  INV_X1 U10910 ( .A(n9148), .ZN(n9149) );
  XNOR2_X1 U10911 ( .A(n9150), .B(n9149), .ZN(n11600) );
  NAND2_X1 U10912 ( .A1(n11600), .A2(n8963), .ZN(n9155) );
  NAND2_X1 U10913 ( .A1(n9165), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9152) );
  XNOR2_X1 U10914 ( .A(n9152), .B(n9151), .ZN(n11601) );
  OAI22_X1 U10915 ( .A1(n9078), .A2(n11603), .B1(n9345), .B2(n11601), .ZN(
        n9153) );
  INV_X1 U10916 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U10917 ( .A1(n9277), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9162) );
  INV_X1 U10918 ( .A(n9171), .ZN(n9158) );
  NAND2_X1 U10919 ( .A1(n9156), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U10920 ( .A1(n9158), .A2(n9157), .ZN(n13556) );
  NAND2_X1 U10921 ( .A1(n9326), .A2(n13556), .ZN(n9161) );
  NAND2_X1 U10922 ( .A1(n9031), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9160) );
  INV_X1 U10923 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n10902) );
  OR2_X1 U10924 ( .A1(n12679), .A2(n10902), .ZN(n9159) );
  NAND4_X1 U10925 ( .A1(n9162), .A2(n9161), .A3(n9160), .A4(n9159), .ZN(n14205) );
  XNOR2_X1 U10926 ( .A(n14886), .B(n14805), .ZN(n13542) );
  NAND2_X1 U10927 ( .A1(n14886), .A2(n14205), .ZN(n9163) );
  XNOR2_X1 U10928 ( .A(n9164), .B(n7625), .ZN(n11751) );
  NAND2_X1 U10929 ( .A1(n11751), .A2(n8963), .ZN(n9170) );
  NAND2_X1 U10930 ( .A1(n9197), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U10931 ( .A1(n9167), .A2(n9166), .ZN(n9181) );
  OAI22_X1 U10932 ( .A1(n9323), .A2(n11753), .B1(n9345), .B2(n14553), .ZN(
        n9168) );
  INV_X1 U10933 ( .A(n9168), .ZN(n9169) );
  NAND2_X1 U10934 ( .A1(n9170), .A2(n9169), .ZN(n14882) );
  NAND2_X1 U10935 ( .A1(n9277), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U10936 ( .A1(n9031), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9176) );
  NOR2_X1 U10937 ( .A1(n9171), .A2(n9662), .ZN(n9172) );
  OR2_X1 U10938 ( .A1(n9186), .A2(n9172), .ZN(n14807) );
  NAND2_X1 U10939 ( .A1(n9326), .A2(n14807), .ZN(n9175) );
  INV_X1 U10940 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n9173) );
  OR2_X1 U10941 ( .A1(n12679), .A2(n9173), .ZN(n9174) );
  NAND4_X1 U10942 ( .A1(n9177), .A2(n9176), .A3(n9175), .A4(n9174), .ZN(n14227) );
  INV_X1 U10943 ( .A(n14227), .ZN(n14787) );
  OR2_X1 U10944 ( .A1(n14882), .A2(n14787), .ZN(n14350) );
  NAND2_X1 U10945 ( .A1(n14882), .A2(n14787), .ZN(n14343) );
  INV_X1 U10946 ( .A(n14785), .ZN(n9192) );
  INV_X1 U10947 ( .A(n9178), .ZN(n9179) );
  XNOR2_X1 U10948 ( .A(n9180), .B(n9179), .ZN(n11804) );
  NAND2_X1 U10949 ( .A1(n11804), .A2(n8963), .ZN(n9185) );
  INV_X1 U10950 ( .A(SI_17_), .ZN(n11807) );
  NAND2_X1 U10951 ( .A1(n9181), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9182) );
  XNOR2_X1 U10952 ( .A(n9182), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14579) );
  OAI22_X1 U10953 ( .A1(n9323), .A2(n11807), .B1(n8994), .B2(n11805), .ZN(
        n9183) );
  INV_X1 U10954 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U10955 ( .A1(n9277), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9191) );
  OR2_X1 U10956 ( .A1(n9186), .A2(n9670), .ZN(n9187) );
  NAND2_X1 U10957 ( .A1(n9206), .A2(n9187), .ZN(n14791) );
  NAND2_X1 U10958 ( .A1(n9326), .A2(n14791), .ZN(n9190) );
  NAND2_X1 U10959 ( .A1(n9031), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9189) );
  INV_X1 U10960 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14794) );
  OR2_X1 U10961 ( .A1(n12679), .A2(n14794), .ZN(n9188) );
  NAND4_X1 U10962 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(n14778) );
  XNOR2_X1 U10963 ( .A(n14796), .B(n14778), .ZN(n14797) );
  NAND2_X1 U10964 ( .A1(n14796), .A2(n14778), .ZN(n9193) );
  INV_X1 U10965 ( .A(n9194), .ZN(n9195) );
  XNOR2_X1 U10966 ( .A(n9196), .B(n9195), .ZN(n11894) );
  NAND2_X1 U10967 ( .A1(n11894), .A2(n8963), .ZN(n9205) );
  NOR2_X1 U10968 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), 
        .ZN(n9198) );
  NAND2_X1 U10969 ( .A1(n9200), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9199) );
  MUX2_X1 U10970 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9199), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n9202) );
  NAND2_X1 U10971 ( .A1(n9202), .A2(n9216), .ZN(n14590) );
  OAI22_X1 U10972 ( .A1(n9078), .A2(n11896), .B1(n9345), .B2(n14590), .ZN(
        n9203) );
  INV_X1 U10973 ( .A(n9203), .ZN(n9204) );
  NAND2_X1 U10974 ( .A1(n9277), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U10975 ( .A1(n9031), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9210) );
  NAND2_X1 U10976 ( .A1(n9206), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U10977 ( .A1(n9221), .A2(n9207), .ZN(n14772) );
  NAND2_X1 U10978 ( .A1(n9326), .A2(n14772), .ZN(n9209) );
  INV_X1 U10979 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n14774) );
  OR2_X1 U10980 ( .A1(n12679), .A2(n14774), .ZN(n9208) );
  NAND4_X1 U10981 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n14156) );
  OR2_X1 U10982 ( .A1(n14873), .A2(n14786), .ZN(n14347) );
  NAND2_X1 U10983 ( .A1(n14873), .A2(n14786), .ZN(n14346) );
  NAND2_X1 U10984 ( .A1(n14347), .A2(n14346), .ZN(n14776) );
  INV_X1 U10985 ( .A(n9212), .ZN(n9213) );
  XNOR2_X1 U10986 ( .A(n9214), .B(n9213), .ZN(n12022) );
  NAND2_X1 U10987 ( .A1(n12022), .A2(n8963), .ZN(n9220) );
  INV_X1 U10988 ( .A(SI_19_), .ZN(n12024) );
  NAND2_X1 U10989 ( .A1(n9216), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9215) );
  MUX2_X1 U10990 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9215), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n9217) );
  OAI22_X1 U10991 ( .A1(n9078), .A2(n12024), .B1(n14605), .B2(n9345), .ZN(
        n9218) );
  INV_X1 U10992 ( .A(n9218), .ZN(n9219) );
  NAND2_X1 U10993 ( .A1(n9031), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9227) );
  NAND2_X1 U10994 ( .A1(n9277), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9226) );
  AND2_X1 U10995 ( .A1(n9221), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9222) );
  OR2_X1 U10996 ( .A1(n9222), .A2(n9233), .ZN(n14766) );
  NAND2_X1 U10997 ( .A1(n9326), .A2(n14766), .ZN(n9225) );
  INV_X1 U10998 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n9223) );
  OR2_X1 U10999 ( .A1(n12679), .A2(n9223), .ZN(n9224) );
  NAND4_X1 U11000 ( .A1(n9227), .A2(n9226), .A3(n9225), .A4(n9224), .ZN(n14780) );
  NOR2_X1 U11001 ( .A1(n14160), .A2(n14780), .ZN(n9228) );
  XNOR2_X1 U11002 ( .A(n9229), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U11003 ( .A1(n12465), .A2(n8963), .ZN(n9231) );
  INV_X1 U11004 ( .A(SI_20_), .ZN(n12466) );
  NAND2_X1 U11005 ( .A1(n9031), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9239) );
  NOR2_X1 U11006 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  OR2_X1 U11007 ( .A1(n9246), .A2(n9234), .ZN(n14755) );
  NAND2_X1 U11008 ( .A1(n14755), .A2(n9326), .ZN(n9238) );
  NAND2_X1 U11009 ( .A1(n9277), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9237) );
  INV_X1 U11010 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n9235) );
  OR2_X1 U11011 ( .A1(n12679), .A2(n9235), .ZN(n9236) );
  NAND4_X1 U11012 ( .A1(n9239), .A2(n9238), .A3(n9237), .A4(n9236), .ZN(n14187) );
  NAND2_X1 U11013 ( .A1(n14934), .A2(n14187), .ZN(n14435) );
  INV_X1 U11014 ( .A(n14934), .ZN(n9240) );
  INV_X1 U11015 ( .A(n14187), .ZN(n14763) );
  NAND2_X1 U11016 ( .A1(n9240), .A2(n14763), .ZN(n14434) );
  NAND2_X1 U11017 ( .A1(n14435), .A2(n14434), .ZN(n14746) );
  NAND2_X1 U11018 ( .A1(n14747), .A2(n14746), .ZN(n14731) );
  NAND2_X1 U11019 ( .A1(n9240), .A2(n14187), .ZN(n14730) );
  INV_X1 U11020 ( .A(n14730), .ZN(n9254) );
  INV_X1 U11021 ( .A(n9241), .ZN(n9242) );
  XNOR2_X1 U11022 ( .A(n9243), .B(n9242), .ZN(n12562) );
  NAND2_X1 U11023 ( .A1(n12562), .A2(n8963), .ZN(n9245) );
  INV_X1 U11024 ( .A(SI_21_), .ZN(n12564) );
  OR2_X1 U11025 ( .A1(n9078), .A2(n12564), .ZN(n9244) );
  OR2_X1 U11026 ( .A1(n9246), .A2(n9485), .ZN(n9247) );
  NAND2_X1 U11027 ( .A1(n9261), .A2(n9247), .ZN(n14741) );
  NAND2_X1 U11028 ( .A1(n14741), .A2(n9326), .ZN(n9252) );
  NAND2_X1 U11029 ( .A1(n9031), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11030 ( .A1(n9277), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9250) );
  INV_X1 U11031 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9248) );
  OR2_X1 U11032 ( .A1(n12679), .A2(n9248), .ZN(n9249) );
  NAND4_X1 U11033 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(n14719) );
  AND2_X1 U11034 ( .A1(n14191), .A2(n14719), .ZN(n9253) );
  NOR2_X1 U11035 ( .A1(n9254), .A2(n9253), .ZN(n9255) );
  NAND2_X1 U11036 ( .A1(n14731), .A2(n9255), .ZN(n14715) );
  NAND2_X1 U11037 ( .A1(n14930), .A2(n14751), .ZN(n14714) );
  INV_X1 U11038 ( .A(n14714), .ZN(n9267) );
  INV_X1 U11039 ( .A(n9256), .ZN(n9257) );
  XNOR2_X1 U11040 ( .A(n9258), .B(n9257), .ZN(n12724) );
  NAND2_X1 U11041 ( .A1(n12724), .A2(n8963), .ZN(n9260) );
  OR2_X1 U11042 ( .A1(n9078), .A2(n10343), .ZN(n9259) );
  NAND2_X1 U11043 ( .A1(n9261), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11044 ( .A1(n9275), .A2(n9262), .ZN(n14723) );
  NAND2_X1 U11045 ( .A1(n14723), .A2(n9326), .ZN(n9265) );
  AOI22_X1 U11046 ( .A1(n9031), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n9277), .B2(
        P3_REG0_REG_22__SCAN_IN), .ZN(n9264) );
  INV_X1 U11047 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n14725) );
  OR2_X1 U11048 ( .A1(n12679), .A2(n14725), .ZN(n9263) );
  NOR2_X1 U11049 ( .A1(n14854), .A2(n14267), .ZN(n9266) );
  NOR2_X1 U11050 ( .A1(n9267), .A2(n9266), .ZN(n9268) );
  NAND2_X1 U11051 ( .A1(n14715), .A2(n9268), .ZN(n9270) );
  NAND2_X1 U11052 ( .A1(n14854), .A2(n14267), .ZN(n9269) );
  NAND2_X1 U11053 ( .A1(n9270), .A2(n9269), .ZN(n14701) );
  XNOR2_X1 U11054 ( .A(n9272), .B(n9271), .ZN(n12875) );
  NAND2_X1 U11055 ( .A1(n12875), .A2(n8963), .ZN(n9274) );
  OR2_X1 U11056 ( .A1(n9078), .A2(n9618), .ZN(n9273) );
  INV_X1 U11057 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11058 ( .A1(n9275), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11059 ( .A1(n9283), .A2(n9276), .ZN(n14707) );
  NAND2_X1 U11060 ( .A1(n14707), .A2(n9326), .ZN(n9279) );
  AOI22_X1 U11061 ( .A1(n9031), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n9277), .B2(
        P3_REG0_REG_23__SCAN_IN), .ZN(n9278) );
  XNOR2_X1 U11062 ( .A(n14323), .B(n14720), .ZN(n14700) );
  INV_X1 U11063 ( .A(n14700), .ZN(n14705) );
  NAND2_X1 U11064 ( .A1(n14323), .A2(n14720), .ZN(n9281) );
  NAND2_X1 U11065 ( .A1(n9283), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11066 ( .A1(n9309), .A2(n9284), .ZN(n14695) );
  NAND2_X1 U11067 ( .A1(n14695), .A2(n9326), .ZN(n9289) );
  INV_X1 U11068 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14847) );
  NAND2_X1 U11069 ( .A1(n9328), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11070 ( .A1(n9277), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9285) );
  OAI211_X1 U11071 ( .C1(n9332), .C2(n14847), .A(n9286), .B(n9285), .ZN(n9287)
         );
  INV_X1 U11072 ( .A(n9287), .ZN(n9288) );
  XOR2_X1 U11073 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9290), .Z(n9291) );
  XNOR2_X1 U11074 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9291), .ZN(n13305) );
  MUX2_X1 U11075 ( .A(n13305), .B(SI_24_), .S(n10674), .Z(n9292) );
  NOR2_X1 U11076 ( .A1(n14702), .A2(n14918), .ZN(n9293) );
  XNOR2_X1 U11077 ( .A(n9295), .B(n7775), .ZN(n13301) );
  NAND2_X1 U11078 ( .A1(n13301), .A2(n8963), .ZN(n9297) );
  XNOR2_X1 U11079 ( .A(n9309), .B(P3_REG3_REG_25__SCAN_IN), .ZN(n14677) );
  NAND2_X1 U11080 ( .A1(n14677), .A2(n9326), .ZN(n9303) );
  INV_X1 U11081 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11082 ( .A1(n9328), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11083 ( .A1(n9277), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9298) );
  OAI211_X1 U11084 ( .C1(n9332), .C2(n9300), .A(n9299), .B(n9298), .ZN(n9301)
         );
  INV_X1 U11085 ( .A(n9301), .ZN(n9302) );
  XNOR2_X1 U11086 ( .A(n14681), .B(n14325), .ZN(n14682) );
  INV_X1 U11087 ( .A(n9304), .ZN(n9305) );
  XNOR2_X1 U11088 ( .A(n9306), .B(n9305), .ZN(n14966) );
  NAND2_X1 U11089 ( .A1(n14966), .A2(n8963), .ZN(n9308) );
  INV_X1 U11090 ( .A(SI_26_), .ZN(n14969) );
  OAI21_X1 U11091 ( .B1(n9309), .B2(P3_REG3_REG_25__SCAN_IN), .A(
        P3_REG3_REG_26__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11092 ( .A1(n9311), .A2(n9310), .ZN(n14665) );
  NAND2_X1 U11093 ( .A1(n14665), .A2(n9326), .ZN(n9317) );
  INV_X1 U11094 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11095 ( .A1(n9031), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U11096 ( .A1(n9277), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9312) );
  OAI211_X1 U11097 ( .C1(n9314), .C2(n12679), .A(n9313), .B(n9312), .ZN(n9315)
         );
  INV_X1 U11098 ( .A(n9315), .ZN(n9316) );
  NAND2_X1 U11099 ( .A1(n14660), .A2(n9318), .ZN(n9319) );
  NAND2_X1 U11100 ( .A1(n14638), .A2(n14647), .ZN(n14445) );
  OAI21_X1 U11101 ( .B1(n14647), .B2(n14902), .A(n14628), .ZN(n9336) );
  INV_X1 U11102 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14300) );
  INV_X1 U11103 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n15610) );
  OAI22_X1 U11104 ( .A1(n14300), .A2(n15610), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14298) );
  INV_X1 U11105 ( .A(n14298), .ZN(n9322) );
  XNOR2_X1 U11106 ( .A(n14299), .B(n9322), .ZN(n14958) );
  NAND2_X1 U11107 ( .A1(n14958), .A2(n8963), .ZN(n9325) );
  OR2_X1 U11108 ( .A1(n9078), .A2(n14960), .ZN(n9324) );
  NAND2_X1 U11109 ( .A1(n9325), .A2(n9324), .ZN(n14624) );
  INV_X1 U11110 ( .A(n14615), .ZN(n9327) );
  NAND2_X1 U11111 ( .A1(n9327), .A2(n9326), .ZN(n12683) );
  INV_X1 U11112 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U11113 ( .A1(n9277), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U11114 ( .A1(n9328), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9329) );
  OAI211_X1 U11115 ( .C1(n9332), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9333)
         );
  INV_X1 U11116 ( .A(n9333), .ZN(n9334) );
  OR2_X1 U11117 ( .A1(n14624), .A2(n14632), .ZN(n14452) );
  NAND2_X1 U11118 ( .A1(n14624), .A2(n14632), .ZN(n14454) );
  NAND2_X1 U11119 ( .A1(n14452), .A2(n14454), .ZN(n14495) );
  INV_X1 U11120 ( .A(n14495), .ZN(n9335) );
  XNOR2_X1 U11121 ( .A(n9336), .B(n9335), .ZN(n9354) );
  NAND2_X1 U11122 ( .A1(n9337), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9339) );
  INV_X1 U11123 ( .A(n12468), .ZN(n9340) );
  NAND2_X1 U11124 ( .A1(n14357), .A2(n9340), .ZN(n14322) );
  NAND2_X1 U11125 ( .A1(n9382), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9341) );
  MUX2_X1 U11126 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9341), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9344) );
  NAND2_X1 U11127 ( .A1(n14500), .A2(n14512), .ZN(n9406) );
  OR2_X1 U11128 ( .A1(n14510), .A2(n10915), .ZN(n10904) );
  NAND2_X1 U11129 ( .A1(n9345), .A2(n10904), .ZN(n12276) );
  INV_X1 U11130 ( .A(n12276), .ZN(n9346) );
  INV_X1 U11131 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U11132 ( .A1(n9277), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11133 ( .A1(n9031), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9347) );
  OAI211_X1 U11134 ( .C1(n9349), .C2(n12679), .A(n9348), .B(n9347), .ZN(n9350)
         );
  INV_X1 U11135 ( .A(n9350), .ZN(n9351) );
  AND2_X1 U11136 ( .A1(n12683), .A2(n9351), .ZN(n14317) );
  INV_X1 U11137 ( .A(P3_B_REG_SCAN_IN), .ZN(n9352) );
  OAI21_X1 U11138 ( .B1(n14510), .B2(n9352), .A(n14779), .ZN(n14613) );
  OAI22_X1 U11139 ( .A1(n14647), .A2(n16495), .B1(n14317), .B2(n14613), .ZN(
        n9353) );
  NAND2_X1 U11140 ( .A1(n9355), .A2(n12078), .ZN(n12708) );
  NAND2_X1 U11141 ( .A1(n14363), .A2(n12708), .ZN(n9356) );
  NAND2_X1 U11142 ( .A1(n9356), .A2(n14356), .ZN(n16490) );
  INV_X1 U11143 ( .A(n16491), .ZN(n12267) );
  NAND2_X1 U11144 ( .A1(n12544), .A2(n12267), .ZN(n9357) );
  INV_X1 U11145 ( .A(n12776), .ZN(n14468) );
  INV_X1 U11146 ( .A(n12833), .ZN(n14470) );
  NAND2_X1 U11147 ( .A1(n12836), .A2(n14470), .ZN(n12835) );
  NAND2_X1 U11148 ( .A1(n12835), .A2(n14375), .ZN(n12593) );
  NAND2_X1 U11149 ( .A1(n12593), .A2(n14473), .ZN(n12592) );
  NAND2_X1 U11150 ( .A1(n12592), .A2(n14379), .ZN(n12760) );
  NAND2_X1 U11151 ( .A1(n12760), .A2(n14474), .ZN(n12759) );
  NAND2_X1 U11152 ( .A1(n12759), .A2(n14383), .ZN(n12809) );
  NAND2_X1 U11153 ( .A1(n12809), .A2(n14475), .ZN(n12808) );
  NAND2_X1 U11154 ( .A1(n12808), .A2(n14387), .ZN(n12965) );
  NAND2_X1 U11155 ( .A1(n12907), .A2(n12970), .ZN(n14393) );
  NOR2_X1 U11156 ( .A1(n14398), .A2(n14397), .ZN(n13209) );
  NAND2_X1 U11157 ( .A1(n14398), .A2(n14397), .ZN(n13208) );
  INV_X1 U11158 ( .A(n14403), .ZN(n9358) );
  NAND2_X1 U11159 ( .A1(n14815), .A2(n13250), .ZN(n14353) );
  NAND2_X1 U11160 ( .A1(n14133), .A2(n16664), .ZN(n14406) );
  NAND2_X1 U11161 ( .A1(n13526), .A2(n16673), .ZN(n14411) );
  INV_X1 U11162 ( .A(n16673), .ZN(n9359) );
  NAND2_X1 U11163 ( .A1(n14254), .A2(n9359), .ZN(n14410) );
  NAND2_X1 U11164 ( .A1(n9360), .A2(n14411), .ZN(n13453) );
  NAND2_X1 U11165 ( .A1(n13453), .A2(n14483), .ZN(n9361) );
  OR2_X1 U11166 ( .A1(n14898), .A2(n14416), .ZN(n14418) );
  NAND2_X1 U11167 ( .A1(n9361), .A2(n14418), .ZN(n13517) );
  INV_X1 U11168 ( .A(n14484), .ZN(n14420) );
  NAND2_X1 U11169 ( .A1(n13517), .A2(n14420), .ZN(n9362) );
  NAND2_X1 U11170 ( .A1(n9362), .A2(n14423), .ZN(n13539) );
  NAND2_X1 U11171 ( .A1(n14886), .A2(n14805), .ZN(n14426) );
  INV_X1 U11172 ( .A(n14778), .ZN(n14806) );
  INV_X1 U11173 ( .A(n14776), .ZN(n9363) );
  NAND2_X1 U11174 ( .A1(n14771), .A2(n9363), .ZN(n9364) );
  AND2_X1 U11175 ( .A1(n14160), .A2(n14750), .ZN(n14342) );
  OR2_X1 U11176 ( .A1(n14191), .A2(n14751), .ZN(n14439) );
  NAND2_X1 U11177 ( .A1(n14191), .A2(n14751), .ZN(n14438) );
  NAND2_X1 U11178 ( .A1(n14854), .A2(n14737), .ZN(n14341) );
  NOR2_X1 U11179 ( .A1(n14918), .A2(n14673), .ZN(n14332) );
  NAND2_X1 U11180 ( .A1(n14918), .A2(n14673), .ZN(n14335) );
  INV_X1 U11181 ( .A(n14335), .ZN(n9366) );
  NOR2_X1 U11182 ( .A1(n14332), .A2(n9366), .ZN(n14687) );
  NAND2_X1 U11183 ( .A1(n9367), .A2(n14335), .ZN(n14683) );
  NAND2_X1 U11184 ( .A1(n14683), .A2(n14682), .ZN(n9369) );
  OR2_X1 U11185 ( .A1(n14681), .A2(n14690), .ZN(n9368) );
  NAND2_X1 U11186 ( .A1(n14293), .A2(n14646), .ZN(n14324) );
  INV_X1 U11187 ( .A(n9371), .ZN(n14446) );
  XNOR2_X1 U11188 ( .A(n14316), .B(n14495), .ZN(n14627) );
  INV_X1 U11189 ( .A(n14627), .ZN(n9376) );
  NAND2_X1 U11190 ( .A1(n12563), .A2(n12468), .ZN(n10600) );
  XNOR2_X1 U11191 ( .A(n10600), .B(n14512), .ZN(n9373) );
  NAND2_X1 U11192 ( .A1(n12563), .A2(n14605), .ZN(n9372) );
  NAND2_X1 U11193 ( .A1(n9373), .A2(n9372), .ZN(n12127) );
  NAND2_X1 U11194 ( .A1(n12468), .A2(n14605), .ZN(n14507) );
  INV_X1 U11195 ( .A(n14507), .ZN(n10597) );
  AND2_X1 U11196 ( .A1(n16663), .A2(n10597), .ZN(n9374) );
  NAND2_X1 U11197 ( .A1(n12127), .A2(n9374), .ZN(n9375) );
  NAND2_X1 U11198 ( .A1(n14507), .A2(n9406), .ZN(n10599) );
  OR2_X1 U11199 ( .A1(n10599), .A2(n12722), .ZN(n10596) );
  OR2_X1 U11200 ( .A1(n16509), .A2(n14512), .ZN(n16676) );
  NAND2_X1 U11201 ( .A1(n14621), .A2(n9377), .ZN(n10605) );
  XNOR2_X1 U11202 ( .A(n9393), .B(P3_B_REG_SCAN_IN), .ZN(n9381) );
  NAND2_X1 U11203 ( .A1(n9381), .A2(n13304), .ZN(n9390) );
  AND2_X1 U11204 ( .A1(n9343), .A2(n9383), .ZN(n9384) );
  NOR2_X1 U11205 ( .A1(n9384), .A2(n9386), .ZN(n9385) );
  MUX2_X1 U11206 ( .A(n9386), .B(n9385), .S(P3_IR_REG_26__SCAN_IN), .Z(n9389)
         );
  INV_X1 U11207 ( .A(n9411), .ZN(n14970) );
  NAND2_X1 U11208 ( .A1(n13304), .A2(n14970), .ZN(n9391) );
  INV_X1 U11209 ( .A(n14946), .ZN(n12663) );
  NAND2_X1 U11210 ( .A1(n14970), .A2(n9393), .ZN(n9394) );
  NOR2_X1 U11211 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9399) );
  NOR4_X1 U11212 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9398) );
  NOR4_X1 U11213 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9397) );
  NOR4_X1 U11214 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9396) );
  NAND4_X1 U11215 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n9405)
         );
  NOR4_X1 U11216 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9403) );
  NOR4_X1 U11217 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9402) );
  NOR4_X1 U11218 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9401) );
  NOR4_X1 U11219 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9400) );
  NAND4_X1 U11220 ( .A1(n9403), .A2(n9402), .A3(n9401), .A4(n9400), .ZN(n9404)
         );
  NAND3_X1 U11221 ( .A1(n12663), .A2(n12266), .A3(n10593), .ZN(n12131) );
  INV_X1 U11222 ( .A(n12127), .ZN(n12120) );
  INV_X1 U11223 ( .A(n12266), .ZN(n14948) );
  INV_X1 U11224 ( .A(n12265), .ZN(n14503) );
  INV_X1 U11225 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U11226 ( .A1(n14503), .A2(n9407), .ZN(n12129) );
  OR2_X1 U11227 ( .A1(n14451), .A2(n14507), .ZN(n12123) );
  NAND2_X1 U11228 ( .A1(n12129), .A2(n12123), .ZN(n9408) );
  NAND2_X1 U11229 ( .A1(n12134), .A2(n9408), .ZN(n9409) );
  OAI21_X1 U11230 ( .B1(n12131), .B2(n12120), .A(n9409), .ZN(n9416) );
  INV_X1 U11231 ( .A(n13304), .ZN(n9412) );
  INV_X1 U11232 ( .A(n9393), .ZN(n9410) );
  NAND2_X1 U11233 ( .A1(n9413), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U11234 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9414), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9415) );
  NOR2_X1 U11235 ( .A1(n16727), .A2(n9417), .ZN(n9419) );
  INV_X1 U11236 ( .A(n14624), .ZN(n10606) );
  INV_X1 U11237 ( .A(n16663), .ZN(n16672) );
  INV_X1 U11238 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U11239 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_247), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_248), .ZN(n9422) );
  OAI221_X1 U11240 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_247), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_248), .A(n9422), .ZN(n9587) );
  INV_X1 U11241 ( .A(keyinput_246), .ZN(n9586) );
  INV_X1 U11242 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9768) );
  INV_X1 U11243 ( .A(keyinput_218), .ZN(n9543) );
  INV_X1 U11244 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n11661) );
  INV_X1 U11245 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n12038) );
  XNOR2_X1 U11246 ( .A(n12038), .B(keyinput_214), .ZN(n9541) );
  INV_X1 U11247 ( .A(keyinput_213), .ZN(n9537) );
  INV_X1 U11248 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n12036) );
  INV_X1 U11249 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n12056) );
  INV_X1 U11250 ( .A(keyinput_207), .ZN(n9531) );
  INV_X1 U11251 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n12052) );
  INV_X1 U11252 ( .A(keyinput_206), .ZN(n9530) );
  INV_X1 U11253 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n12026) );
  XNOR2_X1 U11254 ( .A(n12026), .B(keyinput_201), .ZN(n9528) );
  INV_X1 U11255 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n12193) );
  INV_X1 U11256 ( .A(keyinput_199), .ZN(n9518) );
  INV_X1 U11257 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n12380) );
  INV_X1 U11258 ( .A(keyinput_189), .ZN(n9506) );
  INV_X1 U11259 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9689) );
  INV_X1 U11260 ( .A(keyinput_188), .ZN(n9505) );
  XNOR2_X1 U11261 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n9504)
         );
  INV_X1 U11262 ( .A(keyinput_181), .ZN(n9494) );
  OAI22_X1 U11263 ( .A1(n9670), .A2(keyinput_178), .B1(keyinput_179), .B2(
        P3_REG3_REG_24__SCAN_IN), .ZN(n9423) );
  AOI221_X1 U11264 ( .B1(n9670), .B2(keyinput_178), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_179), .A(n9423), .ZN(n9491) );
  INV_X1 U11265 ( .A(keyinput_177), .ZN(n9489) );
  INV_X1 U11266 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n14166) );
  OAI22_X1 U11267 ( .A1(n14166), .A2(keyinput_170), .B1(keyinput_171), .B2(
        P3_REG3_REG_8__SCAN_IN), .ZN(n9424) );
  AOI221_X1 U11268 ( .B1(n14166), .B2(keyinput_170), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_171), .A(n9424), .ZN(n9482) );
  INV_X1 U11269 ( .A(keyinput_168), .ZN(n9480) );
  INV_X1 U11270 ( .A(keyinput_141), .ZN(n9447) );
  XNOR2_X1 U11271 ( .A(SI_24_), .B(keyinput_136), .ZN(n9446) );
  INV_X1 U11272 ( .A(keyinput_134), .ZN(n9436) );
  INV_X1 U11273 ( .A(keyinput_132), .ZN(n9433) );
  INV_X1 U11274 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9428) );
  INV_X1 U11275 ( .A(keyinput_128), .ZN(n9427) );
  AOI221_X1 U11276 ( .B1(SI_30_), .B2(keyinput_130), .C1(keyinput_129), .C2(
        SI_31_), .A(n9425), .ZN(n9426) );
  OAI221_X1 U11277 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_128), .C1(n9428), 
        .C2(n9427), .A(n9426), .ZN(n9432) );
  INV_X1 U11278 ( .A(keyinput_131), .ZN(n9429) );
  INV_X1 U11279 ( .A(keyinput_133), .ZN(n9434) );
  INV_X1 U11280 ( .A(keyinput_135), .ZN(n9437) );
  INV_X1 U11281 ( .A(SI_23_), .ZN(n9618) );
  AOI22_X1 U11282 ( .A1(n9618), .A2(keyinput_137), .B1(keyinput_139), .B2(
        n12564), .ZN(n9441) );
  OAI221_X1 U11283 ( .B1(n9618), .B2(keyinput_137), .C1(n12564), .C2(
        keyinput_139), .A(n9441), .ZN(n9444) );
  AOI22_X1 U11284 ( .A1(SI_20_), .A2(keyinput_140), .B1(SI_22_), .B2(
        keyinput_138), .ZN(n9442) );
  OAI221_X1 U11285 ( .B1(SI_20_), .B2(keyinput_140), .C1(SI_22_), .C2(
        keyinput_138), .A(n9442), .ZN(n9443) );
  AOI22_X1 U11286 ( .A1(SI_15_), .A2(keyinput_145), .B1(SI_18_), .B2(
        keyinput_142), .ZN(n9448) );
  OAI221_X1 U11287 ( .B1(SI_15_), .B2(keyinput_145), .C1(SI_18_), .C2(
        keyinput_142), .A(n9448), .ZN(n9453) );
  AOI22_X1 U11288 ( .A1(n11807), .A2(keyinput_143), .B1(keyinput_144), .B2(
        n11753), .ZN(n9449) );
  OAI221_X1 U11289 ( .B1(n11807), .B2(keyinput_143), .C1(n11753), .C2(
        keyinput_144), .A(n9449), .ZN(n9452) );
  AOI22_X1 U11290 ( .A1(n11532), .A2(keyinput_146), .B1(keyinput_147), .B2(
        n11452), .ZN(n9450) );
  OAI221_X1 U11291 ( .B1(n11532), .B2(keyinput_146), .C1(n11452), .C2(
        keyinput_147), .A(n9450), .ZN(n9451) );
  INV_X1 U11292 ( .A(SI_7_), .ZN(n11298) );
  AOI22_X1 U11293 ( .A1(SI_8_), .A2(keyinput_152), .B1(n11298), .B2(
        keyinput_153), .ZN(n9454) );
  OAI221_X1 U11294 ( .B1(SI_8_), .B2(keyinput_152), .C1(n11298), .C2(
        keyinput_153), .A(n9454), .ZN(n9455) );
  INV_X1 U11295 ( .A(n9455), .ZN(n9461) );
  AOI22_X1 U11296 ( .A1(SI_10_), .A2(keyinput_150), .B1(n11307), .B2(
        keyinput_149), .ZN(n9456) );
  OAI221_X1 U11297 ( .B1(SI_10_), .B2(keyinput_150), .C1(n11307), .C2(
        keyinput_149), .A(n9456), .ZN(n9457) );
  INV_X1 U11298 ( .A(n9457), .ZN(n9460) );
  XNOR2_X1 U11299 ( .A(SI_9_), .B(keyinput_151), .ZN(n9459) );
  XNOR2_X1 U11300 ( .A(SI_12_), .B(keyinput_148), .ZN(n9458) );
  NAND4_X1 U11301 ( .A1(n9461), .A2(n9460), .A3(n9459), .A4(n9458), .ZN(n9462)
         );
  AOI22_X1 U11302 ( .A1(SI_5_), .A2(keyinput_155), .B1(n11267), .B2(
        keyinput_154), .ZN(n9463) );
  OAI221_X1 U11303 ( .B1(SI_5_), .B2(keyinput_155), .C1(n11267), .C2(
        keyinput_154), .A(n9463), .ZN(n9464) );
  OAI22_X1 U11304 ( .A1(n9465), .A2(n9464), .B1(SI_4_), .B2(keyinput_156), 
        .ZN(n9468) );
  INV_X1 U11305 ( .A(SI_3_), .ZN(n11260) );
  OAI22_X1 U11306 ( .A1(n11260), .A2(keyinput_157), .B1(keyinput_158), .B2(
        SI_2_), .ZN(n9466) );
  AOI221_X1 U11307 ( .B1(n11260), .B2(keyinput_157), .C1(SI_2_), .C2(
        keyinput_158), .A(n9466), .ZN(n9467) );
  OAI221_X1 U11308 ( .B1(n9468), .B2(keyinput_156), .C1(n9468), .C2(SI_4_), 
        .A(n9467), .ZN(n9471) );
  OAI22_X1 U11309 ( .A1(n11271), .A2(keyinput_159), .B1(keyinput_160), .B2(
        SI_0_), .ZN(n9469) );
  AOI221_X1 U11310 ( .B1(n11271), .B2(keyinput_159), .C1(SI_0_), .C2(
        keyinput_160), .A(n9469), .ZN(n9470) );
  INV_X1 U11311 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U11312 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_161), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_162), .ZN(n9473) );
  OAI221_X1 U11313 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_161), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_162), .A(n9473), .ZN(n9474) );
  OAI22_X1 U11314 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_164), .B1(
        keyinput_166), .B2(P3_REG3_REG_23__SCAN_IN), .ZN(n9475) );
  AOI221_X1 U11315 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_164), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_166), .A(n9475), .ZN(n9476) );
  OAI21_X1 U11316 ( .B1(keyinput_167), .B2(P3_REG3_REG_10__SCAN_IN), .A(n9478), 
        .ZN(n9479) );
  OAI221_X1 U11317 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_168), .C1(
        n14146), .C2(n9480), .A(n9479), .ZN(n9481) );
  XNOR2_X1 U11318 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n9488)
         );
  INV_X1 U11319 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13058) );
  OAI22_X1 U11320 ( .A1(n9662), .A2(keyinput_176), .B1(n13058), .B2(
        keyinput_174), .ZN(n9483) );
  AOI221_X1 U11321 ( .B1(n9662), .B2(keyinput_176), .C1(keyinput_174), .C2(
        n13058), .A(n9483), .ZN(n9487) );
  OAI22_X1 U11322 ( .A1(n9485), .A2(keyinput_173), .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_175), .ZN(n9484) );
  AOI221_X1 U11323 ( .B1(n9485), .B2(keyinput_173), .C1(keyinput_175), .C2(
        P3_REG3_REG_25__SCAN_IN), .A(n9484), .ZN(n9486) );
  AOI22_X1 U11324 ( .A1(n9491), .A2(n9490), .B1(keyinput_180), .B2(
        P3_REG3_REG_4__SCAN_IN), .ZN(n9492) );
  OAI21_X1 U11325 ( .B1(keyinput_180), .B2(P3_REG3_REG_4__SCAN_IN), .A(n9492), 
        .ZN(n9493) );
  OAI221_X1 U11326 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_181), .C1(n9047), .C2(n9494), .A(n9493), .ZN(n9498) );
  INV_X1 U11327 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9678) );
  INV_X1 U11328 ( .A(keyinput_182), .ZN(n9495) );
  OAI22_X1 U11329 ( .A1(n9678), .A2(n9495), .B1(P3_REG3_REG_0__SCAN_IN), .B2(
        keyinput_182), .ZN(n9496) );
  INV_X1 U11330 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U11331 ( .A1(n12749), .A2(keyinput_186), .B1(n9126), .B2(
        keyinput_184), .ZN(n9499) );
  OAI221_X1 U11332 ( .B1(n12749), .B2(keyinput_186), .C1(n9126), .C2(
        keyinput_184), .A(n9499), .ZN(n9502) );
  AOI22_X1 U11333 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_187), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_185), .ZN(n9500) );
  OAI221_X1 U11334 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_187), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_185), .A(n9500), .ZN(n9501) );
  INV_X1 U11335 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n12685) );
  INV_X1 U11336 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U11337 ( .A1(n12685), .A2(keyinput_193), .B1(n9508), .B2(
        keyinput_190), .ZN(n9507) );
  OAI221_X1 U11338 ( .B1(n12685), .B2(keyinput_193), .C1(n9508), .C2(
        keyinput_190), .A(n9507), .ZN(n9511) );
  INV_X1 U11339 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U11340 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_192), .B1(n10908), 
        .B2(keyinput_191), .ZN(n9509) );
  OAI221_X1 U11341 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_192), .C1(n10908), 
        .C2(keyinput_191), .A(n9509), .ZN(n9510) );
  INV_X1 U11342 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n12743) );
  INV_X1 U11343 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U11344 ( .A1(n12743), .A2(keyinput_196), .B1(keyinput_195), .B2(
        n12771), .ZN(n9512) );
  OAI221_X1 U11345 ( .B1(n12743), .B2(keyinput_196), .C1(n12771), .C2(
        keyinput_195), .A(n9512), .ZN(n9515) );
  INV_X1 U11346 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n12591) );
  INV_X1 U11347 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n12470) );
  OAI22_X1 U11348 ( .A1(n12591), .A2(keyinput_197), .B1(n12470), .B2(
        keyinput_198), .ZN(n9513) );
  AOI221_X1 U11349 ( .B1(n12591), .B2(keyinput_197), .C1(keyinput_198), .C2(
        n12470), .A(n9513), .ZN(n9514) );
  OAI21_X1 U11350 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(n9517) );
  OAI221_X1 U11351 ( .B1(P3_DATAO_REG_25__SCAN_IN), .B2(keyinput_199), .C1(
        n12193), .C2(n9518), .A(n9517), .ZN(n9522) );
  INV_X1 U11352 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n12263) );
  INV_X1 U11353 ( .A(keyinput_200), .ZN(n9519) );
  INV_X1 U11354 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n12050) );
  INV_X1 U11355 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U11356 ( .A1(n12050), .A2(keyinput_205), .B1(keyinput_204), .B2(
        n12048), .ZN(n9523) );
  OAI221_X1 U11357 ( .B1(n12050), .B2(keyinput_205), .C1(n12048), .C2(
        keyinput_204), .A(n9523), .ZN(n9526) );
  AOI22_X1 U11358 ( .A1(P3_DATAO_REG_22__SCAN_IN), .A2(keyinput_202), .B1(
        P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_203), .ZN(n9524) );
  OAI221_X1 U11359 ( .B1(P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_202), .C1(
        P3_DATAO_REG_21__SCAN_IN), .C2(keyinput_203), .A(n9524), .ZN(n9525) );
  AOI211_X1 U11360 ( .C1(n9528), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9529)
         );
  INV_X1 U11361 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U11362 ( .A1(keyinput_208), .A2(P3_DATAO_REG_16__SCAN_IN), .B1(
        n12058), .B2(keyinput_209), .ZN(n9532) );
  OAI221_X1 U11363 ( .B1(keyinput_208), .B2(P3_DATAO_REG_16__SCAN_IN), .C1(
        n12058), .C2(keyinput_209), .A(n9532), .ZN(n9536) );
  INV_X1 U11364 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n12032) );
  OAI22_X1 U11365 ( .A1(n12032), .A2(keyinput_212), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_210), .ZN(n9533) );
  AOI221_X1 U11366 ( .B1(n12032), .B2(keyinput_212), .C1(keyinput_210), .C2(
        P3_DATAO_REG_14__SCAN_IN), .A(n9533), .ZN(n9535) );
  XNOR2_X1 U11367 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n9534)
         );
  INV_X1 U11368 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n12028) );
  XNOR2_X1 U11369 ( .A(n12028), .B(keyinput_216), .ZN(n9540) );
  AOI22_X1 U11370 ( .A1(P3_DATAO_REG_7__SCAN_IN), .A2(keyinput_217), .B1(
        P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_215), .ZN(n9538) );
  OAI221_X1 U11371 ( .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_217), .C1(
        P3_DATAO_REG_9__SCAN_IN), .C2(keyinput_215), .A(n9538), .ZN(n9539) );
  AOI211_X1 U11372 ( .C1(n9541), .C2(n7560), .A(n9540), .B(n9539), .ZN(n9542)
         );
  AOI221_X1 U11373 ( .B1(P3_DATAO_REG_6__SCAN_IN), .B2(n9543), .C1(n11661), 
        .C2(keyinput_218), .A(n9542), .ZN(n9550) );
  AOI22_X1 U11374 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_220), .B1(
        P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_219), .ZN(n9544) );
  OAI221_X1 U11375 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput_220), .C1(
        P3_DATAO_REG_5__SCAN_IN), .C2(keyinput_219), .A(n9544), .ZN(n9549) );
  OAI22_X1 U11376 ( .A1(n16310), .A2(keyinput_225), .B1(
        P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_222), .ZN(n9545) );
  AOI221_X1 U11377 ( .B1(n16310), .B2(keyinput_225), .C1(keyinput_222), .C2(
        P3_DATAO_REG_2__SCAN_IN), .A(n9545), .ZN(n9548) );
  INV_X1 U11378 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n12044) );
  INV_X1 U11379 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n12064) );
  OAI22_X1 U11380 ( .A1(n12044), .A2(keyinput_221), .B1(n12064), .B2(
        keyinput_224), .ZN(n9546) );
  AOI221_X1 U11381 ( .B1(n12044), .B2(keyinput_221), .C1(keyinput_224), .C2(
        n12064), .A(n9546), .ZN(n9547) );
  OAI211_X1 U11382 ( .C1(n9550), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9557)
         );
  OAI22_X1 U11383 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_227), .B1(
        P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_228), .ZN(n9551) );
  AOI221_X1 U11384 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_227), .C1(
        keyinput_228), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n9551), .ZN(n9556) );
  AOI22_X1 U11385 ( .A1(P3_DATAO_REG_1__SCAN_IN), .A2(keyinput_223), .B1(
        P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_226), .ZN(n9552) );
  OAI221_X1 U11386 ( .B1(P3_DATAO_REG_1__SCAN_IN), .B2(keyinput_223), .C1(
        P3_ADDR_REG_1__SCAN_IN), .C2(keyinput_226), .A(n9552), .ZN(n9555) );
  AOI22_X1 U11387 ( .A1(keyinput_231), .A2(P3_ADDR_REG_6__SCAN_IN), .B1(n16335), .B2(keyinput_229), .ZN(n9553) );
  OAI221_X1 U11388 ( .B1(keyinput_231), .B2(P3_ADDR_REG_6__SCAN_IN), .C1(
        n16335), .C2(keyinput_229), .A(n9553), .ZN(n9554) );
  AOI221_X1 U11389 ( .B1(n9557), .B2(n9556), .C1(n9555), .C2(n9556), .A(n9554), 
        .ZN(n9565) );
  XNOR2_X1 U11390 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_230), .ZN(n9564)
         );
  INV_X1 U11391 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U11392 ( .A1(n16366), .A2(keyinput_233), .B1(keyinput_232), .B2(
        n9559), .ZN(n9558) );
  OAI221_X1 U11393 ( .B1(n16366), .B2(keyinput_233), .C1(n9559), .C2(
        keyinput_232), .A(n9558), .ZN(n9563) );
  XOR2_X1 U11394 ( .A(n16376), .B(keyinput_234), .Z(n9561) );
  XNOR2_X1 U11395 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_235), .ZN(n9560) );
  NAND2_X1 U11396 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  AOI211_X1 U11397 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9562), .ZN(n9569)
         );
  INV_X1 U11398 ( .A(keyinput_236), .ZN(n9566) );
  INV_X1 U11399 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9752) );
  AOI22_X1 U11400 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(n9566), .B1(keyinput_236), 
        .B2(n9752), .ZN(n9567) );
  INV_X1 U11401 ( .A(n9567), .ZN(n9568) );
  XNOR2_X1 U11402 ( .A(n10620), .B(keyinput_237), .ZN(n9571) );
  XNOR2_X1 U11403 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .ZN(n9570) );
  NAND2_X1 U11404 ( .A1(n9571), .A2(n9570), .ZN(n9575) );
  XOR2_X1 U11405 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .Z(n9574) );
  XOR2_X1 U11406 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .Z(n9573) );
  XNOR2_X1 U11407 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_240), .ZN(n9572) );
  INV_X1 U11408 ( .A(keyinput_242), .ZN(n9577) );
  INV_X1 U11409 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9765) );
  OR2_X1 U11410 ( .A1(n9577), .A2(n9765), .ZN(n9578) );
  OAI211_X1 U11411 ( .C1(P1_IR_REG_7__SCAN_IN), .C2(keyinput_242), .A(n9579), 
        .B(n9578), .ZN(n9585) );
  XNOR2_X1 U11412 ( .A(n10611), .B(keyinput_243), .ZN(n9581) );
  XNOR2_X1 U11413 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n9580) );
  NOR2_X1 U11414 ( .A1(n9581), .A2(n9580), .ZN(n9584) );
  AND2_X1 U11415 ( .A1(keyinput_245), .A2(n10610), .ZN(n9583) );
  NOR2_X1 U11416 ( .A1(n10610), .A2(keyinput_245), .ZN(n9582) );
  INV_X1 U11417 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9588) );
  XOR2_X1 U11418 ( .A(keyinput_251), .B(n9588), .Z(n9590) );
  XNOR2_X1 U11419 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_250), .ZN(n9589) );
  NAND2_X1 U11420 ( .A1(n9590), .A2(n9589), .ZN(n9594) );
  XNOR2_X1 U11421 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .ZN(n9593) );
  OAI22_X1 U11422 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_254), .B1(
        keyinput_252), .B2(P1_IR_REG_17__SCAN_IN), .ZN(n9591) );
  AOI221_X1 U11423 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_254), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_252), .A(n9591), .ZN(n9592) );
  OAI211_X1 U11424 ( .C1(n9595), .C2(n9594), .A(n9593), .B(n9592), .ZN(n9597)
         );
  AOI21_X1 U11425 ( .B1(n9597), .B2(keyinput_255), .A(keyinput_127), .ZN(n9599) );
  INV_X1 U11426 ( .A(keyinput_255), .ZN(n9596) );
  AOI21_X1 U11427 ( .B1(n9597), .B2(n9596), .A(P1_IR_REG_20__SCAN_IN), .ZN(
        n9598) );
  AOI22_X1 U11428 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(n9599), .B1(keyinput_127), 
        .B2(n9598), .ZN(n9782) );
  INV_X1 U11429 ( .A(keyinput_118), .ZN(n9769) );
  AOI22_X1 U11430 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_115), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_116), .ZN(n9600) );
  OAI221_X1 U11431 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_115), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_116), .A(n9600), .ZN(n9767) );
  INV_X1 U11432 ( .A(keyinput_114), .ZN(n9766) );
  INV_X1 U11433 ( .A(keyinput_85), .ZN(n9721) );
  INV_X1 U11434 ( .A(keyinput_79), .ZN(n9713) );
  INV_X1 U11435 ( .A(keyinput_78), .ZN(n9712) );
  INV_X1 U11436 ( .A(keyinput_72), .ZN(n9707) );
  INV_X1 U11437 ( .A(keyinput_61), .ZN(n9691) );
  INV_X1 U11438 ( .A(keyinput_60), .ZN(n9690) );
  XOR2_X1 U11439 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .Z(n9688) );
  INV_X1 U11440 ( .A(keyinput_53), .ZN(n9676) );
  INV_X1 U11441 ( .A(keyinput_49), .ZN(n9668) );
  INV_X1 U11442 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n14155) );
  OAI22_X1 U11443 ( .A1(n14155), .A2(keyinput_41), .B1(keyinput_42), .B2(
        P3_REG3_REG_28__SCAN_IN), .ZN(n9601) );
  AOI221_X1 U11444 ( .B1(n14155), .B2(keyinput_41), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_42), .A(n9601), .ZN(n9660) );
  INV_X1 U11445 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n12507) );
  INV_X1 U11446 ( .A(keyinput_39), .ZN(n9654) );
  OAI22_X1 U11447 ( .A1(SI_1_), .A2(keyinput_31), .B1(SI_0_), .B2(keyinput_32), 
        .ZN(n9602) );
  AOI221_X1 U11448 ( .B1(SI_1_), .B2(keyinput_31), .C1(keyinput_32), .C2(SI_0_), .A(n9602), .ZN(n9650) );
  INV_X1 U11449 ( .A(keyinput_13), .ZN(n9624) );
  XNOR2_X1 U11450 ( .A(keyinput_8), .B(n13307), .ZN(n9623) );
  INV_X1 U11451 ( .A(keyinput_7), .ZN(n9616) );
  INV_X1 U11452 ( .A(keyinput_5), .ZN(n9610) );
  INV_X1 U11453 ( .A(keyinput_3), .ZN(n9605) );
  INV_X1 U11454 ( .A(keyinput_1), .ZN(n9604) );
  OAI22_X1 U11455 ( .A1(SI_30_), .A2(keyinput_2), .B1(keyinput_0), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n9603) );
  INV_X1 U11456 ( .A(keyinput_4), .ZN(n9606) );
  OAI221_X1 U11457 ( .B1(SI_27_), .B2(n9610), .C1(n14964), .C2(keyinput_5), 
        .A(n9609), .ZN(n9614) );
  INV_X1 U11458 ( .A(keyinput_6), .ZN(n9611) );
  OAI221_X1 U11459 ( .B1(SI_25_), .B2(n9616), .C1(n13303), .C2(keyinput_7), 
        .A(n9615), .ZN(n9622) );
  AOI22_X1 U11460 ( .A1(n10343), .A2(keyinput_10), .B1(n9618), .B2(keyinput_9), 
        .ZN(n9617) );
  OAI221_X1 U11461 ( .B1(n10343), .B2(keyinput_10), .C1(n9618), .C2(keyinput_9), .A(n9617), .ZN(n9621) );
  AOI22_X1 U11462 ( .A1(SI_21_), .A2(keyinput_11), .B1(n12466), .B2(
        keyinput_12), .ZN(n9619) );
  OAI221_X1 U11463 ( .B1(SI_21_), .B2(keyinput_11), .C1(n12466), .C2(
        keyinput_12), .A(n9619), .ZN(n9620) );
  AOI22_X1 U11464 ( .A1(SI_15_), .A2(keyinput_17), .B1(SI_18_), .B2(
        keyinput_14), .ZN(n9625) );
  OAI221_X1 U11465 ( .B1(SI_15_), .B2(keyinput_17), .C1(SI_18_), .C2(
        keyinput_14), .A(n9625), .ZN(n9630) );
  AOI22_X1 U11466 ( .A1(SI_16_), .A2(keyinput_16), .B1(SI_17_), .B2(
        keyinput_15), .ZN(n9626) );
  OAI221_X1 U11467 ( .B1(SI_16_), .B2(keyinput_16), .C1(SI_17_), .C2(
        keyinput_15), .A(n9626), .ZN(n9629) );
  AOI22_X1 U11468 ( .A1(n11452), .A2(keyinput_19), .B1(n11532), .B2(
        keyinput_18), .ZN(n9627) );
  OAI221_X1 U11469 ( .B1(n11452), .B2(keyinput_19), .C1(n11532), .C2(
        keyinput_18), .A(n9627), .ZN(n9628) );
  AOI22_X1 U11470 ( .A1(n11319), .A2(keyinput_20), .B1(keyinput_21), .B2(
        n11307), .ZN(n9631) );
  OAI221_X1 U11471 ( .B1(n11319), .B2(keyinput_20), .C1(n11307), .C2(
        keyinput_21), .A(n9631), .ZN(n9632) );
  INV_X1 U11472 ( .A(n9632), .ZN(n9639) );
  AOI22_X1 U11473 ( .A1(SI_7_), .A2(keyinput_25), .B1(SI_8_), .B2(keyinput_24), 
        .ZN(n9633) );
  OAI221_X1 U11474 ( .B1(SI_7_), .B2(keyinput_25), .C1(SI_8_), .C2(keyinput_24), .A(n9633), .ZN(n9634) );
  INV_X1 U11475 ( .A(n9634), .ZN(n9638) );
  INV_X1 U11476 ( .A(keyinput_22), .ZN(n9635) );
  XNOR2_X1 U11477 ( .A(n9635), .B(SI_10_), .ZN(n9637) );
  XNOR2_X1 U11478 ( .A(SI_9_), .B(keyinput_23), .ZN(n9636) );
  NAND4_X1 U11479 ( .A1(n9639), .A2(n9638), .A3(n9637), .A4(n9636), .ZN(n9640)
         );
  AOI22_X1 U11480 ( .A1(n11267), .A2(keyinput_26), .B1(keyinput_27), .B2(n9940), .ZN(n9641) );
  OAI221_X1 U11481 ( .B1(n11267), .B2(keyinput_26), .C1(n9940), .C2(
        keyinput_27), .A(n9641), .ZN(n9642) );
  INV_X1 U11482 ( .A(SI_4_), .ZN(n11263) );
  OAI22_X1 U11483 ( .A1(n9643), .A2(n9642), .B1(keyinput_28), .B2(n11263), 
        .ZN(n9646) );
  OAI22_X1 U11484 ( .A1(SI_3_), .A2(keyinput_29), .B1(SI_2_), .B2(keyinput_30), 
        .ZN(n9644) );
  AOI221_X1 U11485 ( .B1(SI_3_), .B2(keyinput_29), .C1(keyinput_30), .C2(SI_2_), .A(n9644), .ZN(n9645) );
  XOR2_X1 U11486 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .Z(n9649) );
  AOI22_X1 U11487 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_34), .ZN(n9647) );
  OAI221_X1 U11488 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_34), .A(n9647), .ZN(n9648) );
  INV_X1 U11489 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U11490 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(n13533), .B2(keyinput_37), .ZN(n9651) );
  OAI221_X1 U11491 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        n13533), .C2(keyinput_37), .A(n9651), .ZN(n9652) );
  OAI221_X1 U11492 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        n12507), .C2(n9654), .A(n9653), .ZN(n9658) );
  INV_X1 U11493 ( .A(keyinput_40), .ZN(n9655) );
  XOR2_X1 U11494 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9667) );
  INV_X1 U11495 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9663) );
  OAI22_X1 U11496 ( .A1(n9663), .A2(keyinput_47), .B1(n9662), .B2(keyinput_48), 
        .ZN(n9661) );
  AOI221_X1 U11497 ( .B1(n9663), .B2(keyinput_47), .C1(keyinput_48), .C2(n9662), .A(n9661), .ZN(n9666) );
  OAI22_X1 U11498 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .ZN(n9664) );
  AOI221_X1 U11499 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        keyinput_46), .C2(P3_REG3_REG_12__SCAN_IN), .A(n9664), .ZN(n9665) );
  OAI22_X1 U11500 ( .A1(n9670), .A2(keyinput_50), .B1(keyinput_51), .B2(
        P3_REG3_REG_24__SCAN_IN), .ZN(n9669) );
  AOI221_X1 U11501 ( .B1(n9670), .B2(keyinput_50), .C1(P3_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n9669), .ZN(n9672) );
  OAI221_X1 U11502 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n9047), 
        .C2(n9676), .A(n9675), .ZN(n9681) );
  INV_X1 U11503 ( .A(keyinput_54), .ZN(n9677) );
  INV_X1 U11504 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9683) );
  AOI22_X1 U11505 ( .A1(n9126), .A2(keyinput_56), .B1(n9683), .B2(keyinput_57), 
        .ZN(n9682) );
  OAI221_X1 U11506 ( .B1(n9126), .B2(keyinput_56), .C1(n9683), .C2(keyinput_57), .A(n9682), .ZN(n9687) );
  INV_X1 U11507 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9685) );
  AOI22_X1 U11508 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_58), .B1(n9685), 
        .B2(keyinput_59), .ZN(n9684) );
  OAI221_X1 U11509 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .C1(n9685), .C2(keyinput_59), .A(n9684), .ZN(n9686) );
  AOI22_X1 U11510 ( .A1(n10908), .A2(keyinput_63), .B1(keyinput_65), .B2(
        n12685), .ZN(n9692) );
  OAI221_X1 U11511 ( .B1(n10908), .B2(keyinput_63), .C1(n12685), .C2(
        keyinput_65), .A(n9692), .ZN(n9695) );
  INV_X1 U11512 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U11513 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_64), .B1(n12740), .B2(
        keyinput_66), .ZN(n9693) );
  OAI221_X1 U11514 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_64), .C1(n12740), 
        .C2(keyinput_66), .A(n9693), .ZN(n9694) );
  AOI211_X1 U11515 ( .C1(keyinput_62), .C2(P3_REG3_REG_26__SCAN_IN), .A(n9695), 
        .B(n9694), .ZN(n9696) );
  OAI21_X1 U11516 ( .B1(keyinput_62), .B2(P3_REG3_REG_26__SCAN_IN), .A(n9696), 
        .ZN(n9699) );
  OAI22_X1 U11517 ( .A1(n12771), .A2(keyinput_67), .B1(
        P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_68), .ZN(n9697) );
  AOI221_X1 U11518 ( .B1(n12771), .B2(keyinput_67), .C1(keyinput_68), .C2(
        P3_DATAO_REG_28__SCAN_IN), .A(n9697), .ZN(n9698) );
  OAI21_X1 U11519 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9704) );
  OAI22_X1 U11520 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput_69), .B1(
        P3_DATAO_REG_26__SCAN_IN), .B2(keyinput_70), .ZN(n9701) );
  AOI221_X1 U11521 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_69), .C1(
        keyinput_70), .C2(P3_DATAO_REG_26__SCAN_IN), .A(n9701), .ZN(n9703) );
  INV_X1 U11522 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U11523 ( .A1(n12048), .A2(keyinput_76), .B1(n12060), .B2(
        keyinput_75), .ZN(n9708) );
  OAI221_X1 U11524 ( .B1(n12048), .B2(keyinput_76), .C1(n12060), .C2(
        keyinput_75), .A(n9708), .ZN(n9711) );
  AOI22_X1 U11525 ( .A1(P3_DATAO_REG_19__SCAN_IN), .A2(keyinput_77), .B1(
        P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_74), .ZN(n9709) );
  OAI221_X1 U11526 ( .B1(P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_77), .C1(
        P3_DATAO_REG_22__SCAN_IN), .C2(keyinput_74), .A(n9709), .ZN(n9710) );
  AOI22_X1 U11527 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput_80), .B1(
        n12058), .B2(keyinput_81), .ZN(n9714) );
  OAI221_X1 U11528 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_80), .C1(
        n12058), .C2(keyinput_81), .A(n9714), .ZN(n9718) );
  INV_X1 U11529 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n12040) );
  OAI22_X1 U11530 ( .A1(n12040), .A2(keyinput_83), .B1(keyinput_84), .B2(
        P3_DATAO_REG_12__SCAN_IN), .ZN(n9715) );
  AOI221_X1 U11531 ( .B1(n12040), .B2(keyinput_83), .C1(
        P3_DATAO_REG_12__SCAN_IN), .C2(keyinput_84), .A(n9715), .ZN(n9717) );
  INV_X1 U11532 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n12054) );
  XOR2_X1 U11533 ( .A(n12054), .B(keyinput_82), .Z(n9716) );
  OAI211_X1 U11534 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9720)
         );
  OAI221_X1 U11535 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_85), .C1(
        n12036), .C2(n9721), .A(n9720), .ZN(n9723) );
  XOR2_X1 U11536 ( .A(n12038), .B(keyinput_86), .Z(n9722) );
  OAI22_X1 U11537 ( .A1(P3_DATAO_REG_7__SCAN_IN), .A2(keyinput_89), .B1(
        P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_88), .ZN(n9724) );
  AOI221_X1 U11538 ( .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_89), .C1(
        keyinput_88), .C2(P3_DATAO_REG_8__SCAN_IN), .A(n9724), .ZN(n9725) );
  INV_X1 U11539 ( .A(keyinput_90), .ZN(n9729) );
  AOI22_X1 U11540 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_92), .B1(
        P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_91), .ZN(n9726) );
  OAI221_X1 U11541 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput_92), .C1(
        P3_DATAO_REG_5__SCAN_IN), .C2(keyinput_91), .A(n9726), .ZN(n9727) );
  INV_X1 U11542 ( .A(n9727), .ZN(n9728) );
  INV_X1 U11543 ( .A(n9730), .ZN(n9737) );
  AOI22_X1 U11544 ( .A1(P3_DATAO_REG_3__SCAN_IN), .A2(keyinput_93), .B1(
        P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_97), .ZN(n9731) );
  OAI221_X1 U11545 ( .B1(P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_93), .C1(
        P3_ADDR_REG_0__SCAN_IN), .C2(keyinput_97), .A(n9731), .ZN(n9736) );
  AOI22_X1 U11546 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput_94), .B1(
        P3_DATAO_REG_1__SCAN_IN), .B2(keyinput_95), .ZN(n9732) );
  OAI221_X1 U11547 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_94), .C1(
        P3_DATAO_REG_1__SCAN_IN), .C2(keyinput_95), .A(n9732), .ZN(n9735) );
  AOI22_X1 U11548 ( .A1(n12064), .A2(keyinput_96), .B1(n16308), .B2(
        keyinput_98), .ZN(n9733) );
  OAI221_X1 U11549 ( .B1(n12064), .B2(keyinput_96), .C1(n16308), .C2(
        keyinput_98), .A(n9733), .ZN(n9734) );
  NOR4_X1 U11550 ( .A1(n9737), .A2(n9736), .A3(n9735), .A4(n9734), .ZN(n9740)
         );
  AOI22_X1 U11551 ( .A1(n16317), .A2(keyinput_99), .B1(keyinput_100), .B2(
        n16322), .ZN(n9738) );
  OAI221_X1 U11552 ( .B1(n16317), .B2(keyinput_99), .C1(n16322), .C2(
        keyinput_100), .A(n9738), .ZN(n9739) );
  AOI22_X1 U11553 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput_103), .B1(n16341), .B2(keyinput_102), .ZN(n9741) );
  OAI221_X1 U11554 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_103), .C1(
        n16341), .C2(keyinput_102), .A(n9741), .ZN(n9744) );
  NAND2_X1 U11555 ( .A1(keyinput_101), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n9742)
         );
  OAI22_X1 U11556 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(keyinput_105), .B1(
        P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_104), .ZN(n9746) );
  AOI221_X1 U11557 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(keyinput_105), .C1(
        keyinput_104), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n9746), .ZN(n9750) );
  INV_X1 U11558 ( .A(keyinput_106), .ZN(n9747) );
  XNOR2_X1 U11559 ( .A(n9747), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n9749) );
  XNOR2_X1 U11560 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_107), .ZN(n9748) );
  NAND3_X1 U11561 ( .A1(n9750), .A2(n9749), .A3(n9748), .ZN(n9755) );
  INV_X1 U11562 ( .A(keyinput_108), .ZN(n9751) );
  OAI22_X1 U11563 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_108), .B1(n9752), 
        .B2(n9751), .ZN(n9753) );
  INV_X1 U11564 ( .A(n9753), .ZN(n9754) );
  OAI21_X1 U11565 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9763) );
  OAI22_X1 U11566 ( .A1(n10620), .A2(keyinput_109), .B1(keyinput_110), .B2(
        P1_IR_REG_3__SCAN_IN), .ZN(n9757) );
  AOI221_X1 U11567 ( .B1(n10620), .B2(keyinput_109), .C1(P1_IR_REG_3__SCAN_IN), 
        .C2(keyinput_110), .A(n9757), .ZN(n9762) );
  XOR2_X1 U11568 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .Z(n9761) );
  XOR2_X1 U11569 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_113), .Z(n9759) );
  XNOR2_X1 U11570 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_112), .ZN(n9758) );
  NAND2_X1 U11571 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  AOI211_X1 U11572 ( .C1(n9763), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9764)
         );
  XOR2_X1 U11573 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_119), .Z(n9771) );
  XNOR2_X1 U11574 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_120), .ZN(n9770) );
  NAND2_X1 U11575 ( .A1(n9771), .A2(n9770), .ZN(n9773) );
  XOR2_X1 U11576 ( .A(n11100), .B(keyinput_121), .Z(n9772) );
  XOR2_X1 U11577 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .Z(n9776) );
  XNOR2_X1 U11578 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_122), .ZN(n9775) );
  INV_X1 U11579 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9778) );
  XOR2_X1 U11580 ( .A(n9778), .B(keyinput_125), .Z(n9781) );
  XNOR2_X1 U11581 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_124), .ZN(n9780) );
  XNOR2_X1 U11582 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_126), .ZN(n9779) );
  INV_X1 U11583 ( .A(n12116), .ZN(n9784) );
  OR2_X1 U11584 ( .A1(n14451), .A2(n9784), .ZN(n9783) );
  NAND2_X1 U11585 ( .A1(n9783), .A2(n9345), .ZN(n10870) );
  NAND2_X1 U11586 ( .A1(n9784), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14515) );
  INV_X1 U11587 ( .A(n14515), .ZN(n9785) );
  NAND2_X1 U11588 ( .A1(n14572), .A2(n10875), .ZN(n9786) );
  INV_X1 U11589 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9792) );
  INV_X1 U11590 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9791) );
  INV_X1 U11592 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12095) );
  OR2_X1 U11593 ( .A1(n9890), .A2(n12095), .ZN(n9801) );
  AND2_X2 U11594 ( .A1(n13918), .A2(n9863), .ZN(n9837) );
  NAND2_X2 U11595 ( .A1(n15612), .A2(n13918), .ZN(n9888) );
  INV_X1 U11596 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9798) );
  INV_X1 U11597 ( .A(n11723), .ZN(n15097) );
  NOR2_X1 U11598 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n9804) );
  NAND4_X1 U11599 ( .A1(n9804), .A2(n9803), .A3(n9802), .A4(n9792), .ZN(n9805)
         );
  INV_X1 U11600 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U11601 ( .A1(n9807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U11602 ( .A1(n9808), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U11603 ( .A1(n9814), .A2(n15605), .ZN(n9815) );
  NAND2_X1 U11604 ( .A1(n9815), .A2(n9790), .ZN(n9810) );
  INV_X1 U11605 ( .A(n9815), .ZN(n9816) );
  XNOR2_X2 U11606 ( .A(n9816), .B(P2_IR_REG_21__SCAN_IN), .ZN(n11248) );
  NAND2_X1 U11607 ( .A1(n15097), .A2(n10540), .ZN(n9836) );
  INV_X1 U11608 ( .A(n9819), .ZN(n9818) );
  NAND2_X1 U11609 ( .A1(n9848), .A2(n9821), .ZN(n9907) );
  NAND2_X1 U11610 ( .A1(n9907), .A2(SI_2_), .ZN(n9899) );
  OAI21_X1 U11611 ( .B1(n9907), .B2(SI_2_), .A(n9899), .ZN(n9823) );
  INV_X1 U11612 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n11329) );
  MUX2_X1 U11613 ( .A(n9822), .B(n11329), .S(n9895), .Z(n9903) );
  NAND2_X1 U11614 ( .A1(n9823), .A2(n9903), .ZN(n9824) );
  NAND2_X1 U11615 ( .A1(n9827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9828) );
  INV_X2 U11616 ( .A(n10101), .ZN(n9944) );
  INV_X1 U11617 ( .A(n9831), .ZN(n9832) );
  NAND2_X1 U11618 ( .A1(n9832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9833) );
  XNOR2_X1 U11619 ( .A(n9833), .B(P2_IR_REG_2__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U11620 ( .A1(n9944), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9909), .B2(
        n16228), .ZN(n9834) );
  INV_X1 U11621 ( .A(n16521), .ZN(n12101) );
  INV_X1 U11622 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9838) );
  OR2_X1 U11623 ( .A1(n9888), .A2(n9838), .ZN(n9843) );
  INV_X1 U11624 ( .A(n9887), .ZN(n9839) );
  NAND2_X1 U11625 ( .A1(n9839), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U11626 ( .A1(n9840), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9841) );
  NAND4_X2 U11627 ( .A1(n9844), .A2(n9843), .A3(n9842), .A4(n9841), .ZN(n9875)
         );
  NAND2_X1 U11628 ( .A1(n9875), .A2(n9986), .ZN(n9850) );
  INV_X1 U11629 ( .A(n9845), .ZN(n9846) );
  NAND2_X1 U11630 ( .A1(n7530), .A2(n9846), .ZN(n9847) );
  NAND2_X1 U11631 ( .A1(n9848), .A2(n9847), .ZN(n11318) );
  NAND2_X1 U11632 ( .A1(n9876), .A2(n10540), .ZN(n9849) );
  NAND2_X1 U11633 ( .A1(n9850), .A2(n9849), .ZN(n9879) );
  AOI22_X1 U11634 ( .A1(n9857), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n9855) );
  INV_X1 U11635 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U11636 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_30__SCAN_IN), 
        .ZN(n9851) );
  OAI21_X1 U11637 ( .B1(n9852), .B2(P2_IR_REG_30__SCAN_IN), .A(n9851), .ZN(
        n9853) );
  NAND2_X1 U11638 ( .A1(n9860), .A2(n9853), .ZN(n9854) );
  OAI21_X1 U11639 ( .B1(n9860), .B2(n9855), .A(n9854), .ZN(n9856) );
  NAND2_X1 U11640 ( .A1(n9856), .A2(n15612), .ZN(n9866) );
  AOI22_X1 U11641 ( .A1(n9857), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n9862) );
  INV_X1 U11642 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U11643 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n9858) );
  OAI21_X1 U11644 ( .B1(n11524), .B2(P2_IR_REG_30__SCAN_IN), .A(n9858), .ZN(
        n9859) );
  NAND2_X1 U11645 ( .A1(n9860), .A2(n9859), .ZN(n9861) );
  OAI21_X1 U11646 ( .B1(n9860), .B2(n9862), .A(n9861), .ZN(n9864) );
  NAND2_X1 U11647 ( .A1(n9864), .A2(n9863), .ZN(n9865) );
  NAND2_X1 U11648 ( .A1(n15099), .A2(n11662), .ZN(n9871) );
  INV_X1 U11649 ( .A(SI_0_), .ZN(n9867) );
  NOR2_X1 U11650 ( .A1(n11277), .A2(n9867), .ZN(n9869) );
  XNOR2_X1 U11651 ( .A(n9869), .B(n9868), .ZN(n15629) );
  MUX2_X1 U11652 ( .A(P2_IR_REG_0__SCAN_IN), .B(n15629), .S(n9870), .Z(n11919)
         );
  NAND2_X1 U11653 ( .A1(n9871), .A2(n11919), .ZN(n9872) );
  OAI211_X1 U11654 ( .C1(n15099), .C2(n11662), .A(n9872), .B(n9986), .ZN(n9874) );
  INV_X1 U11655 ( .A(n11919), .ZN(n11668) );
  NAND2_X1 U11656 ( .A1(n11668), .A2(n15099), .ZN(n11735) );
  NAND2_X1 U11657 ( .A1(n11735), .A2(n9977), .ZN(n9873) );
  NAND2_X1 U11658 ( .A1(n9874), .A2(n9873), .ZN(n9880) );
  NAND2_X1 U11659 ( .A1(n9879), .A2(n9880), .ZN(n9878) );
  OAI22_X1 U11660 ( .A1(n10575), .A2(n9986), .B1(n10540), .B2(n14066), .ZN(
        n9877) );
  NAND2_X1 U11661 ( .A1(n9878), .A2(n9877), .ZN(n9884) );
  INV_X1 U11662 ( .A(n9879), .ZN(n9882) );
  INV_X1 U11663 ( .A(n9880), .ZN(n9881) );
  NAND2_X1 U11664 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  OAI22_X1 U11665 ( .A1(n11723), .A2(n10540), .B1(n16521), .B2(n10499), .ZN(
        n9885) );
  OAI21_X1 U11666 ( .B1(n7451), .B2(n7561), .A(n9885), .ZN(n9886) );
  NAND2_X1 U11667 ( .A1(n9837), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9894) );
  INV_X1 U11668 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11470) );
  OR2_X1 U11669 ( .A1(n9887), .A2(n11470), .ZN(n9893) );
  INV_X1 U11670 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9889) );
  OR2_X1 U11671 ( .A1(n9888), .A2(n9889), .ZN(n9892) );
  OR2_X1 U11672 ( .A1(n10463), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9891) );
  AND4_X2 U11673 ( .A1(n9894), .A2(n9893), .A3(n9892), .A4(n9891), .ZN(n11832)
         );
  NAND2_X1 U11674 ( .A1(n9896), .A2(SI_3_), .ZN(n9921) );
  INV_X1 U11675 ( .A(n9896), .ZN(n9897) );
  NAND2_X1 U11676 ( .A1(n9897), .A2(n11260), .ZN(n9898) );
  NAND2_X1 U11677 ( .A1(n9921), .A2(n9898), .ZN(n9902) );
  NAND3_X1 U11678 ( .A1(n9900), .A2(n9902), .A3(n9899), .ZN(n9908) );
  INV_X1 U11679 ( .A(n9903), .ZN(n9901) );
  AND2_X1 U11680 ( .A1(n9901), .A2(SI_2_), .ZN(n9906) );
  INV_X1 U11681 ( .A(n9902), .ZN(n9905) );
  INV_X1 U11682 ( .A(SI_2_), .ZN(n11301) );
  NAND2_X1 U11683 ( .A1(n9903), .A2(n11301), .ZN(n9904) );
  OAI211_X1 U11684 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9922)
         );
  AND2_X1 U11685 ( .A1(n9908), .A2(n9922), .ZN(n11278) );
  NAND2_X1 U11686 ( .A1(n11278), .A2(n10511), .ZN(n9913) );
  INV_X1 U11687 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U11688 ( .A1(n9831), .A2(n9910), .ZN(n9927) );
  NAND2_X1 U11689 ( .A1(n9927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9911) );
  XNOR2_X1 U11690 ( .A(n9911), .B(P2_IR_REG_3__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U11691 ( .A1(n9944), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9909), .B2(
        n11485), .ZN(n9912) );
  OAI22_X1 U11692 ( .A1(n10540), .A2(n11832), .B1(n12282), .B2(n10499), .ZN(
        n9914) );
  INV_X1 U11693 ( .A(n9986), .ZN(n9977) );
  OAI22_X1 U11694 ( .A1(n11832), .A2(n10499), .B1(n12282), .B2(n10540), .ZN(
        n9915) );
  INV_X2 U11695 ( .A(n9888), .ZN(n9950) );
  NAND2_X1 U11696 ( .A1(n9950), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9920) );
  INV_X1 U11697 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n12107) );
  OR2_X1 U11698 ( .A1(n9887), .A2(n12107), .ZN(n9919) );
  NAND2_X1 U11699 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9953) );
  OAI21_X1 U11700 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n9953), .ZN(n12108) );
  OR2_X1 U11701 ( .A1(n10463), .A2(n12108), .ZN(n9918) );
  INV_X4 U11702 ( .A(n9837), .ZN(n10494) );
  INV_X1 U11703 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9916) );
  OR2_X1 U11704 ( .A1(n10494), .A2(n9916), .ZN(n9917) );
  AND4_X2 U11705 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), .ZN(n11942)
         );
  NAND2_X1 U11706 ( .A1(n9922), .A2(n9921), .ZN(n9925) );
  NAND2_X1 U11707 ( .A1(n9923), .A2(SI_4_), .ZN(n9937) );
  OR2_X1 U11708 ( .A1(n9925), .A2(n9924), .ZN(n9926) );
  NAND2_X1 U11709 ( .A1(n11312), .A2(n10511), .ZN(n9934) );
  NAND2_X1 U11710 ( .A1(n9929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9928) );
  MUX2_X1 U11711 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9928), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9932) );
  INV_X1 U11712 ( .A(n9929), .ZN(n9931) );
  INV_X1 U11713 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U11714 ( .A1(n9931), .A2(n9930), .ZN(n9946) );
  NAND2_X1 U11715 ( .A1(n9932), .A2(n9946), .ZN(n11500) );
  INV_X1 U11716 ( .A(n11500), .ZN(n11495) );
  AOI22_X1 U11717 ( .A1(n9944), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9909), .B2(
        n11495), .ZN(n9933) );
  OAI22_X1 U11718 ( .A1(n11942), .A2(n10499), .B1(n12109), .B2(n10540), .ZN(
        n9935) );
  OAI22_X1 U11719 ( .A1(n10540), .A2(n11942), .B1(n12109), .B2(n10499), .ZN(
        n9936) );
  INV_X1 U11720 ( .A(n9962), .ZN(n9959) );
  NAND2_X1 U11721 ( .A1(n9938), .A2(n9937), .ZN(n9942) );
  NAND2_X1 U11722 ( .A1(n9939), .A2(SI_5_), .ZN(n9966) );
  INV_X1 U11723 ( .A(SI_5_), .ZN(n9940) );
  NAND2_X1 U11724 ( .A1(n9942), .A2(n9941), .ZN(n9967) );
  OR2_X1 U11725 ( .A1(n9942), .A2(n9941), .ZN(n9943) );
  NAND2_X1 U11726 ( .A1(n9967), .A2(n9943), .ZN(n11326) );
  OR2_X1 U11727 ( .A1(n11326), .A2(n10208), .ZN(n9949) );
  NAND2_X1 U11728 ( .A1(n9946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9945) );
  MUX2_X1 U11729 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9945), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9947) );
  AOI22_X1 U11730 ( .A1(n9944), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9909), .B2(
        n11520), .ZN(n9948) );
  NAND2_X1 U11731 ( .A1(n9950), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9958) );
  INV_X1 U11732 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11501) );
  OR2_X1 U11733 ( .A1(n9887), .A2(n11501), .ZN(n9957) );
  INV_X1 U11734 ( .A(n9953), .ZN(n9951) );
  NAND2_X1 U11735 ( .A1(n9951), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9980) );
  INV_X1 U11736 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U11737 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  NAND2_X1 U11738 ( .A1(n9980), .A2(n9954), .ZN(n12082) );
  OR2_X1 U11739 ( .A1(n10463), .A2(n12082), .ZN(n9956) );
  INV_X1 U11740 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11496) );
  OR2_X1 U11741 ( .A1(n10494), .A2(n11496), .ZN(n9955) );
  OAI22_X1 U11742 ( .A1(n11968), .A2(n10220), .B1(n10540), .B2(n11969), .ZN(
        n9960) );
  NAND2_X1 U11743 ( .A1(n9959), .A2(n9960), .ZN(n9965) );
  OAI22_X1 U11744 ( .A1(n11968), .A2(n7420), .B1(n11969), .B2(n10220), .ZN(
        n9964) );
  INV_X1 U11745 ( .A(n9960), .ZN(n9961) );
  AND2_X1 U11746 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  MUX2_X1 U11747 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n11277), .Z(n9968) );
  NAND2_X1 U11748 ( .A1(n9968), .A2(SI_6_), .ZN(n9989) );
  INV_X1 U11749 ( .A(n9968), .ZN(n9969) );
  NAND2_X1 U11750 ( .A1(n9969), .A2(n11267), .ZN(n9970) );
  NAND2_X1 U11751 ( .A1(n9972), .A2(n9971), .ZN(n9990) );
  OR2_X1 U11752 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  NAND2_X1 U11753 ( .A1(n9990), .A2(n9973), .ZN(n11311) );
  OR2_X1 U11754 ( .A1(n11311), .A2(n10208), .ZN(n9976) );
  NAND2_X1 U11755 ( .A1(n9997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9974) );
  XNOR2_X1 U11756 ( .A(n9974), .B(P2_IR_REG_6__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U11757 ( .A1(n9944), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9909), .B2(
        n11547), .ZN(n9975) );
  NAND2_X1 U11758 ( .A1(n9976), .A2(n9975), .ZN(n12296) );
  NAND2_X1 U11759 ( .A1(n9950), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U11760 ( .A1(n9837), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9984) );
  INV_X1 U11761 ( .A(n9980), .ZN(n9978) );
  NAND2_X1 U11762 ( .A1(n9978), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10004) );
  INV_X1 U11763 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U11764 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NAND2_X1 U11765 ( .A1(n10004), .A2(n9981), .ZN(n12144) );
  OR2_X1 U11766 ( .A1(n10463), .A2(n12144), .ZN(n9983) );
  INV_X1 U11767 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n12142) );
  OR2_X1 U11768 ( .A1(n9887), .A2(n12142), .ZN(n9982) );
  NAND4_X1 U11769 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n15093) );
  AOI22_X1 U11770 ( .A1(n12296), .A2(n10499), .B1(n7420), .B2(n15093), .ZN(
        n9987) );
  INV_X1 U11771 ( .A(n15093), .ZN(n12295) );
  OAI22_X1 U11772 ( .A1(n8301), .A2(n10220), .B1(n7420), .B2(n12295), .ZN(
        n9988) );
  MUX2_X1 U11773 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n11277), .Z(n9991) );
  NAND2_X1 U11774 ( .A1(n9991), .A2(SI_7_), .ZN(n10012) );
  INV_X1 U11775 ( .A(n9991), .ZN(n9992) );
  NAND2_X1 U11776 ( .A1(n9992), .A2(n11298), .ZN(n9993) );
  OR2_X1 U11777 ( .A1(n9995), .A2(n9994), .ZN(n9996) );
  NAND2_X1 U11778 ( .A1(n10013), .A2(n9996), .ZN(n11315) );
  OR2_X1 U11779 ( .A1(n11315), .A2(n10208), .ZN(n10001) );
  INV_X1 U11780 ( .A(n9997), .ZN(n9999) );
  INV_X1 U11781 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U11782 ( .A1(n9999), .A2(n9998), .ZN(n10079) );
  NAND2_X1 U11783 ( .A1(n10079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10021) );
  XNOR2_X1 U11784 ( .A(n10021), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U11785 ( .A1(n9944), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9909), .B2(
        n11740), .ZN(n10000) );
  NAND2_X1 U11786 ( .A1(n9950), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U11787 ( .A1(n10514), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10008) );
  INV_X1 U11788 ( .A(n10004), .ZN(n10002) );
  NAND2_X1 U11789 ( .A1(n10002), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10027) );
  INV_X1 U11790 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U11791 ( .A1(n10004), .A2(n10003), .ZN(n10005) );
  NAND2_X1 U11792 ( .A1(n10027), .A2(n10005), .ZN(n12304) );
  OR2_X1 U11793 ( .A1(n10463), .A2(n12304), .ZN(n10007) );
  INV_X1 U11794 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11548) );
  OR2_X1 U11795 ( .A1(n10494), .A2(n11548), .ZN(n10006) );
  NAND4_X1 U11796 ( .A1(n10009), .A2(n10008), .A3(n10007), .A4(n10006), .ZN(
        n15092) );
  AOI22_X1 U11797 ( .A1(n12488), .A2(n7420), .B1(n10499), .B2(n15092), .ZN(
        n10011) );
  INV_X1 U11798 ( .A(n12488), .ZN(n12314) );
  INV_X1 U11799 ( .A(n15092), .ZN(n12487) );
  OAI22_X1 U11800 ( .A1(n12314), .A2(n7420), .B1(n12487), .B2(n10499), .ZN(
        n10010) );
  MUX2_X1 U11801 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n8230), .Z(n10014) );
  NAND2_X1 U11802 ( .A1(n10014), .A2(SI_8_), .ZN(n10042) );
  INV_X1 U11803 ( .A(n10014), .ZN(n10015) );
  NAND2_X1 U11804 ( .A1(n10015), .A2(n11274), .ZN(n10016) );
  OR2_X1 U11805 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  NAND2_X1 U11806 ( .A1(n10043), .A2(n10019), .ZN(n11324) );
  OR2_X1 U11807 ( .A1(n11324), .A2(n10208), .ZN(n10024) );
  INV_X1 U11808 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10020) );
  NAND2_X1 U11809 ( .A1(n10021), .A2(n10020), .ZN(n10022) );
  NAND2_X1 U11810 ( .A1(n10022), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10048) );
  XNOR2_X1 U11811 ( .A(n10048), .B(P2_IR_REG_8__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U11812 ( .A1(n9909), .A2(n11853), .B1(n9944), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U11813 ( .A1(n9837), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10033) );
  INV_X1 U11814 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12494) );
  OR2_X1 U11815 ( .A1(n9887), .A2(n12494), .ZN(n10032) );
  INV_X1 U11816 ( .A(n10027), .ZN(n10025) );
  NAND2_X1 U11817 ( .A1(n10025), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10053) );
  INV_X1 U11818 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U11819 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  NAND2_X1 U11820 ( .A1(n10053), .A2(n10028), .ZN(n12497) );
  OR2_X1 U11821 ( .A1(n10463), .A2(n12497), .ZN(n10031) );
  INV_X1 U11822 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10029) );
  OR2_X1 U11823 ( .A1(n9888), .A2(n10029), .ZN(n10030) );
  OAI22_X1 U11824 ( .A1(n12615), .A2(n10220), .B1(n7420), .B2(n12611), .ZN(
        n10034) );
  NAND2_X1 U11825 ( .A1(n10035), .A2(n10034), .ZN(n10041) );
  INV_X1 U11826 ( .A(n10036), .ZN(n10039) );
  INV_X1 U11827 ( .A(n10037), .ZN(n10038) );
  NAND2_X1 U11828 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  NAND2_X1 U11829 ( .A1(n10075), .A2(SI_9_), .ZN(n10066) );
  MUX2_X1 U11830 ( .A(n11449), .B(n10044), .S(n8230), .Z(n10069) );
  NAND2_X1 U11831 ( .A1(n10045), .A2(n10069), .ZN(n10046) );
  INV_X1 U11832 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U11833 ( .A1(n10048), .A2(n10047), .ZN(n10049) );
  NAND2_X1 U11834 ( .A1(n10049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10050) );
  XNOR2_X1 U11835 ( .A(n10050), .B(P2_IR_REG_9__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U11836 ( .A1(n12534), .A2(n9909), .B1(n9944), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U11837 ( .A1(n10514), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10059) );
  INV_X1 U11838 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11848) );
  OR2_X1 U11839 ( .A1(n10494), .A2(n11848), .ZN(n10058) );
  NAND2_X1 U11840 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  NAND2_X1 U11841 ( .A1(n10088), .A2(n10054), .ZN(n12644) );
  OR2_X1 U11842 ( .A1(n10463), .A2(n12644), .ZN(n10057) );
  INV_X1 U11843 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10055) );
  OR2_X1 U11844 ( .A1(n9888), .A2(n10055), .ZN(n10056) );
  OAI22_X1 U11845 ( .A1(n12789), .A2(n10220), .B1(n7420), .B2(n12621), .ZN(
        n10060) );
  OAI22_X1 U11846 ( .A1(n12789), .A2(n7420), .B1(n12621), .B2(n10220), .ZN(
        n10062) );
  INV_X1 U11847 ( .A(n10060), .ZN(n10061) );
  MUX2_X1 U11848 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n11277), .Z(n10063) );
  NAND2_X1 U11849 ( .A1(n10063), .A2(SI_10_), .ZN(n10096) );
  INV_X1 U11850 ( .A(n10063), .ZN(n10064) );
  NAND2_X1 U11851 ( .A1(n10064), .A2(n11296), .ZN(n10065) );
  NAND2_X1 U11852 ( .A1(n10096), .A2(n10065), .ZN(n10070) );
  AND2_X1 U11853 ( .A1(n10066), .A2(n10070), .ZN(n10067) );
  NAND2_X1 U11854 ( .A1(n10068), .A2(n10067), .ZN(n10076) );
  INV_X1 U11855 ( .A(n10069), .ZN(n10071) );
  AND2_X1 U11856 ( .A1(n10071), .A2(SI_9_), .ZN(n10074) );
  INV_X1 U11857 ( .A(n10070), .ZN(n10073) );
  NAND2_X1 U11858 ( .A1(n10076), .A2(n10097), .ZN(n11454) );
  OR2_X1 U11859 ( .A1(n11454), .A2(n10208), .ZN(n10086) );
  INV_X1 U11860 ( .A(n10077), .ZN(n10078) );
  NAND2_X1 U11861 ( .A1(n10081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U11862 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10080), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n10084) );
  INV_X1 U11863 ( .A(n10081), .ZN(n10083) );
  INV_X1 U11864 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U11865 ( .A1(n10083), .A2(n10082), .ZN(n10098) );
  NAND2_X1 U11866 ( .A1(n10084), .A2(n10098), .ZN(n12535) );
  AOI22_X1 U11867 ( .A1(n16269), .A2(n9909), .B1(n9944), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n10085) );
  AND2_X2 U11868 ( .A1(n10086), .A2(n10085), .ZN(n12917) );
  NAND2_X1 U11869 ( .A1(n9950), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10093) );
  INV_X1 U11870 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n12628) );
  OR2_X1 U11871 ( .A1(n9887), .A2(n12628), .ZN(n10092) );
  INV_X1 U11872 ( .A(n10088), .ZN(n10087) );
  NAND2_X1 U11873 ( .A1(n10087), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10106) );
  INV_X1 U11874 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n16262) );
  NAND2_X1 U11875 ( .A1(n10088), .A2(n16262), .ZN(n10089) );
  NAND2_X1 U11876 ( .A1(n10106), .A2(n10089), .ZN(n12734) );
  OR2_X1 U11877 ( .A1(n10463), .A2(n12734), .ZN(n10091) );
  INV_X1 U11878 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n12536) );
  OR2_X1 U11879 ( .A1(n10494), .A2(n12536), .ZN(n10090) );
  OAI22_X1 U11880 ( .A1(n12917), .A2(n7420), .B1(n12921), .B2(n10220), .ZN(
        n10094) );
  OAI22_X1 U11881 ( .A1(n12917), .A2(n10220), .B1(n7420), .B2(n12921), .ZN(
        n10095) );
  MUX2_X1 U11882 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n11277), .Z(n10118) );
  XNOR2_X1 U11883 ( .A(n10118), .B(SI_11_), .ZN(n10121) );
  XNOR2_X1 U11884 ( .A(n10122), .B(n10121), .ZN(n11541) );
  NAND2_X1 U11885 ( .A1(n11541), .A2(n10511), .ZN(n10104) );
  NAND2_X1 U11886 ( .A1(n10098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U11887 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10099), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n10100) );
  NAND2_X1 U11888 ( .A1(n10100), .A2(n10149), .ZN(n12537) );
  OAI22_X1 U11889 ( .A1(n12537), .A2(n9870), .B1(n10101), .B2(n11542), .ZN(
        n10102) );
  INV_X1 U11890 ( .A(n10102), .ZN(n10103) );
  NAND2_X1 U11891 ( .A1(n9950), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U11892 ( .A1(n10514), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U11893 ( .A1(n10106), .A2(n10105), .ZN(n10107) );
  NAND2_X1 U11894 ( .A1(n10128), .A2(n10107), .ZN(n13030) );
  OR2_X1 U11895 ( .A1(n10463), .A2(n13030), .ZN(n10110) );
  INV_X1 U11896 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10108) );
  OR2_X1 U11897 ( .A1(n10494), .A2(n10108), .ZN(n10109) );
  NAND4_X1 U11898 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n15088) );
  AOI22_X1 U11899 ( .A1(n13052), .A2(n7420), .B1(n10499), .B2(n15088), .ZN(
        n10113) );
  INV_X1 U11900 ( .A(n13052), .ZN(n12927) );
  INV_X1 U11901 ( .A(n15088), .ZN(n13072) );
  OAI22_X1 U11902 ( .A1(n12927), .A2(n7420), .B1(n13072), .B2(n10220), .ZN(
        n10116) );
  INV_X1 U11903 ( .A(n10118), .ZN(n10119) );
  NAND2_X1 U11904 ( .A1(n10119), .A2(n11307), .ZN(n10120) );
  MUX2_X1 U11905 ( .A(n11634), .B(n11636), .S(n11277), .Z(n10140) );
  XNOR2_X1 U11906 ( .A(n10140), .B(SI_12_), .ZN(n10138) );
  XNOR2_X1 U11907 ( .A(n10139), .B(n10138), .ZN(n11633) );
  NAND2_X1 U11908 ( .A1(n11633), .A2(n10511), .ZN(n10125) );
  NAND2_X1 U11909 ( .A1(n10149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10123) );
  XNOR2_X1 U11910 ( .A(n10123), .B(P2_IR_REG_12__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U11911 ( .A1(n9944), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9909), 
        .B2(n12946), .ZN(n10124) );
  NAND2_X1 U11912 ( .A1(n9950), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U11913 ( .A1(n10514), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10132) );
  INV_X1 U11914 ( .A(n10128), .ZN(n10126) );
  NAND2_X1 U11915 ( .A1(n10126), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10171) );
  INV_X1 U11916 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U11917 ( .A1(n10128), .A2(n10127), .ZN(n10129) );
  NAND2_X1 U11918 ( .A1(n10171), .A2(n10129), .ZN(n12984) );
  OR2_X1 U11919 ( .A1(n10463), .A2(n12984), .ZN(n10131) );
  INV_X1 U11920 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12652) );
  OR2_X1 U11921 ( .A1(n10494), .A2(n12652), .ZN(n10130) );
  NAND4_X1 U11922 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n15087) );
  AOI22_X1 U11923 ( .A1(n13191), .A2(n10220), .B1(n7420), .B2(n15087), .ZN(
        n10136) );
  AOI22_X1 U11924 ( .A1(n13191), .A2(n7420), .B1(n10220), .B2(n15087), .ZN(
        n10134) );
  INV_X1 U11925 ( .A(n10134), .ZN(n10135) );
  NAND2_X1 U11926 ( .A1(n10140), .A2(n11319), .ZN(n10141) );
  MUX2_X1 U11927 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n11277), .Z(n10143) );
  NAND2_X1 U11928 ( .A1(n10143), .A2(SI_13_), .ZN(n10162) );
  INV_X1 U11929 ( .A(n10143), .ZN(n10144) );
  NAND2_X1 U11930 ( .A1(n10144), .A2(n11452), .ZN(n10145) );
  NAND2_X1 U11931 ( .A1(n10162), .A2(n10145), .ZN(n10146) );
  NAND2_X1 U11932 ( .A1(n10147), .A2(n10146), .ZN(n10148) );
  NAND2_X1 U11933 ( .A1(n10163), .A2(n10148), .ZN(n11699) );
  OR2_X1 U11934 ( .A1(n11699), .A2(n10208), .ZN(n10153) );
  NOR2_X1 U11935 ( .A1(n10149), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n10164) );
  INV_X1 U11936 ( .A(n10164), .ZN(n10150) );
  NAND2_X1 U11937 ( .A1(n10150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10151) );
  XNOR2_X1 U11938 ( .A(n10151), .B(P2_IR_REG_13__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U11939 ( .A1(n9944), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9909), 
        .B2(n13105), .ZN(n10152) );
  NAND2_X1 U11940 ( .A1(n9950), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10158) );
  INV_X1 U11941 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13130) );
  OR2_X1 U11942 ( .A1(n9887), .A2(n13130), .ZN(n10157) );
  XNOR2_X1 U11943 ( .A(n10171), .B(n13181), .ZN(n13180) );
  OR2_X1 U11944 ( .A1(n13180), .A2(n10463), .ZN(n10156) );
  INV_X1 U11945 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10154) );
  OR2_X1 U11946 ( .A1(n10494), .A2(n10154), .ZN(n10155) );
  OAI22_X1 U11947 ( .A1(n13240), .A2(n10220), .B1(n7420), .B2(n13284), .ZN(
        n10160) );
  OAI22_X1 U11948 ( .A1(n13240), .A2(n7420), .B1(n13284), .B2(n10220), .ZN(
        n10159) );
  INV_X1 U11949 ( .A(n10160), .ZN(n10161) );
  MUX2_X1 U11950 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n11277), .Z(n10184) );
  XNOR2_X1 U11951 ( .A(n10184), .B(SI_14_), .ZN(n10182) );
  XNOR2_X1 U11952 ( .A(n10183), .B(n10182), .ZN(n11842) );
  NAND2_X1 U11953 ( .A1(n11842), .A2(n10511), .ZN(n10169) );
  NAND2_X1 U11954 ( .A1(n10164), .A2(n7660), .ZN(n10166) );
  NAND2_X1 U11955 ( .A1(n10166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10165) );
  MUX2_X1 U11956 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10165), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n10167) );
  AND2_X1 U11957 ( .A1(n10167), .A2(n10209), .ZN(n13436) );
  AOI22_X1 U11958 ( .A1(n9944), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9909), 
        .B2(n13436), .ZN(n10168) );
  INV_X1 U11959 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10170) );
  OAI21_X1 U11960 ( .B1(n10171), .B2(n13181), .A(n10170), .ZN(n10172) );
  AND2_X1 U11961 ( .A1(n10172), .A2(n10191), .ZN(n13288) );
  NAND2_X1 U11962 ( .A1(n13288), .A2(n9840), .ZN(n10176) );
  NAND2_X1 U11963 ( .A1(n10514), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U11964 ( .A1(n9837), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U11965 ( .A1(n9950), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10173) );
  OAI22_X1 U11966 ( .A1(n13348), .A2(n10540), .B1(n13352), .B2(n10220), .ZN(
        n10178) );
  OAI22_X1 U11967 ( .A1(n13348), .A2(n10220), .B1(n7420), .B2(n13352), .ZN(
        n10180) );
  INV_X1 U11968 ( .A(n10177), .ZN(n10179) );
  INV_X1 U11969 ( .A(n10184), .ZN(n10185) );
  NAND2_X1 U11970 ( .A1(n10185), .A2(n11532), .ZN(n10186) );
  MUX2_X1 U11971 ( .A(n11995), .B(n8568), .S(n11277), .Z(n10203) );
  XNOR2_X1 U11972 ( .A(n10203), .B(SI_15_), .ZN(n10201) );
  XNOR2_X1 U11973 ( .A(n10202), .B(n10201), .ZN(n11993) );
  NAND2_X1 U11974 ( .A1(n11993), .A2(n10511), .ZN(n10189) );
  NAND2_X1 U11975 ( .A1(n10209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10187) );
  XNOR2_X1 U11976 ( .A(n10187), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15117) );
  AOI22_X1 U11977 ( .A1(n9944), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9909), 
        .B2(n15117), .ZN(n10188) );
  INV_X1 U11978 ( .A(n10191), .ZN(n10190) );
  INV_X1 U11979 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13438) );
  NAND2_X1 U11980 ( .A1(n10191), .A2(n13438), .ZN(n10192) );
  NAND2_X1 U11981 ( .A1(n10233), .A2(n10192), .ZN(n13458) );
  OR2_X1 U11982 ( .A1(n13458), .A2(n10463), .ZN(n10197) );
  INV_X1 U11983 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13357) );
  OR2_X1 U11984 ( .A1(n9887), .A2(n13357), .ZN(n10194) );
  INV_X1 U11985 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13497) );
  OR2_X1 U11986 ( .A1(n9888), .A2(n13497), .ZN(n10193) );
  AND2_X1 U11987 ( .A1(n10194), .A2(n10193), .ZN(n10196) );
  INV_X1 U11988 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13494) );
  OR2_X1 U11989 ( .A1(n10494), .A2(n13494), .ZN(n10195) );
  OAI22_X1 U11990 ( .A1(n15197), .A2(n10220), .B1(n7420), .B2(n15172), .ZN(
        n10198) );
  OAI22_X1 U11991 ( .A1(n15197), .A2(n10540), .B1(n15172), .B2(n10220), .ZN(
        n10200) );
  INV_X1 U11992 ( .A(n10198), .ZN(n10199) );
  MUX2_X1 U11993 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n11277), .Z(n10206) );
  NAND2_X1 U11994 ( .A1(n7527), .A2(n8644), .ZN(n10207) );
  NAND2_X1 U11995 ( .A1(n10227), .A2(n10207), .ZN(n12320) );
  OR2_X1 U11996 ( .A1(n12320), .A2(n10208), .ZN(n10214) );
  INV_X1 U11997 ( .A(n10209), .ZN(n10210) );
  NAND2_X1 U11998 ( .A1(n10210), .A2(n7662), .ZN(n10257) );
  NAND2_X1 U11999 ( .A1(n10257), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U12000 ( .A1(n10211), .A2(n10255), .ZN(n10228) );
  OR2_X1 U12001 ( .A1(n10211), .A2(n10255), .ZN(n10212) );
  AOI22_X1 U12002 ( .A1(n9944), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n16243), 
        .B2(n9909), .ZN(n10213) );
  XNOR2_X1 U12003 ( .A(n10233), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n15453) );
  NAND2_X1 U12004 ( .A1(n15453), .A2(n9840), .ZN(n10219) );
  INV_X1 U12005 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n15114) );
  NAND2_X1 U12006 ( .A1(n9950), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12007 ( .A1(n9837), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n10215) );
  OAI211_X1 U12008 ( .C1(n9887), .C2(n15114), .A(n10216), .B(n10215), .ZN(
        n10217) );
  INV_X1 U12009 ( .A(n10217), .ZN(n10218) );
  NAND2_X1 U12010 ( .A1(n10219), .A2(n10218), .ZN(n15175) );
  AOI22_X1 U12011 ( .A1(n15539), .A2(n10220), .B1(n7420), .B2(n15175), .ZN(
        n10221) );
  OR2_X1 U12012 ( .A1(n10222), .A2(n10221), .ZN(n10225) );
  INV_X1 U12013 ( .A(n15539), .ZN(n15457) );
  INV_X1 U12014 ( .A(n15175), .ZN(n15200) );
  OAI22_X1 U12015 ( .A1(n15457), .A2(n10220), .B1(n7420), .B2(n15200), .ZN(
        n10224) );
  MUX2_X1 U12016 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n11277), .Z(n10247) );
  XNOR2_X1 U12017 ( .A(n10247), .B(SI_17_), .ZN(n10246) );
  XNOR2_X1 U12018 ( .A(n10245), .B(n10246), .ZN(n12566) );
  NAND2_X1 U12019 ( .A1(n12566), .A2(n10511), .ZN(n10231) );
  NAND2_X1 U12020 ( .A1(n10228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10229) );
  XNOR2_X1 U12021 ( .A(n10229), .B(P2_IR_REG_17__SCAN_IN), .ZN(n16255) );
  AOI22_X1 U12022 ( .A1(n16255), .A2(n9909), .B1(n9944), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n10230) );
  INV_X1 U12023 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10239) );
  INV_X1 U12024 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13406) );
  INV_X1 U12025 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10232) );
  OAI21_X1 U12026 ( .B1(n10233), .B2(n13406), .A(n10232), .ZN(n10236) );
  INV_X1 U12027 ( .A(n10233), .ZN(n10235) );
  NAND2_X1 U12028 ( .A1(n10235), .A2(n10234), .ZN(n10261) );
  NAND2_X1 U12029 ( .A1(n10236), .A2(n10261), .ZN(n15428) );
  OR2_X1 U12030 ( .A1(n15428), .A2(n10463), .ZN(n10238) );
  AOI22_X1 U12031 ( .A1(n10514), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9950), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n10237) );
  OAI211_X1 U12032 ( .C1(n10494), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n15177) );
  AOI22_X1 U12033 ( .A1(n15598), .A2(n7420), .B1(n10220), .B2(n15177), .ZN(
        n10241) );
  INV_X1 U12034 ( .A(n15598), .ZN(n15430) );
  INV_X1 U12035 ( .A(n15177), .ZN(n15202) );
  OAI22_X1 U12036 ( .A1(n15430), .A2(n10540), .B1(n15202), .B2(n10220), .ZN(
        n10240) );
  OAI21_X1 U12037 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(n10244) );
  NAND2_X1 U12038 ( .A1(n10244), .A2(n10243), .ZN(n10268) );
  INV_X1 U12039 ( .A(n10246), .ZN(n10249) );
  NOR2_X1 U12040 ( .A1(n10247), .A2(SI_17_), .ZN(n10248) );
  NAND2_X1 U12041 ( .A1(n10251), .A2(SI_18_), .ZN(n10274) );
  MUX2_X1 U12042 ( .A(n12878), .B(n8554), .S(n11277), .Z(n10254) );
  NAND2_X1 U12043 ( .A1(n12847), .A2(n10511), .ZN(n10260) );
  NAND2_X1 U12044 ( .A1(n10255), .A2(n9791), .ZN(n10256) );
  OAI21_X1 U12045 ( .B1(n10257), .B2(n10256), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n10258) );
  XNOR2_X1 U12046 ( .A(n10258), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U12047 ( .A1(n15123), .A2(n9909), .B1(n9944), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12048 ( .A1(n10261), .A2(n15127), .ZN(n10262) );
  AND2_X1 U12049 ( .A1(n10280), .A2(n10262), .ZN(n15410) );
  NAND2_X1 U12050 ( .A1(n15410), .A2(n9840), .ZN(n10265) );
  AOI22_X1 U12051 ( .A1(n10514), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9950), 
        .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n10264) );
  NAND2_X1 U12052 ( .A1(n9837), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U12053 ( .A1(n10268), .A2(n10269), .ZN(n10267) );
  OAI22_X1 U12054 ( .A1(n15595), .A2(n10499), .B1(n7420), .B2(n15203), .ZN(
        n10266) );
  NAND2_X1 U12055 ( .A1(n10267), .A2(n10266), .ZN(n10273) );
  INV_X1 U12056 ( .A(n10268), .ZN(n10271) );
  INV_X1 U12057 ( .A(n10269), .ZN(n10270) );
  NAND2_X1 U12058 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  NAND2_X1 U12059 ( .A1(n10273), .A2(n10272), .ZN(n10289) );
  MUX2_X1 U12060 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n11277), .Z(n10295) );
  XNOR2_X1 U12061 ( .A(n10295), .B(SI_19_), .ZN(n10296) );
  XNOR2_X1 U12062 ( .A(n10297), .B(n10296), .ZN(n13025) );
  NAND2_X1 U12063 ( .A1(n13025), .A2(n10511), .ZN(n10277) );
  AOI22_X1 U12064 ( .A1(n9944), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10515), 
        .B2(n9909), .ZN(n10276) );
  INV_X1 U12065 ( .A(n10280), .ZN(n10278) );
  NAND2_X1 U12066 ( .A1(n10278), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n10301) );
  INV_X1 U12067 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U12068 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  NAND2_X1 U12069 ( .A1(n10301), .A2(n10281), .ZN(n15387) );
  OR2_X1 U12070 ( .A1(n15387), .A2(n10463), .ZN(n10286) );
  INV_X1 U12071 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n15388) );
  NAND2_X1 U12072 ( .A1(n9950), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12073 ( .A1(n9837), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n10282) );
  OAI211_X1 U12074 ( .C1(n9887), .C2(n15388), .A(n10283), .B(n10282), .ZN(
        n10284) );
  INV_X1 U12075 ( .A(n10284), .ZN(n10285) );
  OAI22_X1 U12076 ( .A1(n15590), .A2(n10499), .B1(n7420), .B2(n15181), .ZN(
        n10290) );
  NAND2_X1 U12077 ( .A1(n10289), .A2(n10290), .ZN(n10288) );
  OAI22_X1 U12078 ( .A1(n15590), .A2(n10540), .B1(n15181), .B2(n10499), .ZN(
        n10287) );
  NAND2_X1 U12079 ( .A1(n10288), .A2(n10287), .ZN(n10294) );
  INV_X1 U12080 ( .A(n10289), .ZN(n10292) );
  INV_X1 U12081 ( .A(n10290), .ZN(n10291) );
  NAND2_X1 U12082 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  NAND2_X1 U12083 ( .A1(n10294), .A2(n10293), .ZN(n10311) );
  MUX2_X1 U12084 ( .A(n13118), .B(n13167), .S(n11277), .Z(n10312) );
  XNOR2_X1 U12085 ( .A(n10312), .B(SI_20_), .ZN(n10298) );
  XNOR2_X1 U12086 ( .A(n10314), .B(n10298), .ZN(n13116) );
  NAND2_X1 U12087 ( .A1(n13116), .A2(n10511), .ZN(n10300) );
  NAND2_X1 U12088 ( .A1(n9944), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n10299) );
  AND2_X2 U12089 ( .A1(n10300), .A2(n10299), .ZN(n15585) );
  INV_X1 U12090 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U12091 ( .A1(n10301), .A2(n15044), .ZN(n10302) );
  AND2_X1 U12092 ( .A1(n10318), .A2(n10302), .ZN(n15373) );
  NAND2_X1 U12093 ( .A1(n15373), .A2(n9840), .ZN(n10308) );
  INV_X1 U12094 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12095 ( .A1(n9950), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12096 ( .A1(n10514), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n10303) );
  OAI211_X1 U12097 ( .C1(n10305), .C2(n10494), .A(n10304), .B(n10303), .ZN(
        n10306) );
  INV_X1 U12098 ( .A(n10306), .ZN(n10307) );
  OAI22_X1 U12099 ( .A1(n15585), .A2(n10540), .B1(n15183), .B2(n10220), .ZN(
        n10310) );
  OAI22_X1 U12100 ( .A1(n15585), .A2(n10499), .B1(n10540), .B2(n15183), .ZN(
        n10309) );
  MUX2_X1 U12101 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n11277), .Z(n10330) );
  XNOR2_X1 U12102 ( .A(n10330), .B(SI_21_), .ZN(n10328) );
  XNOR2_X1 U12103 ( .A(n10329), .B(n10328), .ZN(n13703) );
  NAND2_X1 U12104 ( .A1(n13703), .A2(n10511), .ZN(n10316) );
  NAND2_X1 U12105 ( .A1(n9944), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n10315) );
  INV_X1 U12106 ( .A(n10318), .ZN(n10317) );
  NAND2_X1 U12107 ( .A1(n10317), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n10333) );
  INV_X1 U12108 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14999) );
  NAND2_X1 U12109 ( .A1(n10318), .A2(n14999), .ZN(n10319) );
  NAND2_X1 U12110 ( .A1(n10333), .A2(n10319), .ZN(n14998) );
  OR2_X1 U12111 ( .A1(n14998), .A2(n10463), .ZN(n10325) );
  INV_X1 U12112 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U12113 ( .A1(n10514), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U12114 ( .A1(n9950), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n10320) );
  OAI211_X1 U12115 ( .C1(n10494), .C2(n10322), .A(n10321), .B(n10320), .ZN(
        n10323) );
  INV_X1 U12116 ( .A(n10323), .ZN(n10324) );
  OAI22_X1 U12117 ( .A1(n15360), .A2(n10220), .B1(n7420), .B2(n15184), .ZN(
        n10326) );
  OAI22_X1 U12118 ( .A1(n15360), .A2(n10540), .B1(n15184), .B2(n10220), .ZN(
        n10327) );
  XNOR2_X1 U12119 ( .A(n10346), .B(SI_22_), .ZN(n13710) );
  MUX2_X1 U12120 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n11277), .Z(n10347) );
  XNOR2_X1 U12121 ( .A(n13710), .B(n10347), .ZN(n13430) );
  NAND2_X1 U12122 ( .A1(n13430), .A2(n10511), .ZN(n10332) );
  NAND2_X1 U12123 ( .A1(n9944), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n10331) );
  INV_X1 U12124 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n15053) );
  NAND2_X1 U12125 ( .A1(n10333), .A2(n15053), .ZN(n10334) );
  NAND2_X1 U12126 ( .A1(n10359), .A2(n10334), .ZN(n15343) );
  OR2_X1 U12127 ( .A1(n15343), .A2(n10463), .ZN(n10339) );
  INV_X1 U12128 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15508) );
  NAND2_X1 U12129 ( .A1(n9950), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U12130 ( .A1(n10514), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n10335) );
  OAI211_X1 U12131 ( .C1(n15508), .C2(n10494), .A(n10336), .B(n10335), .ZN(
        n10337) );
  INV_X1 U12132 ( .A(n10337), .ZN(n10338) );
  NAND2_X1 U12133 ( .A1(n10339), .A2(n10338), .ZN(n15215) );
  AOI22_X1 U12134 ( .A1(n15342), .A2(n10220), .B1(n7420), .B2(n15215), .ZN(
        n10341) );
  INV_X1 U12135 ( .A(n15215), .ZN(n15214) );
  OAI22_X1 U12136 ( .A1(n15580), .A2(n10499), .B1(n10540), .B2(n15214), .ZN(
        n10340) );
  INV_X1 U12137 ( .A(n10347), .ZN(n10344) );
  NAND2_X1 U12138 ( .A1(n10344), .A2(n10343), .ZN(n10345) );
  NAND2_X1 U12139 ( .A1(n10346), .A2(n10345), .ZN(n10349) );
  NAND2_X1 U12140 ( .A1(n10347), .A2(SI_22_), .ZN(n10348) );
  MUX2_X1 U12141 ( .A(n13339), .B(n13730), .S(n11277), .Z(n10350) );
  NAND2_X1 U12142 ( .A1(n10350), .A2(n9618), .ZN(n10369) );
  INV_X1 U12143 ( .A(n10350), .ZN(n10351) );
  NAND2_X1 U12144 ( .A1(n10351), .A2(SI_23_), .ZN(n10352) );
  NAND2_X1 U12145 ( .A1(n10369), .A2(n10352), .ZN(n10353) );
  NAND2_X1 U12146 ( .A1(n10354), .A2(n10353), .ZN(n10355) );
  NAND2_X1 U12147 ( .A1(n10370), .A2(n10355), .ZN(n13729) );
  NAND2_X1 U12148 ( .A1(n13729), .A2(n10511), .ZN(n10357) );
  NAND2_X1 U12149 ( .A1(n9944), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n10356) );
  AND2_X2 U12150 ( .A1(n10357), .A2(n10356), .ZN(n15576) );
  NAND2_X1 U12151 ( .A1(n10359), .A2(n10358), .ZN(n10360) );
  AND2_X1 U12152 ( .A1(n10375), .A2(n10360), .ZN(n15329) );
  NAND2_X1 U12153 ( .A1(n15329), .A2(n9840), .ZN(n10366) );
  INV_X1 U12154 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10363) );
  NAND2_X1 U12155 ( .A1(n9950), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U12156 ( .A1(n10514), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n10361) );
  OAI211_X1 U12157 ( .C1(n10363), .C2(n10494), .A(n10362), .B(n10361), .ZN(
        n10364) );
  INV_X1 U12158 ( .A(n10364), .ZN(n10365) );
  INV_X1 U12159 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13514) );
  MUX2_X1 U12160 ( .A(n13514), .B(n13750), .S(n11277), .Z(n10388) );
  XNOR2_X1 U12161 ( .A(n10388), .B(SI_24_), .ZN(n10371) );
  XNOR2_X1 U12162 ( .A(n10391), .B(n10371), .ZN(n13749) );
  NAND2_X1 U12163 ( .A1(n13749), .A2(n7423), .ZN(n10373) );
  NAND2_X1 U12164 ( .A1(n9944), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n10372) );
  INV_X1 U12165 ( .A(n10375), .ZN(n10374) );
  NAND2_X1 U12166 ( .A1(n10374), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n10399) );
  INV_X1 U12167 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15031) );
  NAND2_X1 U12168 ( .A1(n10375), .A2(n15031), .ZN(n10376) );
  NAND2_X1 U12169 ( .A1(n10399), .A2(n10376), .ZN(n15314) );
  OR2_X1 U12170 ( .A1(n15314), .A2(n10463), .ZN(n10382) );
  INV_X1 U12171 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U12172 ( .A1(n9950), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U12173 ( .A1(n10514), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n10377) );
  OAI211_X1 U12174 ( .C1(n10379), .C2(n10494), .A(n10378), .B(n10377), .ZN(
        n10380) );
  INV_X1 U12175 ( .A(n10380), .ZN(n10381) );
  NAND2_X1 U12176 ( .A1(n10382), .A2(n10381), .ZN(n15191) );
  AOI22_X1 U12177 ( .A1(n15496), .A2(n10220), .B1(n7420), .B2(n15191), .ZN(
        n10384) );
  INV_X1 U12178 ( .A(n15191), .ZN(n15010) );
  OAI22_X1 U12179 ( .A1(n15572), .A2(n10499), .B1(n10540), .B2(n15010), .ZN(
        n10383) );
  OAI21_X1 U12180 ( .B1(n10385), .B2(n10384), .A(n10383), .ZN(n10387) );
  NAND2_X1 U12181 ( .A1(n10387), .A2(n10386), .ZN(n10409) );
  INV_X1 U12182 ( .A(n10388), .ZN(n10389) );
  NAND2_X1 U12183 ( .A1(n10390), .A2(n10389), .ZN(n10392) );
  MUX2_X1 U12184 ( .A(n15627), .B(n16179), .S(n11277), .Z(n10393) );
  NAND2_X1 U12185 ( .A1(n10393), .A2(n13303), .ZN(n10414) );
  INV_X1 U12186 ( .A(n10393), .ZN(n10394) );
  NAND2_X1 U12187 ( .A1(n10394), .A2(SI_25_), .ZN(n10395) );
  NAND2_X1 U12188 ( .A1(n10414), .A2(n10395), .ZN(n10411) );
  XNOR2_X1 U12189 ( .A(n10410), .B(n10411), .ZN(n15624) );
  NAND2_X1 U12190 ( .A1(n15624), .A2(n7423), .ZN(n10397) );
  NAND2_X1 U12191 ( .A1(n9944), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10396) );
  INV_X1 U12192 ( .A(n10399), .ZN(n10398) );
  NAND2_X1 U12193 ( .A1(n10398), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n10419) );
  INV_X1 U12194 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U12195 ( .A1(n10399), .A2(n15011), .ZN(n10400) );
  NAND2_X1 U12196 ( .A1(n10419), .A2(n10400), .ZN(n15297) );
  OR2_X1 U12197 ( .A1(n15297), .A2(n10463), .ZN(n10405) );
  INV_X1 U12198 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15490) );
  NAND2_X1 U12199 ( .A1(n10514), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U12200 ( .A1(n9950), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10401) );
  OAI211_X1 U12201 ( .C1(n15490), .C2(n10494), .A(n10402), .B(n10401), .ZN(
        n10403) );
  INV_X1 U12202 ( .A(n10403), .ZN(n10404) );
  NAND2_X1 U12203 ( .A1(n10405), .A2(n10404), .ZN(n15084) );
  AOI22_X1 U12204 ( .A1(n15299), .A2(n7420), .B1(n15084), .B2(n10220), .ZN(
        n10408) );
  INV_X1 U12205 ( .A(n10408), .ZN(n10407) );
  AOI22_X1 U12206 ( .A1(n15299), .A2(n10220), .B1(n7420), .B2(n15084), .ZN(
        n10406) );
  INV_X1 U12207 ( .A(n10410), .ZN(n10413) );
  INV_X1 U12208 ( .A(n10411), .ZN(n10412) );
  NAND2_X1 U12209 ( .A1(n10413), .A2(n10412), .ZN(n10415) );
  MUX2_X1 U12210 ( .A(n15623), .B(n8126), .S(n11277), .Z(n10428) );
  XNOR2_X1 U12211 ( .A(n10428), .B(SI_26_), .ZN(n10427) );
  XNOR2_X1 U12212 ( .A(n10432), .B(n10427), .ZN(n15621) );
  NAND2_X1 U12213 ( .A1(n15621), .A2(n10511), .ZN(n10417) );
  NAND2_X1 U12214 ( .A1(n9944), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10416) );
  INV_X1 U12215 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U12216 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  NAND2_X1 U12217 ( .A1(n15281), .A2(n9840), .ZN(n10426) );
  INV_X1 U12218 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10423) );
  NAND2_X1 U12219 ( .A1(n9950), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U12220 ( .A1(n10514), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n10421) );
  OAI211_X1 U12221 ( .C1(n10423), .C2(n10494), .A(n10422), .B(n10421), .ZN(
        n10424) );
  INV_X1 U12222 ( .A(n10424), .ZN(n10425) );
  AOI22_X1 U12223 ( .A1(n15483), .A2(n7420), .B1(n10220), .B2(n15219), .ZN(
        n10504) );
  OAI22_X1 U12224 ( .A1(n15284), .A2(n10540), .B1(n15192), .B2(n10499), .ZN(
        n10503) );
  INV_X1 U12225 ( .A(n10427), .ZN(n10431) );
  INV_X1 U12226 ( .A(n10428), .ZN(n10429) );
  NAND2_X1 U12227 ( .A1(n10429), .A2(SI_26_), .ZN(n10430) );
  MUX2_X1 U12228 ( .A(n15620), .B(n16172), .S(n11277), .Z(n10433) );
  NAND2_X1 U12229 ( .A1(n10433), .A2(n14964), .ZN(n10436) );
  INV_X1 U12230 ( .A(n10433), .ZN(n10434) );
  NAND2_X1 U12231 ( .A1(n10434), .A2(SI_27_), .ZN(n10435) );
  NAND2_X1 U12232 ( .A1(n10436), .A2(n10435), .ZN(n10487) );
  MUX2_X1 U12233 ( .A(n15616), .B(n13802), .S(n11277), .Z(n10437) );
  NAND2_X1 U12234 ( .A1(n10437), .A2(n13916), .ZN(n10459) );
  INV_X1 U12235 ( .A(n10437), .ZN(n10438) );
  NAND2_X1 U12236 ( .A1(n10438), .A2(SI_28_), .ZN(n10439) );
  INV_X1 U12237 ( .A(n10440), .ZN(n10441) );
  NAND2_X1 U12238 ( .A1(n10441), .A2(n7634), .ZN(n10442) );
  NAND2_X1 U12239 ( .A1(n15613), .A2(n7423), .ZN(n10444) );
  NAND2_X1 U12240 ( .A1(n9944), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10443) );
  INV_X1 U12241 ( .A(n10491), .ZN(n10446) );
  AND2_X1 U12242 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n10445) );
  NAND2_X1 U12243 ( .A1(n10446), .A2(n10445), .ZN(n15234) );
  INV_X1 U12244 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10448) );
  INV_X1 U12245 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10447) );
  OAI21_X1 U12246 ( .B1(n10491), .B2(n10448), .A(n10447), .ZN(n10449) );
  NAND2_X1 U12247 ( .A1(n15234), .A2(n10449), .ZN(n15255) );
  OR2_X1 U12248 ( .A1(n15255), .A2(n10463), .ZN(n10455) );
  INV_X1 U12249 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12250 ( .A1(n9950), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U12251 ( .A1(n10514), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n10450) );
  OAI211_X1 U12252 ( .C1(n10452), .C2(n10494), .A(n10451), .B(n10450), .ZN(
        n10453) );
  INV_X1 U12253 ( .A(n10453), .ZN(n10454) );
  AND2_X1 U12254 ( .A1(n15226), .A2(n10499), .ZN(n10456) );
  AOI21_X1 U12255 ( .B1(n15474), .B2(n7420), .A(n10456), .ZN(n10526) );
  NAND2_X1 U12256 ( .A1(n15474), .A2(n10499), .ZN(n10458) );
  NAND2_X1 U12257 ( .A1(n15226), .A2(n7420), .ZN(n10457) );
  NAND2_X1 U12258 ( .A1(n10458), .A2(n10457), .ZN(n10525) );
  MUX2_X1 U12259 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n11277), .Z(n10473) );
  XNOR2_X1 U12260 ( .A(n10473), .B(n14960), .ZN(n10471) );
  XNOR2_X1 U12261 ( .A(n10472), .B(n10471), .ZN(n13567) );
  NAND2_X1 U12262 ( .A1(n13567), .A2(n7423), .ZN(n10462) );
  NAND2_X1 U12263 ( .A1(n9944), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10461) );
  OR2_X1 U12264 ( .A1(n15234), .A2(n10463), .ZN(n10469) );
  INV_X1 U12265 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U12266 ( .A1(n9950), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U12267 ( .A1(n10514), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10464) );
  OAI211_X1 U12268 ( .C1(n10466), .C2(n10494), .A(n10465), .B(n10464), .ZN(
        n10467) );
  INV_X1 U12269 ( .A(n10467), .ZN(n10468) );
  AND2_X1 U12270 ( .A1(n10469), .A2(n10468), .ZN(n10470) );
  OAI22_X1 U12271 ( .A1(n15470), .A2(n10499), .B1(n7420), .B2(n10470), .ZN(
        n10519) );
  AOI22_X1 U12272 ( .A1(n15236), .A2(n10220), .B1(n7420), .B2(n15083), .ZN(
        n10520) );
  NOR2_X1 U12273 ( .A1(n10519), .A2(n10520), .ZN(n10527) );
  INV_X1 U12274 ( .A(n10473), .ZN(n10474) );
  NAND2_X1 U12275 ( .A1(n10474), .A2(n14960), .ZN(n10475) );
  MUX2_X1 U12276 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n11277), .Z(n10476) );
  NAND2_X1 U12277 ( .A1(n10476), .A2(SI_30_), .ZN(n10479) );
  INV_X1 U12278 ( .A(n10476), .ZN(n10477) );
  INV_X1 U12279 ( .A(SI_30_), .ZN(n14955) );
  NAND2_X1 U12280 ( .A1(n10477), .A2(n14955), .ZN(n10478) );
  NAND2_X1 U12281 ( .A1(n10479), .A2(n10478), .ZN(n10507) );
  MUX2_X1 U12282 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n11277), .Z(n10480) );
  XNOR2_X1 U12283 ( .A(n10480), .B(SI_31_), .ZN(n10481) );
  NAND2_X1 U12284 ( .A1(n9944), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n10482) );
  INV_X1 U12285 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10483) );
  OR2_X1 U12286 ( .A1(n10494), .A2(n10483), .ZN(n10486) );
  INV_X1 U12287 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n15158) );
  OR2_X1 U12288 ( .A1(n9887), .A2(n15158), .ZN(n10485) );
  INV_X1 U12289 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n15554) );
  OR2_X1 U12290 ( .A1(n9888), .A2(n15554), .ZN(n10484) );
  AND3_X1 U12291 ( .A1(n10486), .A2(n10485), .A3(n10484), .ZN(n10524) );
  NAND2_X1 U12292 ( .A1(n16169), .A2(n7423), .ZN(n10490) );
  NAND2_X1 U12293 ( .A1(n9944), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10489) );
  XNOR2_X1 U12294 ( .A(n10491), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n15264) );
  NAND2_X1 U12295 ( .A1(n15264), .A2(n9840), .ZN(n10498) );
  INV_X1 U12296 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10495) );
  NAND2_X1 U12297 ( .A1(n9950), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10493) );
  NAND2_X1 U12298 ( .A1(n10514), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n10492) );
  OAI211_X1 U12299 ( .C1(n10495), .C2(n10494), .A(n10493), .B(n10492), .ZN(
        n10496) );
  INV_X1 U12300 ( .A(n10496), .ZN(n10497) );
  AND2_X1 U12301 ( .A1(n15193), .A2(n10499), .ZN(n10500) );
  AOI21_X1 U12302 ( .B1(n15478), .B2(n7420), .A(n10500), .ZN(n10528) );
  NAND2_X1 U12303 ( .A1(n15478), .A2(n10220), .ZN(n10502) );
  NAND2_X1 U12304 ( .A1(n15193), .A2(n7420), .ZN(n10501) );
  NAND2_X1 U12305 ( .A1(n10502), .A2(n10501), .ZN(n10529) );
  AOI22_X1 U12306 ( .A1(n10528), .A2(n10529), .B1(n10504), .B2(n10503), .ZN(
        n10505) );
  NAND2_X1 U12307 ( .A1(n10508), .A2(n10507), .ZN(n10509) );
  NAND2_X1 U12308 ( .A1(n13919), .A2(n10511), .ZN(n10513) );
  NAND2_X1 U12309 ( .A1(n9944), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10512) );
  AOI222_X1 U12310 ( .A1(n9837), .A2(P2_REG1_REG_30__SCAN_IN), .B1(n10514), 
        .B2(P2_REG2_REG_30__SCAN_IN), .C1(n9950), .C2(P2_REG0_REG_30__SCAN_IN), 
        .ZN(n10570) );
  OAI22_X1 U12311 ( .A1(n15560), .A2(n7420), .B1(n10570), .B2(n10499), .ZN(
        n10537) );
  INV_X1 U12312 ( .A(n10570), .ZN(n15228) );
  NAND2_X1 U12313 ( .A1(n15163), .A2(n10499), .ZN(n10541) );
  NAND2_X1 U12314 ( .A1(n11922), .A2(n13431), .ZN(n10551) );
  NAND3_X1 U12315 ( .A1(n10541), .A2(n10517), .A3(n10551), .ZN(n10518) );
  AOI22_X1 U12316 ( .A1(n15467), .A2(n7420), .B1(n15228), .B2(n10518), .ZN(
        n10536) );
  INV_X1 U12317 ( .A(n10519), .ZN(n10522) );
  INV_X1 U12318 ( .A(n10520), .ZN(n10521) );
  OAI22_X1 U12319 ( .A1(n10537), .A2(n10536), .B1(n10522), .B2(n10521), .ZN(
        n10535) );
  MUX2_X1 U12320 ( .A(n15163), .B(n10540), .S(n15552), .Z(n10523) );
  OAI21_X1 U12321 ( .B1(n10524), .B2(n10220), .A(n10523), .ZN(n10534) );
  NOR4_X1 U12322 ( .A1(n10571), .A2(n10527), .A3(n10526), .A4(n10525), .ZN(
        n10533) );
  INV_X1 U12323 ( .A(n10528), .ZN(n10531) );
  INV_X1 U12324 ( .A(n10529), .ZN(n10530) );
  NAND2_X1 U12325 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  NAND2_X1 U12326 ( .A1(n15163), .A2(n10540), .ZN(n10543) );
  NAND2_X1 U12327 ( .A1(n10541), .A2(n10220), .ZN(n10542) );
  MUX2_X1 U12328 ( .A(n10543), .B(n10542), .S(n15552), .Z(n10544) );
  INV_X1 U12329 ( .A(n11685), .ZN(n10567) );
  NOR2_X1 U12330 ( .A1(n11662), .A2(n13431), .ZN(n10546) );
  AOI211_X1 U12331 ( .C1(n11248), .C2(n13027), .A(n10567), .B(n10546), .ZN(
        n10547) );
  NAND2_X1 U12332 ( .A1(n10556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U12333 ( .A1(n10607), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13337) );
  INV_X1 U12334 ( .A(n13337), .ZN(n10555) );
  INV_X1 U12335 ( .A(n10551), .ZN(n10553) );
  INV_X1 U12336 ( .A(n11248), .ZN(n13257) );
  NOR3_X1 U12337 ( .A1(n13117), .A2(n13257), .A3(n13027), .ZN(n10552) );
  NOR2_X1 U12338 ( .A1(n10553), .A2(n10552), .ZN(n10554) );
  NAND2_X1 U12339 ( .A1(n10565), .A2(n10564), .ZN(n10557) );
  INV_X1 U12340 ( .A(n15160), .ZN(n11467) );
  INV_X1 U12341 ( .A(n10566), .ZN(n11463) );
  NAND4_X1 U12342 ( .A1(n16223), .A2(n10567), .A3(n11467), .A4(n15225), .ZN(
        n10568) );
  OAI211_X1 U12343 ( .C1(n13431), .C2(n13337), .A(n10568), .B(P2_B_REG_SCAN_IN), .ZN(n10592) );
  XOR2_X1 U12344 ( .A(n15467), .B(n10570), .Z(n10588) );
  INV_X1 U12345 ( .A(n10571), .ZN(n10587) );
  INV_X1 U12346 ( .A(n15474), .ZN(n15248) );
  NAND2_X1 U12347 ( .A1(n15248), .A2(n15226), .ZN(n15221) );
  INV_X1 U12348 ( .A(n15226), .ZN(n10572) );
  NAND2_X1 U12349 ( .A1(n15474), .A2(n10572), .ZN(n10573) );
  NAND2_X1 U12350 ( .A1(n15221), .A2(n10573), .ZN(n15241) );
  XNOR2_X1 U12351 ( .A(n15478), .B(n15220), .ZN(n15268) );
  XNOR2_X1 U12352 ( .A(n15483), .B(n15192), .ZN(n15276) );
  XNOR2_X1 U12353 ( .A(n15299), .B(n15084), .ZN(n15289) );
  NAND2_X1 U12354 ( .A1(n15496), .A2(n15010), .ZN(n15217) );
  OR2_X1 U12355 ( .A1(n15496), .A2(n15010), .ZN(n10574) );
  NAND2_X1 U12356 ( .A1(n15217), .A2(n10574), .ZN(n15306) );
  XNOR2_X1 U12357 ( .A(n15503), .B(n15188), .ZN(n15333) );
  XNOR2_X1 U12358 ( .A(n8227), .B(n15184), .ZN(n15362) );
  INV_X1 U12359 ( .A(n15585), .ZN(n15518) );
  INV_X1 U12360 ( .A(n15183), .ZN(n15210) );
  XNOR2_X1 U12361 ( .A(n15518), .B(n15210), .ZN(n15375) );
  XNOR2_X1 U12362 ( .A(n15598), .B(n15202), .ZN(n15418) );
  XNOR2_X1 U12363 ( .A(n15539), .B(n15200), .ZN(n15437) );
  XNOR2_X1 U12364 ( .A(n13463), .B(n15172), .ZN(n13350) );
  XNOR2_X1 U12365 ( .A(n15545), .B(n15085), .ZN(n13232) );
  XNOR2_X1 U12366 ( .A(n12853), .B(n12921), .ZN(n12913) );
  XNOR2_X1 U12367 ( .A(n13052), .B(n13072), .ZN(n12978) );
  XNOR2_X1 U12368 ( .A(n12521), .B(n15091), .ZN(n12608) );
  INV_X1 U12369 ( .A(n11942), .ZN(n15095) );
  NAND2_X1 U12370 ( .A1(n11968), .A2(n11969), .ZN(n11949) );
  INV_X1 U12371 ( .A(n11968), .ZN(n15022) );
  INV_X1 U12372 ( .A(n11969), .ZN(n15094) );
  NAND2_X1 U12373 ( .A1(n15022), .A2(n15094), .ZN(n11952) );
  NAND2_X1 U12374 ( .A1(n11949), .A2(n11952), .ZN(n11941) );
  NAND2_X1 U12375 ( .A1(n9875), .A2(n14066), .ZN(n10576) );
  INV_X1 U12376 ( .A(n15099), .ZN(n11227) );
  NAND2_X1 U12377 ( .A1(n11227), .A2(n11919), .ZN(n11224) );
  NAND4_X1 U12378 ( .A1(n11941), .A2(n11716), .A3(n12204), .A4(n10569), .ZN(
        n10577) );
  INV_X1 U12379 ( .A(n11832), .ZN(n15096) );
  NOR4_X1 U12380 ( .A1(n11935), .A2(n12102), .A3(n10577), .A4(n11827), .ZN(
        n10578) );
  XNOR2_X1 U12381 ( .A(n12488), .B(n15092), .ZN(n12298) );
  XNOR2_X1 U12382 ( .A(n12296), .B(n15093), .ZN(n12293) );
  NAND4_X1 U12383 ( .A1(n12608), .A2(n10578), .A3(n12298), .A4(n12293), .ZN(
        n10579) );
  NOR4_X1 U12384 ( .A1(n12913), .A2(n12978), .A3(n12638), .A4(n10579), .ZN(
        n10580) );
  XNOR2_X1 U12385 ( .A(n13191), .B(n15087), .ZN(n12982) );
  XNOR2_X1 U12386 ( .A(n13274), .B(n15086), .ZN(n13237) );
  NAND4_X1 U12387 ( .A1(n13232), .A2(n10580), .A3(n12982), .A4(n13237), .ZN(
        n10581) );
  NOR4_X1 U12388 ( .A1(n15418), .A2(n15437), .A3(n13350), .A4(n10581), .ZN(
        n10582) );
  INV_X1 U12389 ( .A(n15590), .ZN(n15386) );
  INV_X1 U12390 ( .A(n15181), .ZN(n15208) );
  XNOR2_X1 U12391 ( .A(n15386), .B(n15208), .ZN(n15391) );
  INV_X1 U12392 ( .A(n15595), .ZN(n15409) );
  INV_X1 U12393 ( .A(n15203), .ZN(n15205) );
  XNOR2_X1 U12394 ( .A(n15409), .B(n15205), .ZN(n15403) );
  NAND4_X1 U12395 ( .A1(n15375), .A2(n10582), .A3(n15391), .A4(n15403), .ZN(
        n10583) );
  NOR4_X1 U12396 ( .A1(n15306), .A2(n15333), .A3(n15362), .A4(n10583), .ZN(
        n10584) );
  XNOR2_X1 U12397 ( .A(n15342), .B(n15215), .ZN(n15348) );
  NAND3_X1 U12398 ( .A1(n15289), .A2(n10584), .A3(n15348), .ZN(n10585) );
  NOR4_X1 U12399 ( .A1(n15241), .A2(n15268), .A3(n15276), .A4(n10585), .ZN(
        n10586) );
  XNOR2_X1 U12400 ( .A(n15236), .B(n15083), .ZN(n15222) );
  NAND4_X1 U12401 ( .A1(n10588), .A2(n10587), .A3(n10586), .A4(n15222), .ZN(
        n10589) );
  XOR2_X1 U12402 ( .A(n10515), .B(n10589), .Z(n10590) );
  NOR3_X1 U12403 ( .A1(n10590), .A2(n11248), .A3(n13337), .ZN(n10591) );
  XNOR2_X1 U12404 ( .A(n14946), .B(n12266), .ZN(n10595) );
  AND2_X1 U12405 ( .A1(n10593), .A2(n12135), .ZN(n10594) );
  AND2_X1 U12406 ( .A1(n10595), .A2(n10594), .ZN(n12670) );
  NAND2_X1 U12407 ( .A1(n10596), .A2(n14451), .ZN(n12665) );
  OR2_X1 U12408 ( .A1(n14451), .A2(n10597), .ZN(n12664) );
  NAND2_X1 U12409 ( .A1(n12665), .A2(n12664), .ZN(n10598) );
  NAND2_X1 U12410 ( .A1(n14946), .A2(n10598), .ZN(n10603) );
  AOI22_X1 U12411 ( .A1(n12722), .A2(n10600), .B1(n10599), .B2(n12563), .ZN(
        n10601) );
  NAND2_X1 U12412 ( .A1(n10601), .A2(n12663), .ZN(n10602) );
  NOR2_X1 U12413 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n10612) );
  NOR2_X1 U12414 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n10619) );
  NOR2_X1 U12415 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n10618) );
  NOR2_X1 U12416 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n10617) );
  NOR2_X1 U12417 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n10616) );
  NAND2_X1 U12418 ( .A1(n10626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10627) );
  NAND2_X1 U12419 ( .A1(n7523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10630) );
  INV_X1 U12420 ( .A(n11015), .ZN(n10637) );
  NAND3_X1 U12421 ( .A1(n10633), .A2(n10632), .A3(n10638), .ZN(n10634) );
  NOR2_X1 U12422 ( .A1(n10639), .A2(n10634), .ZN(n10635) );
  INV_X1 U12423 ( .A(n10639), .ZN(n10640) );
  NAND2_X1 U12424 ( .A1(n11106), .A2(n10640), .ZN(n10645) );
  NAND2_X1 U12425 ( .A1(n10642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10643) );
  AND2_X2 U12426 ( .A1(n13850), .A2(n13849), .ZN(n13587) );
  NAND2_X1 U12427 ( .A1(n10645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10646) );
  NOR2_X1 U12428 ( .A1(n13839), .A2(n10650), .ZN(n10647) );
  NAND2_X1 U12429 ( .A1(n13587), .A2(n16180), .ZN(n10649) );
  XNOR2_X2 U12430 ( .A(n10653), .B(P1_IR_REG_30__SCAN_IN), .ZN(n10659) );
  INV_X1 U12431 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10656) );
  INV_X1 U12432 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10657) );
  OR2_X1 U12433 ( .A1(n10700), .A2(n10657), .ZN(n10662) );
  INV_X1 U12434 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n11016) );
  OR2_X1 U12435 ( .A1(n10679), .A2(n11016), .ZN(n10661) );
  NAND2_X1 U12436 ( .A1(n13829), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10660) );
  INV_X1 U12437 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n16281) );
  NAND2_X1 U12438 ( .A1(n11277), .A2(SI_0_), .ZN(n10663) );
  XNOR2_X1 U12439 ( .A(n10663), .B(n8375), .ZN(n16182) );
  NAND2_X1 U12440 ( .A1(n10651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10665) );
  MUX2_X1 U12441 ( .A(n16281), .B(n16182), .S(n13712), .Z(n16474) );
  INV_X1 U12442 ( .A(n16474), .ZN(n13584) );
  NAND2_X1 U12443 ( .A1(n13829), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10670) );
  INV_X1 U12444 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n12423) );
  INV_X1 U12445 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10668) );
  INV_X1 U12446 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U12447 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10671) );
  MUX2_X1 U12448 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10671), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n10673) );
  INV_X1 U12449 ( .A(n10672), .ZN(n10683) );
  NAND2_X1 U12450 ( .A1(n10673), .A2(n10683), .ZN(n11341) );
  INV_X1 U12451 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n11317) );
  INV_X1 U12452 ( .A(n13854), .ZN(n10676) );
  NAND2_X1 U12453 ( .A1(n13829), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10682) );
  INV_X1 U12454 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10678) );
  OR2_X1 U12455 ( .A1(n10677), .A2(n10678), .ZN(n10681) );
  INV_X1 U12456 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n12458) );
  OR2_X1 U12457 ( .A1(n10700), .A2(n12458), .ZN(n10680) );
  INV_X1 U12458 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n11350) );
  INV_X2 U12459 ( .A(n13712), .ZN(n11177) );
  NAND2_X1 U12460 ( .A1(n10683), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10684) );
  MUX2_X1 U12461 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10684), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n10685) );
  NAND2_X1 U12462 ( .A1(n10685), .A2(n10695), .ZN(n11349) );
  INV_X1 U12463 ( .A(n11349), .ZN(n15769) );
  AOI22_X1 U12464 ( .A1(n11178), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n11177), 
        .B2(n15769), .ZN(n10687) );
  NAND2_X1 U12465 ( .A1(n11290), .A2(n13838), .ZN(n10686) );
  NAND2_X1 U12466 ( .A1(n11774), .A2(n11777), .ZN(n11773) );
  INV_X1 U12467 ( .A(n8105), .ZN(n13580) );
  NAND2_X1 U12468 ( .A1(n13581), .A2(n13580), .ZN(n10688) );
  NAND2_X1 U12469 ( .A1(n13805), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10694) );
  INV_X1 U12470 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10689) );
  OR2_X1 U12471 ( .A1(n13807), .A2(n10689), .ZN(n10693) );
  INV_X1 U12472 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10690) );
  OR2_X1 U12473 ( .A1(n13810), .A2(n10690), .ZN(n10692) );
  OR2_X1 U12474 ( .A1(n10700), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U12475 ( .A1(n11278), .A2(n13838), .ZN(n10698) );
  NAND2_X1 U12476 ( .A1(n10695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10696) );
  XNOR2_X1 U12477 ( .A(n10696), .B(P1_IR_REG_3__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U12478 ( .A1(n11178), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11177), 
        .B2(n11390), .ZN(n10697) );
  INV_X1 U12479 ( .A(n15755), .ZN(n11775) );
  INV_X1 U12480 ( .A(n13607), .ZN(n13608) );
  NAND2_X1 U12481 ( .A1(n11775), .A2(n13608), .ZN(n10699) );
  NAND2_X1 U12482 ( .A1(n13830), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10704) );
  INV_X1 U12483 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11342) );
  OR2_X1 U12484 ( .A1(n13807), .A2(n11342), .ZN(n10703) );
  INV_X1 U12485 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11359) );
  OR2_X1 U12486 ( .A1(n10679), .A2(n11359), .ZN(n10702) );
  AND2_X1 U12487 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10711) );
  INV_X1 U12488 ( .A(n10711), .ZN(n10713) );
  OAI21_X1 U12489 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n10713), .ZN(n12449) );
  OR2_X1 U12490 ( .A1(n10700), .A2(n12449), .ZN(n10701) );
  NAND2_X1 U12491 ( .A1(n11312), .A2(n13838), .ZN(n10708) );
  NAND2_X1 U12492 ( .A1(n10705), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10706) );
  XNOR2_X1 U12493 ( .A(n10706), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U12494 ( .A1(n11178), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11177), 
        .B2(n15782), .ZN(n10707) );
  NAND2_X1 U12495 ( .A1(n10708), .A2(n10707), .ZN(n13611) );
  INV_X1 U12496 ( .A(n15754), .ZN(n10772) );
  NAND2_X1 U12497 ( .A1(n10772), .A2(n16546), .ZN(n10709) );
  NAND2_X1 U12498 ( .A1(n13829), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10719) );
  INV_X1 U12499 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10710) );
  OR2_X1 U12500 ( .A1(n13810), .A2(n10710), .ZN(n10718) );
  NAND2_X1 U12501 ( .A1(n10711), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10730) );
  INV_X1 U12502 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10712) );
  NAND2_X1 U12503 ( .A1(n10713), .A2(n10712), .ZN(n10714) );
  NAND2_X1 U12504 ( .A1(n10730), .A2(n10714), .ZN(n12475) );
  OR2_X1 U12505 ( .A1(n10700), .A2(n12475), .ZN(n10717) );
  INV_X1 U12506 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10715) );
  OR2_X1 U12507 ( .A1(n10679), .A2(n10715), .ZN(n10716) );
  NAND4_X1 U12508 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n15753) );
  INV_X1 U12509 ( .A(n15753), .ZN(n11903) );
  OR2_X1 U12510 ( .A1(n11326), .A2(n11123), .ZN(n10724) );
  INV_X1 U12511 ( .A(n10720), .ZN(n10721) );
  NAND2_X1 U12512 ( .A1(n10721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10722) );
  XNOR2_X1 U12513 ( .A(n10722), .B(P1_IR_REG_5__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U12514 ( .A1(n11178), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11177), 
        .B2(n11403), .ZN(n10723) );
  NAND2_X1 U12515 ( .A1(n10724), .A2(n10723), .ZN(n13619) );
  XNOR2_X1 U12516 ( .A(n11903), .B(n13619), .ZN(n13858) );
  INV_X1 U12517 ( .A(n13619), .ZN(n12476) );
  NAND2_X1 U12518 ( .A1(n12476), .A2(n11903), .ZN(n10725) );
  OR2_X1 U12519 ( .A1(n11311), .A2(n11123), .ZN(n10728) );
  INV_X1 U12520 ( .A(n11106), .ZN(n10740) );
  NAND2_X1 U12521 ( .A1(n10740), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10726) );
  XNOR2_X1 U12522 ( .A(n10726), .B(P1_IR_REG_6__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U12523 ( .A1(n11178), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11177), 
        .B2(n11364), .ZN(n10727) );
  NAND2_X1 U12524 ( .A1(n10728), .A2(n10727), .ZN(n13628) );
  NAND2_X1 U12525 ( .A1(n13805), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10736) );
  INV_X1 U12526 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n12341) );
  OR2_X1 U12527 ( .A1(n13807), .A2(n12341), .ZN(n10735) );
  INV_X1 U12528 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10729) );
  NOR2_X1 U12529 ( .A1(n10730), .A2(n10729), .ZN(n10744) );
  INV_X1 U12530 ( .A(n10744), .ZN(n10746) );
  NAND2_X1 U12531 ( .A1(n10730), .A2(n10729), .ZN(n10731) );
  NAND2_X1 U12532 ( .A1(n10746), .A2(n10731), .ZN(n12344) );
  OR2_X1 U12533 ( .A1(n10700), .A2(n12344), .ZN(n10734) );
  INV_X1 U12534 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10732) );
  OR2_X1 U12535 ( .A1(n13810), .A2(n10732), .ZN(n10733) );
  NAND4_X1 U12536 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        n15752) );
  NAND2_X1 U12537 ( .A1(n13628), .A2(n15752), .ZN(n10737) );
  NAND2_X1 U12538 ( .A1(n12335), .A2(n10737), .ZN(n10739) );
  OR2_X1 U12539 ( .A1(n13628), .A2(n15752), .ZN(n10738) );
  OR2_X1 U12540 ( .A1(n11315), .A2(n11123), .ZN(n10742) );
  OAI21_X1 U12541 ( .B1(n10740), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10755) );
  XNOR2_X1 U12542 ( .A(n10755), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U12543 ( .A1(n11178), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11177), 
        .B2(n11420), .ZN(n10741) );
  NAND2_X1 U12544 ( .A1(n13805), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10752) );
  INV_X1 U12545 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10743) );
  OR2_X1 U12546 ( .A1(n13807), .A2(n10743), .ZN(n10751) );
  NAND2_X1 U12547 ( .A1(n10744), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10761) );
  INV_X1 U12548 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U12549 ( .A1(n10746), .A2(n10745), .ZN(n10747) );
  NAND2_X1 U12550 ( .A1(n10761), .A2(n10747), .ZN(n16583) );
  OR2_X1 U12551 ( .A1(n10700), .A2(n16583), .ZN(n10750) );
  INV_X1 U12552 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10748) );
  OR2_X1 U12553 ( .A1(n13810), .A2(n10748), .ZN(n10749) );
  NAND4_X1 U12554 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n15751) );
  XNOR2_X1 U12555 ( .A(n13633), .B(n15751), .ZN(n16574) );
  INV_X1 U12556 ( .A(n16574), .ZN(n16569) );
  OR2_X1 U12557 ( .A1(n13633), .A2(n15751), .ZN(n10753) );
  OR2_X1 U12558 ( .A1(n11324), .A2(n11123), .ZN(n10758) );
  NAND2_X1 U12559 ( .A1(n10755), .A2(n9765), .ZN(n10756) );
  NAND2_X1 U12560 ( .A1(n10756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10995) );
  XNOR2_X1 U12561 ( .A(n10995), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U12562 ( .A1(n11178), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11177), 
        .B2(n11436), .ZN(n10757) );
  NAND2_X1 U12563 ( .A1(n10758), .A2(n10757), .ZN(n13637) );
  NAND2_X1 U12564 ( .A1(n13830), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10766) );
  INV_X1 U12565 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10759) );
  OR2_X1 U12566 ( .A1(n10679), .A2(n10759), .ZN(n10765) );
  INV_X1 U12567 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11414) );
  OR2_X1 U12568 ( .A1(n13807), .A2(n11414), .ZN(n10764) );
  NAND2_X1 U12569 ( .A1(n10761), .A2(n10760), .ZN(n10762) );
  NAND2_X1 U12570 ( .A1(n10788), .A2(n10762), .ZN(n12574) );
  OR2_X1 U12571 ( .A1(n10700), .A2(n12574), .ZN(n10763) );
  NAND4_X1 U12572 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n15750) );
  XNOR2_X1 U12573 ( .A(n13637), .B(n12896), .ZN(n13863) );
  NAND2_X1 U12574 ( .A1(n10767), .A2(n10780), .ZN(n10768) );
  NAND2_X1 U12575 ( .A1(n12879), .A2(n10768), .ZN(n16603) );
  NAND2_X1 U12576 ( .A1(n10675), .A2(n13599), .ZN(n11776) );
  NAND2_X1 U12577 ( .A1(n11778), .A2(n11776), .ZN(n10769) );
  NAND2_X1 U12578 ( .A1(n10769), .A2(n13855), .ZN(n11780) );
  NAND2_X1 U12579 ( .A1(n13581), .A2(n8105), .ZN(n10770) );
  NAND2_X1 U12580 ( .A1(n11790), .A2(n13607), .ZN(n10771) );
  NAND2_X1 U12581 ( .A1(n10772), .A2(n13611), .ZN(n10773) );
  NAND2_X1 U12582 ( .A1(n10774), .A2(n10773), .ZN(n11931) );
  NAND2_X1 U12583 ( .A1(n12476), .A2(n15753), .ZN(n10776) );
  XNOR2_X1 U12584 ( .A(n13628), .B(n15752), .ZN(n13860) );
  INV_X1 U12585 ( .A(n13628), .ZN(n16555) );
  NAND2_X1 U12586 ( .A1(n16555), .A2(n15752), .ZN(n10777) );
  INV_X1 U12587 ( .A(n15751), .ZN(n12575) );
  NAND2_X1 U12588 ( .A1(n13633), .A2(n12575), .ZN(n10779) );
  NOR2_X1 U12589 ( .A1(n13633), .A2(n12575), .ZN(n10778) );
  XNOR2_X1 U12590 ( .A(n12883), .B(n10780), .ZN(n10783) );
  INV_X1 U12591 ( .A(n13850), .ZN(n10781) );
  NAND2_X1 U12592 ( .A1(n10650), .A2(n16180), .ZN(n13578) );
  INV_X1 U12593 ( .A(n13578), .ZN(n10782) );
  NAND2_X1 U12594 ( .A1(n10783), .A2(n16623), .ZN(n10795) );
  NAND2_X1 U12595 ( .A1(n16180), .A2(n13849), .ZN(n13840) );
  NAND2_X1 U12596 ( .A1(n13830), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10793) );
  INV_X1 U12597 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10785) );
  OR2_X1 U12598 ( .A1(n10679), .A2(n10785), .ZN(n10792) );
  INV_X1 U12599 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10786) );
  OR2_X1 U12600 ( .A1(n13807), .A2(n10786), .ZN(n10791) );
  NOR2_X1 U12601 ( .A1(n10788), .A2(n10787), .ZN(n10940) );
  INV_X1 U12602 ( .A(n10940), .ZN(n11064) );
  NAND2_X1 U12603 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  NAND2_X1 U12604 ( .A1(n11064), .A2(n10789), .ZN(n16629) );
  OR2_X1 U12605 ( .A1(n10700), .A2(n16629), .ZN(n10790) );
  NAND4_X1 U12606 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n15749) );
  INV_X1 U12607 ( .A(n13840), .ZN(n10808) );
  AOI22_X1 U12608 ( .A1(n15956), .A2(n15749), .B1(n15751), .B2(n15955), .ZN(
        n10794) );
  OAI211_X1 U12609 ( .C1(n16619), .C2(n16603), .A(n10795), .B(n10794), .ZN(
        n16607) );
  NAND2_X1 U12610 ( .A1(n16176), .A2(P1_B_REG_SCAN_IN), .ZN(n10796) );
  MUX2_X1 U12611 ( .A(P1_B_REG_SCAN_IN), .B(n10796), .S(n13516), .Z(n10797) );
  NAND2_X1 U12612 ( .A1(n10797), .A2(n10810), .ZN(n11281) );
  NOR4_X1 U12613 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10806) );
  NOR4_X1 U12614 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10805) );
  INV_X1 U12615 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n16213) );
  INV_X1 U12616 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n16212) );
  INV_X1 U12617 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n16211) );
  INV_X1 U12618 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n16210) );
  NAND4_X1 U12619 ( .A1(n16213), .A2(n16212), .A3(n16211), .A4(n16210), .ZN(
        n10803) );
  NOR4_X1 U12620 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10801) );
  NOR4_X1 U12621 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10800) );
  NOR4_X1 U12622 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10799) );
  NOR4_X1 U12623 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U12624 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10802) );
  NOR4_X1 U12625 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n10803), .A4(n10802), .ZN(n10804) );
  AND3_X1 U12626 ( .A1(n10806), .A2(n10805), .A3(n10804), .ZN(n10807) );
  NOR2_X1 U12627 ( .A1(n11281), .A2(n10807), .ZN(n11570) );
  NAND2_X1 U12628 ( .A1(n13850), .A2(n16033), .ZN(n11200) );
  NAND2_X1 U12629 ( .A1(n11200), .A2(n10808), .ZN(n10809) );
  INV_X1 U12630 ( .A(n11304), .ZN(n11282) );
  NAND3_X1 U12631 ( .A1(n10809), .A2(n11282), .A3(n11015), .ZN(n11569) );
  NOR2_X1 U12632 ( .A1(n11570), .A2(n11569), .ZN(n10812) );
  NAND2_X1 U12633 ( .A1(n16175), .A2(n16176), .ZN(n10811) );
  OAI21_X1 U12634 ( .B1(n11281), .B2(P1_D_REG_1__SCAN_IN), .A(n10811), .ZN(
        n11571) );
  INV_X1 U12635 ( .A(n11571), .ZN(n11197) );
  NAND2_X1 U12636 ( .A1(n10812), .A2(n11197), .ZN(n11208) );
  NAND2_X1 U12637 ( .A1(n16175), .A2(n13516), .ZN(n10813) );
  NAND2_X1 U12638 ( .A1(n11218), .A2(n11770), .ZN(n14035) );
  MUX2_X1 U12639 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n16607), .S(n16014), .Z(
        n10820) );
  OR2_X1 U12640 ( .A1(n10947), .A2(n16033), .ZN(n13843) );
  NOR2_X1 U12641 ( .A1(n16603), .A2(n16006), .ZN(n10819) );
  NAND2_X1 U12642 ( .A1(n12448), .A2(n16546), .ZN(n12447) );
  OR2_X1 U12643 ( .A1(n12447), .A2(n13619), .ZN(n12343) );
  OR2_X1 U12644 ( .A1(n12343), .A2(n13628), .ZN(n12342) );
  OAI211_X1 U12645 ( .C1(n16571), .C2(n8041), .A(n16698), .B(n16613), .ZN(
        n16604) );
  NOR2_X1 U12646 ( .A1(n16604), .A2(n15825), .ZN(n10818) );
  NOR2_X1 U12647 ( .A1(n13850), .A2(n10815), .ZN(n11204) );
  INV_X1 U12648 ( .A(n11204), .ZN(n10816) );
  OR2_X2 U12649 ( .A1(n16642), .A2(n10816), .ZN(n16587) );
  OAI22_X1 U12650 ( .A1(n8041), .A2(n16587), .B1(n12574), .B2(n16036), .ZN(
        n10817) );
  MUX2_X1 U12651 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n10915), .Z(n10841) );
  MUX2_X1 U12652 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n10915), .Z(n10840) );
  INV_X1 U12653 ( .A(n13070), .ZN(n11321) );
  MUX2_X1 U12654 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n10915), .Z(n10838) );
  MUX2_X1 U12655 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n10837), .Z(n10821) );
  XNOR2_X1 U12656 ( .A(n10821), .B(n12166), .ZN(n12164) );
  INV_X1 U12657 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10844) );
  MUX2_X1 U12658 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n10837), .Z(n10822) );
  XNOR2_X1 U12659 ( .A(n10822), .B(n10878), .ZN(n12016) );
  INV_X1 U12660 ( .A(n10822), .ZN(n10823) );
  MUX2_X1 U12661 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n10837), .Z(n10824) );
  XOR2_X1 U12662 ( .A(n12161), .B(n10824), .Z(n12152) );
  INV_X1 U12663 ( .A(n12161), .ZN(n11262) );
  OAI22_X1 U12664 ( .A1(n12151), .A2(n12152), .B1(n10824), .B2(n11262), .ZN(
        n12394) );
  MUX2_X1 U12665 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n10915), .Z(n10825) );
  XNOR2_X1 U12666 ( .A(n10825), .B(n12412), .ZN(n12395) );
  INV_X1 U12667 ( .A(n10825), .ZN(n10826) );
  AOI22_X1 U12668 ( .A1(n12394), .A2(n12395), .B1(n12412), .B2(n10826), .ZN(
        n12180) );
  MUX2_X1 U12669 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n10915), .Z(n10827) );
  XOR2_X1 U12670 ( .A(n12189), .B(n10827), .Z(n12181) );
  INV_X1 U12671 ( .A(n12189), .ZN(n11259) );
  OAI22_X1 U12672 ( .A1(n12180), .A2(n12181), .B1(n10827), .B2(n11259), .ZN(
        n12372) );
  MUX2_X1 U12673 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n10915), .Z(n10828) );
  XOR2_X1 U12674 ( .A(n11269), .B(n10828), .Z(n12373) );
  INV_X1 U12675 ( .A(n11269), .ZN(n12391) );
  INV_X1 U12676 ( .A(n10828), .ZN(n10829) );
  AOI22_X1 U12677 ( .A1(n12372), .A2(n12373), .B1(n12391), .B2(n10829), .ZN(
        n12247) );
  MUX2_X1 U12678 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n10915), .Z(n10830) );
  XOR2_X1 U12679 ( .A(n12259), .B(n10830), .Z(n12248) );
  MUX2_X1 U12680 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n10915), .Z(n10831) );
  XOR2_X1 U12681 ( .A(n11276), .B(n10831), .Z(n12227) );
  INV_X1 U12682 ( .A(n11276), .ZN(n12236) );
  INV_X1 U12683 ( .A(n10831), .ZN(n10832) );
  AOI22_X1 U12684 ( .A1(n12226), .A2(n12227), .B1(n12236), .B2(n10832), .ZN(
        n12361) );
  MUX2_X1 U12685 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n10915), .Z(n10833) );
  XOR2_X1 U12686 ( .A(n12368), .B(n10833), .Z(n12360) );
  INV_X1 U12687 ( .A(n12368), .ZN(n11289) );
  OAI22_X1 U12688 ( .A1(n12361), .A2(n12360), .B1(n10833), .B2(n11289), .ZN(
        n12502) );
  MUX2_X1 U12689 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n10915), .Z(n10834) );
  XNOR2_X1 U12690 ( .A(n10834), .B(n12515), .ZN(n12503) );
  INV_X1 U12691 ( .A(n10834), .ZN(n10835) );
  AOI22_X1 U12692 ( .A1(n12502), .A2(n12503), .B1(n12515), .B2(n10835), .ZN(
        n12744) );
  MUX2_X1 U12693 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n10915), .Z(n10836) );
  XOR2_X1 U12694 ( .A(n12756), .B(n10836), .Z(n12745) );
  INV_X1 U12695 ( .A(n12756), .ZN(n11309) );
  XOR2_X1 U12696 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n13070), .Z(n13057) );
  XOR2_X1 U12697 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n13070), .Z(n13061) );
  INV_X1 U12698 ( .A(n10837), .ZN(n14594) );
  MUX2_X1 U12699 ( .A(n13057), .B(n13061), .S(n14594), .Z(n13067) );
  XNOR2_X1 U12700 ( .A(n10840), .B(n10839), .ZN(n14517) );
  OAI21_X1 U12701 ( .B1(n10840), .B2(n14531), .A(n14516), .ZN(n14543) );
  XNOR2_X1 U12702 ( .A(n10841), .B(n11534), .ZN(n14544) );
  INV_X1 U12703 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n10868) );
  MUX2_X1 U12704 ( .A(n10902), .B(n10868), .S(n10915), .Z(n10842) );
  INV_X1 U12705 ( .A(n14510), .ZN(n10874) );
  AOI211_X1 U12706 ( .C1(n10843), .C2(n10842), .A(n14574), .B(n10917), .ZN(
        n10914) );
  INV_X1 U12707 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16680) );
  OR2_X1 U12708 ( .A1(n13070), .A2(n16680), .ZN(n10862) );
  INV_X1 U12709 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n16505) );
  NAND2_X1 U12710 ( .A1(n8952), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10845) );
  OAI21_X1 U12711 ( .B1(n12166), .B2(n11998), .A(n10845), .ZN(n12169) );
  INV_X1 U12712 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n16485) );
  OR2_X1 U12713 ( .A1(n12169), .A2(n16485), .ZN(n12167) );
  NAND2_X1 U12714 ( .A1(n12167), .A2(n10845), .ZN(n12007) );
  INV_X1 U12715 ( .A(n10878), .ZN(n12021) );
  NAND2_X1 U12716 ( .A1(n12021), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10846) );
  NAND2_X1 U12717 ( .A1(n10847), .A2(n11262), .ZN(n12397) );
  OAI21_X1 U12718 ( .B1(n10847), .B2(n11262), .A(n12397), .ZN(n12154) );
  INV_X1 U12719 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n16534) );
  NAND2_X1 U12720 ( .A1(n12153), .A2(n12397), .ZN(n10848) );
  INV_X1 U12721 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n16541) );
  MUX2_X1 U12722 ( .A(n16541), .B(P3_REG1_REG_4__SCAN_IN), .S(n12412), .Z(
        n12399) );
  NAND2_X1 U12723 ( .A1(n10848), .A2(n12399), .ZN(n12396) );
  OR2_X1 U12724 ( .A1(n12412), .A2(n16541), .ZN(n10849) );
  NAND2_X1 U12725 ( .A1(n12396), .A2(n10849), .ZN(n10850) );
  INV_X1 U12726 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n12600) );
  INV_X1 U12727 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n12765) );
  MUX2_X1 U12728 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n12765), .S(n11269), .Z(
        n12377) );
  NAND2_X1 U12729 ( .A1(n10851), .A2(n12377), .ZN(n12374) );
  NAND2_X1 U12730 ( .A1(n11269), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U12731 ( .A1(n10853), .A2(n7705), .ZN(n12230) );
  INV_X1 U12732 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n16566) );
  INV_X1 U12733 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n16599) );
  MUX2_X1 U12734 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n16599), .S(n11276), .Z(
        n12229) );
  NAND2_X1 U12735 ( .A1(n11276), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10854) );
  NAND2_X1 U12736 ( .A1(n12233), .A2(n10854), .ZN(n10856) );
  INV_X1 U12737 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n13226) );
  OAI21_X1 U12738 ( .B1(n10856), .B2(n11289), .A(n10855), .ZN(n12364) );
  NAND2_X1 U12739 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11297), .ZN(n10857) );
  OAI21_X1 U12740 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11297), .A(n10857), 
        .ZN(n12511) );
  NAND2_X1 U12741 ( .A1(n10859), .A2(n11309), .ZN(n10858) );
  INV_X1 U12742 ( .A(n10858), .ZN(n10860) );
  INV_X1 U12743 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16668) );
  OAI21_X1 U12744 ( .B1(n10859), .B2(n11309), .A(n10858), .ZN(n12752) );
  NAND2_X1 U12745 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n11534), .ZN(n10865) );
  OAI21_X1 U12746 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n11534), .A(n10865), 
        .ZN(n14533) );
  NOR2_X1 U12747 ( .A1(n14534), .A2(n14533), .ZN(n14532) );
  AND2_X1 U12748 ( .A1(n11534), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n10866) );
  OAI21_X1 U12749 ( .B1(n10867), .B2(n11601), .A(n10928), .ZN(n10869) );
  AOI21_X1 U12750 ( .B1(n10869), .B2(n10868), .A(n10929), .ZN(n10873) );
  INV_X1 U12751 ( .A(n10870), .ZN(n10872) );
  NOR2_X1 U12752 ( .A1(n10873), .A2(n14611), .ZN(n10913) );
  MUX2_X1 U12753 ( .A(n10876), .B(n10875), .S(n10874), .Z(n14606) );
  NOR2_X1 U12754 ( .A1(n14606), .A2(n11601), .ZN(n10912) );
  INV_X1 U12755 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n16422) );
  NAND2_X1 U12756 ( .A1(n11534), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n10900) );
  NAND2_X1 U12757 ( .A1(n11297), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10895) );
  MUX2_X1 U12758 ( .A(n8944), .B(P3_REG2_REG_2__SCAN_IN), .S(n10878), .Z(
        n12011) );
  NAND2_X1 U12759 ( .A1(n8952), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10880) );
  OAI21_X1 U12760 ( .B1(n12166), .B2(n12002), .A(n10880), .ZN(n12172) );
  NAND2_X1 U12761 ( .A1(n12174), .A2(n10880), .ZN(n12010) );
  NAND2_X1 U12762 ( .A1(n12021), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10881) );
  MUX2_X1 U12763 ( .A(n10884), .B(P3_REG2_REG_4__SCAN_IN), .S(n12412), .Z(
        n12404) );
  OR2_X1 U12764 ( .A1(n12412), .A2(n10884), .ZN(n10885) );
  NAND2_X1 U12765 ( .A1(n12409), .A2(n10885), .ZN(n10886) );
  NAND2_X1 U12766 ( .A1(n10886), .A2(n11259), .ZN(n12384) );
  OAI21_X1 U12767 ( .B1(n10886), .B2(n11259), .A(n12384), .ZN(n12185) );
  NAND2_X1 U12768 ( .A1(n12386), .A2(n12384), .ZN(n10887) );
  MUX2_X1 U12769 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n9003), .S(n11269), .Z(
        n12383) );
  NAND2_X1 U12770 ( .A1(n10887), .A2(n12383), .ZN(n12388) );
  NAND2_X1 U12771 ( .A1(n11269), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U12772 ( .A1(n12237), .A2(n12238), .ZN(n10889) );
  MUX2_X1 U12773 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n9034), .S(n11276), .Z(
        n12240) );
  NAND2_X1 U12774 ( .A1(n11276), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10890) );
  OAI21_X1 U12775 ( .B1(n10892), .B2(n11289), .A(n10891), .ZN(n12359) );
  OAI21_X1 U12776 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11297), .A(n10895), 
        .ZN(n12506) );
  NOR2_X1 U12777 ( .A1(n13060), .A2(n13061), .ZN(n13059) );
  OAI21_X1 U12778 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n11534), .A(n10900), 
        .ZN(n14537) );
  AND2_X1 U12779 ( .A1(n10903), .A2(n10902), .ZN(n10907) );
  INV_X1 U12780 ( .A(n10904), .ZN(n10905) );
  OAI21_X1 U12781 ( .B1(n7562), .B2(n10907), .A(n14603), .ZN(n10910) );
  NOR2_X1 U12782 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10908), .ZN(n13555) );
  INV_X1 U12783 ( .A(n13555), .ZN(n10909) );
  OAI211_X1 U12784 ( .C1(n16422), .C2(n14572), .A(n10910), .B(n10909), .ZN(
        n10911) );
  INV_X4 U12785 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X2 U12786 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  MUX2_X1 U12787 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n10915), .Z(n10922) );
  MUX2_X1 U12788 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n10915), .Z(n10920) );
  MUX2_X1 U12789 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n10915), .Z(n10919) );
  INV_X1 U12790 ( .A(n10916), .ZN(n10918) );
  XNOR2_X1 U12791 ( .A(n10919), .B(n14553), .ZN(n14562) );
  NOR2_X1 U12792 ( .A1(n14563), .A2(n14562), .ZN(n14561) );
  XNOR2_X1 U12793 ( .A(n10920), .B(n11805), .ZN(n14575) );
  NOR2_X1 U12794 ( .A1(n10921), .A2(n10922), .ZN(n14591) );
  AOI21_X1 U12795 ( .B1(n10922), .B2(n10921), .A(n14591), .ZN(n10927) );
  NAND2_X1 U12796 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14553), .ZN(n10923) );
  OAI21_X1 U12797 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n14553), .A(n10923), 
        .ZN(n14555) );
  NAND2_X1 U12798 ( .A1(n14590), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n14597) );
  OAI21_X1 U12799 ( .B1(n14590), .B2(P3_REG2_REG_18__SCAN_IN), .A(n14597), 
        .ZN(n10926) );
  NAND2_X1 U12800 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14553), .ZN(n10930) );
  OAI21_X1 U12801 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n14553), .A(n10930), 
        .ZN(n14551) );
  NOR2_X1 U12802 ( .A1(n14579), .A2(n7500), .ZN(n10931) );
  INV_X1 U12803 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U12804 ( .A1(n14590), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n14587) );
  OAI21_X1 U12805 ( .B1(n14590), .B2(P3_REG1_REG_18__SCAN_IN), .A(n14587), 
        .ZN(n10932) );
  NAND2_X1 U12806 ( .A1(n10933), .A2(n10932), .ZN(n10934) );
  NOR2_X1 U12807 ( .A1(n14606), .A2(n14590), .ZN(n10936) );
  INV_X1 U12808 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n16460) );
  NAND2_X1 U12809 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14277)
         );
  OAI21_X1 U12810 ( .B1(n14572), .B2(n16460), .A(n14277), .ZN(n10935) );
  NAND2_X1 U12811 ( .A1(n13116), .A2(n13838), .ZN(n10939) );
  OR2_X1 U12812 ( .A1(n10937), .A2(n13167), .ZN(n10938) );
  NAND2_X1 U12813 ( .A1(n11062), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11085) );
  INV_X1 U12814 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U12815 ( .A1(n10961), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U12816 ( .A1(n11145), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11182) );
  INV_X1 U12817 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11181) );
  INV_X1 U12818 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n11209) );
  AND2_X1 U12819 ( .A1(n11184), .A2(n11209), .ZN(n10941) );
  OR2_X1 U12820 ( .A1(n10941), .A2(n11210), .ZN(n15959) );
  INV_X1 U12821 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U12822 ( .A1(n13829), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n10943) );
  NAND2_X1 U12823 ( .A1(n13830), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n10942) );
  OAI211_X1 U12824 ( .C1(n10944), .C2(n10679), .A(n10943), .B(n10942), .ZN(
        n10945) );
  INV_X1 U12825 ( .A(n10945), .ZN(n10946) );
  AND2_X1 U12826 ( .A1(n15739), .A2(n14012), .ZN(n10948) );
  AOI21_X1 U12827 ( .B1(n15958), .B2(n14013), .A(n10948), .ZN(n13960) );
  NAND2_X1 U12828 ( .A1(n15958), .A2(n8750), .ZN(n10950) );
  NAND2_X1 U12829 ( .A1(n15739), .A2(n14013), .ZN(n10949) );
  NAND2_X1 U12830 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  XNOR2_X1 U12831 ( .A(n10951), .B(n13999), .ZN(n13962) );
  XOR2_X1 U12832 ( .A(n13960), .B(n13962), .Z(n11203) );
  NAND2_X1 U12833 ( .A1(n11842), .A2(n13838), .ZN(n10960) );
  NAND2_X1 U12834 ( .A1(n11103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U12835 ( .A1(n10995), .A2(n10952), .ZN(n11079) );
  NAND2_X1 U12836 ( .A1(n10953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10982) );
  INV_X1 U12837 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U12838 ( .A1(n10982), .A2(n10954), .ZN(n10955) );
  NAND2_X1 U12839 ( .A1(n10955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10969) );
  INV_X1 U12840 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U12841 ( .A1(n10969), .A2(n10956), .ZN(n10957) );
  NAND2_X1 U12842 ( .A1(n10957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10958) );
  XNOR2_X1 U12843 ( .A(n10958), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U12844 ( .A1(n12695), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10959) );
  INV_X4 U12845 ( .A(n13967), .ZN(n14001) );
  INV_X1 U12846 ( .A(n10961), .ZN(n11111) );
  NAND2_X1 U12847 ( .A1(n10974), .A2(n10962), .ZN(n10963) );
  NAND2_X1 U12848 ( .A1(n11111), .A2(n10963), .ZN(n15642) );
  OR2_X1 U12849 ( .A1(n15642), .A2(n10700), .ZN(n10967) );
  NAND2_X1 U12850 ( .A1(n13829), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U12851 ( .A1(n13830), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10965) );
  INV_X1 U12852 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11882) );
  OR2_X1 U12853 ( .A1(n10679), .A2(n11882), .ZN(n10964) );
  NAND4_X1 U12854 ( .A1(n10967), .A2(n10966), .A3(n10965), .A4(n10964), .ZN(
        n15744) );
  AOI22_X1 U12855 ( .A1(n16137), .A2(n14013), .B1(n14001), .B2(n15744), .ZN(
        n11099) );
  INV_X2 U12856 ( .A(n13968), .ZN(n14013) );
  AOI22_X1 U12857 ( .A1(n16137), .A2(n8750), .B1(n14013), .B2(n15744), .ZN(
        n10968) );
  XNOR2_X1 U12858 ( .A(n10968), .B(n11072), .ZN(n11098) );
  OR2_X1 U12859 ( .A1(n11699), .A2(n11123), .ZN(n10971) );
  XNOR2_X1 U12860 ( .A(n10969), .B(P1_IR_REG_13__SCAN_IN), .ZN(n15804) );
  AOI22_X1 U12861 ( .A1(n15804), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U12862 ( .A1(n10988), .A2(n10972), .ZN(n10973) );
  NAND2_X1 U12863 ( .A1(n10974), .A2(n10973), .ZN(n13484) );
  OR2_X1 U12864 ( .A1(n13484), .A2(n10700), .ZN(n10979) );
  INV_X1 U12865 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15805) );
  OR2_X1 U12866 ( .A1(n10679), .A2(n15805), .ZN(n10978) );
  INV_X1 U12867 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11875) );
  OR2_X1 U12868 ( .A1(n13807), .A2(n11875), .ZN(n10977) );
  INV_X1 U12869 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10975) );
  OR2_X1 U12870 ( .A1(n13810), .A2(n10975), .ZN(n10976) );
  NAND4_X1 U12871 ( .A1(n10979), .A2(n10978), .A3(n10977), .A4(n10976), .ZN(
        n15745) );
  AND2_X1 U12872 ( .A1(n15745), .A2(n14012), .ZN(n10980) );
  AOI21_X1 U12873 ( .B1(n16697), .B2(n14013), .A(n10980), .ZN(n11097) );
  AOI22_X1 U12874 ( .A1(n16697), .A2(n8750), .B1(n14013), .B2(n15745), .ZN(
        n10981) );
  XNOR2_X1 U12875 ( .A(n10981), .B(n11072), .ZN(n11096) );
  NAND2_X1 U12876 ( .A1(n11633), .A2(n13838), .ZN(n10984) );
  XNOR2_X1 U12877 ( .A(n10982), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U12878 ( .A1(n11883), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10983) );
  NAND2_X1 U12879 ( .A1(n13830), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10992) );
  INV_X1 U12880 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10985) );
  OR2_X1 U12881 ( .A1(n10679), .A2(n10985), .ZN(n10991) );
  INV_X1 U12882 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11637) );
  OR2_X1 U12883 ( .A1(n13807), .A2(n11637), .ZN(n10990) );
  NAND2_X1 U12884 ( .A1(n11085), .A2(n10986), .ZN(n10987) );
  NAND2_X1 U12885 ( .A1(n10988), .A2(n10987), .ZN(n13326) );
  OR2_X1 U12886 ( .A1(n10700), .A2(n13326), .ZN(n10989) );
  NAND4_X1 U12887 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n15746) );
  AND2_X1 U12888 ( .A1(n15746), .A2(n14012), .ZN(n10993) );
  AOI21_X1 U12889 ( .B1(n13659), .B2(n14013), .A(n10993), .ZN(n11095) );
  AOI22_X1 U12890 ( .A1(n13659), .A2(n8750), .B1(n14013), .B2(n15746), .ZN(
        n10994) );
  XNOR2_X1 U12891 ( .A(n10994), .B(n11072), .ZN(n11094) );
  OR2_X1 U12892 ( .A1(n11450), .A2(n11123), .ZN(n11000) );
  NAND2_X1 U12893 ( .A1(n10995), .A2(n10611), .ZN(n10996) );
  NAND2_X1 U12894 ( .A1(n10996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U12895 ( .A1(n10997), .A2(n10609), .ZN(n11058) );
  OR2_X1 U12896 ( .A1(n10997), .A2(n10609), .ZN(n10998) );
  AOI22_X1 U12897 ( .A1(n11587), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n10999) );
  AND2_X1 U12898 ( .A1(n15749), .A2(n14012), .ZN(n11001) );
  AOI21_X1 U12899 ( .B1(n16633), .B2(n14013), .A(n11001), .ZN(n11057) );
  AOI22_X1 U12900 ( .A1(n16633), .A2(n8750), .B1(n14013), .B2(n15749), .ZN(
        n11002) );
  XNOR2_X1 U12901 ( .A(n11002), .B(n11072), .ZN(n11056) );
  AND2_X1 U12902 ( .A1(n15752), .A2(n14012), .ZN(n11003) );
  AOI21_X1 U12903 ( .B1(n13628), .B2(n14013), .A(n11003), .ZN(n11047) );
  NAND2_X1 U12904 ( .A1(n13628), .A2(n8750), .ZN(n11005) );
  NAND2_X1 U12905 ( .A1(n15752), .A2(n14005), .ZN(n11004) );
  NAND2_X1 U12906 ( .A1(n11005), .A2(n11004), .ZN(n11006) );
  XNOR2_X1 U12907 ( .A(n11006), .B(n11072), .ZN(n11046) );
  AOI22_X1 U12908 ( .A1(n15755), .A2(n14001), .B1(n14013), .B2(n13607), .ZN(
        n11032) );
  NAND2_X1 U12909 ( .A1(n15755), .A2(n14005), .ZN(n11008) );
  NAND2_X1 U12910 ( .A1(n13607), .A2(n8750), .ZN(n11007) );
  NAND2_X1 U12911 ( .A1(n11008), .A2(n11007), .ZN(n11009) );
  XNOR2_X1 U12912 ( .A(n11009), .B(n10648), .ZN(n11031) );
  NAND2_X1 U12913 ( .A1(n15757), .A2(n14005), .ZN(n11011) );
  NAND2_X1 U12914 ( .A1(n8750), .A2(n13599), .ZN(n11010) );
  NAND2_X1 U12915 ( .A1(n11011), .A2(n11010), .ZN(n11012) );
  AND2_X1 U12916 ( .A1(n13599), .A2(n14013), .ZN(n11013) );
  AOI21_X1 U12917 ( .B1(n15757), .B2(n14001), .A(n11013), .ZN(n11021) );
  XNOR2_X1 U12918 ( .A(n11020), .B(n11021), .ZN(n11613) );
  OAI22_X1 U12919 ( .A1(n16474), .A2(n13968), .B1(n16281), .B2(n11015), .ZN(
        n11014) );
  AOI21_X1 U12920 ( .B1(n8099), .B2(n14001), .A(n11014), .ZN(n11535) );
  NAND2_X1 U12921 ( .A1(n8099), .A2(n14005), .ZN(n11019) );
  OAI22_X1 U12922 ( .A1(n16474), .A2(n13969), .B1(n11016), .B2(n11015), .ZN(
        n11017) );
  INV_X1 U12923 ( .A(n11017), .ZN(n11018) );
  NAND2_X1 U12924 ( .A1(n11019), .A2(n11018), .ZN(n11536) );
  MUX2_X1 U12925 ( .A(n11072), .B(n11535), .S(n11536), .Z(n11612) );
  INV_X1 U12926 ( .A(n11020), .ZN(n11022) );
  NAND2_X1 U12927 ( .A1(n11022), .A2(n11021), .ZN(n11023) );
  NAND2_X1 U12928 ( .A1(n11611), .A2(n11023), .ZN(n11605) );
  NAND2_X1 U12929 ( .A1(n15756), .A2(n14005), .ZN(n11025) );
  NAND2_X1 U12930 ( .A1(n13582), .A2(n8750), .ZN(n11024) );
  NAND2_X1 U12931 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  XNOR2_X1 U12932 ( .A(n11026), .B(n11072), .ZN(n11027) );
  AOI22_X1 U12933 ( .A1(n15756), .A2(n14001), .B1(n14013), .B2(n8105), .ZN(
        n11028) );
  XNOR2_X1 U12934 ( .A(n11028), .B(n11027), .ZN(n11606) );
  INV_X1 U12935 ( .A(n11027), .ZN(n11029) );
  NAND2_X1 U12936 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  XNOR2_X1 U12937 ( .A(n11031), .B(n11032), .ZN(n11869) );
  NAND2_X1 U12938 ( .A1(n15754), .A2(n14001), .ZN(n11034) );
  NAND2_X1 U12939 ( .A1(n13611), .A2(n14005), .ZN(n11033) );
  NAND2_X1 U12940 ( .A1(n11034), .A2(n11033), .ZN(n11038) );
  NAND2_X1 U12941 ( .A1(n11039), .A2(n11038), .ZN(n11899) );
  NAND2_X1 U12942 ( .A1(n15754), .A2(n14005), .ZN(n11036) );
  NAND2_X1 U12943 ( .A1(n13611), .A2(n8750), .ZN(n11035) );
  NAND2_X1 U12944 ( .A1(n11036), .A2(n11035), .ZN(n11037) );
  XNOR2_X1 U12945 ( .A(n11037), .B(n10648), .ZN(n11898) );
  NAND2_X1 U12946 ( .A1(n11899), .A2(n11898), .ZN(n11897) );
  NAND2_X1 U12947 ( .A1(n13619), .A2(n8750), .ZN(n11041) );
  NAND2_X1 U12948 ( .A1(n15753), .A2(n14013), .ZN(n11040) );
  NAND2_X1 U12949 ( .A1(n11041), .A2(n11040), .ZN(n11042) );
  XNOR2_X1 U12950 ( .A(n11042), .B(n13999), .ZN(n11043) );
  AOI22_X1 U12951 ( .A1(n13619), .A2(n14013), .B1(n15753), .B2(n14001), .ZN(
        n11044) );
  XNOR2_X1 U12952 ( .A(n11043), .B(n11044), .ZN(n11986) );
  INV_X1 U12953 ( .A(n11043), .ZN(n11045) );
  XNOR2_X1 U12954 ( .A(n11046), .B(n11047), .ZN(n12068) );
  AND2_X1 U12955 ( .A1(n15751), .A2(n14012), .ZN(n11048) );
  AOI21_X1 U12956 ( .B1(n13633), .B2(n14013), .A(n11048), .ZN(n11050) );
  AOI22_X1 U12957 ( .A1(n13633), .A2(n8750), .B1(n14013), .B2(n15751), .ZN(
        n11049) );
  XNOR2_X1 U12958 ( .A(n11049), .B(n11072), .ZN(n11051) );
  XOR2_X1 U12959 ( .A(n11050), .B(n11051), .Z(n12416) );
  AOI22_X1 U12960 ( .A1(n13637), .A2(n8750), .B1(n14013), .B2(n15750), .ZN(
        n11053) );
  XNOR2_X1 U12961 ( .A(n11053), .B(n11072), .ZN(n11055) );
  AOI22_X1 U12962 ( .A1(n13637), .A2(n14013), .B1(n14012), .B2(n15750), .ZN(
        n11054) );
  XNOR2_X1 U12963 ( .A(n11055), .B(n11054), .ZN(n12572) );
  XOR2_X1 U12964 ( .A(n11057), .B(n11056), .Z(n12895) );
  OR2_X1 U12965 ( .A1(n11454), .A2(n11123), .ZN(n11061) );
  NAND2_X1 U12966 ( .A1(n11058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11059) );
  XNOR2_X1 U12967 ( .A(n11059), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U12968 ( .A1(n11588), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U12969 ( .A1(n13805), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11070) );
  INV_X1 U12970 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12886) );
  OR2_X1 U12971 ( .A1(n13807), .A2(n12886), .ZN(n11069) );
  INV_X1 U12972 ( .A(n11062), .ZN(n11083) );
  INV_X1 U12973 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U12974 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U12975 ( .A1(n11083), .A2(n11065), .ZN(n13017) );
  OR2_X1 U12976 ( .A1(n10700), .A2(n13017), .ZN(n11068) );
  INV_X1 U12977 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11066) );
  OR2_X1 U12978 ( .A1(n13810), .A2(n11066), .ZN(n11067) );
  NAND4_X1 U12979 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n15748) );
  AND2_X1 U12980 ( .A1(n15748), .A2(n14012), .ZN(n11071) );
  AOI21_X1 U12981 ( .B1(n13649), .B2(n14013), .A(n11071), .ZN(n11075) );
  AOI22_X1 U12982 ( .A1(n13649), .A2(n8750), .B1(n14013), .B2(n15748), .ZN(
        n11073) );
  XNOR2_X1 U12983 ( .A(n11073), .B(n11072), .ZN(n11074) );
  XOR2_X1 U12984 ( .A(n11075), .B(n11074), .Z(n13015) );
  INV_X1 U12985 ( .A(n11074), .ZN(n11077) );
  NAND2_X1 U12986 ( .A1(n11541), .A2(n13838), .ZN(n11081) );
  XNOR2_X1 U12987 ( .A(n11079), .B(n9768), .ZN(n11645) );
  AOI22_X1 U12988 ( .A1(n11178), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11645), 
        .B2(n11177), .ZN(n11080) );
  NAND2_X1 U12989 ( .A1(n13829), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11090) );
  INV_X1 U12990 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11082) );
  OR2_X1 U12991 ( .A1(n10679), .A2(n11082), .ZN(n11089) );
  INV_X1 U12992 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n13218) );
  NAND2_X1 U12993 ( .A1(n11083), .A2(n13218), .ZN(n11084) );
  NAND2_X1 U12994 ( .A1(n11085), .A2(n11084), .ZN(n13219) );
  OR2_X1 U12995 ( .A1(n10700), .A2(n13219), .ZN(n11088) );
  INV_X1 U12996 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11086) );
  OR2_X1 U12997 ( .A1(n13810), .A2(n11086), .ZN(n11087) );
  NAND4_X1 U12998 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n15747) );
  AOI22_X1 U12999 ( .A1(n13656), .A2(n8750), .B1(n14013), .B2(n15747), .ZN(
        n11091) );
  XNOR2_X1 U13000 ( .A(n11091), .B(n11072), .ZN(n11093) );
  AOI22_X1 U13001 ( .A1(n13656), .A2(n14013), .B1(n14012), .B2(n15747), .ZN(
        n11092) );
  XNOR2_X1 U13002 ( .A(n11093), .B(n11092), .ZN(n13217) );
  XOR2_X1 U13003 ( .A(n11095), .B(n11094), .Z(n13324) );
  XOR2_X1 U13004 ( .A(n11097), .B(n11096), .Z(n13482) );
  XNOR2_X1 U13005 ( .A(n11098), .B(n11099), .ZN(n15640) );
  NAND2_X1 U13006 ( .A1(n11993), .A2(n13838), .ZN(n11109) );
  NAND4_X1 U13007 ( .A1(n11102), .A2(n11101), .A3(n9768), .A4(n11100), .ZN(
        n11104) );
  NOR2_X1 U13008 ( .A1(n11104), .A2(n11103), .ZN(n11105) );
  NAND2_X1 U13009 ( .A1(n11106), .A2(n11105), .ZN(n11124) );
  NAND2_X1 U13010 ( .A1(n11124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11107) );
  XNOR2_X1 U13011 ( .A(n11107), .B(P1_IR_REG_15__SCAN_IN), .ZN(n16293) );
  AOI22_X1 U13012 ( .A1(n11178), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11177), 
        .B2(n16293), .ZN(n11108) );
  NAND2_X1 U13013 ( .A1(n16718), .A2(n8750), .ZN(n11120) );
  INV_X1 U13014 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11118) );
  INV_X1 U13015 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U13016 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  NAND2_X1 U13017 ( .A1(n11129), .A2(n11112), .ZN(n16722) );
  OR2_X1 U13018 ( .A1(n16722), .A2(n10700), .ZN(n11117) );
  INV_X1 U13019 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11113) );
  OR2_X1 U13020 ( .A1(n10679), .A2(n11113), .ZN(n11115) );
  INV_X1 U13021 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n13509) );
  OR2_X1 U13022 ( .A1(n13807), .A2(n13509), .ZN(n11114) );
  AND2_X1 U13023 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  OAI211_X1 U13024 ( .C1(n13810), .C2(n11118), .A(n11117), .B(n11116), .ZN(
        n15743) );
  NAND2_X1 U13025 ( .A1(n15743), .A2(n14013), .ZN(n11119) );
  NAND2_X1 U13026 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  XNOR2_X1 U13027 ( .A(n11121), .B(n11072), .ZN(n11122) );
  AOI22_X1 U13028 ( .A1(n16718), .A2(n14005), .B1(n14012), .B2(n15743), .ZN(
        n16712) );
  NAND2_X1 U13029 ( .A1(n11139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11125) );
  XNOR2_X1 U13030 ( .A(n11125), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U13031 ( .A1(n11178), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11177), 
        .B2(n12859), .ZN(n11126) );
  NAND2_X1 U13032 ( .A1(n16129), .A2(n8750), .ZN(n11134) );
  NAND2_X1 U13033 ( .A1(n11129), .A2(n11128), .ZN(n11130) );
  NAND2_X1 U13034 ( .A1(n11147), .A2(n11130), .ZN(n16035) );
  AOI22_X1 U13035 ( .A1(n13805), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n13829), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U13036 ( .A1(n13830), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11131) );
  OAI211_X1 U13037 ( .C1(n16035), .C2(n10700), .A(n11132), .B(n11131), .ZN(
        n15742) );
  NAND2_X1 U13038 ( .A1(n15742), .A2(n14005), .ZN(n11133) );
  NAND2_X1 U13039 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  XNOR2_X1 U13040 ( .A(n11135), .B(n13999), .ZN(n11136) );
  AOI22_X1 U13041 ( .A1(n16129), .A2(n14013), .B1(n14012), .B2(n15742), .ZN(
        n11137) );
  XNOR2_X1 U13042 ( .A(n11136), .B(n11137), .ZN(n15681) );
  INV_X1 U13043 ( .A(n11136), .ZN(n11138) );
  NAND2_X1 U13044 ( .A1(n12566), .A2(n13838), .ZN(n11144) );
  NAND2_X1 U13045 ( .A1(n11158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11141) );
  INV_X1 U13046 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n11140) );
  XNOR2_X1 U13047 ( .A(n11141), .B(n11140), .ZN(n13158) );
  INV_X1 U13048 ( .A(n13158), .ZN(n11142) );
  AOI22_X1 U13049 ( .A1(n11142), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n11143) );
  INV_X1 U13050 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n11151) );
  INV_X1 U13051 ( .A(n11145), .ZN(n11163) );
  NAND2_X1 U13052 ( .A1(n11147), .A2(n11146), .ZN(n11148) );
  NAND2_X1 U13053 ( .A1(n11163), .A2(n11148), .ZN(n16013) );
  OR2_X1 U13054 ( .A1(n16013), .A2(n10700), .ZN(n11150) );
  AOI22_X1 U13055 ( .A1(n13805), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n13829), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n11149) );
  OAI211_X1 U13056 ( .C1(n13810), .C2(n11151), .A(n11150), .B(n11149), .ZN(
        n15741) );
  AOI22_X1 U13057 ( .A1(n16123), .A2(n14005), .B1(n14012), .B2(n15741), .ZN(
        n11155) );
  NAND2_X1 U13058 ( .A1(n16123), .A2(n8750), .ZN(n11153) );
  NAND2_X1 U13059 ( .A1(n15741), .A2(n14013), .ZN(n11152) );
  NAND2_X1 U13060 ( .A1(n11153), .A2(n11152), .ZN(n11154) );
  XNOR2_X1 U13061 ( .A(n11154), .B(n13999), .ZN(n11157) );
  XOR2_X1 U13062 ( .A(n11155), .B(n11157), .Z(n15687) );
  INV_X1 U13063 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U13064 ( .A1(n12847), .A2(n13838), .ZN(n11161) );
  OAI21_X1 U13065 ( .B1(n11158), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n11159) );
  XNOR2_X1 U13066 ( .A(n11159), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U13067 ( .A1(n13378), .A2(n11177), .B1(n11178), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n11160) );
  NAND2_X1 U13068 ( .A1(n16118), .A2(n8750), .ZN(n11172) );
  INV_X1 U13069 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U13070 ( .A1(n11163), .A2(n11162), .ZN(n11164) );
  NAND2_X1 U13071 ( .A1(n11182), .A2(n11164), .ZN(n16000) );
  OR2_X1 U13072 ( .A1(n16000), .A2(n10700), .ZN(n11170) );
  INV_X1 U13073 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U13074 ( .A1(n13830), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11166) );
  INV_X1 U13075 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n16001) );
  OR2_X1 U13076 ( .A1(n13807), .A2(n16001), .ZN(n11165) );
  OAI211_X1 U13077 ( .C1(n10679), .C2(n11167), .A(n11166), .B(n11165), .ZN(
        n11168) );
  INV_X1 U13078 ( .A(n11168), .ZN(n11169) );
  NAND2_X1 U13079 ( .A1(n15740), .A2(n14013), .ZN(n11171) );
  NAND2_X1 U13080 ( .A1(n11172), .A2(n11171), .ZN(n11173) );
  XNOR2_X1 U13081 ( .A(n11173), .B(n13999), .ZN(n11174) );
  AOI22_X1 U13082 ( .A1(n16118), .A2(n14013), .B1(n14012), .B2(n15740), .ZN(
        n11175) );
  XNOR2_X1 U13083 ( .A(n11174), .B(n11175), .ZN(n15714) );
  INV_X1 U13084 ( .A(n11174), .ZN(n11176) );
  NAND2_X1 U13085 ( .A1(n13025), .A2(n13838), .ZN(n11180) );
  AOI22_X1 U13086 ( .A1(n11178), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11177), 
        .B2(n10650), .ZN(n11179) );
  NAND2_X1 U13087 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  NAND2_X1 U13088 ( .A1(n11184), .A2(n11183), .ZN(n15979) );
  OR2_X1 U13089 ( .A1(n15979), .A2(n10700), .ZN(n11189) );
  INV_X1 U13090 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13382) );
  NAND2_X1 U13091 ( .A1(n13830), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U13092 ( .A1(n13829), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11185) );
  OAI211_X1 U13093 ( .C1(n10679), .C2(n13382), .A(n11186), .B(n11185), .ZN(
        n11187) );
  INV_X1 U13094 ( .A(n11187), .ZN(n11188) );
  AOI22_X1 U13095 ( .A1(n16111), .A2(n14013), .B1(n14001), .B2(n15954), .ZN(
        n11193) );
  NAND2_X1 U13096 ( .A1(n16111), .A2(n8750), .ZN(n11191) );
  NAND2_X1 U13097 ( .A1(n15954), .A2(n14005), .ZN(n11190) );
  NAND2_X1 U13098 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  XNOR2_X1 U13099 ( .A(n11192), .B(n13999), .ZN(n11195) );
  XOR2_X1 U13100 ( .A(n11193), .B(n11195), .Z(n15655) );
  INV_X1 U13101 ( .A(n11193), .ZN(n11194) );
  INV_X1 U13102 ( .A(n11770), .ZN(n11574) );
  INV_X1 U13103 ( .A(n11303), .ZN(n11196) );
  NOR2_X1 U13104 ( .A1(n11570), .A2(n11196), .ZN(n11198) );
  AND3_X1 U13105 ( .A1(n11574), .A2(n11198), .A3(n11197), .ZN(n11205) );
  AND2_X1 U13106 ( .A1(n16684), .A2(n13840), .ZN(n11201) );
  AOI211_X1 U13107 ( .C1(n11203), .C2(n11202), .A(n15729), .B(n7506), .ZN(
        n11222) );
  INV_X1 U13108 ( .A(n15958), .ZN(n16104) );
  NAND2_X1 U13109 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  INV_X1 U13110 ( .A(n16719), .ZN(n15712) );
  NOR2_X1 U13111 ( .A1(n16104), .A2(n15712), .ZN(n11221) );
  INV_X1 U13112 ( .A(n11207), .ZN(n11573) );
  OAI22_X1 U13113 ( .A1(n11208), .A2(n11770), .B1(n11569), .B2(n11573), .ZN(
        n11537) );
  OAI22_X1 U13114 ( .A1(n15959), .A2(n16723), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11209), .ZN(n11220) );
  OR2_X1 U13115 ( .A1(n11210), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U13116 ( .A1(n11210), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n13571) );
  NAND2_X1 U13117 ( .A1(n11211), .A2(n13571), .ZN(n15942) );
  OR2_X1 U13118 ( .A1(n15942), .A2(n10700), .ZN(n11217) );
  INV_X1 U13119 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U13120 ( .A1(n13830), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U13121 ( .A1(n13829), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11212) );
  OAI211_X1 U13122 ( .C1(n10679), .C2(n11214), .A(n11213), .B(n11212), .ZN(
        n11215) );
  INV_X1 U13123 ( .A(n11215), .ZN(n11216) );
  NAND2_X1 U13124 ( .A1(n11218), .A2(n11574), .ZN(n15691) );
  INV_X1 U13125 ( .A(n15954), .ZN(n15996) );
  OR2_X1 U13126 ( .A1(n15691), .A2(n16031), .ZN(n15716) );
  OAI22_X1 U13127 ( .A1(n8149), .A2(n15717), .B1(n15996), .B2(n15716), .ZN(
        n11219) );
  AND2_X1 U13128 ( .A1(n11919), .A2(n15099), .ZN(n11715) );
  XNOR2_X1 U13129 ( .A(n11716), .B(n8283), .ZN(n11754) );
  INV_X1 U13130 ( .A(n11224), .ZN(n11225) );
  OAI21_X1 U13131 ( .B1(n11716), .B2(n11225), .A(n11722), .ZN(n11228) );
  NAND2_X1 U13132 ( .A1(n11682), .A2(n10566), .ZN(n15162) );
  INV_X1 U13133 ( .A(n15225), .ZN(n15043) );
  OAI22_X1 U13134 ( .A1(n11723), .A2(n15162), .B1(n11227), .B2(n15043), .ZN(
        n14059) );
  AOI21_X1 U13135 ( .B1(n11228), .B2(n15446), .A(n14059), .ZN(n11229) );
  OAI21_X1 U13136 ( .B1(n11754), .B2(n15443), .A(n11229), .ZN(n11755) );
  NAND2_X1 U13137 ( .A1(n11918), .A2(n11922), .ZN(n11709) );
  INV_X1 U13138 ( .A(n11709), .ZN(n11230) );
  NAND2_X1 U13139 ( .A1(n11682), .A2(n11685), .ZN(n11710) );
  XNOR2_X1 U13140 ( .A(P2_B_REG_SCAN_IN), .B(n13513), .ZN(n11231) );
  AND2_X1 U13141 ( .A1(n15625), .A2(n11231), .ZN(n11232) );
  OR2_X1 U13142 ( .A1(n15622), .A2(n11232), .ZN(n11234) );
  NAND2_X1 U13143 ( .A1(n15622), .A2(n13513), .ZN(n11233) );
  INV_X1 U13144 ( .A(n11234), .ZN(n16218) );
  INV_X1 U13145 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n16217) );
  AOI22_X1 U13146 ( .A1(n16218), .A2(n16217), .B1(n15622), .B2(n15625), .ZN(
        n11708) );
  NOR4_X1 U13147 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n11238) );
  NOR4_X1 U13148 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n11237) );
  NOR4_X1 U13149 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n11236) );
  NOR4_X1 U13150 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n11235) );
  NAND4_X1 U13151 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11244) );
  NOR2_X1 U13152 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n11242) );
  NOR4_X1 U13153 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n11241) );
  NOR4_X1 U13154 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n11240) );
  NOR4_X1 U13155 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U13156 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11243) );
  OAI21_X1 U13157 ( .B1(n11244), .B2(n11243), .A(n16218), .ZN(n11711) );
  NAND2_X1 U13158 ( .A1(n11708), .A2(n11711), .ZN(n11680) );
  INV_X1 U13159 ( .A(n11680), .ZN(n11245) );
  NAND4_X1 U13160 ( .A1(n16223), .A2(n11710), .A3(n16222), .A4(n11245), .ZN(
        n11246) );
  MUX2_X1 U13161 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11755), .S(n15429), .Z(
        n11255) );
  NOR2_X1 U13162 ( .A1(n11250), .A2(n13117), .ZN(n11686) );
  INV_X1 U13163 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11247) );
  OAI22_X1 U13164 ( .A1(n15456), .A2(n14066), .B1(n11247), .B2(n15427), .ZN(
        n11254) );
  NAND2_X1 U13165 ( .A1(n11922), .A2(n11248), .ZN(n12080) );
  INV_X1 U13166 ( .A(n12080), .ZN(n11249) );
  NAND2_X1 U13167 ( .A1(n15429), .A2(n11249), .ZN(n15458) );
  OAI21_X1 U13168 ( .B1(n11668), .B2(n14066), .A(n15232), .ZN(n11251) );
  AND2_X1 U13169 ( .A1(n11668), .A2(n14066), .ZN(n12098) );
  NOR2_X1 U13170 ( .A1(n11251), .A2(n12098), .ZN(n11756) );
  INV_X1 U13171 ( .A(n11756), .ZN(n11252) );
  OAI22_X1 U13172 ( .A1(n11754), .A2(n15458), .B1(n15318), .B2(n11252), .ZN(
        n11253) );
  OR3_X1 U13173 ( .A1(n11255), .A2(n11254), .A3(n11253), .ZN(P2_U3264) );
  INV_X2 U13174 ( .A(n15608), .ZN(n15628) );
  OR2_X2 U13175 ( .A1(n8230), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15626) );
  INV_X1 U13176 ( .A(n15100), .ZN(n11256) );
  OAI222_X1 U13177 ( .A1(n15628), .A2(n11257), .B1(n15626), .B2(n11318), .C1(
        P2_U3088), .C2(n11256), .ZN(P2_U3326) );
  INV_X2 U13178 ( .A(n12874), .ZN(n14968) );
  NOR2_X1 U13179 ( .A1(n11277), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14952) );
  OAI222_X1 U13180 ( .A1(P3_U3151), .A2(n11259), .B1(n14968), .B2(n11258), 
        .C1(n14959), .C2(n9940), .ZN(P3_U3290) );
  OAI222_X1 U13181 ( .A1(P3_U3151), .A2(n11262), .B1(n14968), .B2(n11261), 
        .C1(n14959), .C2(n11260), .ZN(P3_U3292) );
  INV_X1 U13182 ( .A(n12412), .ZN(n11265) );
  OAI222_X1 U13183 ( .A1(n11265), .A2(P3_U3151), .B1(n14968), .B2(n11264), 
        .C1(n11263), .C2(n14959), .ZN(P3_U3291) );
  INV_X1 U13184 ( .A(n11266), .ZN(n11268) );
  OAI222_X1 U13185 ( .A1(P3_U3151), .A2(n11269), .B1(n14968), .B2(n11268), 
        .C1(n11267), .C2(n14959), .ZN(P3_U3289) );
  INV_X1 U13186 ( .A(n11270), .ZN(n11272) );
  OAI222_X1 U13187 ( .A1(n12166), .A2(P3_U3151), .B1(n14968), .B2(n11272), 
        .C1(n11271), .C2(n14959), .ZN(P3_U3294) );
  INV_X1 U13188 ( .A(n11273), .ZN(n11275) );
  OAI222_X1 U13189 ( .A1(n11276), .A2(P3_U3151), .B1(n14968), .B2(n11275), 
        .C1(n11274), .C2(n14959), .ZN(P3_U3287) );
  OR2_X2 U13190 ( .A1(n11277), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16174) );
  INV_X1 U13191 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n11279) );
  INV_X1 U13192 ( .A(n11278), .ZN(n11293) );
  INV_X1 U13193 ( .A(n11390), .ZN(n11397) );
  OAI222_X1 U13194 ( .A1(n16174), .A2(n11279), .B1(n13259), .B2(n11293), .C1(
        n11397), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U13195 ( .A(n11364), .ZN(n11386) );
  OAI222_X1 U13196 ( .A1(n16174), .A2(n11280), .B1(n13259), .B2(n11311), .C1(
        n11386), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U13197 ( .A(n13516), .ZN(n11283) );
  NAND3_X1 U13198 ( .A1(n16175), .A2(P1_STATE_REG_SCAN_IN), .A3(n11282), .ZN(
        n11285) );
  OAI22_X1 U13199 ( .A1(n16214), .A2(P1_D_REG_0__SCAN_IN), .B1(n11283), .B2(
        n11285), .ZN(n11284) );
  INV_X1 U13200 ( .A(n11284), .ZN(P1_U3445) );
  INV_X1 U13201 ( .A(n16176), .ZN(n11286) );
  OAI22_X1 U13202 ( .A1(n16214), .A2(P1_D_REG_1__SCAN_IN), .B1(n11286), .B2(
        n11285), .ZN(n11287) );
  INV_X1 U13203 ( .A(n11287), .ZN(P1_U3446) );
  OAI222_X1 U13204 ( .A1(n11289), .A2(P3_U3151), .B1(n14968), .B2(n11288), 
        .C1(n8112), .C2(n14959), .ZN(P3_U3286) );
  INV_X1 U13205 ( .A(n11290), .ZN(n11328) );
  AOI22_X1 U13206 ( .A1(n16228), .A2(P2_STATE_REG_SCAN_IN), .B1(n15608), .B2(
        P1_DATAO_REG_2__SCAN_IN), .ZN(n11291) );
  OAI21_X1 U13207 ( .B1(n11328), .B2(n15626), .A(n11291), .ZN(P2_U3325) );
  AOI22_X1 U13208 ( .A1(n11485), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n15608), .ZN(n11292) );
  OAI21_X1 U13209 ( .B1(n11293), .B2(n15626), .A(n11292), .ZN(P2_U3324) );
  AOI22_X1 U13210 ( .A1(n11520), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n15608), .ZN(n11294) );
  OAI21_X1 U13211 ( .B1(n11326), .B2(n15626), .A(n11294), .ZN(P2_U3322) );
  OAI222_X1 U13212 ( .A1(P3_U3151), .A2(n11297), .B1(n14959), .B2(n11296), 
        .C1(n14968), .C2(n11295), .ZN(P3_U3285) );
  OAI222_X1 U13213 ( .A1(n14968), .A2(n11299), .B1(n14959), .B2(n11298), .C1(
        n7705), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U13214 ( .A(n11420), .ZN(n11413) );
  OAI222_X1 U13215 ( .A1(n16174), .A2(n11300), .B1(n13259), .B2(n11315), .C1(
        n11413), .C2(P1_U3086), .ZN(P1_U3348) );
  OAI222_X1 U13216 ( .A1(n12021), .A2(P3_U3151), .B1(n14968), .B2(n11302), 
        .C1(n11301), .C2(n14959), .ZN(P3_U3293) );
  NAND2_X1 U13217 ( .A1(n11304), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13908) );
  INV_X1 U13218 ( .A(n13908), .ZN(n13889) );
  OR2_X1 U13219 ( .A1(n11303), .A2(n13889), .ZN(n11331) );
  OR2_X1 U13220 ( .A1(n13840), .A2(n11304), .ZN(n11305) );
  INV_X1 U13221 ( .A(n11330), .ZN(n11306) );
  AND2_X1 U13222 ( .A1(n11331), .A2(n11306), .ZN(n16283) );
  NOR2_X1 U13223 ( .A1(n16283), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U13224 ( .A1(P3_U3151), .A2(n11309), .B1(n14968), .B2(n11308), 
        .C1(n14959), .C2(n11307), .ZN(P3_U3284) );
  INV_X1 U13225 ( .A(n11547), .ZN(n11551) );
  OAI222_X1 U13226 ( .A1(P2_U3088), .A2(n11551), .B1(n15626), .B2(n11311), 
        .C1(n11310), .C2(n15628), .ZN(P2_U3321) );
  INV_X1 U13227 ( .A(n11312), .ZN(n11322) );
  OAI222_X1 U13228 ( .A1(n15628), .A2(n11313), .B1(n15626), .B2(n11322), .C1(
        P2_U3088), .C2(n11500), .ZN(P2_U3323) );
  INV_X1 U13229 ( .A(n11740), .ZN(n11560) );
  INV_X1 U13230 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n11314) );
  OAI222_X1 U13231 ( .A1(P2_U3088), .A2(n11560), .B1(n15626), .B2(n11315), 
        .C1(n11314), .C2(n15628), .ZN(P2_U3320) );
  INV_X1 U13232 ( .A(n11853), .ZN(n11746) );
  OAI222_X1 U13233 ( .A1(P2_U3088), .A2(n11746), .B1(n15626), .B2(n11324), 
        .C1(n11316), .C2(n15628), .ZN(P2_U3319) );
  INV_X1 U13234 ( .A(n13335), .ZN(n16178) );
  OAI222_X1 U13235 ( .A1(n16178), .A2(n11318), .B1(n16174), .B2(n11317), .C1(
        P1_U3086), .C2(n11341), .ZN(P1_U3354) );
  OAI222_X1 U13236 ( .A1(P3_U3151), .A2(n11321), .B1(n14968), .B2(n11320), 
        .C1(n14959), .C2(n11319), .ZN(P3_U3283) );
  INV_X1 U13237 ( .A(n15782), .ZN(n15790) );
  OAI222_X1 U13238 ( .A1(P1_U3086), .A2(n15790), .B1(n16178), .B2(n11322), 
        .C1(n8115), .C2(n16174), .ZN(P1_U3351) );
  INV_X1 U13239 ( .A(n11436), .ZN(n11323) );
  OAI222_X1 U13240 ( .A1(n16174), .A2(n11325), .B1(n16178), .B2(n11324), .C1(
        n11323), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U13241 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n11327) );
  INV_X1 U13242 ( .A(n11403), .ZN(n11344) );
  OAI222_X1 U13243 ( .A1(n16174), .A2(n11327), .B1(n16178), .B2(n11326), .C1(
        n11344), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U13244 ( .A1(n16174), .A2(n11329), .B1(n16178), .B2(n11328), .C1(
        n11349), .C2(P1_U3086), .ZN(P1_U3353) );
  NAND2_X1 U13245 ( .A1(n11331), .A2(n11330), .ZN(n16285) );
  INV_X1 U13246 ( .A(n16285), .ZN(n11332) );
  NAND2_X1 U13247 ( .A1(n11332), .A2(n16170), .ZN(n16297) );
  XNOR2_X1 U13248 ( .A(n11341), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n11352) );
  AND2_X1 U13249 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n11351) );
  XNOR2_X1 U13250 ( .A(n11352), .B(n11351), .ZN(n11339) );
  INV_X1 U13251 ( .A(n11341), .ZN(n11353) );
  INV_X1 U13252 ( .A(n16283), .ZN(n16301) );
  OAI22_X1 U13253 ( .A1(n16301), .A2(n11333), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12423), .ZN(n11334) );
  AOI21_X1 U13254 ( .B1(n11353), .B2(n16294), .A(n11334), .ZN(n11338) );
  INV_X1 U13255 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15758) );
  NOR2_X1 U13256 ( .A1(n16281), .A2(n15758), .ZN(n15759) );
  INV_X1 U13257 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11335) );
  MUX2_X1 U13258 ( .A(n11335), .B(P1_REG2_REG_1__SCAN_IN), .S(n11341), .Z(
        n11336) );
  NOR2_X1 U13259 ( .A1(n16285), .A2(n16170), .ZN(n13387) );
  NAND3_X1 U13260 ( .A1(n11336), .A2(P1_REG2_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n11340) );
  OAI211_X1 U13261 ( .C1(n15759), .C2(n11336), .A(n15797), .B(n11340), .ZN(
        n11337) );
  OAI211_X1 U13262 ( .C1(n16297), .C2(n11339), .A(n11338), .B(n11337), .ZN(
        P1_U3244) );
  OAI21_X1 U13263 ( .B1(n11335), .B2(n11341), .A(n11340), .ZN(n15765) );
  XNOR2_X1 U13264 ( .A(n11349), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U13265 ( .A1(n15765), .A2(n15764), .B1(n15769), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n11389) );
  MUX2_X1 U13266 ( .A(n10689), .B(P1_REG2_REG_3__SCAN_IN), .S(n11390), .Z(
        n11388) );
  NOR2_X1 U13267 ( .A1(n11389), .A2(n11388), .ZN(n15779) );
  NOR2_X1 U13268 ( .A1(n11397), .A2(n10689), .ZN(n15778) );
  MUX2_X1 U13269 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11342), .S(n15782), .Z(
        n15777) );
  OAI21_X1 U13270 ( .B1(n15779), .B2(n15778), .A(n15777), .ZN(n15776) );
  NAND2_X1 U13271 ( .A1(n15782), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n11406) );
  INV_X1 U13272 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11343) );
  MUX2_X1 U13273 ( .A(n11343), .B(P1_REG2_REG_5__SCAN_IN), .S(n11403), .Z(
        n11405) );
  AOI21_X1 U13274 ( .B1(n15776), .B2(n11406), .A(n11405), .ZN(n11408) );
  NOR2_X1 U13275 ( .A1(n11344), .A2(n11343), .ZN(n11375) );
  MUX2_X1 U13276 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n12341), .S(n11364), .Z(
        n11374) );
  OAI21_X1 U13277 ( .B1(n11408), .B2(n11375), .A(n11374), .ZN(n11377) );
  NAND2_X1 U13278 ( .A1(n11364), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11346) );
  MUX2_X1 U13279 ( .A(n10743), .B(P1_REG2_REG_7__SCAN_IN), .S(n11420), .Z(
        n11345) );
  AOI21_X1 U13280 ( .B1(n11377), .B2(n11346), .A(n11345), .ZN(n11442) );
  NAND3_X1 U13281 ( .A1(n11377), .A2(n11346), .A3(n11345), .ZN(n11347) );
  NAND2_X1 U13282 ( .A1(n15797), .A2(n11347), .ZN(n11373) );
  AND2_X1 U13283 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n12420) );
  NOR2_X1 U13284 ( .A1(n16301), .A2(n16358), .ZN(n11348) );
  AOI211_X1 U13285 ( .C1(n16294), .C2(n11420), .A(n12420), .B(n11348), .ZN(
        n11372) );
  MUX2_X1 U13286 ( .A(n11350), .B(P1_REG1_REG_2__SCAN_IN), .S(n11349), .Z(
        n15768) );
  NAND2_X1 U13287 ( .A1(n11352), .A2(n11351), .ZN(n11355) );
  NAND2_X1 U13288 ( .A1(n11353), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11354) );
  NAND2_X1 U13289 ( .A1(n11355), .A2(n11354), .ZN(n15767) );
  NAND2_X1 U13290 ( .A1(n15768), .A2(n15767), .ZN(n15766) );
  NAND2_X1 U13291 ( .A1(n15769), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U13292 ( .A1(n15766), .A2(n11391), .ZN(n11358) );
  INV_X1 U13293 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11356) );
  MUX2_X1 U13294 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n11356), .S(n11390), .Z(
        n11357) );
  NAND2_X1 U13295 ( .A1(n11358), .A2(n11357), .ZN(n15785) );
  NAND2_X1 U13296 ( .A1(n11390), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15784) );
  NAND2_X1 U13297 ( .A1(n15785), .A2(n15784), .ZN(n11361) );
  MUX2_X1 U13298 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n11359), .S(n15782), .Z(
        n11360) );
  NAND2_X1 U13299 ( .A1(n11361), .A2(n11360), .ZN(n15787) );
  NAND2_X1 U13300 ( .A1(n15782), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n11362) );
  AND2_X1 U13301 ( .A1(n15787), .A2(n11362), .ZN(n11401) );
  MUX2_X1 U13302 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10715), .S(n11403), .Z(
        n11402) );
  NAND2_X1 U13303 ( .A1(n11401), .A2(n11402), .ZN(n11400) );
  OR2_X1 U13304 ( .A1(n11403), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U13305 ( .A1(n11400), .A2(n11363), .ZN(n11378) );
  INV_X1 U13306 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n16560) );
  MUX2_X1 U13307 ( .A(n16560), .B(P1_REG1_REG_6__SCAN_IN), .S(n11364), .Z(
        n11379) );
  OR2_X1 U13308 ( .A1(n11378), .A2(n11379), .ZN(n11380) );
  NAND2_X1 U13309 ( .A1(n11364), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U13310 ( .A1(n11380), .A2(n11369), .ZN(n11367) );
  INV_X1 U13311 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11365) );
  MUX2_X1 U13312 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n11365), .S(n11420), .Z(
        n11366) );
  NAND2_X1 U13313 ( .A1(n11367), .A2(n11366), .ZN(n11422) );
  MUX2_X1 U13314 ( .A(n11365), .B(P1_REG1_REG_7__SCAN_IN), .S(n11420), .Z(
        n11368) );
  NAND3_X1 U13315 ( .A1(n11380), .A2(n11369), .A3(n11368), .ZN(n11370) );
  NAND3_X1 U13316 ( .A1(n15807), .A2(n11422), .A3(n11370), .ZN(n11371) );
  OAI211_X1 U13317 ( .C1(n11442), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        P1_U3250) );
  INV_X1 U13318 ( .A(n16294), .ZN(n15791) );
  OR3_X1 U13319 ( .A1(n11408), .A2(n11375), .A3(n11374), .ZN(n11376) );
  NAND3_X1 U13320 ( .A1(n15797), .A2(n11377), .A3(n11376), .ZN(n11385) );
  NAND2_X1 U13321 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n12070) );
  AOI21_X1 U13322 ( .B1(n11379), .B2(n11378), .A(n16297), .ZN(n11381) );
  NAND2_X1 U13323 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  NAND2_X1 U13324 ( .A1(n12070), .A2(n11382), .ZN(n11383) );
  AOI21_X1 U13325 ( .B1(n16283), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11383), .ZN(
        n11384) );
  OAI211_X1 U13326 ( .C1(n15791), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        P1_U3249) );
  AOI22_X1 U13327 ( .A1(n11587), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n12848), .ZN(n11387) );
  OAI21_X1 U13328 ( .B1(n11450), .B2(n13259), .A(n11387), .ZN(P1_U3346) );
  AOI211_X1 U13329 ( .C1(n11389), .C2(n11388), .A(n15779), .B(n16291), .ZN(
        n11399) );
  MUX2_X1 U13330 ( .A(n11356), .B(P1_REG1_REG_3__SCAN_IN), .S(n11390), .Z(
        n11392) );
  NAND3_X1 U13331 ( .A1(n15766), .A2(n11392), .A3(n11391), .ZN(n11393) );
  NAND3_X1 U13332 ( .A1(n15807), .A2(n15785), .A3(n11393), .ZN(n11396) );
  NAND2_X1 U13333 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n11864) );
  INV_X1 U13334 ( .A(n11864), .ZN(n11394) );
  AOI21_X1 U13335 ( .B1(n16283), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n11394), .ZN(
        n11395) );
  OAI211_X1 U13336 ( .C1(n15791), .C2(n11397), .A(n11396), .B(n11395), .ZN(
        n11398) );
  OR2_X1 U13337 ( .A1(n11399), .A2(n11398), .ZN(P1_U3246) );
  OAI21_X1 U13338 ( .B1(n11402), .B2(n11401), .A(n11400), .ZN(n11411) );
  INV_X1 U13339 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n16340) );
  NAND2_X1 U13340 ( .A1(n16294), .A2(n11403), .ZN(n11404) );
  NAND2_X1 U13341 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11988) );
  OAI211_X1 U13342 ( .C1(n16340), .C2(n16301), .A(n11404), .B(n11988), .ZN(
        n11410) );
  AND3_X1 U13343 ( .A1(n15776), .A2(n11406), .A3(n11405), .ZN(n11407) );
  NOR3_X1 U13344 ( .A1(n16291), .A2(n11408), .A3(n11407), .ZN(n11409) );
  AOI211_X1 U13345 ( .C1(n15807), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        n11412) );
  INV_X1 U13346 ( .A(n11412), .ZN(P1_U3248) );
  NOR2_X1 U13347 ( .A1(n11413), .A2(n10743), .ZN(n11441) );
  MUX2_X1 U13348 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11414), .S(n11436), .Z(
        n11440) );
  OAI21_X1 U13349 ( .B1(n11442), .B2(n11441), .A(n11440), .ZN(n11439) );
  NAND2_X1 U13350 ( .A1(n11436), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11416) );
  MUX2_X1 U13351 ( .A(n10786), .B(P1_REG2_REG_9__SCAN_IN), .S(n11587), .Z(
        n11415) );
  AOI21_X1 U13352 ( .B1(n11439), .B2(n11416), .A(n11415), .ZN(n11586) );
  NAND3_X1 U13353 ( .A1(n11439), .A2(n11416), .A3(n11415), .ZN(n11417) );
  NAND2_X1 U13354 ( .A1(n11417), .A2(n15797), .ZN(n11432) );
  AND2_X1 U13355 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12898) );
  INV_X1 U13356 ( .A(n11587), .ZN(n11418) );
  NOR2_X1 U13357 ( .A1(n15791), .A2(n11418), .ZN(n11419) );
  AOI211_X1 U13358 ( .C1(n16283), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n12898), .B(
        n11419), .ZN(n11431) );
  NAND2_X1 U13359 ( .A1(n11420), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11421) );
  AND2_X1 U13360 ( .A1(n11422), .A2(n11421), .ZN(n11434) );
  MUX2_X1 U13361 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10759), .S(n11436), .Z(
        n11435) );
  NAND2_X1 U13362 ( .A1(n11434), .A2(n11435), .ZN(n11433) );
  INV_X1 U13363 ( .A(n11433), .ZN(n11424) );
  MUX2_X1 U13364 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10785), .S(n11587), .Z(
        n11426) );
  OR2_X1 U13365 ( .A1(n11436), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11425) );
  INV_X1 U13366 ( .A(n11425), .ZN(n11423) );
  NOR3_X1 U13367 ( .A1(n11424), .A2(n11426), .A3(n11423), .ZN(n11429) );
  NAND2_X1 U13368 ( .A1(n11433), .A2(n11425), .ZN(n11427) );
  NAND2_X1 U13369 ( .A1(n11427), .A2(n11426), .ZN(n11582) );
  INV_X1 U13370 ( .A(n11582), .ZN(n11428) );
  OAI21_X1 U13371 ( .B1(n11429), .B2(n11428), .A(n15807), .ZN(n11430) );
  OAI211_X1 U13372 ( .C1(n11586), .C2(n11432), .A(n11431), .B(n11430), .ZN(
        P1_U3252) );
  OAI21_X1 U13373 ( .B1(n11435), .B2(n11434), .A(n11433), .ZN(n11447) );
  INV_X1 U13374 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U13375 ( .A1(n16294), .A2(n11436), .ZN(n11437) );
  NAND2_X1 U13376 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12573) );
  OAI211_X1 U13377 ( .C1(n11438), .C2(n16301), .A(n11437), .B(n12573), .ZN(
        n11446) );
  INV_X1 U13378 ( .A(n11439), .ZN(n11444) );
  NOR3_X1 U13379 ( .A1(n11442), .A2(n11441), .A3(n11440), .ZN(n11443) );
  NOR3_X1 U13380 ( .A1(n11444), .A2(n11443), .A3(n16291), .ZN(n11445) );
  AOI211_X1 U13381 ( .C1(n15807), .C2(n11447), .A(n11446), .B(n11445), .ZN(
        n11448) );
  INV_X1 U13382 ( .A(n11448), .ZN(P1_U3251) );
  INV_X1 U13383 ( .A(n12534), .ZN(n11858) );
  OAI222_X1 U13384 ( .A1(P2_U3088), .A2(n11858), .B1(n15626), .B2(n11450), 
        .C1(n11449), .C2(n15628), .ZN(P2_U3318) );
  OAI222_X1 U13385 ( .A1(P3_U3151), .A2(n14531), .B1(n14959), .B2(n11452), 
        .C1(n14968), .C2(n11451), .ZN(P3_U3282) );
  INV_X1 U13386 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n11453) );
  OAI222_X1 U13387 ( .A1(P2_U3088), .A2(n12535), .B1(n15626), .B2(n11454), 
        .C1(n11453), .C2(n15628), .ZN(P2_U3317) );
  INV_X1 U13388 ( .A(n11588), .ZN(n11631) );
  OAI222_X1 U13389 ( .A1(n16174), .A2(n11455), .B1(n13259), .B2(n11454), .C1(
        n11631), .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U13390 ( .A1(n11682), .A2(n11456), .ZN(n11457) );
  AND2_X1 U13391 ( .A1(n11457), .A2(n9870), .ZN(n11458) );
  OR2_X1 U13392 ( .A1(n11459), .A2(n11458), .ZN(n11478) );
  NOR2_X1 U13393 ( .A1(n11478), .A2(P2_U3088), .ZN(n16224) );
  INV_X1 U13394 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n11481) );
  INV_X1 U13395 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11460) );
  AND2_X1 U13396 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15107) );
  NAND2_X1 U13397 ( .A1(n15108), .A2(n15107), .ZN(n15106) );
  NAND2_X1 U13398 ( .A1(n15100), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U13399 ( .A1(n15106), .A2(n11461), .ZN(n16225) );
  INV_X1 U13400 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11462) );
  XNOR2_X1 U13401 ( .A(n16228), .B(n11462), .ZN(n16226) );
  XNOR2_X1 U13402 ( .A(n11485), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n11465) );
  NOR2_X1 U13403 ( .A1(n11466), .A2(n11465), .ZN(n11482) );
  NAND2_X1 U13404 ( .A1(n11463), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15614) );
  NOR2_X1 U13405 ( .A1(n15614), .A2(n11467), .ZN(n11464) );
  AOI211_X1 U13406 ( .C1(n11466), .C2(n11465), .A(n11482), .B(n16264), .ZN(
        n11476) );
  NAND2_X1 U13407 ( .A1(n11467), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15618) );
  NOR2_X1 U13408 ( .A1(n15618), .A2(n10566), .ZN(n11468) );
  INV_X1 U13409 ( .A(n16257), .ZN(n16272) );
  INV_X1 U13410 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11469) );
  MUX2_X1 U13411 ( .A(n11469), .B(P2_REG2_REG_1__SCAN_IN), .S(n15100), .Z(
        n15102) );
  INV_X1 U13412 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11525) );
  NOR3_X1 U13413 ( .A1(n15102), .A2(n11525), .A3(n15103), .ZN(n15101) );
  AOI21_X1 U13414 ( .B1(n15100), .B2(P2_REG2_REG_1__SCAN_IN), .A(n15101), .ZN(
        n16233) );
  INV_X1 U13415 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n12096) );
  MUX2_X1 U13416 ( .A(n12096), .B(P2_REG2_REG_2__SCAN_IN), .S(n16228), .Z(
        n16232) );
  NOR2_X1 U13417 ( .A1(n16233), .A2(n16232), .ZN(n16231) );
  AND2_X1 U13418 ( .A1(n16228), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11472) );
  MUX2_X1 U13419 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11470), .S(n11485), .Z(
        n11471) );
  OAI21_X1 U13420 ( .B1(n16231), .B2(n11472), .A(n11471), .ZN(n11488) );
  INV_X1 U13421 ( .A(n11488), .ZN(n11474) );
  NOR3_X1 U13422 ( .A1(n16231), .A2(n11472), .A3(n11471), .ZN(n11473) );
  NOR3_X1 U13423 ( .A1(n16272), .A2(n11474), .A3(n11473), .ZN(n11475) );
  NOR2_X1 U13424 ( .A1(n11476), .A2(n11475), .ZN(n11480) );
  AND2_X1 U13425 ( .A1(n10566), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11477) );
  AOI22_X1 U13426 ( .A1(n16270), .A2(n11485), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11479) );
  OAI211_X1 U13427 ( .C1(n16278), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        P2_U3217) );
  AOI21_X1 U13428 ( .B1(n11485), .B2(P2_REG1_REG_3__SCAN_IN), .A(n11482), .ZN(
        n11484) );
  XNOR2_X1 U13429 ( .A(n11495), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n11483) );
  NOR2_X1 U13430 ( .A1(n11484), .A2(n11483), .ZN(n11494) );
  AOI211_X1 U13431 ( .C1(n11484), .C2(n11483), .A(n11494), .B(n16264), .ZN(
        n11491) );
  NAND2_X1 U13432 ( .A1(n11485), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n11487) );
  MUX2_X1 U13433 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n12107), .S(n11500), .Z(
        n11486) );
  AOI21_X1 U13434 ( .B1(n11488), .B2(n11487), .A(n11486), .ZN(n11515) );
  AND3_X1 U13435 ( .A1(n11488), .A2(n11487), .A3(n11486), .ZN(n11489) );
  NOR3_X1 U13436 ( .A1(n16272), .A2(n11515), .A3(n11489), .ZN(n11490) );
  NOR2_X1 U13437 ( .A1(n11491), .A2(n11490), .ZN(n11493) );
  AND2_X1 U13438 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n11824) );
  AOI21_X1 U13439 ( .B1(n16270), .B2(n11495), .A(n11824), .ZN(n11492) );
  OAI211_X1 U13440 ( .C1(n16278), .C2(n8590), .A(n11493), .B(n11492), .ZN(
        P2_U3218) );
  INV_X1 U13441 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n11508) );
  AND2_X1 U13442 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n11978) );
  MUX2_X1 U13443 ( .A(n11496), .B(P2_REG1_REG_5__SCAN_IN), .S(n11520), .Z(
        n11510) );
  XNOR2_X1 U13444 ( .A(n11547), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n11497) );
  AOI211_X1 U13445 ( .C1(n11498), .C2(n11497), .A(n16264), .B(n11546), .ZN(
        n11499) );
  AOI211_X1 U13446 ( .C1(n16270), .C2(n11547), .A(n11978), .B(n11499), .ZN(
        n11507) );
  NOR2_X1 U13447 ( .A1(n11500), .A2(n12107), .ZN(n11514) );
  MUX2_X1 U13448 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11501), .S(n11520), .Z(
        n11513) );
  OAI21_X1 U13449 ( .B1(n11515), .B2(n11514), .A(n11513), .ZN(n11512) );
  NAND2_X1 U13450 ( .A1(n11520), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11503) );
  MUX2_X1 U13451 ( .A(n12142), .B(P2_REG2_REG_6__SCAN_IN), .S(n11547), .Z(
        n11502) );
  AOI21_X1 U13452 ( .B1(n11512), .B2(n11503), .A(n11502), .ZN(n11555) );
  INV_X1 U13453 ( .A(n11555), .ZN(n11505) );
  NAND3_X1 U13454 ( .A1(n11512), .A2(n11503), .A3(n11502), .ZN(n11504) );
  NAND3_X1 U13455 ( .A1(n11505), .A2(n16257), .A3(n11504), .ZN(n11506) );
  OAI211_X1 U13456 ( .C1(n11508), .C2(n16278), .A(n11507), .B(n11506), .ZN(
        P2_U3220) );
  INV_X1 U13457 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n11523) );
  AOI211_X1 U13458 ( .C1(n11511), .C2(n11510), .A(n16264), .B(n11509), .ZN(
        n11519) );
  INV_X1 U13459 ( .A(n11512), .ZN(n11517) );
  NOR3_X1 U13460 ( .A1(n11515), .A2(n11514), .A3(n11513), .ZN(n11516) );
  NOR3_X1 U13461 ( .A1(n16272), .A2(n11517), .A3(n11516), .ZN(n11518) );
  NOR2_X1 U13462 ( .A1(n11519), .A2(n11518), .ZN(n11522) );
  AND2_X1 U13463 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15019) );
  AOI21_X1 U13464 ( .B1(n16270), .B2(n11520), .A(n15019), .ZN(n11521) );
  OAI211_X1 U13465 ( .C1(n16278), .C2(n11523), .A(n11522), .B(n11521), .ZN(
        P2_U3219) );
  OAI22_X1 U13466 ( .A1(n16272), .A2(n11525), .B1(n11524), .B2(n16264), .ZN(
        n11528) );
  INV_X1 U13467 ( .A(n16270), .ZN(n15128) );
  NAND2_X1 U13468 ( .A1(n16257), .A2(n11525), .ZN(n11526) );
  OAI211_X1 U13469 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n16264), .A(n15128), .B(
        n11526), .ZN(n11527) );
  MUX2_X1 U13470 ( .A(n11528), .B(n11527), .S(P2_IR_REG_0__SCAN_IN), .Z(n11529) );
  INV_X1 U13471 ( .A(n11529), .ZN(n11531) );
  AOI22_X1 U13472 ( .A1(n16224), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11530) );
  NAND2_X1 U13473 ( .A1(n11531), .A2(n11530), .ZN(P2_U3214) );
  OAI222_X1 U13474 ( .A1(P3_U3151), .A2(n11534), .B1(n14968), .B2(n11533), 
        .C1(n14959), .C2(n11532), .ZN(P3_U3281) );
  XOR2_X1 U13475 ( .A(n11536), .B(n11535), .Z(n15760) );
  INV_X1 U13476 ( .A(n15691), .ZN(n16716) );
  AND2_X1 U13477 ( .A1(n15757), .A2(n15956), .ZN(n11577) );
  AOI22_X1 U13478 ( .A1(n16716), .A2(n11577), .B1(n13584), .B2(n16719), .ZN(
        n11540) );
  AND2_X1 U13479 ( .A1(n11537), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11614) );
  INV_X1 U13480 ( .A(n11614), .ZN(n11538) );
  NAND2_X1 U13481 ( .A1(n11538), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n11539) );
  OAI211_X1 U13482 ( .C1(n15760), .C2(n15729), .A(n11540), .B(n11539), .ZN(
        P1_U3232) );
  INV_X1 U13483 ( .A(n11541), .ZN(n11543) );
  OAI222_X1 U13484 ( .A1(n12537), .A2(P2_U3088), .B1(n15626), .B2(n11543), 
        .C1(n11542), .C2(n15628), .ZN(P2_U3316) );
  INV_X1 U13485 ( .A(n11645), .ZN(n11640) );
  OAI222_X1 U13486 ( .A1(n11544), .A2(n16174), .B1(P1_U3086), .B2(n11640), 
        .C1(n16178), .C2(n11543), .ZN(P1_U3344) );
  AND2_X1 U13487 ( .A1(n11750), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13488 ( .A1(n11750), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13489 ( .A1(n11750), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13490 ( .A1(n11750), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13491 ( .A1(n11750), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13492 ( .A1(n11750), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13493 ( .A1(n11750), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13494 ( .A1(n11750), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13495 ( .A1(n11750), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13496 ( .A1(n11750), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13497 ( .A1(n11750), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13498 ( .A1(n11750), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13499 ( .A1(n11750), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13500 ( .A1(n11750), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13501 ( .A1(n11750), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13502 ( .A1(n11750), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  MUX2_X1 U13503 ( .A(n11548), .B(P2_REG1_REG_7__SCAN_IN), .S(n11740), .Z(
        n11549) );
  NOR2_X1 U13504 ( .A1(n11550), .A2(n11549), .ZN(n11736) );
  AOI211_X1 U13505 ( .C1(n11550), .C2(n11549), .A(n16264), .B(n11736), .ZN(
        n11562) );
  NOR2_X1 U13506 ( .A1(n11551), .A2(n12142), .ZN(n11554) );
  INV_X1 U13507 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11552) );
  MUX2_X1 U13508 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11552), .S(n11740), .Z(
        n11553) );
  OAI21_X1 U13509 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n11743) );
  INV_X1 U13510 ( .A(n11743), .ZN(n11557) );
  NOR3_X1 U13511 ( .A1(n11555), .A2(n11554), .A3(n11553), .ZN(n11556) );
  NOR3_X1 U13512 ( .A1(n11557), .A2(n11556), .A3(n16272), .ZN(n11558) );
  AOI21_X1 U13513 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(n16224), .A(n11558), .ZN(
        n11559) );
  NAND2_X1 U13514 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n12222) );
  OAI211_X1 U13515 ( .C1(n11560), .C2(n15128), .A(n11559), .B(n12222), .ZN(
        n11561) );
  OR2_X1 U13516 ( .A1(n11562), .A2(n11561), .ZN(P2_U3221) );
  INV_X1 U13517 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14303) );
  INV_X1 U13518 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U13519 ( .A1(n13829), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11564) );
  NAND2_X1 U13520 ( .A1(n13830), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11563) );
  OAI211_X1 U13521 ( .C1(n10679), .C2(n11565), .A(n11564), .B(n11563), .ZN(
        n15815) );
  NAND2_X1 U13522 ( .A1(n15815), .A2(P1_U4016), .ZN(n11566) );
  OAI21_X1 U13523 ( .B1(P1_U4016), .B2(n14303), .A(n11566), .ZN(P1_U3591) );
  NAND2_X1 U13524 ( .A1(n15954), .A2(P1_U4016), .ZN(n11567) );
  OAI21_X1 U13525 ( .B1(P1_U4016), .B2(n11568), .A(n11567), .ZN(P1_U3579) );
  NOR2_X1 U13526 ( .A1(n11569), .A2(P1_U3086), .ZN(n13902) );
  INV_X1 U13527 ( .A(n11570), .ZN(n11572) );
  NAND4_X1 U13528 ( .A1(n13902), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11771) );
  INV_X2 U13529 ( .A(n16709), .ZN(n16694) );
  NAND2_X1 U13530 ( .A1(n8099), .A2(n16474), .ZN(n11575) );
  AND2_X1 U13531 ( .A1(n11576), .A2(n11575), .ZN(n16473) );
  AOI21_X1 U13532 ( .B1(n16702), .B2(n16619), .A(n16473), .ZN(n11578) );
  NOR2_X1 U13533 ( .A1(n11578), .A2(n11577), .ZN(n16480) );
  NAND3_X1 U13534 ( .A1(n13850), .A2(n10650), .A3(n13839), .ZN(n16602) );
  OR2_X1 U13535 ( .A1(n16473), .A2(n16602), .ZN(n11579) );
  OAI211_X1 U13536 ( .C1(n10815), .C2(n16474), .A(n16480), .B(n11579), .ZN(
        n16143) );
  NAND2_X1 U13537 ( .A1(n16143), .A2(n16694), .ZN(n11580) );
  OAI21_X1 U13538 ( .B1(n16694), .B2(n10656), .A(n11580), .ZN(P1_U3459) );
  MUX2_X1 U13539 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11082), .S(n11645), .Z(
        n11585) );
  OR2_X1 U13540 ( .A1(n11587), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U13541 ( .A1(n11582), .A2(n11581), .ZN(n11620) );
  INV_X1 U13542 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n16660) );
  MUX2_X1 U13543 ( .A(n16660), .B(P1_REG1_REG_10__SCAN_IN), .S(n11588), .Z(
        n11619) );
  OR2_X1 U13544 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U13545 ( .A1(n11588), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11583) );
  AND2_X1 U13546 ( .A1(n11621), .A2(n11583), .ZN(n11584) );
  NAND2_X1 U13547 ( .A1(n11584), .A2(n11585), .ZN(n11649) );
  OAI21_X1 U13548 ( .B1(n11585), .B2(n11584), .A(n11649), .ZN(n11598) );
  AOI21_X1 U13549 ( .B1(n11587), .B2(P1_REG2_REG_9__SCAN_IN), .A(n11586), .ZN(
        n11625) );
  MUX2_X1 U13550 ( .A(n12886), .B(P1_REG2_REG_10__SCAN_IN), .S(n11588), .Z(
        n11624) );
  NOR2_X1 U13551 ( .A1(n11625), .A2(n11624), .ZN(n11623) );
  NOR2_X1 U13552 ( .A1(n11631), .A2(n12886), .ZN(n11592) );
  INV_X1 U13553 ( .A(n11592), .ZN(n11590) );
  INV_X1 U13554 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11639) );
  MUX2_X1 U13555 ( .A(n11639), .B(P1_REG2_REG_11__SCAN_IN), .S(n11645), .Z(
        n11589) );
  NAND2_X1 U13556 ( .A1(n11590), .A2(n11589), .ZN(n11593) );
  MUX2_X1 U13557 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11639), .S(n11645), .Z(
        n11591) );
  OAI21_X1 U13558 ( .B1(n11623), .B2(n11592), .A(n11591), .ZN(n11638) );
  OAI211_X1 U13559 ( .C1(n11623), .C2(n11593), .A(n11638), .B(n15797), .ZN(
        n11596) );
  NOR2_X1 U13560 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13218), .ZN(n11594) );
  AOI21_X1 U13561 ( .B1(n16283), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n11594), 
        .ZN(n11595) );
  OAI211_X1 U13562 ( .C1(n11640), .C2(n15791), .A(n11596), .B(n11595), .ZN(
        n11597) );
  AOI21_X1 U13563 ( .B1(n15807), .B2(n11598), .A(n11597), .ZN(n11599) );
  INV_X1 U13564 ( .A(n11599), .ZN(P1_U3254) );
  INV_X1 U13565 ( .A(n11600), .ZN(n11602) );
  OAI222_X1 U13566 ( .A1(n14959), .A2(n11603), .B1(n14968), .B2(n11602), .C1(
        P3_U3151), .C2(n11601), .ZN(P3_U3280) );
  OAI21_X1 U13567 ( .B1(n11606), .B2(n11605), .A(n11604), .ZN(n11609) );
  OAI22_X1 U13568 ( .A1(n11614), .A2(n12458), .B1(n15712), .B2(n13580), .ZN(
        n11608) );
  OAI22_X1 U13569 ( .A1(n11775), .A2(n15717), .B1(n15716), .B2(n10675), .ZN(
        n11607) );
  AOI211_X1 U13570 ( .C1(n11609), .C2(n16714), .A(n11608), .B(n11607), .ZN(
        n11610) );
  INV_X1 U13571 ( .A(n11610), .ZN(P1_U3237) );
  OAI21_X1 U13572 ( .B1(n11613), .B2(n11612), .A(n11611), .ZN(n11617) );
  OAI22_X1 U13573 ( .A1(n11614), .A2(n12423), .B1(n15712), .B2(n11762), .ZN(
        n11616) );
  OAI22_X1 U13574 ( .A1(n11764), .A2(n15716), .B1(n15717), .B2(n13581), .ZN(
        n11615) );
  AOI211_X1 U13575 ( .C1(n11617), .C2(n16714), .A(n11616), .B(n11615), .ZN(
        n11618) );
  INV_X1 U13576 ( .A(n11618), .ZN(P1_U3222) );
  AOI21_X1 U13577 ( .B1(n11620), .B2(n11619), .A(n16297), .ZN(n11622) );
  NAND2_X1 U13578 ( .A1(n11622), .A2(n11621), .ZN(n11630) );
  NAND2_X1 U13579 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n13018)
         );
  AOI211_X1 U13580 ( .C1(n11625), .C2(n11624), .A(n11623), .B(n16291), .ZN(
        n11626) );
  INV_X1 U13581 ( .A(n11626), .ZN(n11627) );
  NAND2_X1 U13582 ( .A1(n13018), .A2(n11627), .ZN(n11628) );
  AOI21_X1 U13583 ( .B1(n16283), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11628), 
        .ZN(n11629) );
  OAI211_X1 U13584 ( .C1(n15791), .C2(n11631), .A(n11630), .B(n11629), .ZN(
        P1_U3253) );
  AOI22_X1 U13585 ( .A1(n15804), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n12848), .ZN(n11632) );
  OAI21_X1 U13586 ( .B1(n11699), .B2(n13259), .A(n11632), .ZN(P1_U3342) );
  INV_X1 U13587 ( .A(n12946), .ZN(n12950) );
  INV_X1 U13588 ( .A(n11633), .ZN(n11635) );
  OAI222_X1 U13589 ( .A1(P2_U3088), .A2(n12950), .B1(n15626), .B2(n11635), 
        .C1(n11634), .C2(n15628), .ZN(P2_U3315) );
  INV_X1 U13590 ( .A(n11883), .ZN(n11874) );
  OAI222_X1 U13591 ( .A1(n16174), .A2(n11636), .B1(n13259), .B2(n11635), .C1(
        n11874), .C2(P1_U3086), .ZN(P1_U3343) );
  MUX2_X1 U13592 ( .A(n11637), .B(P1_REG2_REG_12__SCAN_IN), .S(n11883), .Z(
        n11642) );
  OAI21_X1 U13593 ( .B1(n11640), .B2(n11639), .A(n11638), .ZN(n11641) );
  NOR2_X1 U13594 ( .A1(n11641), .A2(n11642), .ZN(n11873) );
  AOI21_X1 U13595 ( .B1(n11642), .B2(n11641), .A(n11873), .ZN(n11656) );
  INV_X1 U13596 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11643) );
  NAND2_X1 U13597 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n13327)
         );
  OAI21_X1 U13598 ( .B1(n16301), .B2(n11643), .A(n13327), .ZN(n11644) );
  AOI21_X1 U13599 ( .B1(n11883), .B2(n16294), .A(n11644), .ZN(n11655) );
  INV_X1 U13600 ( .A(n11649), .ZN(n11647) );
  MUX2_X1 U13601 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10985), .S(n11883), .Z(
        n11650) );
  OR2_X1 U13602 ( .A1(n11645), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11648) );
  INV_X1 U13603 ( .A(n11648), .ZN(n11646) );
  NOR3_X1 U13604 ( .A1(n11647), .A2(n11650), .A3(n11646), .ZN(n11653) );
  NAND2_X1 U13605 ( .A1(n11649), .A2(n11648), .ZN(n11651) );
  NAND2_X1 U13606 ( .A1(n11651), .A2(n11650), .ZN(n11885) );
  INV_X1 U13607 ( .A(n11885), .ZN(n11652) );
  OAI21_X1 U13608 ( .B1(n11653), .B2(n11652), .A(n15807), .ZN(n11654) );
  OAI211_X1 U13609 ( .C1(n11656), .C2(n16291), .A(n11655), .B(n11654), .ZN(
        P1_U3255) );
  NAND2_X1 U13610 ( .A1(n15215), .A2(P2_U3947), .ZN(n11657) );
  OAI21_X1 U13611 ( .B1(n8577), .B2(P2_U3947), .A(n11657), .ZN(P2_U3553) );
  INV_X1 U13612 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n11659) );
  NAND2_X1 U13613 ( .A1(n14216), .A2(P3_U3897), .ZN(n11658) );
  OAI21_X1 U13614 ( .B1(P3_U3897), .B2(n11659), .A(n11658), .ZN(P3_U3495) );
  NAND2_X1 U13615 ( .A1(n14217), .A2(P3_U3897), .ZN(n11660) );
  OAI21_X1 U13616 ( .B1(P3_U3897), .B2(n11661), .A(n11660), .ZN(P3_U3497) );
  NOR2_X1 U13617 ( .A1(n10575), .A2(n15232), .ZN(n11663) );
  NAND2_X1 U13618 ( .A1(n11663), .A2(n11664), .ZN(n11667) );
  INV_X1 U13619 ( .A(n11663), .ZN(n11666) );
  INV_X1 U13620 ( .A(n11664), .ZN(n11665) );
  NAND2_X1 U13621 ( .A1(n11666), .A2(n11665), .ZN(n11671) );
  NAND2_X1 U13622 ( .A1(n11715), .A2(n7418), .ZN(n11670) );
  NAND2_X1 U13623 ( .A1(n11668), .A2(n11672), .ZN(n11669) );
  AND2_X1 U13624 ( .A1(n11670), .A2(n11669), .ZN(n14062) );
  NAND2_X1 U13625 ( .A1(n14060), .A2(n11671), .ZN(n11702) );
  INV_X2 U13626 ( .A(n7460), .ZN(n15232) );
  NOR2_X1 U13627 ( .A1(n11723), .A2(n15232), .ZN(n11674) );
  XNOR2_X1 U13628 ( .A(n16521), .B(n11672), .ZN(n11673) );
  NAND2_X1 U13629 ( .A1(n11674), .A2(n11673), .ZN(n11677) );
  INV_X1 U13630 ( .A(n11673), .ZN(n11676) );
  INV_X1 U13631 ( .A(n11674), .ZN(n11675) );
  NAND2_X1 U13632 ( .A1(n11676), .A2(n11675), .ZN(n11678) );
  AND2_X1 U13633 ( .A1(n11677), .A2(n11678), .ZN(n11703) );
  NAND2_X1 U13634 ( .A1(n11702), .A2(n11703), .ZN(n11701) );
  NAND2_X1 U13635 ( .A1(n11701), .A2(n11678), .ZN(n11808) );
  XNOR2_X1 U13636 ( .A(n12282), .B(n11679), .ZN(n11810) );
  OR2_X1 U13637 ( .A1(n11832), .A2(n15232), .ZN(n11811) );
  XNOR2_X1 U13638 ( .A(n11810), .B(n11811), .ZN(n11809) );
  XNOR2_X1 U13639 ( .A(n11808), .B(n11809), .ZN(n11697) );
  OR2_X1 U13640 ( .A1(n16222), .A2(n11680), .ZN(n11690) );
  INV_X1 U13641 ( .A(n11690), .ZN(n11681) );
  NAND2_X1 U13642 ( .A1(n11681), .A2(n16223), .ZN(n11688) );
  INV_X1 U13643 ( .A(n11682), .ZN(n11683) );
  NAND2_X1 U13644 ( .A1(n16520), .A2(n11683), .ZN(n11684) );
  OR2_X1 U13645 ( .A1(n11688), .A2(n11685), .ZN(n15076) );
  OAI22_X1 U13646 ( .A1(n11942), .A2(n15162), .B1(n11723), .B2(n15043), .ZN(
        n11725) );
  INV_X1 U13647 ( .A(n11686), .ZN(n11687) );
  OR2_X1 U13648 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  INV_X1 U13649 ( .A(n12282), .ZN(n11833) );
  AOI22_X1 U13650 ( .A1(n15033), .A2(n11725), .B1(n15080), .B2(n11833), .ZN(
        n11696) );
  NAND2_X1 U13651 ( .A1(n11690), .A2(n11709), .ZN(n11691) );
  NAND2_X1 U13652 ( .A1(n11691), .A2(n11710), .ZN(n11705) );
  INV_X1 U13653 ( .A(n11692), .ZN(n11693) );
  OR2_X1 U13654 ( .A1(n11705), .A2(n11693), .ZN(n11694) );
  INV_X1 U13655 ( .A(n15074), .ZN(n15052) );
  MUX2_X1 U13656 ( .A(n15052), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n11695) );
  OAI211_X1 U13657 ( .C1(n11697), .C2(n15077), .A(n11696), .B(n11695), .ZN(
        P2_U3190) );
  INV_X1 U13658 ( .A(n13105), .ZN(n11700) );
  INV_X1 U13659 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11698) );
  OAI222_X1 U13660 ( .A1(P2_U3088), .A2(n11700), .B1(n15626), .B2(n11699), 
        .C1(n11698), .C2(n15628), .ZN(P2_U3314) );
  INV_X1 U13661 ( .A(n15080), .ZN(n15066) );
  OAI21_X1 U13662 ( .B1(n11703), .B2(n11702), .A(n11701), .ZN(n11704) );
  NAND2_X1 U13663 ( .A1(n11704), .A2(n15070), .ZN(n11707) );
  OAI22_X1 U13664 ( .A1(n11832), .A2(n15162), .B1(n10575), .B2(n15043), .ZN(
        n12093) );
  INV_X1 U13665 ( .A(n16223), .ZN(n16220) );
  OR2_X1 U13666 ( .A1(n11705), .A2(n16220), .ZN(n14058) );
  AOI22_X1 U13667 ( .A1(n15033), .A2(n12093), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14058), .ZN(n11706) );
  OAI211_X1 U13668 ( .C1(n16521), .C2(n15066), .A(n11707), .B(n11706), .ZN(
        P2_U3209) );
  OR2_X1 U13669 ( .A1(n11708), .A2(n16220), .ZN(n16215) );
  NAND3_X1 U13670 ( .A1(n11711), .A2(n11710), .A3(n11709), .ZN(n11712) );
  INV_X1 U13671 ( .A(n16222), .ZN(n11713) );
  INV_X1 U13672 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11731) );
  INV_X1 U13673 ( .A(n11714), .ZN(n15543) );
  NAND2_X1 U13674 ( .A1(n10575), .A2(n14066), .ZN(n11717) );
  NAND2_X1 U13675 ( .A1(n11718), .A2(n11717), .ZN(n12103) );
  NAND2_X1 U13676 ( .A1(n12103), .A2(n12102), .ZN(n11720) );
  NAND2_X1 U13677 ( .A1(n11723), .A2(n16521), .ZN(n11719) );
  NAND2_X1 U13678 ( .A1(n11720), .A2(n11719), .ZN(n11828) );
  INV_X1 U13679 ( .A(n11827), .ZN(n11830) );
  XNOR2_X1 U13680 ( .A(n11828), .B(n11830), .ZN(n12286) );
  NAND2_X1 U13681 ( .A1(n11722), .A2(n11721), .ZN(n12092) );
  NAND2_X1 U13682 ( .A1(n11723), .A2(n12101), .ZN(n11724) );
  NAND2_X1 U13683 ( .A1(n12090), .A2(n11724), .ZN(n11831) );
  XNOR2_X1 U13684 ( .A(n11831), .B(n11830), .ZN(n11726) );
  AOI21_X1 U13685 ( .B1(n11726), .B2(n15446), .A(n11725), .ZN(n12289) );
  AND2_X1 U13686 ( .A1(n16521), .A2(n12098), .ZN(n11727) );
  INV_X1 U13687 ( .A(n11727), .ZN(n12097) );
  NAND2_X1 U13688 ( .A1(n11727), .A2(n12282), .ZN(n11839) );
  INV_X1 U13689 ( .A(n11839), .ZN(n11728) );
  AOI211_X1 U13690 ( .C1(n11833), .C2(n12097), .A(n7418), .B(n11728), .ZN(
        n12285) );
  AOI21_X1 U13691 ( .B1(n15546), .B2(n11833), .A(n12285), .ZN(n11729) );
  OAI211_X1 U13692 ( .C1(n15550), .C2(n12286), .A(n12289), .B(n11729), .ZN(
        n12200) );
  NAND2_X1 U13693 ( .A1(n12200), .A2(n16526), .ZN(n11730) );
  OAI21_X1 U13694 ( .B1(n16526), .B2(n11731), .A(n11730), .ZN(P2_U3502) );
  NAND2_X1 U13695 ( .A1(n15070), .A2(n7418), .ZN(n15067) );
  AOI21_X1 U13696 ( .B1(n15099), .B2(n7418), .A(n15077), .ZN(n11732) );
  OAI21_X1 U13697 ( .B1(n11732), .B2(n15080), .A(n11919), .ZN(n11734) );
  NOR2_X1 U13698 ( .A1(n10575), .A2(n15162), .ZN(n11921) );
  AOI22_X1 U13699 ( .A1(n15033), .A2(n11921), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14058), .ZN(n11733) );
  OAI211_X1 U13700 ( .C1(n15067), .C2(n11735), .A(n11734), .B(n11733), .ZN(
        P2_U3204) );
  INV_X1 U13701 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11737) );
  MUX2_X1 U13702 ( .A(n11737), .B(P2_REG1_REG_8__SCAN_IN), .S(n11853), .Z(
        n11738) );
  AOI211_X1 U13703 ( .C1(n11739), .C2(n11738), .A(n16264), .B(n11847), .ZN(
        n11749) );
  NAND2_X1 U13704 ( .A1(n11740), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11742) );
  MUX2_X1 U13705 ( .A(n12494), .B(P2_REG2_REG_8__SCAN_IN), .S(n11853), .Z(
        n11741) );
  AOI21_X1 U13706 ( .B1(n11743), .B2(n11742), .A(n11741), .ZN(n11852) );
  AND3_X1 U13707 ( .A1(n11743), .A2(n11742), .A3(n11741), .ZN(n11744) );
  NOR3_X1 U13708 ( .A1(n11852), .A2(n11744), .A3(n16272), .ZN(n11748) );
  NAND2_X1 U13709 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U13710 ( .A1(n16224), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n11745) );
  OAI211_X1 U13711 ( .C1(n15128), .C2(n11746), .A(n12330), .B(n11745), .ZN(
        n11747) );
  OR3_X1 U13712 ( .A1(n11749), .A2(n11748), .A3(n11747), .ZN(P2_U3222) );
  AND2_X1 U13713 ( .A1(n11750), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13714 ( .A1(n11750), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13715 ( .A1(n11750), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13716 ( .A1(n11750), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13717 ( .A1(n11750), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13718 ( .A1(n11750), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13719 ( .A1(n11750), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13720 ( .A1(n11750), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13721 ( .A1(n11750), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13722 ( .A1(n11750), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13723 ( .A1(n11750), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13724 ( .A1(n11750), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13725 ( .A1(n11750), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13726 ( .A1(n11750), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  INV_X1 U13727 ( .A(n11751), .ZN(n11752) );
  OAI222_X1 U13728 ( .A1(P3_U3151), .A2(n14553), .B1(n14959), .B2(n11753), 
        .C1(n14968), .C2(n11752), .ZN(P3_U3279) );
  INV_X1 U13729 ( .A(n11754), .ZN(n11757) );
  AOI211_X1 U13730 ( .C1(n11714), .C2(n11757), .A(n11756), .B(n11755), .ZN(
        n11911) );
  AOI22_X1 U13731 ( .A1(n15536), .A2(n9876), .B1(n16525), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n11758) );
  OAI21_X1 U13732 ( .B1(n11911), .B2(n16525), .A(n11758), .ZN(P2_U3500) );
  INV_X1 U13733 ( .A(n16602), .ZN(n16691) );
  INV_X1 U13734 ( .A(n11759), .ZN(n11760) );
  INV_X1 U13735 ( .A(n11768), .ZN(n12428) );
  OAI211_X1 U13736 ( .C1(n11762), .C2(n16474), .A(n16698), .B(n11784), .ZN(
        n12424) );
  OAI21_X1 U13737 ( .B1(n11762), .B2(n16684), .A(n12424), .ZN(n11769) );
  OAI22_X1 U13738 ( .A1(n11764), .A2(n16031), .B1(n13581), .B2(n16029), .ZN(
        n11765) );
  AOI21_X1 U13739 ( .B1(n11766), .B2(n16623), .A(n11765), .ZN(n11767) );
  OAI21_X1 U13740 ( .B1(n11768), .B2(n16619), .A(n11767), .ZN(n12427) );
  AOI211_X1 U13741 ( .C1(n16691), .C2(n12428), .A(n11769), .B(n12427), .ZN(
        n16488) );
  NAND2_X1 U13742 ( .A1(n16707), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11772) );
  OAI21_X1 U13743 ( .B1(n16488), .B2(n16707), .A(n11772), .ZN(P1_U3529) );
  OAI21_X1 U13744 ( .B1(n11774), .B2(n11777), .A(n11773), .ZN(n11783) );
  INV_X1 U13745 ( .A(n11783), .ZN(n12460) );
  INV_X1 U13746 ( .A(n16619), .ZN(n16579) );
  OAI22_X1 U13747 ( .A1(n11775), .A2(n16029), .B1(n10675), .B2(n16031), .ZN(
        n11782) );
  NAND3_X1 U13748 ( .A1(n11778), .A2(n11777), .A3(n11776), .ZN(n11779) );
  AOI21_X1 U13749 ( .B1(n11780), .B2(n11779), .A(n16702), .ZN(n11781) );
  AOI211_X1 U13750 ( .C1(n16579), .C2(n11783), .A(n11782), .B(n11781), .ZN(
        n12464) );
  AOI21_X1 U13751 ( .B1(n11784), .B2(n8105), .A(n16686), .ZN(n11785) );
  AND2_X1 U13752 ( .A1(n11785), .A2(n11793), .ZN(n12457) );
  AOI21_X1 U13753 ( .B1(n16696), .B2(n8105), .A(n12457), .ZN(n11786) );
  OAI211_X1 U13754 ( .C1(n12460), .C2(n16602), .A(n12464), .B(n11786), .ZN(
        n11788) );
  NAND2_X1 U13755 ( .A1(n11788), .A2(n16694), .ZN(n11787) );
  OAI21_X1 U13756 ( .B1(n16694), .B2(n10678), .A(n11787), .ZN(P1_U3465) );
  NAND2_X1 U13757 ( .A1(n11788), .A2(n16708), .ZN(n11789) );
  OAI21_X1 U13758 ( .B1(n16708), .B2(n11350), .A(n11789), .ZN(P1_U3530) );
  XNOR2_X1 U13759 ( .A(n11790), .B(n11797), .ZN(n12445) );
  NAND2_X1 U13760 ( .A1(n15754), .A2(n15956), .ZN(n11792) );
  NAND2_X1 U13761 ( .A1(n15756), .A2(n15955), .ZN(n11791) );
  NAND2_X1 U13762 ( .A1(n11792), .A2(n11791), .ZN(n12434) );
  NAND2_X1 U13763 ( .A1(n11793), .A2(n13607), .ZN(n11794) );
  NAND2_X1 U13764 ( .A1(n11794), .A2(n16698), .ZN(n11795) );
  NOR2_X1 U13765 ( .A1(n12448), .A2(n11795), .ZN(n12433) );
  AOI211_X1 U13766 ( .C1(n16696), .C2(n13607), .A(n12434), .B(n12433), .ZN(
        n11800) );
  OAI21_X1 U13767 ( .B1(n11798), .B2(n11797), .A(n11796), .ZN(n12443) );
  NAND2_X1 U13768 ( .A1(n12443), .A2(n16705), .ZN(n11799) );
  OAI211_X1 U13769 ( .C1(n12445), .C2(n16702), .A(n11800), .B(n11799), .ZN(
        n11802) );
  NAND2_X1 U13770 ( .A1(n11802), .A2(n16694), .ZN(n11801) );
  OAI21_X1 U13771 ( .B1(n16694), .B2(n10690), .A(n11801), .ZN(P1_U3468) );
  NAND2_X1 U13772 ( .A1(n11802), .A2(n16708), .ZN(n11803) );
  OAI21_X1 U13773 ( .B1(n16708), .B2(n11356), .A(n11803), .ZN(P1_U3531) );
  INV_X1 U13774 ( .A(n11804), .ZN(n11806) );
  OAI222_X1 U13775 ( .A1(n14959), .A2(n11807), .B1(n14968), .B2(n11806), .C1(
        n11805), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13776 ( .A(n11810), .ZN(n11813) );
  INV_X1 U13777 ( .A(n11811), .ZN(n11812) );
  XNOR2_X1 U13778 ( .A(n12109), .B(n11679), .ZN(n11814) );
  OR2_X1 U13779 ( .A1(n11942), .A2(n15232), .ZN(n11815) );
  NAND2_X1 U13780 ( .A1(n11814), .A2(n11815), .ZN(n11966) );
  INV_X1 U13781 ( .A(n11814), .ZN(n11817) );
  INV_X1 U13782 ( .A(n11815), .ZN(n11816) );
  NAND2_X1 U13783 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  AND2_X1 U13784 ( .A1(n11966), .A2(n11818), .ZN(n11819) );
  OAI21_X1 U13785 ( .B1(n11820), .B2(n11819), .A(n11967), .ZN(n11821) );
  NAND2_X1 U13786 ( .A1(n11821), .A2(n15070), .ZN(n11826) );
  OR2_X1 U13787 ( .A1(n11969), .A2(n15162), .ZN(n11822) );
  OAI21_X1 U13788 ( .B1(n11832), .B2(n15043), .A(n11822), .ZN(n11837) );
  NOR2_X1 U13789 ( .A1(n15066), .A2(n12109), .ZN(n11823) );
  AOI211_X1 U13790 ( .C1(n15033), .C2(n11837), .A(n11824), .B(n11823), .ZN(
        n11825) );
  OAI211_X1 U13791 ( .C1(n15052), .C2(n12108), .A(n11826), .B(n11825), .ZN(
        P2_U3202) );
  NAND2_X1 U13792 ( .A1(n11832), .A2(n12282), .ZN(n11829) );
  XNOR2_X1 U13793 ( .A(n11936), .B(n8281), .ZN(n12114) );
  NAND2_X1 U13794 ( .A1(n11831), .A2(n11830), .ZN(n11835) );
  NAND2_X1 U13795 ( .A1(n11833), .A2(n11832), .ZN(n11834) );
  NAND2_X1 U13796 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  NAND2_X1 U13797 ( .A1(n11836), .A2(n8281), .ZN(n11940) );
  OAI21_X1 U13798 ( .B1(n11836), .B2(n8281), .A(n11940), .ZN(n11838) );
  AOI21_X1 U13799 ( .B1(n11838), .B2(n15446), .A(n11837), .ZN(n12106) );
  INV_X1 U13800 ( .A(n12109), .ZN(n11938) );
  AOI211_X1 U13801 ( .C1(n11938), .C2(n11839), .A(n7418), .B(n11937), .ZN(
        n12111) );
  AOI21_X1 U13802 ( .B1(n15546), .B2(n11938), .A(n12111), .ZN(n11840) );
  OAI211_X1 U13803 ( .C1(n15550), .C2(n12114), .A(n12106), .B(n11840), .ZN(
        n12194) );
  NAND2_X1 U13804 ( .A1(n12194), .A2(n16526), .ZN(n11841) );
  OAI21_X1 U13805 ( .B1(n16526), .B2(n9916), .A(n11841), .ZN(P2_U3503) );
  INV_X1 U13806 ( .A(n13436), .ZN(n11844) );
  INV_X1 U13807 ( .A(n11842), .ZN(n11845) );
  OAI222_X1 U13808 ( .A1(n11844), .A2(P2_U3088), .B1(n15626), .B2(n11845), 
        .C1(n11843), .C2(n15628), .ZN(P2_U3313) );
  INV_X1 U13809 ( .A(n12695), .ZN(n12688) );
  OAI222_X1 U13810 ( .A1(n16174), .A2(n11846), .B1(n13259), .B2(n11845), .C1(
        P1_U3086), .C2(n12688), .ZN(P1_U3341) );
  MUX2_X1 U13811 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11848), .S(n12534), .Z(
        n11849) );
  OAI21_X1 U13812 ( .B1(n11850), .B2(n11849), .A(n12533), .ZN(n11851) );
  INV_X1 U13813 ( .A(n16264), .ZN(n16230) );
  NAND2_X1 U13814 ( .A1(n11851), .A2(n16230), .ZN(n11862) );
  AOI21_X1 U13815 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n11853), .A(n11852), .ZN(
        n11856) );
  INV_X1 U13816 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11854) );
  MUX2_X1 U13817 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11854), .S(n12534), .Z(
        n11855) );
  NAND2_X1 U13818 ( .A1(n11856), .A2(n11855), .ZN(n12526) );
  OAI21_X1 U13819 ( .B1(n11856), .B2(n11855), .A(n12526), .ZN(n11860) );
  NAND2_X1 U13820 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U13821 ( .A1(n16224), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11857) );
  OAI211_X1 U13822 ( .C1(n15128), .C2(n11858), .A(n12585), .B(n11857), .ZN(
        n11859) );
  AOI21_X1 U13823 ( .B1(n11860), .B2(n16257), .A(n11859), .ZN(n11861) );
  NAND2_X1 U13824 ( .A1(n11862), .A2(n11861), .ZN(P2_U3223) );
  NAND2_X1 U13825 ( .A1(n15191), .A2(P2_U3947), .ZN(n11863) );
  OAI21_X1 U13826 ( .B1(n13750), .B2(P2_U3947), .A(n11863), .ZN(P2_U3555) );
  INV_X1 U13827 ( .A(n16723), .ZN(n13331) );
  INV_X1 U13828 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n12435) );
  NAND2_X1 U13829 ( .A1(n16716), .A2(n12434), .ZN(n11865) );
  OAI211_X1 U13830 ( .C1(n15712), .C2(n13608), .A(n11865), .B(n11864), .ZN(
        n11871) );
  INV_X1 U13831 ( .A(n11866), .ZN(n11867) );
  AOI211_X1 U13832 ( .C1(n11869), .C2(n11868), .A(n15729), .B(n11867), .ZN(
        n11870) );
  AOI211_X1 U13833 ( .C1(n13331), .C2(n12435), .A(n11871), .B(n11870), .ZN(
        n11872) );
  INV_X1 U13834 ( .A(n11872), .ZN(P1_U3218) );
  AOI21_X1 U13835 ( .B1(n11637), .B2(n11874), .A(n11873), .ZN(n15800) );
  MUX2_X1 U13836 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11875), .S(n15804), .Z(
        n15799) );
  NAND2_X1 U13837 ( .A1(n15800), .A2(n15799), .ZN(n15798) );
  NAND2_X1 U13838 ( .A1(n15804), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11877) );
  INV_X1 U13839 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11876) );
  MUX2_X1 U13840 ( .A(n11876), .B(P1_REG2_REG_14__SCAN_IN), .S(n12695), .Z(
        n11878) );
  AOI21_X1 U13841 ( .B1(n15798), .B2(n11877), .A(n11878), .ZN(n12686) );
  INV_X1 U13842 ( .A(n15798), .ZN(n11880) );
  NAND2_X1 U13843 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  OAI21_X1 U13844 ( .B1(n11880), .B2(n11879), .A(n15797), .ZN(n11893) );
  NAND2_X1 U13845 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15641)
         );
  OAI21_X1 U13846 ( .B1(n16301), .B2(n16421), .A(n15641), .ZN(n11881) );
  AOI21_X1 U13847 ( .B1(n12695), .B2(n16294), .A(n11881), .ZN(n11892) );
  XNOR2_X1 U13848 ( .A(n12695), .B(n11882), .ZN(n11889) );
  OR2_X1 U13849 ( .A1(n11883), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U13850 ( .A1(n11885), .A2(n11884), .ZN(n15803) );
  MUX2_X1 U13851 ( .A(n15805), .B(P1_REG1_REG_13__SCAN_IN), .S(n15804), .Z(
        n11886) );
  OR2_X1 U13852 ( .A1(n15803), .A2(n11886), .ZN(n15806) );
  NAND2_X1 U13853 ( .A1(n15804), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11887) );
  AND2_X1 U13854 ( .A1(n15806), .A2(n11887), .ZN(n11888) );
  NAND2_X1 U13855 ( .A1(n11888), .A2(n11889), .ZN(n12697) );
  OAI21_X1 U13856 ( .B1(n11889), .B2(n11888), .A(n12697), .ZN(n11890) );
  NAND2_X1 U13857 ( .A1(n11890), .A2(n15807), .ZN(n11891) );
  OAI211_X1 U13858 ( .C1(n12686), .C2(n11893), .A(n11892), .B(n11891), .ZN(
        P1_U3257) );
  INV_X1 U13859 ( .A(n11894), .ZN(n11895) );
  OAI222_X1 U13860 ( .A1(P3_U3151), .A2(n14590), .B1(n14959), .B2(n11896), 
        .C1(n14968), .C2(n11895), .ZN(P3_U3277) );
  INV_X1 U13861 ( .A(n11897), .ZN(n11902) );
  AOI21_X1 U13862 ( .B1(n11899), .B2(n11901), .A(n11898), .ZN(n11900) );
  AOI21_X1 U13863 ( .B1(n11902), .B2(n11901), .A(n11900), .ZN(n11907) );
  INV_X1 U13864 ( .A(n15716), .ZN(n12073) );
  NAND2_X1 U13865 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15788) );
  OAI21_X1 U13866 ( .B1(n15712), .B2(n16546), .A(n15788), .ZN(n11905) );
  OAI22_X1 U13867 ( .A1(n15717), .A2(n11903), .B1(n16723), .B2(n12449), .ZN(
        n11904) );
  AOI211_X1 U13868 ( .C1(n12073), .C2(n15755), .A(n11905), .B(n11904), .ZN(
        n11906) );
  OAI21_X1 U13869 ( .B1(n11907), .B2(n15729), .A(n11906), .ZN(P1_U3230) );
  OAI22_X1 U13870 ( .A1(n15594), .A2(n14066), .B1(n15586), .B2(n9838), .ZN(
        n11909) );
  INV_X1 U13871 ( .A(n11909), .ZN(n11910) );
  OAI21_X1 U13872 ( .B1(n11911), .B2(n16527), .A(n11910), .ZN(P2_U3433) );
  INV_X1 U13873 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n11913) );
  NAND2_X1 U13874 ( .A1(n14398), .A2(P3_U3897), .ZN(n11912) );
  OAI21_X1 U13875 ( .B1(P3_U3897), .B2(n11913), .A(n11912), .ZN(P3_U3500) );
  INV_X1 U13876 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U13877 ( .A1(n14366), .A2(P3_U3897), .ZN(n11914) );
  OAI21_X1 U13878 ( .B1(P3_U3897), .B2(n11915), .A(n11914), .ZN(P3_U3493) );
  INV_X1 U13879 ( .A(n15458), .ZN(n11917) );
  INV_X1 U13880 ( .A(n12204), .ZN(n11916) );
  NAND2_X1 U13881 ( .A1(n11917), .A2(n11916), .ZN(n11925) );
  NAND2_X1 U13882 ( .A1(n11919), .A2(n11918), .ZN(n12202) );
  AOI21_X1 U13883 ( .B1(n11226), .B2(n15443), .A(n12204), .ZN(n11920) );
  NOR2_X1 U13884 ( .A1(n11921), .A2(n11920), .ZN(n12203) );
  OAI21_X1 U13885 ( .B1(n11922), .B2(n12202), .A(n12203), .ZN(n11923) );
  INV_X1 U13886 ( .A(n15427), .ZN(n15452) );
  AOI22_X1 U13887 ( .A1(n11923), .A2(n15429), .B1(n15452), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n11924) );
  OAI211_X1 U13888 ( .C1(n11525), .C2(n15429), .A(n11925), .B(n11924), .ZN(
        P2_U3265) );
  OAI21_X1 U13889 ( .B1(n11927), .B2(n13858), .A(n11926), .ZN(n12471) );
  AOI21_X1 U13890 ( .B1(n12447), .B2(n13619), .A(n16686), .ZN(n11928) );
  NAND2_X1 U13891 ( .A1(n11928), .A2(n12343), .ZN(n12472) );
  NAND2_X1 U13892 ( .A1(n15752), .A2(n15956), .ZN(n11930) );
  NAND2_X1 U13893 ( .A1(n15754), .A2(n15955), .ZN(n11929) );
  AND2_X1 U13894 ( .A1(n11930), .A2(n11929), .ZN(n12473) );
  OAI211_X1 U13895 ( .C1(n12476), .C2(n16684), .A(n12472), .B(n12473), .ZN(
        n11933) );
  NAND2_X1 U13896 ( .A1(n11931), .A2(n13858), .ZN(n12480) );
  AND3_X1 U13897 ( .A1(n12481), .A2(n16623), .A3(n12480), .ZN(n11932) );
  AOI211_X1 U13898 ( .C1(n16705), .C2(n12471), .A(n11933), .B(n11932), .ZN(
        n12061) );
  NAND2_X1 U13899 ( .A1(n16707), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11934) );
  OAI21_X1 U13900 ( .B1(n12061), .B2(n16707), .A(n11934), .ZN(P1_U3533) );
  XOR2_X1 U13901 ( .A(n11941), .B(n11951), .Z(n12088) );
  OAI211_X1 U13902 ( .C1(n11937), .C2(n11968), .A(n11961), .B(n15232), .ZN(
        n12084) );
  OAI21_X1 U13903 ( .B1(n11968), .B2(n16520), .A(n12084), .ZN(n11947) );
  NAND2_X1 U13904 ( .A1(n11938), .A2(n11942), .ZN(n11939) );
  NAND2_X1 U13905 ( .A1(n11940), .A2(n11939), .ZN(n11955) );
  XOR2_X1 U13906 ( .A(n11955), .B(n11941), .Z(n11946) );
  OR2_X1 U13907 ( .A1(n11942), .A2(n15043), .ZN(n11944) );
  NAND2_X1 U13908 ( .A1(n15093), .A2(n15073), .ZN(n11943) );
  NAND2_X1 U13909 ( .A1(n11944), .A2(n11943), .ZN(n15020) );
  INV_X1 U13910 ( .A(n15020), .ZN(n11945) );
  OAI21_X1 U13911 ( .B1(n11946), .B2(n11226), .A(n11945), .ZN(n12085) );
  AOI211_X1 U13912 ( .C1(n12088), .C2(n16523), .A(n11947), .B(n12085), .ZN(
        n12197) );
  NAND2_X1 U13913 ( .A1(n16525), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11948) );
  OAI21_X1 U13914 ( .B1(n12197), .B2(n16525), .A(n11948), .ZN(P2_U3504) );
  INV_X1 U13915 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11965) );
  INV_X1 U13916 ( .A(n11949), .ZN(n11950) );
  OR2_X1 U13917 ( .A1(n11951), .A2(n11950), .ZN(n11953) );
  XOR2_X1 U13918 ( .A(n12293), .B(n12290), .Z(n12149) );
  NAND2_X1 U13919 ( .A1(n11968), .A2(n15094), .ZN(n11954) );
  NAND2_X1 U13920 ( .A1(n11955), .A2(n11954), .ZN(n11957) );
  NAND2_X1 U13921 ( .A1(n15022), .A2(n11969), .ZN(n11956) );
  NAND2_X1 U13922 ( .A1(n11957), .A2(n11956), .ZN(n12294) );
  XNOR2_X1 U13923 ( .A(n12294), .B(n12293), .ZN(n11960) );
  OR2_X1 U13924 ( .A1(n11969), .A2(n15043), .ZN(n11959) );
  NAND2_X1 U13925 ( .A1(n15092), .A2(n15073), .ZN(n11958) );
  NAND2_X1 U13926 ( .A1(n11959), .A2(n11958), .ZN(n11979) );
  AOI21_X1 U13927 ( .B1(n11960), .B2(n15446), .A(n11979), .ZN(n12141) );
  AOI21_X1 U13928 ( .B1(n11961), .B2(n12296), .A(n7418), .ZN(n11962) );
  NAND2_X1 U13929 ( .A1(n11962), .A2(n12303), .ZN(n12143) );
  OAI211_X1 U13930 ( .C1(n12149), .C2(n15550), .A(n12141), .B(n12143), .ZN(
        n11984) );
  NAND2_X1 U13931 ( .A1(n11984), .A2(n16526), .ZN(n11964) );
  NAND2_X1 U13932 ( .A1(n15536), .A2(n12296), .ZN(n11963) );
  OAI211_X1 U13933 ( .C1(n16526), .C2(n11965), .A(n11964), .B(n11963), .ZN(
        P2_U3505) );
  XNOR2_X1 U13934 ( .A(n12296), .B(n7695), .ZN(n12208) );
  NAND2_X1 U13935 ( .A1(n15093), .A2(n7418), .ZN(n12209) );
  XNOR2_X1 U13936 ( .A(n12208), .B(n12209), .ZN(n12207) );
  NAND2_X1 U13937 ( .A1(n11967), .A2(n11966), .ZN(n15016) );
  XNOR2_X1 U13938 ( .A(n11968), .B(n11679), .ZN(n11970) );
  OR2_X1 U13939 ( .A1(n11969), .A2(n15232), .ZN(n11971) );
  NAND2_X1 U13940 ( .A1(n11970), .A2(n11971), .ZN(n11975) );
  INV_X1 U13941 ( .A(n11970), .ZN(n11973) );
  INV_X1 U13942 ( .A(n11971), .ZN(n11972) );
  NAND2_X1 U13943 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  AND2_X1 U13944 ( .A1(n11975), .A2(n11974), .ZN(n15017) );
  XOR2_X1 U13945 ( .A(n12207), .B(n12206), .Z(n11976) );
  NAND2_X1 U13946 ( .A1(n11976), .A2(n15070), .ZN(n11981) );
  NOR2_X1 U13947 ( .A1(n15066), .A2(n8301), .ZN(n11977) );
  AOI211_X1 U13948 ( .C1(n15033), .C2(n11979), .A(n11978), .B(n11977), .ZN(
        n11980) );
  OAI211_X1 U13949 ( .C1(n15052), .C2(n12144), .A(n11981), .B(n11980), .ZN(
        P2_U3211) );
  INV_X1 U13950 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11982) );
  OAI22_X1 U13951 ( .A1(n15594), .A2(n8301), .B1(n15586), .B2(n11982), .ZN(
        n11983) );
  AOI21_X1 U13952 ( .B1(n11984), .B2(n15586), .A(n11983), .ZN(n11985) );
  INV_X1 U13953 ( .A(n11985), .ZN(P2_U3448) );
  XOR2_X1 U13954 ( .A(n11987), .B(n11986), .Z(n11992) );
  OAI21_X1 U13955 ( .B1(n15712), .B2(n12476), .A(n11988), .ZN(n11990) );
  INV_X1 U13956 ( .A(n15752), .ZN(n12418) );
  OAI22_X1 U13957 ( .A1(n15717), .A2(n12418), .B1(n16723), .B2(n12475), .ZN(
        n11989) );
  AOI211_X1 U13958 ( .C1(n12073), .C2(n15754), .A(n11990), .B(n11989), .ZN(
        n11991) );
  OAI21_X1 U13959 ( .B1(n11992), .B2(n15729), .A(n11991), .ZN(P1_U3227) );
  INV_X1 U13960 ( .A(n11993), .ZN(n11994) );
  INV_X1 U13961 ( .A(n16293), .ZN(n12699) );
  OAI222_X1 U13962 ( .A1(n16174), .A2(n8568), .B1(n13259), .B2(n11994), .C1(
        n12699), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13963 ( .A(n15117), .ZN(n15131) );
  OAI222_X1 U13964 ( .A1(n15628), .A2(n11995), .B1(n15626), .B2(n11994), .C1(
        P2_U3088), .C2(n15131), .ZN(P2_U3312) );
  INV_X1 U13965 ( .A(n14611), .ZN(n14528) );
  NOR3_X1 U13966 ( .A1(n14528), .A2(n14603), .A3(n14604), .ZN(n12005) );
  OR2_X1 U13967 ( .A1(n14574), .A2(n11996), .ZN(n11997) );
  INV_X1 U13968 ( .A(n11998), .ZN(n12000) );
  INV_X1 U13969 ( .A(n14572), .ZN(n14609) );
  AOI22_X1 U13970 ( .A1(n14609), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11999) );
  OAI21_X1 U13971 ( .B1(n14611), .B2(n12000), .A(n11999), .ZN(n12001) );
  AOI21_X1 U13972 ( .B1(n14603), .B2(n12002), .A(n12001), .ZN(n12003) );
  OAI211_X1 U13973 ( .C1(n12005), .C2(n12165), .A(n12004), .B(n12003), .ZN(
        P3_U3182) );
  OAI21_X1 U13974 ( .B1(n12008), .B2(n12007), .A(n12006), .ZN(n12015) );
  OAI22_X1 U13975 ( .A1(n14572), .A2(n16317), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9685), .ZN(n12014) );
  OAI21_X1 U13976 ( .B1(n12011), .B2(n12010), .A(n12009), .ZN(n12012) );
  AND2_X1 U13977 ( .A1(n14603), .A2(n12012), .ZN(n12013) );
  AOI211_X1 U13978 ( .C1(n14528), .C2(n12015), .A(n12014), .B(n12013), .ZN(
        n12020) );
  XNOR2_X1 U13979 ( .A(n12017), .B(n12016), .ZN(n12018) );
  NAND2_X1 U13980 ( .A1(n12018), .A2(n14604), .ZN(n12019) );
  OAI211_X1 U13981 ( .C1(n14606), .C2(n12021), .A(n12020), .B(n12019), .ZN(
        P3_U3184) );
  INV_X1 U13982 ( .A(n12022), .ZN(n12023) );
  OAI222_X1 U13983 ( .A1(n14959), .A2(n12024), .B1(P3_U3151), .B2(n14605), 
        .C1(n14968), .C2(n12023), .ZN(P3_U3276) );
  NAND2_X1 U13984 ( .A1(n14720), .A2(P3_U3897), .ZN(n12025) );
  OAI21_X1 U13985 ( .B1(P3_U3897), .B2(n12026), .A(n12025), .ZN(P3_U3514) );
  NAND2_X1 U13986 ( .A1(n14391), .A2(P3_U3897), .ZN(n12027) );
  OAI21_X1 U13987 ( .B1(P3_U3897), .B2(n12028), .A(n12027), .ZN(P3_U3499) );
  INV_X1 U13988 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U13989 ( .A1(n12933), .A2(P3_U3897), .ZN(n12029) );
  OAI21_X1 U13990 ( .B1(P3_U3897), .B2(n12030), .A(n12029), .ZN(P3_U3496) );
  NAND2_X1 U13991 ( .A1(n14254), .A2(P3_U3897), .ZN(n12031) );
  OAI21_X1 U13992 ( .B1(P3_U3897), .B2(n12032), .A(n12031), .ZN(P3_U3503) );
  INV_X1 U13993 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U13994 ( .A1(n14227), .A2(P3_U3897), .ZN(n12033) );
  OAI21_X1 U13995 ( .B1(P3_U3897), .B2(n12034), .A(n12033), .ZN(P3_U3507) );
  NAND2_X1 U13996 ( .A1(n14133), .A2(P3_U3897), .ZN(n12035) );
  OAI21_X1 U13997 ( .B1(P3_U3897), .B2(n12036), .A(n12035), .ZN(P3_U3502) );
  NAND2_X1 U13998 ( .A1(n14403), .A2(P3_U3897), .ZN(n12037) );
  OAI21_X1 U13999 ( .B1(P3_U3897), .B2(n12038), .A(n12037), .ZN(P3_U3501) );
  NAND2_X1 U14000 ( .A1(n14416), .A2(P3_U3897), .ZN(n12039) );
  OAI21_X1 U14001 ( .B1(P3_U3897), .B2(n12040), .A(n12039), .ZN(P3_U3504) );
  INV_X1 U14002 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n12042) );
  NAND2_X1 U14003 ( .A1(n14267), .A2(P3_U3897), .ZN(n12041) );
  OAI21_X1 U14004 ( .B1(P3_U3897), .B2(n12042), .A(n12041), .ZN(P3_U3513) );
  NAND2_X1 U14005 ( .A1(n12556), .A2(P3_U3897), .ZN(n12043) );
  OAI21_X1 U14006 ( .B1(P3_U3897), .B2(n12044), .A(n12043), .ZN(P3_U3494) );
  INV_X1 U14007 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U14008 ( .A1(n12963), .A2(P3_U3897), .ZN(n12045) );
  OAI21_X1 U14009 ( .B1(P3_U3897), .B2(n12046), .A(n12045), .ZN(P3_U3498) );
  NAND2_X1 U14010 ( .A1(n14187), .A2(P3_U3897), .ZN(n12047) );
  OAI21_X1 U14011 ( .B1(P3_U3897), .B2(n12048), .A(n12047), .ZN(P3_U3511) );
  NAND2_X1 U14012 ( .A1(n14780), .A2(P3_U3897), .ZN(n12049) );
  OAI21_X1 U14013 ( .B1(P3_U3897), .B2(n12050), .A(n12049), .ZN(P3_U3510) );
  NAND2_X1 U14014 ( .A1(n14156), .A2(P3_U3897), .ZN(n12051) );
  OAI21_X1 U14015 ( .B1(P3_U3897), .B2(n12052), .A(n12051), .ZN(P3_U3509) );
  NAND2_X1 U14016 ( .A1(n13557), .A2(P3_U3897), .ZN(n12053) );
  OAI21_X1 U14017 ( .B1(P3_U3897), .B2(n12054), .A(n12053), .ZN(P3_U3505) );
  NAND2_X1 U14018 ( .A1(n14778), .A2(P3_U3897), .ZN(n12055) );
  OAI21_X1 U14019 ( .B1(P3_U3897), .B2(n12056), .A(n12055), .ZN(P3_U3508) );
  NAND2_X1 U14020 ( .A1(n14205), .A2(P3_U3897), .ZN(n12057) );
  OAI21_X1 U14021 ( .B1(P3_U3897), .B2(n12058), .A(n12057), .ZN(P3_U3506) );
  NAND2_X1 U14022 ( .A1(n14719), .A2(P3_U3897), .ZN(n12059) );
  OAI21_X1 U14023 ( .B1(P3_U3897), .B2(n12060), .A(n12059), .ZN(P3_U3512) );
  OR2_X1 U14024 ( .A1(n12061), .A2(n16709), .ZN(n12062) );
  OAI21_X1 U14025 ( .B1(n16694), .B2(n10710), .A(n12062), .ZN(P1_U3474) );
  OAI21_X1 U14026 ( .B1(P3_U3897), .B2(n12064), .A(n12063), .ZN(P3_U3491) );
  INV_X1 U14027 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U14028 ( .A1(n12279), .A2(P3_U3897), .ZN(n12065) );
  OAI21_X1 U14029 ( .B1(P3_U3897), .B2(n12066), .A(n12065), .ZN(P3_U3492) );
  OAI211_X1 U14030 ( .C1(n12069), .C2(n12068), .A(n12067), .B(n16714), .ZN(
        n12075) );
  OAI21_X1 U14031 ( .B1(n15712), .B2(n16555), .A(n12070), .ZN(n12072) );
  OAI22_X1 U14032 ( .A1(n15717), .A2(n12575), .B1(n16723), .B2(n12344), .ZN(
        n12071) );
  AOI211_X1 U14033 ( .C1(n12073), .C2(n15753), .A(n12072), .B(n12071), .ZN(
        n12074) );
  NAND2_X1 U14034 ( .A1(n12075), .A2(n12074), .ZN(P1_U3239) );
  INV_X1 U14035 ( .A(n14872), .ZN(n16730) );
  AND2_X1 U14036 ( .A1(n12708), .A2(n14355), .ZN(n14472) );
  NAND2_X1 U14037 ( .A1(n12123), .A2(n16663), .ZN(n12076) );
  OAI22_X1 U14038 ( .A1(n14472), .A2(n12076), .B1(n16496), .B2(n16497), .ZN(
        n12671) );
  MUX2_X1 U14039 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n12671), .S(n16724), .Z(
        n12077) );
  AOI21_X1 U14040 ( .B1(n16730), .B2(n12078), .A(n12077), .ZN(n12079) );
  INV_X1 U14041 ( .A(n12079), .ZN(P3_U3459) );
  NAND2_X1 U14042 ( .A1(n15443), .A2(n12080), .ZN(n12081) );
  INV_X1 U14043 ( .A(n15435), .ZN(n15336) );
  INV_X1 U14044 ( .A(n12082), .ZN(n15021) );
  AOI22_X1 U14045 ( .A1(n15316), .A2(n15022), .B1(n15021), .B2(n15452), .ZN(
        n12083) );
  OAI21_X1 U14046 ( .B1(n15318), .B2(n12084), .A(n12083), .ZN(n12087) );
  MUX2_X1 U14047 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n12085), .S(n15429), .Z(
        n12086) );
  AOI211_X1 U14048 ( .C1(n12088), .C2(n15336), .A(n12087), .B(n12086), .ZN(
        n12089) );
  INV_X1 U14049 ( .A(n12089), .ZN(P2_U3260) );
  OAI21_X1 U14050 ( .B1(n12092), .B2(n12091), .A(n12090), .ZN(n12094) );
  AOI21_X1 U14051 ( .B1(n12094), .B2(n15446), .A(n12093), .ZN(n16519) );
  OAI22_X1 U14052 ( .A1(n15429), .A2(n12096), .B1(n12095), .B2(n15427), .ZN(
        n12100) );
  OAI211_X1 U14053 ( .C1(n16521), .C2(n12098), .A(n12097), .B(n15232), .ZN(
        n16518) );
  NOR2_X1 U14054 ( .A1(n15318), .A2(n16518), .ZN(n12099) );
  AOI211_X1 U14055 ( .C1(n15316), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        n12105) );
  XNOR2_X1 U14056 ( .A(n12103), .B(n12102), .ZN(n16524) );
  NAND2_X1 U14057 ( .A1(n16524), .A2(n15336), .ZN(n12104) );
  OAI211_X1 U14058 ( .C1(n15454), .C2(n16519), .A(n12105), .B(n12104), .ZN(
        P2_U3263) );
  MUX2_X1 U14059 ( .A(n12107), .B(n12106), .S(n15429), .Z(n12113) );
  OAI22_X1 U14060 ( .A1(n15456), .A2(n12109), .B1(n15427), .B2(n12108), .ZN(
        n12110) );
  AOI21_X1 U14061 ( .B1(n15461), .B2(n12111), .A(n12110), .ZN(n12112) );
  OAI211_X1 U14062 ( .C1(n15435), .C2(n12114), .A(n12113), .B(n12112), .ZN(
        P2_U3261) );
  INV_X1 U14063 ( .A(n12129), .ZN(n12115) );
  NAND2_X1 U14064 ( .A1(n12131), .A2(n12115), .ZN(n12119) );
  AND3_X1 U14065 ( .A1(n12664), .A2(n12117), .A3(n12116), .ZN(n12118) );
  OAI211_X1 U14066 ( .C1(n12134), .C2(n12120), .A(n12119), .B(n12118), .ZN(
        n12121) );
  NAND2_X1 U14067 ( .A1(n12121), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12126) );
  INV_X1 U14068 ( .A(n12135), .ZN(n12122) );
  OR2_X1 U14069 ( .A1(n12123), .A2(n12122), .ZN(n14511) );
  INV_X1 U14070 ( .A(n14511), .ZN(n12124) );
  NAND2_X1 U14071 ( .A1(n12131), .A2(n12124), .ZN(n12125) );
  NOR2_X1 U14072 ( .A1(n14287), .A2(P3_U3151), .ZN(n12353) );
  NAND3_X1 U14073 ( .A1(n12134), .A2(n12127), .A3(n16663), .ZN(n12128) );
  OAI21_X1 U14074 ( .B1(n12131), .B2(n12129), .A(n12128), .ZN(n12130) );
  INV_X1 U14075 ( .A(n14472), .ZN(n12139) );
  OR2_X1 U14076 ( .A1(n12131), .A2(n14511), .ZN(n12277) );
  INV_X1 U14077 ( .A(n12277), .ZN(n12132) );
  AND2_X1 U14078 ( .A1(n16672), .A2(n12135), .ZN(n12133) );
  NAND2_X1 U14079 ( .A1(n12134), .A2(n12133), .ZN(n12137) );
  OAI22_X1 U14080 ( .A1(n14290), .A2(n16496), .B1(n14282), .B2(n12674), .ZN(
        n12138) );
  AOI21_X1 U14081 ( .B1(n14273), .B2(n12139), .A(n12138), .ZN(n12140) );
  OAI21_X1 U14082 ( .B1(n12353), .B2(n9678), .A(n12140), .ZN(P3_U3172) );
  MUX2_X1 U14083 ( .A(n12142), .B(n12141), .S(n15429), .Z(n12148) );
  INV_X1 U14084 ( .A(n12143), .ZN(n12146) );
  OAI22_X1 U14085 ( .A1(n15456), .A2(n8301), .B1(n15427), .B2(n12144), .ZN(
        n12145) );
  AOI21_X1 U14086 ( .B1(n15461), .B2(n12146), .A(n12145), .ZN(n12147) );
  OAI211_X1 U14087 ( .C1(n12149), .C2(n15435), .A(n12148), .B(n12147), .ZN(
        P2_U3259) );
  NAND2_X1 U14088 ( .A1(n15219), .A2(P2_U3947), .ZN(n12150) );
  OAI21_X1 U14089 ( .B1(n8126), .B2(P2_U3947), .A(n12150), .ZN(P2_U3557) );
  XOR2_X1 U14090 ( .A(n12152), .B(n12151), .Z(n12163) );
  INV_X1 U14091 ( .A(n12153), .ZN(n12400) );
  AOI21_X1 U14092 ( .B1(n16534), .B2(n12154), .A(n12400), .ZN(n12156) );
  NOR2_X1 U14093 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14146), .ZN(n14144) );
  AOI21_X1 U14094 ( .B1(n14609), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n14144), .ZN(
        n12155) );
  OAI21_X1 U14095 ( .B1(n12156), .B2(n14611), .A(n12155), .ZN(n12160) );
  NAND2_X1 U14096 ( .A1(n12157), .A2(n8955), .ZN(n12158) );
  AOI21_X1 U14097 ( .B1(n12407), .B2(n12158), .A(n14541), .ZN(n12159) );
  AOI211_X1 U14098 ( .C1(n14580), .C2(n12161), .A(n12160), .B(n12159), .ZN(
        n12162) );
  OAI21_X1 U14099 ( .B1(n12163), .B2(n14574), .A(n12162), .ZN(P3_U3185) );
  XOR2_X1 U14100 ( .A(n12165), .B(n12164), .Z(n12179) );
  INV_X1 U14101 ( .A(n12166), .ZN(n12177) );
  INV_X1 U14102 ( .A(n12167), .ZN(n12168) );
  AOI21_X1 U14103 ( .B1(n16485), .B2(n12169), .A(n12168), .ZN(n12171) );
  AOI22_X1 U14104 ( .A1(n14609), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n12170) );
  OAI21_X1 U14105 ( .B1(n12171), .B2(n14611), .A(n12170), .ZN(n12176) );
  NAND2_X1 U14106 ( .A1(n12172), .A2(n8925), .ZN(n12173) );
  AOI21_X1 U14107 ( .B1(n12174), .B2(n12173), .A(n14541), .ZN(n12175) );
  AOI211_X1 U14108 ( .C1(n14580), .C2(n12177), .A(n12176), .B(n12175), .ZN(
        n12178) );
  OAI21_X1 U14109 ( .B1(n14574), .B2(n12179), .A(n12178), .ZN(P3_U3183) );
  XOR2_X1 U14110 ( .A(n12180), .B(n12181), .Z(n12191) );
  AOI21_X1 U14111 ( .B1(n12600), .B2(n12182), .A(n7638), .ZN(n12184) );
  NOR2_X1 U14112 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8984), .ZN(n14214) );
  AOI21_X1 U14113 ( .B1(n14609), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n14214), .ZN(
        n12183) );
  OAI21_X1 U14114 ( .B1(n12184), .B2(n14611), .A(n12183), .ZN(n12188) );
  NAND2_X1 U14115 ( .A1(n12185), .A2(n8986), .ZN(n12186) );
  AOI21_X1 U14116 ( .B1(n12386), .B2(n12186), .A(n14541), .ZN(n12187) );
  AOI211_X1 U14117 ( .C1(n14580), .C2(n12189), .A(n12188), .B(n12187), .ZN(
        n12190) );
  OAI21_X1 U14118 ( .B1(n12191), .B2(n14574), .A(n12190), .ZN(P3_U3187) );
  NAND2_X1 U14119 ( .A1(n14325), .A2(P3_U3897), .ZN(n12192) );
  OAI21_X1 U14120 ( .B1(P3_U3897), .B2(n12193), .A(n12192), .ZN(P3_U3516) );
  INV_X1 U14121 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U14122 ( .A1(n12194), .A2(n15586), .ZN(n12195) );
  OAI21_X1 U14123 ( .B1(n16529), .B2(n12196), .A(n12195), .ZN(P2_U3442) );
  INV_X1 U14124 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n12199) );
  OR2_X1 U14125 ( .A1(n12197), .A2(n16527), .ZN(n12198) );
  OAI21_X1 U14126 ( .B1(n16529), .B2(n12199), .A(n12198), .ZN(P2_U3445) );
  NAND2_X1 U14127 ( .A1(n12200), .A2(n15586), .ZN(n12201) );
  OAI21_X1 U14128 ( .B1(n16529), .B2(n9889), .A(n12201), .ZN(P2_U3439) );
  OAI211_X1 U14129 ( .C1(n12204), .C2(n15543), .A(n12203), .B(n12202), .ZN(
        n15551) );
  NAND2_X1 U14130 ( .A1(n15586), .A2(n15551), .ZN(n12205) );
  OAI21_X1 U14131 ( .B1(n16529), .B2(n9852), .A(n12205), .ZN(P2_U3430) );
  INV_X1 U14132 ( .A(n12208), .ZN(n12211) );
  INV_X1 U14133 ( .A(n12209), .ZN(n12210) );
  XNOR2_X1 U14134 ( .A(n12488), .B(n7695), .ZN(n12212) );
  NAND2_X1 U14135 ( .A1(n15092), .A2(n7418), .ZN(n12213) );
  NAND2_X1 U14136 ( .A1(n12212), .A2(n12213), .ZN(n12324) );
  INV_X1 U14137 ( .A(n12212), .ZN(n12215) );
  INV_X1 U14138 ( .A(n12213), .ZN(n12214) );
  NAND2_X1 U14139 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  AND2_X1 U14140 ( .A1(n12324), .A2(n12216), .ZN(n12217) );
  NAND2_X1 U14141 ( .A1(n12218), .A2(n12217), .ZN(n12325) );
  OAI21_X1 U14142 ( .B1(n12218), .B2(n12217), .A(n12325), .ZN(n12219) );
  NAND2_X1 U14143 ( .A1(n12219), .A2(n15070), .ZN(n12225) );
  OR2_X1 U14144 ( .A1(n12611), .A2(n15162), .ZN(n12221) );
  NAND2_X1 U14145 ( .A1(n15093), .A2(n15225), .ZN(n12220) );
  AND2_X1 U14146 ( .A1(n12221), .A2(n12220), .ZN(n12301) );
  OAI21_X1 U14147 ( .B1(n15076), .B2(n12301), .A(n12222), .ZN(n12223) );
  AOI21_X1 U14148 ( .B1(n12488), .B2(n15080), .A(n12223), .ZN(n12224) );
  OAI211_X1 U14149 ( .C1(n15052), .C2(n12304), .A(n12225), .B(n12224), .ZN(
        P2_U3185) );
  XOR2_X1 U14150 ( .A(n12227), .B(n12226), .Z(n12246) );
  OR2_X1 U14151 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12228), .ZN(n12908) );
  OAI21_X1 U14152 ( .B1(n14572), .B2(n16366), .A(n12908), .ZN(n12235) );
  INV_X1 U14153 ( .A(n12229), .ZN(n12231) );
  NAND3_X1 U14154 ( .A1(n12252), .A2(n12231), .A3(n12230), .ZN(n12232) );
  AOI21_X1 U14155 ( .B1(n12233), .B2(n12232), .A(n14611), .ZN(n12234) );
  AOI211_X1 U14156 ( .C1(n14580), .C2(n12236), .A(n12235), .B(n12234), .ZN(
        n12245) );
  INV_X1 U14157 ( .A(n12237), .ZN(n12250) );
  INV_X1 U14158 ( .A(n12238), .ZN(n12239) );
  NOR3_X1 U14159 ( .A1(n12250), .A2(n12240), .A3(n12239), .ZN(n12243) );
  INV_X1 U14160 ( .A(n12241), .ZN(n12242) );
  OAI21_X1 U14161 ( .B1(n12243), .B2(n12242), .A(n14603), .ZN(n12244) );
  OAI211_X1 U14162 ( .C1(n12246), .C2(n14574), .A(n12245), .B(n12244), .ZN(
        P3_U3190) );
  XOR2_X1 U14163 ( .A(n12248), .B(n12247), .Z(n12261) );
  OR2_X1 U14164 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12249), .ZN(n12801) );
  OAI21_X1 U14165 ( .B1(n14572), .B2(n9559), .A(n12801), .ZN(n12258) );
  AOI21_X1 U14166 ( .B1(n9018), .B2(n12251), .A(n12250), .ZN(n12256) );
  INV_X1 U14167 ( .A(n12252), .ZN(n12253) );
  AOI21_X1 U14168 ( .B1(n16566), .B2(n12254), .A(n12253), .ZN(n12255) );
  OAI22_X1 U14169 ( .A1(n14541), .A2(n12256), .B1(n12255), .B2(n14611), .ZN(
        n12257) );
  AOI211_X1 U14170 ( .C1(n12259), .C2(n14580), .A(n12258), .B(n12257), .ZN(
        n12260) );
  OAI21_X1 U14171 ( .B1(n12261), .B2(n14574), .A(n12260), .ZN(P3_U3189) );
  NAND2_X1 U14172 ( .A1(n14673), .A2(P3_U3897), .ZN(n12262) );
  OAI21_X1 U14173 ( .B1(P3_U3897), .B2(n12263), .A(n12262), .ZN(P3_U3515) );
  OAI21_X1 U14174 ( .B1(n14357), .B2(n14605), .A(n12468), .ZN(n12264) );
  OAI21_X2 U14175 ( .B1(n12266), .B2(n12265), .A(n12264), .ZN(n12268) );
  XNOR2_X1 U14176 ( .A(n12268), .B(n12267), .ZN(n12545) );
  XNOR2_X1 U14177 ( .A(n12545), .B(n14366), .ZN(n12274) );
  XNOR2_X1 U14178 ( .A(n12268), .B(n12709), .ZN(n12269) );
  NAND2_X1 U14179 ( .A1(n12269), .A2(n16496), .ZN(n12272) );
  NAND2_X1 U14180 ( .A1(n12272), .A2(n12270), .ZN(n12350) );
  NAND2_X1 U14181 ( .A1(n12268), .A2(n12674), .ZN(n12271) );
  NAND2_X1 U14182 ( .A1(n12711), .A2(n12271), .ZN(n12351) );
  OAI21_X1 U14183 ( .B1(n12274), .B2(n12273), .A(n14140), .ZN(n12275) );
  NAND2_X1 U14184 ( .A1(n12275), .A2(n14273), .ZN(n12281) );
  OR2_X1 U14185 ( .A1(n12277), .A2(n12276), .ZN(n14167) );
  OAI22_X1 U14186 ( .A1(n14290), .A2(n16498), .B1(n14282), .B2(n16491), .ZN(
        n12278) );
  AOI21_X1 U14187 ( .B1(n7422), .B2(n12279), .A(n12278), .ZN(n12280) );
  OAI211_X1 U14188 ( .C1(n12353), .C2(n9685), .A(n12281), .B(n12280), .ZN(
        P3_U3177) );
  OAI22_X1 U14189 ( .A1(n15429), .A2(n11470), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15427), .ZN(n12284) );
  NOR2_X1 U14190 ( .A1(n15456), .A2(n12282), .ZN(n12283) );
  AOI211_X1 U14191 ( .C1(n12285), .C2(n15461), .A(n12284), .B(n12283), .ZN(
        n12288) );
  OR2_X1 U14192 ( .A1(n12286), .A2(n15435), .ZN(n12287) );
  OAI211_X1 U14193 ( .C1(n15454), .C2(n12289), .A(n12288), .B(n12287), .ZN(
        P2_U3262) );
  NAND2_X1 U14194 ( .A1(n12291), .A2(n12298), .ZN(n12292) );
  NAND2_X1 U14195 ( .A1(n12486), .A2(n12292), .ZN(n12308) );
  NAND2_X1 U14196 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  XNOR2_X1 U14197 ( .A(n12490), .B(n12298), .ZN(n12299) );
  NAND2_X1 U14198 ( .A1(n12299), .A2(n15446), .ZN(n12300) );
  OAI211_X1 U14199 ( .C1(n12308), .C2(n15443), .A(n12301), .B(n12300), .ZN(
        n12309) );
  MUX2_X1 U14200 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n12309), .S(n15429), .Z(
        n12302) );
  INV_X1 U14201 ( .A(n12302), .ZN(n12307) );
  AOI211_X1 U14202 ( .C1(n12488), .C2(n12303), .A(n7418), .B(n12495), .ZN(
        n12310) );
  OAI22_X1 U14203 ( .A1(n15456), .A2(n12314), .B1(n12304), .B2(n15427), .ZN(
        n12305) );
  AOI21_X1 U14204 ( .B1(n12310), .B2(n15461), .A(n12305), .ZN(n12306) );
  OAI211_X1 U14205 ( .C1(n12308), .C2(n15458), .A(n12307), .B(n12306), .ZN(
        P2_U3258) );
  INV_X1 U14206 ( .A(n12308), .ZN(n12311) );
  AOI211_X1 U14207 ( .C1(n12311), .C2(n11714), .A(n12310), .B(n12309), .ZN(
        n12317) );
  AOI22_X1 U14208 ( .A1(n15536), .A2(n12488), .B1(n16525), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n12312) );
  OAI21_X1 U14209 ( .B1(n12317), .B2(n16525), .A(n12312), .ZN(P2_U3506) );
  INV_X1 U14210 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n12313) );
  OAI22_X1 U14211 ( .A1(n15594), .A2(n12314), .B1(n15586), .B2(n12313), .ZN(
        n12315) );
  INV_X1 U14212 ( .A(n12315), .ZN(n12316) );
  OAI21_X1 U14213 ( .B1(n12317), .B2(n16527), .A(n12316), .ZN(P2_U3451) );
  INV_X1 U14214 ( .A(n12859), .ZN(n12866) );
  OAI222_X1 U14215 ( .A1(P1_U3086), .A2(n12866), .B1(n13259), .B2(n12320), 
        .C1(n12318), .C2(n16174), .ZN(P1_U3339) );
  INV_X1 U14216 ( .A(n16243), .ZN(n15120) );
  INV_X1 U14217 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n12319) );
  OAI222_X1 U14218 ( .A1(P2_U3088), .A2(n15120), .B1(n15626), .B2(n12320), 
        .C1(n12319), .C2(n15628), .ZN(P2_U3311) );
  INV_X1 U14219 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12321) );
  NOR2_X1 U14220 ( .A1(n16727), .A2(n12321), .ZN(n12322) );
  AOI21_X1 U14221 ( .B1(n12671), .B2(n16727), .A(n12322), .ZN(n12323) );
  OAI21_X1 U14222 ( .B1(n12674), .B2(n14938), .A(n12323), .ZN(P3_U3390) );
  XNOR2_X1 U14223 ( .A(n12615), .B(n11679), .ZN(n12581) );
  OR2_X1 U14224 ( .A1(n12611), .A2(n15232), .ZN(n12580) );
  XNOR2_X1 U14225 ( .A(n12581), .B(n12580), .ZN(n12326) );
  XNOR2_X1 U14226 ( .A(n12582), .B(n12326), .ZN(n12334) );
  OR2_X1 U14227 ( .A1(n12621), .A2(n15162), .ZN(n12328) );
  NAND2_X1 U14228 ( .A1(n15092), .A2(n15225), .ZN(n12327) );
  AND2_X1 U14229 ( .A1(n12328), .A2(n12327), .ZN(n12491) );
  INV_X1 U14230 ( .A(n12497), .ZN(n12329) );
  NAND2_X1 U14231 ( .A1(n15074), .A2(n12329), .ZN(n12331) );
  OAI211_X1 U14232 ( .C1(n12491), .C2(n15076), .A(n12331), .B(n12330), .ZN(
        n12332) );
  AOI21_X1 U14233 ( .B1(n12521), .B2(n15080), .A(n12332), .ZN(n12333) );
  OAI21_X1 U14234 ( .B1(n12334), .B2(n15077), .A(n12333), .ZN(P2_U3193) );
  XNOR2_X1 U14235 ( .A(n12335), .B(n13860), .ZN(n16553) );
  AOI22_X1 U14236 ( .A1(n15956), .A2(n15751), .B1(n15753), .B2(n15955), .ZN(
        n12339) );
  OAI211_X1 U14237 ( .C1(n12337), .C2(n13860), .A(n12336), .B(n16623), .ZN(
        n12338) );
  OAI211_X1 U14238 ( .C1(n16553), .C2(n16619), .A(n12339), .B(n12338), .ZN(
        n16557) );
  INV_X1 U14239 ( .A(n16557), .ZN(n12340) );
  MUX2_X1 U14240 ( .A(n12341), .B(n12340), .S(n16014), .Z(n12347) );
  INV_X1 U14241 ( .A(n12342), .ZN(n16573) );
  AOI21_X1 U14242 ( .B1(n13628), .B2(n12343), .A(n16573), .ZN(n16554) );
  NOR2_X1 U14243 ( .A1(n15825), .A2(n16686), .ZN(n15987) );
  OAI22_X1 U14244 ( .A1(n16587), .A2(n16555), .B1(n12344), .B2(n16036), .ZN(
        n12345) );
  AOI21_X1 U14245 ( .B1(n16554), .B2(n15987), .A(n12345), .ZN(n12346) );
  OAI211_X1 U14246 ( .C1(n16553), .C2(n16006), .A(n12347), .B(n12346), .ZN(
        P1_U3287) );
  INV_X1 U14247 ( .A(n12348), .ZN(n12349) );
  AOI21_X1 U14248 ( .B1(n12351), .B2(n12350), .A(n12349), .ZN(n12357) );
  OAI22_X1 U14249 ( .A1(n14290), .A2(n12544), .B1(n14282), .B2(n12352), .ZN(
        n12355) );
  INV_X1 U14250 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n12717) );
  NOR2_X1 U14251 ( .A1(n12353), .A2(n12717), .ZN(n12354) );
  OAI21_X1 U14252 ( .B1(n12357), .B2(n14295), .A(n12356), .ZN(P3_U3162) );
  AOI21_X1 U14253 ( .B1(n12359), .B2(n9050), .A(n12358), .ZN(n12371) );
  XNOR2_X1 U14254 ( .A(n12361), .B(n12360), .ZN(n12362) );
  NAND2_X1 U14255 ( .A1(n12362), .A2(n14604), .ZN(n12370) );
  OR2_X1 U14256 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9047), .ZN(n13094) );
  OAI21_X1 U14257 ( .B1(n14572), .B2(n16376), .A(n13094), .ZN(n12367) );
  AOI21_X1 U14258 ( .B1(n12364), .B2(n13226), .A(n12363), .ZN(n12365) );
  NOR2_X1 U14259 ( .A1(n12365), .A2(n14611), .ZN(n12366) );
  AOI211_X1 U14260 ( .C1(n14580), .C2(n12368), .A(n12367), .B(n12366), .ZN(
        n12369) );
  OAI211_X1 U14261 ( .C1(n12371), .C2(n14541), .A(n12370), .B(n12369), .ZN(
        P3_U3191) );
  XOR2_X1 U14262 ( .A(n12373), .B(n12372), .Z(n12393) );
  INV_X1 U14263 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n12382) );
  INV_X1 U14264 ( .A(n12374), .ZN(n12379) );
  INV_X1 U14265 ( .A(n12375), .ZN(n12376) );
  NOR3_X1 U14266 ( .A1(n7638), .A2(n12377), .A3(n12376), .ZN(n12378) );
  OAI21_X1 U14267 ( .B1(n12379), .B2(n12378), .A(n14528), .ZN(n12381) );
  OR2_X1 U14268 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12380), .ZN(n12934) );
  OAI211_X1 U14269 ( .C1(n14572), .C2(n12382), .A(n12381), .B(n12934), .ZN(
        n12390) );
  INV_X1 U14270 ( .A(n12383), .ZN(n12385) );
  NAND3_X1 U14271 ( .A1(n12386), .A2(n12385), .A3(n12384), .ZN(n12387) );
  AOI21_X1 U14272 ( .B1(n12388), .B2(n12387), .A(n14541), .ZN(n12389) );
  AOI211_X1 U14273 ( .C1(n14580), .C2(n12391), .A(n12390), .B(n12389), .ZN(
        n12392) );
  OAI21_X1 U14274 ( .B1(n12393), .B2(n14574), .A(n12392), .ZN(P3_U3188) );
  XOR2_X1 U14275 ( .A(n12394), .B(n12395), .Z(n12414) );
  INV_X1 U14276 ( .A(n12396), .ZN(n12402) );
  INV_X1 U14277 ( .A(n12397), .ZN(n12398) );
  NOR3_X1 U14278 ( .A1(n12400), .A2(n12399), .A3(n12398), .ZN(n12401) );
  OAI21_X1 U14279 ( .B1(n12402), .B2(n12401), .A(n14528), .ZN(n12403) );
  NAND2_X1 U14280 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n12557) );
  OAI211_X1 U14281 ( .C1(n14572), .C2(n16335), .A(n12403), .B(n12557), .ZN(
        n12411) );
  INV_X1 U14282 ( .A(n12404), .ZN(n12406) );
  NAND3_X1 U14283 ( .A1(n12407), .A2(n12406), .A3(n12405), .ZN(n12408) );
  AOI21_X1 U14284 ( .B1(n12409), .B2(n12408), .A(n14541), .ZN(n12410) );
  AOI211_X1 U14285 ( .C1(n14580), .C2(n12412), .A(n12411), .B(n12410), .ZN(
        n12413) );
  OAI21_X1 U14286 ( .B1(n12414), .B2(n14574), .A(n12413), .ZN(P3_U3186) );
  INV_X1 U14287 ( .A(n13633), .ZN(n16586) );
  OAI211_X1 U14288 ( .C1(n12417), .C2(n12416), .A(n12415), .B(n16714), .ZN(
        n12422) );
  OAI22_X1 U14289 ( .A1(n12896), .A2(n16029), .B1(n12418), .B2(n16031), .ZN(
        n16578) );
  NOR2_X1 U14290 ( .A1(n16723), .A2(n16583), .ZN(n12419) );
  AOI211_X1 U14291 ( .C1(n16716), .C2(n16578), .A(n12420), .B(n12419), .ZN(
        n12421) );
  OAI211_X1 U14292 ( .C1(n16586), .C2(n15712), .A(n12422), .B(n12421), .ZN(
        P1_U3213) );
  AND2_X1 U14293 ( .A1(n16642), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n12426) );
  OAI22_X1 U14294 ( .A1(n15825), .A2(n12424), .B1(n12423), .B2(n16036), .ZN(
        n12425) );
  AOI211_X1 U14295 ( .C1(n12427), .C2(n16014), .A(n12426), .B(n12425), .ZN(
        n12430) );
  INV_X1 U14296 ( .A(n16006), .ZN(n16637) );
  AOI22_X1 U14297 ( .A1(n12428), .A2(n16637), .B1(n16632), .B2(n13599), .ZN(
        n12429) );
  NAND2_X1 U14298 ( .A1(n12430), .A2(n12429), .ZN(P1_U3292) );
  INV_X1 U14299 ( .A(n12431), .ZN(n12432) );
  NOR2_X1 U14300 ( .A1(n16587), .A2(n13608), .ZN(n12442) );
  NAND2_X1 U14301 ( .A1(n12433), .A2(n16033), .ZN(n12438) );
  INV_X1 U14302 ( .A(n12434), .ZN(n12437) );
  NAND2_X1 U14303 ( .A1(n16631), .A2(n12435), .ZN(n12436) );
  NAND3_X1 U14304 ( .A1(n12438), .A2(n12437), .A3(n12436), .ZN(n12439) );
  NAND2_X1 U14305 ( .A1(n12439), .A2(n16014), .ZN(n12440) );
  OAI21_X1 U14306 ( .B1(n10689), .B2(n16014), .A(n12440), .ZN(n12441) );
  AOI211_X1 U14307 ( .C1(n15929), .C2(n12443), .A(n12442), .B(n12441), .ZN(
        n12444) );
  OAI21_X1 U14308 ( .B1(n12445), .B2(n15970), .A(n12444), .ZN(P1_U3290) );
  XNOR2_X1 U14309 ( .A(n12446), .B(n13857), .ZN(n16547) );
  OAI211_X1 U14310 ( .C1(n12448), .C2(n16546), .A(n12447), .B(n16698), .ZN(
        n16545) );
  OAI22_X1 U14311 ( .A1(n16545), .A2(n15825), .B1(n12449), .B2(n16036), .ZN(
        n12452) );
  AOI22_X1 U14312 ( .A1(n15956), .A2(n15753), .B1(n15755), .B2(n15955), .ZN(
        n16544) );
  INV_X1 U14313 ( .A(n16544), .ZN(n12450) );
  MUX2_X1 U14314 ( .A(n12450), .B(P1_REG2_REG_4__SCAN_IN), .S(n16642), .Z(
        n12451) );
  AOI211_X1 U14315 ( .C1(n16632), .C2(n13611), .A(n12452), .B(n12451), .ZN(
        n12456) );
  OAI21_X1 U14316 ( .B1(n12454), .B2(n13857), .A(n12453), .ZN(n16550) );
  NAND2_X1 U14317 ( .A1(n16550), .A2(n15929), .ZN(n12455) );
  OAI211_X1 U14318 ( .C1(n16547), .C2(n15970), .A(n12456), .B(n12455), .ZN(
        P1_U3289) );
  INV_X1 U14319 ( .A(n12457), .ZN(n12459) );
  OAI22_X1 U14320 ( .A1(n15825), .A2(n12459), .B1(n12458), .B2(n16036), .ZN(
        n12462) );
  OAI22_X1 U14321 ( .A1(n12460), .A2(n16006), .B1(n13580), .B2(n16587), .ZN(
        n12461) );
  AOI211_X1 U14322 ( .C1(P1_REG2_REG_2__SCAN_IN), .C2(n16642), .A(n12462), .B(
        n12461), .ZN(n12463) );
  OAI21_X1 U14323 ( .B1(n16642), .B2(n12464), .A(n12463), .ZN(P1_U3291) );
  INV_X1 U14324 ( .A(n12465), .ZN(n12467) );
  OAI222_X1 U14325 ( .A1(P3_U3151), .A2(n12468), .B1(n14968), .B2(n12467), 
        .C1(n12466), .C2(n14959), .ZN(P3_U3275) );
  NAND2_X1 U14326 ( .A1(n14674), .A2(P3_U3897), .ZN(n12469) );
  OAI21_X1 U14327 ( .B1(P3_U3897), .B2(n12470), .A(n12469), .ZN(P3_U3517) );
  INV_X1 U14328 ( .A(n12471), .ZN(n12484) );
  AOI21_X1 U14329 ( .B1(n16579), .B2(n16014), .A(n16637), .ZN(n15897) );
  INV_X1 U14330 ( .A(n12472), .ZN(n12479) );
  INV_X1 U14331 ( .A(n12473), .ZN(n12474) );
  MUX2_X1 U14332 ( .A(n12474), .B(P1_REG2_REG_5__SCAN_IN), .S(n16642), .Z(
        n12478) );
  OAI22_X1 U14333 ( .A1(n16587), .A2(n12476), .B1(n16036), .B2(n12475), .ZN(
        n12477) );
  AOI211_X1 U14334 ( .C1(n12479), .C2(n16636), .A(n12478), .B(n12477), .ZN(
        n12483) );
  NAND3_X1 U14335 ( .A1(n12481), .A2(n12480), .A3(n15948), .ZN(n12482) );
  OAI211_X1 U14336 ( .C1(n12484), .C2(n15897), .A(n12483), .B(n12482), .ZN(
        P1_U3288) );
  NAND2_X1 U14337 ( .A1(n12488), .A2(n15092), .ZN(n12485) );
  XNOR2_X1 U14338 ( .A(n12610), .B(n12608), .ZN(n12520) );
  INV_X1 U14339 ( .A(n12520), .ZN(n12501) );
  AND2_X1 U14340 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  XNOR2_X1 U14341 ( .A(n12617), .B(n12608), .ZN(n12492) );
  OAI21_X1 U14342 ( .B1(n12492), .B2(n11226), .A(n12491), .ZN(n12518) );
  INV_X1 U14343 ( .A(n12518), .ZN(n12493) );
  MUX2_X1 U14344 ( .A(n12494), .B(n12493), .S(n15429), .Z(n12500) );
  OAI21_X1 U14345 ( .B1(n12495), .B2(n12615), .A(n15232), .ZN(n12496) );
  NOR2_X1 U14346 ( .A1(n12496), .A2(n12641), .ZN(n12519) );
  OAI22_X1 U14347 ( .A1(n12615), .A2(n15456), .B1(n15427), .B2(n12497), .ZN(
        n12498) );
  AOI21_X1 U14348 ( .B1(n12519), .B2(n15461), .A(n12498), .ZN(n12499) );
  OAI211_X1 U14349 ( .C1(n12501), .C2(n15435), .A(n12500), .B(n12499), .ZN(
        P2_U3257) );
  XOR2_X1 U14350 ( .A(n12503), .B(n12502), .Z(n12517) );
  AOI21_X1 U14351 ( .B1(n12506), .B2(n12505), .A(n12504), .ZN(n12509) );
  NOR2_X1 U14352 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12507), .ZN(n14132) );
  AOI21_X1 U14353 ( .B1(n14609), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n14132), 
        .ZN(n12508) );
  OAI21_X1 U14354 ( .B1(n14541), .B2(n12509), .A(n12508), .ZN(n12514) );
  AOI21_X1 U14355 ( .B1(n7629), .B2(n12511), .A(n12510), .ZN(n12512) );
  NOR2_X1 U14356 ( .A1(n12512), .A2(n14611), .ZN(n12513) );
  AOI211_X1 U14357 ( .C1(n14580), .C2(n12515), .A(n12514), .B(n12513), .ZN(
        n12516) );
  OAI21_X1 U14358 ( .B1(n12517), .B2(n14574), .A(n12516), .ZN(P3_U3192) );
  AOI211_X1 U14359 ( .C1(n16523), .C2(n12520), .A(n12519), .B(n12518), .ZN(
        n12525) );
  AOI22_X1 U14360 ( .A1(n15536), .A2(n12521), .B1(n16525), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n12522) );
  OAI21_X1 U14361 ( .B1(n12525), .B2(n16525), .A(n12522), .ZN(P2_U3507) );
  OAI22_X1 U14362 ( .A1(n15594), .A2(n12615), .B1(n15586), .B2(n10029), .ZN(
        n12523) );
  INV_X1 U14363 ( .A(n12523), .ZN(n12524) );
  OAI21_X1 U14364 ( .B1(n12525), .B2(n16527), .A(n12524), .ZN(P2_U3454) );
  OAI21_X1 U14365 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n12534), .A(n12526), .ZN(
        n16273) );
  MUX2_X1 U14366 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n12628), .S(n12535), .Z(
        n16274) );
  NOR2_X1 U14367 ( .A1(n16273), .A2(n16274), .ZN(n16271) );
  AOI21_X1 U14368 ( .B1(n16269), .B2(P2_REG2_REG_10__SCAN_IN), .A(n16271), 
        .ZN(n12529) );
  INV_X1 U14369 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12527) );
  MUX2_X1 U14370 ( .A(n12527), .B(P2_REG2_REG_11__SCAN_IN), .S(n12537), .Z(
        n12528) );
  NAND2_X1 U14371 ( .A1(n12529), .A2(n12528), .ZN(n12650) );
  OAI21_X1 U14372 ( .B1(n12529), .B2(n12528), .A(n12650), .ZN(n12542) );
  INV_X1 U14373 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n12532) );
  INV_X1 U14374 ( .A(n12537), .ZN(n12654) );
  AND2_X1 U14375 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12530) );
  AOI21_X1 U14376 ( .B1(n16270), .B2(n12654), .A(n12530), .ZN(n12531) );
  OAI21_X1 U14377 ( .B1(n16278), .B2(n12532), .A(n12531), .ZN(n12541) );
  OAI21_X1 U14378 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n12534), .A(n12533), .ZN(
        n16265) );
  MUX2_X1 U14379 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n12536), .S(n12535), .Z(
        n16266) );
  NOR2_X1 U14380 ( .A1(n16265), .A2(n16266), .ZN(n16263) );
  XOR2_X1 U14381 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n12537), .Z(n12538) );
  AOI211_X1 U14382 ( .C1(n12539), .C2(n12538), .A(n16264), .B(n12653), .ZN(
        n12540) );
  AOI211_X1 U14383 ( .C1(n16257), .C2(n12542), .A(n12541), .B(n12540), .ZN(
        n12543) );
  INV_X1 U14384 ( .A(n12543), .ZN(P2_U3225) );
  XNOR2_X1 U14385 ( .A(n12268), .B(n14145), .ZN(n12546) );
  XNOR2_X1 U14386 ( .A(n12546), .B(n12556), .ZN(n14142) );
  NAND2_X1 U14387 ( .A1(n12545), .A2(n12544), .ZN(n14139) );
  INV_X1 U14388 ( .A(n12546), .ZN(n12547) );
  NAND2_X1 U14389 ( .A1(n12547), .A2(n12556), .ZN(n12548) );
  XNOR2_X1 U14390 ( .A(n12268), .B(n12842), .ZN(n12550) );
  NAND2_X1 U14391 ( .A1(n12550), .A2(n12549), .ZN(n12795) );
  INV_X1 U14392 ( .A(n12550), .ZN(n12551) );
  NAND2_X1 U14393 ( .A1(n12551), .A2(n14216), .ZN(n12552) );
  NAND2_X1 U14394 ( .A1(n12795), .A2(n12552), .ZN(n12554) );
  INV_X1 U14395 ( .A(n12796), .ZN(n12553) );
  AOI21_X1 U14396 ( .B1(n12555), .B2(n12554), .A(n12553), .ZN(n12561) );
  INV_X1 U14397 ( .A(n14290), .ZN(n14218) );
  AOI22_X1 U14398 ( .A1(n14218), .A2(n12933), .B1(n7422), .B2(n12556), .ZN(
        n12558) );
  OAI211_X1 U14399 ( .C1(n14282), .C2(n16537), .A(n12558), .B(n12557), .ZN(
        n12559) );
  AOI21_X1 U14400 ( .B1(n12841), .B2(n14287), .A(n12559), .ZN(n12560) );
  OAI21_X1 U14401 ( .B1(n12561), .B2(n14295), .A(n12560), .ZN(P3_U3170) );
  INV_X1 U14402 ( .A(n12562), .ZN(n12565) );
  OAI222_X1 U14403 ( .A1(n14968), .A2(n12565), .B1(n14959), .B2(n12564), .C1(
        P3_U3151), .C2(n12563), .ZN(P3_U3274) );
  INV_X1 U14404 ( .A(n12566), .ZN(n12569) );
  OAI222_X1 U14405 ( .A1(n16174), .A2(n12567), .B1(n13259), .B2(n12569), .C1(
        P1_U3086), .C2(n13158), .ZN(P1_U3338) );
  INV_X1 U14406 ( .A(n16255), .ZN(n15122) );
  INV_X1 U14407 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n12568) );
  OAI222_X1 U14408 ( .A1(n15122), .A2(P2_U3088), .B1(n15626), .B2(n12569), 
        .C1(n12568), .C2(n15628), .ZN(P2_U3310) );
  AOI21_X1 U14409 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(n12579) );
  OAI21_X1 U14410 ( .B1(n16723), .B2(n12574), .A(n12573), .ZN(n12577) );
  INV_X1 U14411 ( .A(n15749), .ZN(n13019) );
  OAI22_X1 U14412 ( .A1(n13019), .A2(n15717), .B1(n15716), .B2(n12575), .ZN(
        n12576) );
  AOI211_X1 U14413 ( .C1(n13637), .C2(n16719), .A(n12577), .B(n12576), .ZN(
        n12578) );
  OAI21_X1 U14414 ( .B1(n12579), .B2(n15729), .A(n12578), .ZN(P1_U3221) );
  NOR2_X1 U14415 ( .A1(n12621), .A2(n15232), .ZN(n12728) );
  XOR2_X1 U14416 ( .A(n12727), .B(n12726), .Z(n12588) );
  OR2_X1 U14417 ( .A1(n12611), .A2(n15043), .ZN(n12583) );
  OAI21_X1 U14418 ( .B1(n12921), .B2(n15162), .A(n12583), .ZN(n12639) );
  NAND2_X1 U14419 ( .A1(n15033), .A2(n12639), .ZN(n12584) );
  OAI211_X1 U14420 ( .C1(n15052), .C2(n12644), .A(n12585), .B(n12584), .ZN(
        n12586) );
  AOI21_X1 U14421 ( .B1(n12792), .B2(n15080), .A(n12586), .ZN(n12587) );
  OAI21_X1 U14422 ( .B1(n12588), .B2(n15077), .A(n12587), .ZN(P2_U3203) );
  INV_X1 U14423 ( .A(n14661), .ZN(n12589) );
  NAND2_X1 U14424 ( .A1(n12589), .A2(P3_U3897), .ZN(n12590) );
  OAI21_X1 U14425 ( .B1(P3_U3897), .B2(n12591), .A(n12590), .ZN(P3_U3518) );
  OAI21_X1 U14426 ( .B1(n12593), .B2(n14473), .A(n12592), .ZN(n12823) );
  INV_X1 U14427 ( .A(n12594), .ZN(n12595) );
  AOI21_X1 U14428 ( .B1(n14473), .B2(n12596), .A(n12595), .ZN(n12599) );
  AOI22_X1 U14429 ( .A1(n14777), .A2(n14216), .B1(n14217), .B2(n14779), .ZN(
        n12598) );
  NAND2_X1 U14430 ( .A1(n12823), .A2(n16678), .ZN(n12597) );
  OAI211_X1 U14431 ( .C1(n12599), .C2(n14817), .A(n12598), .B(n12597), .ZN(
        n12820) );
  AOI21_X1 U14432 ( .B1(n16643), .B2(n12823), .A(n12820), .ZN(n12607) );
  OAI22_X1 U14433 ( .A1(n14872), .A2(n12604), .B1(n16724), .B2(n12600), .ZN(
        n12601) );
  INV_X1 U14434 ( .A(n12601), .ZN(n12602) );
  OAI21_X1 U14435 ( .B1(n12607), .B2(n7821), .A(n12602), .ZN(P3_U3464) );
  INV_X1 U14436 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n12603) );
  OAI22_X1 U14437 ( .A1(n14938), .A2(n12604), .B1(n16727), .B2(n12603), .ZN(
        n12605) );
  INV_X1 U14438 ( .A(n12605), .ZN(n12606) );
  OAI21_X1 U14439 ( .B1(n12607), .B2(n16733), .A(n12606), .ZN(P3_U3405) );
  INV_X1 U14440 ( .A(n12608), .ZN(n12609) );
  NAND2_X1 U14441 ( .A1(n12610), .A2(n12609), .ZN(n12613) );
  OR2_X1 U14442 ( .A1(n12615), .A2(n12611), .ZN(n12612) );
  OR2_X1 U14443 ( .A1(n12789), .A2(n12621), .ZN(n12614) );
  INV_X1 U14444 ( .A(n12913), .ZN(n12619) );
  XNOR2_X1 U14445 ( .A(n12914), .B(n12619), .ZN(n12852) );
  INV_X1 U14446 ( .A(n12852), .ZN(n12633) );
  AND2_X1 U14447 ( .A1(n12615), .A2(n15091), .ZN(n12616) );
  OR2_X2 U14448 ( .A1(n12637), .A2(n12638), .ZN(n12635) );
  INV_X1 U14449 ( .A(n12621), .ZN(n15090) );
  NAND2_X1 U14450 ( .A1(n12789), .A2(n15090), .ZN(n12618) );
  OAI211_X1 U14451 ( .C1(n12620), .C2(n12619), .A(n12919), .B(n15446), .ZN(
        n12625) );
  OR2_X1 U14452 ( .A1(n12621), .A2(n15043), .ZN(n12623) );
  NAND2_X1 U14453 ( .A1(n15088), .A2(n15073), .ZN(n12622) );
  NAND2_X1 U14454 ( .A1(n12623), .A2(n12622), .ZN(n12732) );
  INV_X1 U14455 ( .A(n12732), .ZN(n12624) );
  NAND2_X1 U14456 ( .A1(n12625), .A2(n12624), .ZN(n12850) );
  NAND2_X1 U14457 ( .A1(n12850), .A2(n15429), .ZN(n12632) );
  INV_X1 U14458 ( .A(n12643), .ZN(n12627) );
  INV_X1 U14459 ( .A(n12926), .ZN(n12626) );
  AOI211_X1 U14460 ( .C1(n12853), .C2(n12627), .A(n7418), .B(n12626), .ZN(
        n12851) );
  NOR2_X1 U14461 ( .A1(n12917), .A2(n15456), .ZN(n12630) );
  OAI22_X1 U14462 ( .A1(n15429), .A2(n12628), .B1(n12734), .B2(n15427), .ZN(
        n12629) );
  AOI211_X1 U14463 ( .C1(n12851), .C2(n15461), .A(n12630), .B(n12629), .ZN(
        n12631) );
  OAI211_X1 U14464 ( .C1(n15435), .C2(n12633), .A(n12632), .B(n12631), .ZN(
        P2_U3255) );
  XOR2_X1 U14465 ( .A(n12638), .B(n12634), .Z(n12788) );
  INV_X1 U14466 ( .A(n12788), .ZN(n12649) );
  INV_X1 U14467 ( .A(n12635), .ZN(n12636) );
  AOI211_X1 U14468 ( .C1(n12638), .C2(n12637), .A(n11226), .B(n12636), .ZN(
        n12640) );
  OR2_X1 U14469 ( .A1(n12640), .A2(n12639), .ZN(n12786) );
  OAI21_X1 U14470 ( .B1(n12789), .B2(n12641), .A(n15232), .ZN(n12642) );
  OR2_X1 U14471 ( .A1(n12643), .A2(n12642), .ZN(n12785) );
  OAI22_X1 U14472 ( .A1(n15429), .A2(n11854), .B1(n12644), .B2(n15427), .ZN(
        n12645) );
  AOI21_X1 U14473 ( .B1(n12792), .B2(n15316), .A(n12645), .ZN(n12646) );
  OAI21_X1 U14474 ( .B1(n12785), .B2(n15318), .A(n12646), .ZN(n12647) );
  AOI21_X1 U14475 ( .B1(n12786), .B2(n15429), .A(n12647), .ZN(n12648) );
  OAI21_X1 U14476 ( .B1(n15435), .B2(n12649), .A(n12648), .ZN(P2_U3256) );
  OAI21_X1 U14477 ( .B1(n12654), .B2(P2_REG2_REG_11__SCAN_IN), .A(n12650), 
        .ZN(n12951) );
  XNOR2_X1 U14478 ( .A(n12951), .B(n12950), .ZN(n12651) );
  NOR2_X1 U14479 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n12651), .ZN(n12949) );
  AOI21_X1 U14480 ( .B1(n12651), .B2(P2_REG2_REG_12__SCAN_IN), .A(n12949), 
        .ZN(n12661) );
  XNOR2_X1 U14481 ( .A(n12946), .B(n12652), .ZN(n12656) );
  OAI21_X1 U14482 ( .B1(n12656), .B2(n12655), .A(n12945), .ZN(n12659) );
  NAND2_X1 U14483 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n13076)
         );
  NAND2_X1 U14484 ( .A1(n16224), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n12657) );
  OAI211_X1 U14485 ( .C1(n15128), .C2(n12950), .A(n13076), .B(n12657), .ZN(
        n12658) );
  AOI21_X1 U14486 ( .B1(n12659), .B2(n16230), .A(n12658), .ZN(n12660) );
  OAI21_X1 U14487 ( .B1(n12661), .B2(n16272), .A(n12660), .ZN(P2_U3226) );
  INV_X1 U14488 ( .A(n12665), .ZN(n12662) );
  NAND2_X1 U14489 ( .A1(n12663), .A2(n12662), .ZN(n12668) );
  INV_X1 U14490 ( .A(n12664), .ZN(n12666) );
  OAI21_X1 U14491 ( .B1(n14946), .B2(n12666), .A(n12665), .ZN(n12667) );
  AND2_X1 U14492 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  MUX2_X1 U14493 ( .A(P3_REG2_REG_0__SCAN_IN), .B(n12671), .S(n14819), .Z(
        n12676) );
  INV_X1 U14494 ( .A(n16509), .ZN(n14504) );
  OAI22_X1 U14495 ( .A1(n14809), .A2(n12674), .B1(n14792), .B2(n9678), .ZN(
        n12675) );
  OR2_X1 U14496 ( .A1(n12676), .A2(n12675), .ZN(P3_U3233) );
  INV_X1 U14497 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12680) );
  NAND2_X1 U14498 ( .A1(n9277), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12678) );
  NAND2_X1 U14499 ( .A1(n9031), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12677) );
  OAI211_X1 U14500 ( .C1(n12680), .C2(n12679), .A(n12678), .B(n12677), .ZN(
        n12681) );
  INV_X1 U14501 ( .A(n12681), .ZN(n12682) );
  NAND2_X1 U14502 ( .A1(n12683), .A2(n12682), .ZN(n14313) );
  NAND2_X1 U14503 ( .A1(n14313), .A2(P3_U3897), .ZN(n12684) );
  OAI21_X1 U14504 ( .B1(P3_U3897), .B2(n12685), .A(n12684), .ZN(P3_U3522) );
  INV_X1 U14505 ( .A(n12686), .ZN(n12687) );
  OAI21_X1 U14506 ( .B1(n12688), .B2(n11876), .A(n12687), .ZN(n12689) );
  NOR2_X1 U14507 ( .A1(n16293), .A2(n12689), .ZN(n12690) );
  XNOR2_X1 U14508 ( .A(n12689), .B(n16293), .ZN(n16290) );
  NOR2_X1 U14509 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n16290), .ZN(n16289) );
  NOR2_X1 U14510 ( .A1(n12690), .A2(n16289), .ZN(n12694) );
  INV_X1 U14511 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12691) );
  MUX2_X1 U14512 ( .A(n12691), .B(P1_REG2_REG_16__SCAN_IN), .S(n12859), .Z(
        n12692) );
  INV_X1 U14513 ( .A(n12692), .ZN(n12693) );
  NAND2_X1 U14514 ( .A1(n12693), .A2(n12694), .ZN(n12860) );
  OAI211_X1 U14515 ( .C1(n12694), .C2(n12693), .A(n15797), .B(n12860), .ZN(
        n12705) );
  NAND2_X1 U14516 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15682)
         );
  OR2_X1 U14517 ( .A1(n12695), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U14518 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  XNOR2_X1 U14519 ( .A(n12698), .B(n12699), .ZN(n16288) );
  NOR2_X1 U14520 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n16288), .ZN(n16287) );
  AOI21_X1 U14521 ( .B1(n12699), .B2(n12698), .A(n16287), .ZN(n12701) );
  XNOR2_X1 U14522 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12866), .ZN(n12700) );
  NAND2_X1 U14523 ( .A1(n12700), .A2(n12701), .ZN(n12865) );
  OAI211_X1 U14524 ( .C1(n12701), .C2(n12700), .A(n15807), .B(n12865), .ZN(
        n12702) );
  NAND2_X1 U14525 ( .A1(n15682), .A2(n12702), .ZN(n12703) );
  AOI21_X1 U14526 ( .B1(n16283), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12703), 
        .ZN(n12704) );
  OAI211_X1 U14527 ( .C1(n15791), .C2(n12866), .A(n12705), .B(n12704), .ZN(
        P1_U3259) );
  NAND2_X1 U14528 ( .A1(n14504), .A2(n14357), .ZN(n16512) );
  NAND2_X1 U14529 ( .A1(n16503), .A2(n16512), .ZN(n12706) );
  NAND2_X1 U14530 ( .A1(n14819), .A2(n12706), .ZN(n14813) );
  XNOR2_X1 U14531 ( .A(n12707), .B(n12708), .ZN(n16481) );
  INV_X1 U14532 ( .A(n16481), .ZN(n12721) );
  NAND2_X1 U14533 ( .A1(n12709), .A2(n16672), .ZN(n16483) );
  OR2_X1 U14534 ( .A1(n12707), .A2(n12711), .ZN(n12712) );
  NAND2_X1 U14535 ( .A1(n12710), .A2(n12712), .ZN(n12716) );
  NAND2_X1 U14536 ( .A1(n14366), .A2(n14779), .ZN(n12713) );
  NAND2_X1 U14537 ( .A1(n12714), .A2(n12713), .ZN(n12715) );
  AOI21_X1 U14538 ( .B1(n12716), .B2(n16500), .A(n12715), .ZN(n16484) );
  OAI21_X1 U14539 ( .B1(n14504), .B2(n16483), .A(n16484), .ZN(n12719) );
  OAI22_X1 U14540 ( .A1(n14819), .A2(n8925), .B1(n12717), .B2(n14792), .ZN(
        n12718) );
  AOI21_X1 U14541 ( .B1(n12719), .B2(n14819), .A(n12718), .ZN(n12720) );
  OAI21_X1 U14542 ( .B1(n14813), .B2(n12721), .A(n12720), .ZN(P3_U3232) );
  AOI22_X1 U14543 ( .A1(n12722), .A2(P3_STATE_REG_SCAN_IN), .B1(n10343), .B2(
        n14952), .ZN(n12723) );
  OAI21_X1 U14544 ( .B1(n12724), .B2(n14968), .A(n12723), .ZN(n12725) );
  INV_X1 U14545 ( .A(n12725), .ZN(P3_U3273) );
  INV_X1 U14546 ( .A(n12728), .ZN(n12729) );
  NAND2_X1 U14547 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  XNOR2_X1 U14548 ( .A(n12917), .B(n11679), .ZN(n13039) );
  NOR2_X1 U14549 ( .A1(n12921), .A2(n15232), .ZN(n13037) );
  XNOR2_X1 U14550 ( .A(n13039), .B(n13037), .ZN(n13035) );
  XOR2_X1 U14551 ( .A(n13036), .B(n13035), .Z(n12737) );
  AOI22_X1 U14552 ( .A1(n15033), .A2(n12732), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12733) );
  OAI21_X1 U14553 ( .B1(n15052), .B2(n12734), .A(n12733), .ZN(n12735) );
  AOI21_X1 U14554 ( .B1(n12853), .B2(n15080), .A(n12735), .ZN(n12736) );
  OAI21_X1 U14555 ( .B1(n12737), .B2(n15077), .A(n12736), .ZN(P2_U3189) );
  INV_X1 U14556 ( .A(n14317), .ZN(n12738) );
  NAND2_X1 U14557 ( .A1(n12738), .A2(P3_U3897), .ZN(n12739) );
  OAI21_X1 U14558 ( .B1(P3_U3897), .B2(n12740), .A(n12739), .ZN(P3_U3521) );
  INV_X1 U14559 ( .A(n14647), .ZN(n12741) );
  NAND2_X1 U14560 ( .A1(n12741), .A2(P3_U3897), .ZN(n12742) );
  OAI21_X1 U14561 ( .B1(P3_U3897), .B2(n12743), .A(n12742), .ZN(P3_U3519) );
  XOR2_X1 U14562 ( .A(n12745), .B(n12744), .Z(n12758) );
  INV_X1 U14563 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n16397) );
  NAND2_X1 U14564 ( .A1(n12746), .A2(n9089), .ZN(n12747) );
  NAND2_X1 U14565 ( .A1(n12747), .A2(n7607), .ZN(n12748) );
  NAND2_X1 U14566 ( .A1(n14603), .A2(n12748), .ZN(n12750) );
  OR2_X1 U14567 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12749), .ZN(n13251) );
  OAI211_X1 U14568 ( .C1(n16397), .C2(n14572), .A(n12750), .B(n13251), .ZN(
        n12755) );
  AOI21_X1 U14569 ( .B1(n12752), .B2(n16668), .A(n12751), .ZN(n12753) );
  NOR2_X1 U14570 ( .A1(n12753), .A2(n14611), .ZN(n12754) );
  AOI211_X1 U14571 ( .C1(n14580), .C2(n12756), .A(n12755), .B(n12754), .ZN(
        n12757) );
  OAI21_X1 U14572 ( .B1(n12758), .B2(n14574), .A(n12757), .ZN(P3_U3193) );
  OAI21_X1 U14573 ( .B1(n12760), .B2(n14474), .A(n12759), .ZN(n12830) );
  INV_X1 U14574 ( .A(n12830), .ZN(n12764) );
  AOI22_X1 U14575 ( .A1(n14777), .A2(n12933), .B1(n12963), .B2(n14779), .ZN(
        n12763) );
  OAI211_X1 U14576 ( .C1(n7462), .C2(n9014), .A(n16500), .B(n12761), .ZN(
        n12762) );
  OAI211_X1 U14577 ( .C1(n12764), .C2(n16503), .A(n12763), .B(n12762), .ZN(
        n12826) );
  AOI21_X1 U14578 ( .B1(n16643), .B2(n12830), .A(n12826), .ZN(n12769) );
  OAI22_X1 U14579 ( .A1(n14872), .A2(n12936), .B1(n16724), .B2(n12765), .ZN(
        n12766) );
  INV_X1 U14580 ( .A(n12766), .ZN(n12767) );
  OAI21_X1 U14581 ( .B1(n12769), .B2(n7821), .A(n12767), .ZN(P3_U3465) );
  INV_X1 U14582 ( .A(n14938), .ZN(n16734) );
  AOI22_X1 U14583 ( .A1(n16734), .A2(n12827), .B1(P3_REG0_REG_6__SCAN_IN), 
        .B2(n16733), .ZN(n12768) );
  OAI21_X1 U14584 ( .B1(n12769), .B2(n16733), .A(n12768), .ZN(P3_U3408) );
  INV_X1 U14585 ( .A(n14632), .ZN(n14169) );
  NAND2_X1 U14586 ( .A1(n14169), .A2(P3_U3897), .ZN(n12770) );
  OAI21_X1 U14587 ( .B1(P3_U3897), .B2(n12771), .A(n12770), .ZN(P3_U3520) );
  INV_X1 U14588 ( .A(n16512), .ZN(n12773) );
  OAI21_X1 U14589 ( .B1(n14360), .B2(n14468), .A(n12774), .ZN(n16533) );
  OAI22_X1 U14590 ( .A1(n14809), .A2(n16530), .B1(n14792), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n12783) );
  NAND2_X1 U14591 ( .A1(n12775), .A2(n16500), .ZN(n12781) );
  AOI21_X1 U14592 ( .B1(n16492), .B2(n12777), .A(n12776), .ZN(n12780) );
  AOI22_X1 U14593 ( .A1(n14777), .A2(n14366), .B1(n14216), .B2(n14779), .ZN(
        n12779) );
  NAND2_X1 U14594 ( .A1(n16533), .A2(n16678), .ZN(n12778) );
  OAI211_X1 U14595 ( .C1(n12781), .C2(n12780), .A(n12779), .B(n12778), .ZN(
        n16531) );
  MUX2_X1 U14596 ( .A(n16531), .B(P3_REG2_REG_3__SCAN_IN), .S(n16517), .Z(
        n12782) );
  AOI211_X1 U14597 ( .C1(n14758), .C2(n16533), .A(n12783), .B(n12782), .ZN(
        n12784) );
  INV_X1 U14598 ( .A(n12784), .ZN(P3_U3230) );
  INV_X1 U14599 ( .A(n12785), .ZN(n12787) );
  AOI211_X1 U14600 ( .C1(n16523), .C2(n12788), .A(n12787), .B(n12786), .ZN(
        n12794) );
  OAI22_X1 U14601 ( .A1(n12789), .A2(n15594), .B1(n16529), .B2(n10055), .ZN(
        n12790) );
  INV_X1 U14602 ( .A(n12790), .ZN(n12791) );
  OAI21_X1 U14603 ( .B1(n12794), .B2(n16527), .A(n12791), .ZN(P2_U3457) );
  AOI22_X1 U14604 ( .A1(n12792), .A2(n15536), .B1(n16525), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n12793) );
  OAI21_X1 U14605 ( .B1(n12794), .B2(n16525), .A(n12793), .ZN(P2_U3508) );
  NAND2_X1 U14606 ( .A1(n12796), .A2(n12795), .ZN(n14211) );
  XNOR2_X1 U14607 ( .A(n14163), .B(n14215), .ZN(n12797) );
  XNOR2_X1 U14608 ( .A(n12797), .B(n12933), .ZN(n14212) );
  NAND2_X1 U14609 ( .A1(n12797), .A2(n12837), .ZN(n12798) );
  XNOR2_X1 U14610 ( .A(n14163), .B(n12936), .ZN(n12799) );
  XNOR2_X1 U14611 ( .A(n12799), .B(n14217), .ZN(n12940) );
  NAND2_X1 U14612 ( .A1(n12799), .A2(n14217), .ZN(n12800) );
  XNOR2_X1 U14613 ( .A(n12268), .B(n12815), .ZN(n12903) );
  XNOR2_X1 U14614 ( .A(n12903), .B(n12963), .ZN(n12901) );
  XNOR2_X1 U14615 ( .A(n12902), .B(n12901), .ZN(n12805) );
  AOI22_X1 U14616 ( .A1(n14218), .A2(n14391), .B1(n7422), .B2(n14217), .ZN(
        n12802) );
  OAI211_X1 U14617 ( .C1(n14282), .C2(n16562), .A(n12802), .B(n12801), .ZN(
        n12803) );
  AOI21_X1 U14618 ( .B1(n12814), .B2(n14287), .A(n12803), .ZN(n12804) );
  OAI21_X1 U14619 ( .B1(n12805), .B2(n14295), .A(n12804), .ZN(P3_U3153) );
  XNOR2_X1 U14620 ( .A(n12807), .B(n12806), .ZN(n12813) );
  OAI21_X1 U14621 ( .B1(n12809), .B2(n14475), .A(n12808), .ZN(n16565) );
  OAI22_X1 U14622 ( .A1(n12810), .A2(n16495), .B1(n12907), .B2(n16497), .ZN(
        n12811) );
  AOI21_X1 U14623 ( .B1(n16565), .B2(n16678), .A(n12811), .ZN(n12812) );
  OAI21_X1 U14624 ( .B1(n14817), .B2(n12813), .A(n12812), .ZN(n16563) );
  INV_X1 U14625 ( .A(n16563), .ZN(n12819) );
  AOI22_X1 U14626 ( .A1(n14821), .A2(n12815), .B1(n16508), .B2(n12814), .ZN(
        n12816) );
  OAI21_X1 U14627 ( .B1(n9018), .B2(n14819), .A(n12816), .ZN(n12817) );
  AOI21_X1 U14628 ( .B1(n16565), .B2(n14758), .A(n12817), .ZN(n12818) );
  OAI21_X1 U14629 ( .B1(n12819), .B2(n16517), .A(n12818), .ZN(P3_U3226) );
  INV_X1 U14630 ( .A(n12820), .ZN(n12825) );
  AOI22_X1 U14631 ( .A1(n14821), .A2(n14215), .B1(n16508), .B2(n14219), .ZN(
        n12821) );
  OAI21_X1 U14632 ( .B1(n8986), .B2(n14819), .A(n12821), .ZN(n12822) );
  AOI21_X1 U14633 ( .B1(n12823), .B2(n14758), .A(n12822), .ZN(n12824) );
  OAI21_X1 U14634 ( .B1(n12825), .B2(n16517), .A(n12824), .ZN(P3_U3228) );
  INV_X1 U14635 ( .A(n12826), .ZN(n12832) );
  AOI22_X1 U14636 ( .A1(n14821), .A2(n12827), .B1(n16508), .B2(n12943), .ZN(
        n12828) );
  OAI21_X1 U14637 ( .B1(n9003), .B2(n14819), .A(n12828), .ZN(n12829) );
  AOI21_X1 U14638 ( .B1(n12830), .B2(n14758), .A(n12829), .ZN(n12831) );
  OAI21_X1 U14639 ( .B1(n12832), .B2(n16517), .A(n12831), .ZN(P3_U3227) );
  XNOR2_X1 U14640 ( .A(n12834), .B(n12833), .ZN(n12840) );
  OAI21_X1 U14641 ( .B1(n12836), .B2(n14470), .A(n12835), .ZN(n16540) );
  OAI22_X1 U14642 ( .A1(n16498), .A2(n16495), .B1(n12837), .B2(n16497), .ZN(
        n12838) );
  AOI21_X1 U14643 ( .B1(n16540), .B2(n16678), .A(n12838), .ZN(n12839) );
  OAI21_X1 U14644 ( .B1(n14817), .B2(n12840), .A(n12839), .ZN(n16538) );
  INV_X1 U14645 ( .A(n16538), .ZN(n12846) );
  AOI22_X1 U14646 ( .A1(n14821), .A2(n12842), .B1(n16508), .B2(n12841), .ZN(
        n12843) );
  OAI21_X1 U14647 ( .B1(n10884), .B2(n14819), .A(n12843), .ZN(n12844) );
  AOI21_X1 U14648 ( .B1(n16540), .B2(n14758), .A(n12844), .ZN(n12845) );
  OAI21_X1 U14649 ( .B1(n12846), .B2(n16517), .A(n12845), .ZN(P3_U3229) );
  INV_X1 U14650 ( .A(n12847), .ZN(n12877) );
  AOI22_X1 U14651 ( .A1(n13378), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n12848), .ZN(n12849) );
  OAI21_X1 U14652 ( .B1(n12877), .B2(n16178), .A(n12849), .ZN(P1_U3337) );
  AOI211_X1 U14653 ( .C1(n16523), .C2(n12852), .A(n12851), .B(n12850), .ZN(
        n12858) );
  AOI22_X1 U14654 ( .A1(n12853), .A2(n15536), .B1(n16525), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U14655 ( .B1(n12858), .B2(n16525), .A(n12854), .ZN(P2_U3509) );
  INV_X1 U14656 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n12855) );
  OAI22_X1 U14657 ( .A1(n12917), .A2(n15594), .B1(n15586), .B2(n12855), .ZN(
        n12856) );
  INV_X1 U14658 ( .A(n12856), .ZN(n12857) );
  OAI21_X1 U14659 ( .B1(n12858), .B2(n16527), .A(n12857), .ZN(P2_U3460) );
  NAND2_X1 U14660 ( .A1(n12859), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12861) );
  NAND2_X1 U14661 ( .A1(n12861), .A2(n12860), .ZN(n12864) );
  INV_X1 U14662 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13155) );
  NOR2_X1 U14663 ( .A1(n13158), .A2(n13155), .ZN(n12862) );
  AOI21_X1 U14664 ( .B1(n13155), .B2(n13158), .A(n12862), .ZN(n12863) );
  NAND2_X1 U14665 ( .A1(n12863), .A2(n12864), .ZN(n13154) );
  OAI211_X1 U14666 ( .C1(n12864), .C2(n12863), .A(n15797), .B(n13154), .ZN(
        n12873) );
  NAND2_X1 U14667 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15690)
         );
  XNOR2_X1 U14668 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n13158), .ZN(n12869) );
  INV_X1 U14669 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12867) );
  OAI21_X1 U14670 ( .B1(n12867), .B2(n12866), .A(n12865), .ZN(n12868) );
  NAND2_X1 U14671 ( .A1(n12869), .A2(n12868), .ZN(n13157) );
  OAI211_X1 U14672 ( .C1(n12869), .C2(n12868), .A(n15807), .B(n13157), .ZN(
        n12870) );
  NAND2_X1 U14673 ( .A1(n15690), .A2(n12870), .ZN(n12871) );
  AOI21_X1 U14674 ( .B1(n16283), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12871), 
        .ZN(n12872) );
  OAI211_X1 U14675 ( .C1(n15791), .C2(n13158), .A(n12873), .B(n12872), .ZN(
        P1_U3260) );
  NAND2_X1 U14676 ( .A1(n12875), .A2(n12874), .ZN(n12876) );
  OAI211_X1 U14677 ( .C1(n9618), .C2(n14959), .A(n12876), .B(n14515), .ZN(
        P3_U3272) );
  INV_X1 U14678 ( .A(n15123), .ZN(n15135) );
  OAI222_X1 U14679 ( .A1(n15628), .A2(n12878), .B1(n15626), .B2(n12877), .C1(
        P2_U3088), .C2(n15135), .ZN(P2_U3309) );
  XNOR2_X1 U14680 ( .A(n16633), .B(n15749), .ZN(n16618) );
  OR2_X1 U14681 ( .A1(n16633), .A2(n15749), .ZN(n12882) );
  XNOR2_X1 U14682 ( .A(n13649), .B(n15748), .ZN(n13864) );
  XNOR2_X1 U14683 ( .A(n12991), .B(n13864), .ZN(n16652) );
  OAI211_X1 U14684 ( .C1(n12884), .C2(n13864), .A(n16623), .B(n12996), .ZN(
        n16656) );
  NAND2_X1 U14685 ( .A1(n15749), .A2(n15955), .ZN(n16654) );
  AND2_X1 U14686 ( .A1(n16656), .A2(n16654), .ZN(n12885) );
  MUX2_X1 U14687 ( .A(n12886), .B(n12885), .S(n16014), .Z(n12893) );
  NAND2_X1 U14688 ( .A1(n16614), .A2(n13649), .ZN(n12887) );
  NAND2_X1 U14689 ( .A1(n12887), .A2(n16698), .ZN(n12888) );
  OR2_X1 U14690 ( .A1(n12888), .A2(n7628), .ZN(n12890) );
  NAND2_X1 U14691 ( .A1(n15747), .A2(n15956), .ZN(n12889) );
  NAND2_X1 U14692 ( .A1(n12890), .A2(n12889), .ZN(n16653) );
  OAI22_X1 U14693 ( .A1(n12994), .A2(n16587), .B1(n13017), .B2(n16036), .ZN(
        n12891) );
  AOI21_X1 U14694 ( .B1(n16653), .B2(n16636), .A(n12891), .ZN(n12892) );
  OAI211_X1 U14695 ( .C1(n15897), .C2(n16652), .A(n12893), .B(n12892), .ZN(
        P1_U3283) );
  OAI211_X1 U14696 ( .C1(n7637), .C2(n12895), .A(n12894), .B(n16714), .ZN(
        n12900) );
  INV_X1 U14697 ( .A(n15748), .ZN(n13220) );
  OAI22_X1 U14698 ( .A1(n13220), .A2(n16029), .B1(n12896), .B2(n16031), .ZN(
        n16622) );
  NOR2_X1 U14699 ( .A1(n16723), .A2(n16629), .ZN(n12897) );
  AOI211_X1 U14700 ( .C1(n16716), .C2(n16622), .A(n12898), .B(n12897), .ZN(
        n12899) );
  OAI211_X1 U14701 ( .C1(n16616), .C2(n15712), .A(n12900), .B(n12899), .ZN(
        P1_U3231) );
  NAND2_X1 U14702 ( .A1(n12902), .A2(n12901), .ZN(n12906) );
  INV_X1 U14703 ( .A(n12903), .ZN(n12904) );
  NAND2_X1 U14704 ( .A1(n12904), .A2(n12963), .ZN(n12905) );
  XNOR2_X1 U14705 ( .A(n14163), .B(n16595), .ZN(n13088) );
  XNOR2_X1 U14706 ( .A(n13088), .B(n12907), .ZN(n13086) );
  XNOR2_X1 U14707 ( .A(n13087), .B(n13086), .ZN(n12912) );
  AOI22_X1 U14708 ( .A1(n14218), .A2(n14398), .B1(n7422), .B2(n12963), .ZN(
        n12909) );
  OAI211_X1 U14709 ( .C1(n16595), .C2(n14282), .A(n12909), .B(n12908), .ZN(
        n12910) );
  AOI21_X1 U14710 ( .B1(n12969), .B2(n14287), .A(n12910), .ZN(n12911) );
  OAI21_X1 U14711 ( .B1(n12912), .B2(n14295), .A(n12911), .ZN(P3_U3161) );
  OR2_X1 U14712 ( .A1(n12917), .A2(n12921), .ZN(n12915) );
  NAND2_X1 U14713 ( .A1(n12916), .A2(n12915), .ZN(n12979) );
  XOR2_X1 U14714 ( .A(n12978), .B(n12979), .Z(n13050) );
  INV_X1 U14715 ( .A(n13050), .ZN(n12932) );
  INV_X1 U14716 ( .A(n12921), .ZN(n15089) );
  NAND2_X1 U14717 ( .A1(n12917), .A2(n15089), .ZN(n12918) );
  AOI21_X1 U14718 ( .B1(n12978), .B2(n12920), .A(n7611), .ZN(n12925) );
  OR2_X1 U14719 ( .A1(n12921), .A2(n15043), .ZN(n12923) );
  NAND2_X1 U14720 ( .A1(n15087), .A2(n15073), .ZN(n12922) );
  NAND2_X1 U14721 ( .A1(n12923), .A2(n12922), .ZN(n13028) );
  INV_X1 U14722 ( .A(n13028), .ZN(n12924) );
  OAI21_X1 U14723 ( .B1(n12925), .B2(n11226), .A(n12924), .ZN(n13048) );
  NAND2_X1 U14724 ( .A1(n13048), .A2(n15429), .ZN(n12931) );
  AOI211_X1 U14725 ( .C1(n13052), .C2(n12926), .A(n7418), .B(n7669), .ZN(
        n13049) );
  NOR2_X1 U14726 ( .A1(n12927), .A2(n15456), .ZN(n12929) );
  OAI22_X1 U14727 ( .A1(n15429), .A2(n12527), .B1(n13030), .B2(n15427), .ZN(
        n12928) );
  AOI211_X1 U14728 ( .C1(n13049), .C2(n15461), .A(n12929), .B(n12928), .ZN(
        n12930) );
  OAI211_X1 U14729 ( .C1(n15435), .C2(n12932), .A(n12931), .B(n12930), .ZN(
        P2_U3254) );
  AOI22_X1 U14730 ( .A1(n14218), .A2(n12963), .B1(n7422), .B2(n12933), .ZN(
        n12935) );
  OAI211_X1 U14731 ( .C1(n12936), .C2(n14282), .A(n12935), .B(n12934), .ZN(
        n12942) );
  INV_X1 U14732 ( .A(n12937), .ZN(n12938) );
  AOI211_X1 U14733 ( .C1(n12940), .C2(n12939), .A(n14295), .B(n12938), .ZN(
        n12941) );
  AOI211_X1 U14734 ( .C1(n12943), .C2(n14287), .A(n12942), .B(n12941), .ZN(
        n12944) );
  INV_X1 U14735 ( .A(n12944), .ZN(P3_U3179) );
  XNOR2_X1 U14736 ( .A(n13105), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n12948) );
  OAI21_X1 U14737 ( .B1(n12946), .B2(P2_REG1_REG_12__SCAN_IN), .A(n12945), 
        .ZN(n12947) );
  NOR2_X1 U14738 ( .A1(n12947), .A2(n12948), .ZN(n13099) );
  AOI211_X1 U14739 ( .C1(n12948), .C2(n12947), .A(n16264), .B(n13099), .ZN(
        n12959) );
  INV_X1 U14740 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n12957) );
  AOI21_X1 U14741 ( .B1(n12951), .B2(n12950), .A(n12949), .ZN(n12953) );
  MUX2_X1 U14742 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n13130), .S(n13105), .Z(
        n12952) );
  NAND2_X1 U14743 ( .A1(n12952), .A2(n12953), .ZN(n13103) );
  OAI211_X1 U14744 ( .C1(n12953), .C2(n12952), .A(n13103), .B(n16257), .ZN(
        n12956) );
  AND2_X1 U14745 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n12954) );
  AOI21_X1 U14746 ( .B1(n16270), .B2(n13105), .A(n12954), .ZN(n12955) );
  OAI211_X1 U14747 ( .C1(n16278), .C2(n12957), .A(n12956), .B(n12955), .ZN(
        n12958) );
  OR2_X1 U14748 ( .A1(n12959), .A2(n12958), .ZN(P2_U3227) );
  INV_X1 U14749 ( .A(n12960), .ZN(n12961) );
  AOI21_X1 U14750 ( .B1(n14479), .B2(n12962), .A(n12961), .ZN(n12968) );
  AOI22_X1 U14751 ( .A1(n14779), .A2(n14398), .B1(n12963), .B2(n14777), .ZN(
        n12967) );
  OAI21_X1 U14752 ( .B1(n12965), .B2(n14479), .A(n12964), .ZN(n16598) );
  NAND2_X1 U14753 ( .A1(n16598), .A2(n16678), .ZN(n12966) );
  OAI211_X1 U14754 ( .C1(n12968), .C2(n14817), .A(n12967), .B(n12966), .ZN(
        n16596) );
  INV_X1 U14755 ( .A(n16596), .ZN(n12974) );
  AOI22_X1 U14756 ( .A1(n14821), .A2(n12970), .B1(n16508), .B2(n12969), .ZN(
        n12971) );
  OAI21_X1 U14757 ( .B1(n9034), .B2(n14819), .A(n12971), .ZN(n12972) );
  AOI21_X1 U14758 ( .B1(n16598), .B2(n14758), .A(n12972), .ZN(n12973) );
  OAI21_X1 U14759 ( .B1(n12974), .B2(n16517), .A(n12973), .ZN(P3_U3225) );
  NAND2_X1 U14760 ( .A1(n13052), .A2(n13072), .ZN(n12975) );
  INV_X1 U14761 ( .A(n12982), .ZN(n13119) );
  OAI211_X1 U14762 ( .C1(n7633), .C2(n12982), .A(n15446), .B(n13124), .ZN(
        n12977) );
  AND2_X1 U14763 ( .A1(n15088), .A2(n15225), .ZN(n12976) );
  AOI21_X1 U14764 ( .B1(n15086), .B2(n15073), .A(n12976), .ZN(n13078) );
  NAND2_X1 U14765 ( .A1(n12977), .A2(n13078), .ZN(n13187) );
  INV_X1 U14766 ( .A(n13187), .ZN(n12989) );
  NAND2_X1 U14767 ( .A1(n12979), .A2(n12978), .ZN(n12981) );
  NAND2_X1 U14768 ( .A1(n13052), .A2(n15088), .ZN(n12980) );
  XNOR2_X1 U14769 ( .A(n13120), .B(n12982), .ZN(n13189) );
  AOI211_X1 U14770 ( .C1(n13191), .C2(n12983), .A(n7418), .B(n13129), .ZN(
        n13188) );
  NAND2_X1 U14771 ( .A1(n13188), .A2(n15461), .ZN(n12986) );
  INV_X1 U14772 ( .A(n12984), .ZN(n13075) );
  AOI22_X1 U14773 ( .A1(n15454), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n13075), 
        .B2(n15452), .ZN(n12985) );
  OAI211_X1 U14774 ( .C1(n7668), .C2(n15456), .A(n12986), .B(n12985), .ZN(
        n12987) );
  AOI21_X1 U14775 ( .B1(n15336), .B2(n13189), .A(n12987), .ZN(n12988) );
  OAI21_X1 U14776 ( .B1(n12989), .B2(n15454), .A(n12988), .ZN(P2_U3253) );
  INV_X1 U14777 ( .A(n13864), .ZN(n12990) );
  OR2_X1 U14778 ( .A1(n13649), .A2(n15748), .ZN(n12992) );
  XNOR2_X1 U14779 ( .A(n13656), .B(n15747), .ZN(n13866) );
  XNOR2_X1 U14780 ( .A(n13149), .B(n13866), .ZN(n13010) );
  NAND2_X1 U14781 ( .A1(n12994), .A2(n15748), .ZN(n12995) );
  OAI211_X1 U14782 ( .C1(n12997), .C2(n13866), .A(n13138), .B(n16623), .ZN(
        n12999) );
  AOI22_X1 U14783 ( .A1(n15956), .A2(n15746), .B1(n15748), .B2(n15955), .ZN(
        n12998) );
  AND2_X1 U14784 ( .A1(n12999), .A2(n12998), .ZN(n13009) );
  INV_X1 U14785 ( .A(n13009), .ZN(n13005) );
  OR2_X1 U14786 ( .A1(n7628), .A2(n13136), .ZN(n13000) );
  AND2_X1 U14787 ( .A1(n13201), .A2(n13000), .ZN(n13007) );
  NAND2_X1 U14788 ( .A1(n13007), .A2(n15987), .ZN(n13003) );
  INV_X1 U14789 ( .A(n13219), .ZN(n13001) );
  AOI22_X1 U14790 ( .A1(n16642), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n13001), 
        .B2(n16631), .ZN(n13002) );
  OAI211_X1 U14791 ( .C1(n13136), .C2(n16587), .A(n13003), .B(n13002), .ZN(
        n13004) );
  AOI21_X1 U14792 ( .B1(n13005), .B2(n16014), .A(n13004), .ZN(n13006) );
  OAI21_X1 U14793 ( .B1(n15897), .B2(n13010), .A(n13006), .ZN(P1_U3282) );
  AOI22_X1 U14794 ( .A1(n13007), .A2(n16698), .B1(n16696), .B2(n13656), .ZN(
        n13008) );
  OAI211_X1 U14795 ( .C1(n16142), .C2(n13010), .A(n13009), .B(n13008), .ZN(
        n13012) );
  NAND2_X1 U14796 ( .A1(n13012), .A2(n16694), .ZN(n13011) );
  OAI21_X1 U14797 ( .B1(n16694), .B2(n11086), .A(n13011), .ZN(P1_U3492) );
  NAND2_X1 U14798 ( .A1(n13012), .A2(n16708), .ZN(n13013) );
  OAI21_X1 U14799 ( .B1(n16708), .B2(n11082), .A(n13013), .ZN(P1_U3539) );
  OAI211_X1 U14800 ( .C1(n13016), .C2(n13015), .A(n13014), .B(n16714), .ZN(
        n13024) );
  INV_X1 U14801 ( .A(n13017), .ZN(n13022) );
  INV_X1 U14802 ( .A(n13018), .ZN(n13021) );
  INV_X1 U14803 ( .A(n15747), .ZN(n13328) );
  OAI22_X1 U14804 ( .A1(n13328), .A2(n15717), .B1(n15716), .B2(n13019), .ZN(
        n13020) );
  AOI211_X1 U14805 ( .C1(n13022), .C2(n13331), .A(n13021), .B(n13020), .ZN(
        n13023) );
  OAI211_X1 U14806 ( .C1(n12994), .C2(n15712), .A(n13024), .B(n13023), .ZN(
        P1_U3217) );
  INV_X1 U14807 ( .A(n13025), .ZN(n13026) );
  OAI222_X1 U14808 ( .A1(n16174), .A2(n8551), .B1(n13259), .B2(n13026), .C1(
        n16033), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U14809 ( .A1(n13027), .A2(P2_U3088), .B1(n15626), .B2(n13026), 
        .C1(n11568), .C2(n15628), .ZN(P2_U3308) );
  AOI22_X1 U14810 ( .A1(n15033), .A2(n13028), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13029) );
  OAI21_X1 U14811 ( .B1(n15052), .B2(n13030), .A(n13029), .ZN(n13046) );
  XNOR2_X1 U14812 ( .A(n13052), .B(n11679), .ZN(n13031) );
  AND2_X1 U14813 ( .A1(n15088), .A2(n7418), .ZN(n13032) );
  NAND2_X1 U14814 ( .A1(n13031), .A2(n13032), .ZN(n13079) );
  INV_X1 U14815 ( .A(n13031), .ZN(n13073) );
  INV_X1 U14816 ( .A(n13032), .ZN(n13033) );
  NAND2_X1 U14817 ( .A1(n13073), .A2(n13033), .ZN(n13034) );
  NAND2_X1 U14818 ( .A1(n13079), .A2(n13034), .ZN(n13044) );
  INV_X1 U14819 ( .A(n13037), .ZN(n13038) );
  NAND2_X1 U14820 ( .A1(n13039), .A2(n13038), .ZN(n13040) );
  AOI211_X1 U14821 ( .C1(n13044), .C2(n13043), .A(n15077), .B(n7624), .ZN(
        n13045) );
  AOI211_X1 U14822 ( .C1(n13052), .C2(n15080), .A(n13046), .B(n13045), .ZN(
        n13047) );
  INV_X1 U14823 ( .A(n13047), .ZN(P2_U3208) );
  AOI211_X1 U14824 ( .C1(n16523), .C2(n13050), .A(n13049), .B(n13048), .ZN(
        n13054) );
  INV_X1 U14825 ( .A(n15594), .ZN(n15599) );
  AOI22_X1 U14826 ( .A1(n13052), .A2(n15599), .B1(P2_REG0_REG_11__SCAN_IN), 
        .B2(n16527), .ZN(n13051) );
  OAI21_X1 U14827 ( .B1(n13054), .B2(n16527), .A(n13051), .ZN(P2_U3463) );
  AOI22_X1 U14828 ( .A1(n13052), .A2(n15536), .B1(P2_REG1_REG_11__SCAN_IN), 
        .B2(n16525), .ZN(n13053) );
  OAI21_X1 U14829 ( .B1(n13054), .B2(n16525), .A(n13053), .ZN(P2_U3510) );
  AOI21_X1 U14830 ( .B1(n13057), .B2(n13056), .A(n13055), .ZN(n13065) );
  NOR2_X1 U14831 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13058), .ZN(n13315) );
  AOI21_X1 U14832 ( .B1(n13061), .B2(n13060), .A(n13059), .ZN(n13062) );
  NOR2_X1 U14833 ( .A1(n14541), .A2(n13062), .ZN(n13063) );
  AOI211_X1 U14834 ( .C1(n14609), .C2(P3_ADDR_REG_12__SCAN_IN), .A(n13315), 
        .B(n13063), .ZN(n13064) );
  OAI21_X1 U14835 ( .B1(n13065), .B2(n14611), .A(n13064), .ZN(n13069) );
  AOI211_X1 U14836 ( .C1(n13067), .C2(n13066), .A(n14574), .B(n7630), .ZN(
        n13068) );
  AOI211_X1 U14837 ( .C1(n14580), .C2(n13070), .A(n13069), .B(n13068), .ZN(
        n13071) );
  INV_X1 U14838 ( .A(n13071), .ZN(P3_U3194) );
  NOR3_X1 U14839 ( .A1(n13073), .A2(n13072), .A3(n15067), .ZN(n13074) );
  AOI21_X1 U14840 ( .B1(n7624), .B2(n15070), .A(n13074), .ZN(n13085) );
  XNOR2_X1 U14841 ( .A(n13191), .B(n11679), .ZN(n13172) );
  NAND2_X1 U14842 ( .A1(n15087), .A2(n7418), .ZN(n13173) );
  XNOR2_X1 U14843 ( .A(n13172), .B(n13173), .ZN(n13084) );
  NAND2_X1 U14844 ( .A1(n15074), .A2(n13075), .ZN(n13077) );
  OAI211_X1 U14845 ( .C1(n13078), .C2(n15076), .A(n13077), .B(n13076), .ZN(
        n13082) );
  AND2_X1 U14846 ( .A1(n13084), .A2(n13079), .ZN(n13080) );
  NOR2_X1 U14847 ( .A1(n13176), .A2(n15077), .ZN(n13081) );
  AOI211_X1 U14848 ( .C1(n13191), .C2(n15080), .A(n13082), .B(n13081), .ZN(
        n13083) );
  OAI21_X1 U14849 ( .B1(n13085), .B2(n13084), .A(n13083), .ZN(P2_U3196) );
  XNOR2_X1 U14850 ( .A(n14163), .B(n13213), .ZN(n13246) );
  XNOR2_X1 U14851 ( .A(n13246), .B(n13262), .ZN(n13093) );
  NAND2_X1 U14852 ( .A1(n13088), .A2(n14391), .ZN(n13089) );
  INV_X1 U14853 ( .A(n13093), .ZN(n13090) );
  INV_X1 U14854 ( .A(n14128), .ZN(n13091) );
  AOI21_X1 U14855 ( .B1(n13093), .B2(n13092), .A(n13091), .ZN(n13098) );
  AOI22_X1 U14856 ( .A1(n14218), .A2(n14403), .B1(n7422), .B2(n14391), .ZN(
        n13095) );
  OAI211_X1 U14857 ( .C1(n14282), .C2(n14397), .A(n13095), .B(n13094), .ZN(
        n13096) );
  AOI21_X1 U14858 ( .B1(n13277), .B2(n14287), .A(n13096), .ZN(n13097) );
  OAI21_X1 U14859 ( .B1(n13098), .B2(n14295), .A(n13097), .ZN(P3_U3171) );
  XNOR2_X1 U14860 ( .A(n13436), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n13100) );
  AOI211_X1 U14861 ( .C1(n13101), .C2(n13100), .A(n16264), .B(n13435), .ZN(
        n13115) );
  INV_X1 U14862 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U14863 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n13291)
         );
  INV_X1 U14864 ( .A(n13291), .ZN(n13102) );
  AOI21_X1 U14865 ( .B1(n16270), .B2(n13436), .A(n13102), .ZN(n13112) );
  INV_X1 U14866 ( .A(n13103), .ZN(n13104) );
  AOI21_X1 U14867 ( .B1(n13105), .B2(P2_REG2_REG_13__SCAN_IN), .A(n13104), 
        .ZN(n13107) );
  NAND2_X1 U14868 ( .A1(n13436), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13108) );
  OAI211_X1 U14869 ( .C1(n13436), .C2(P2_REG2_REG_14__SCAN_IN), .A(n13107), 
        .B(n13108), .ZN(n13106) );
  INV_X1 U14870 ( .A(n13106), .ZN(n13440) );
  NOR2_X1 U14871 ( .A1(n13436), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13441) );
  INV_X1 U14872 ( .A(n13441), .ZN(n13109) );
  AOI21_X1 U14873 ( .B1(n13109), .B2(n13108), .A(n13107), .ZN(n13110) );
  OAI21_X1 U14874 ( .B1(n13440), .B2(n13110), .A(n16257), .ZN(n13111) );
  OAI211_X1 U14875 ( .C1(n16278), .C2(n13113), .A(n13112), .B(n13111), .ZN(
        n13114) );
  OR2_X1 U14876 ( .A1(n13115), .A2(n13114), .ZN(P2_U3228) );
  INV_X1 U14877 ( .A(n13116), .ZN(n13166) );
  OAI222_X1 U14878 ( .A1(n15628), .A2(n13118), .B1(P2_U3088), .B2(n13117), 
        .C1(n13166), .C2(n15626), .ZN(P2_U3307) );
  NAND2_X1 U14879 ( .A1(n13191), .A2(n15087), .ZN(n13121) );
  XNOR2_X1 U14880 ( .A(n13239), .B(n13237), .ZN(n13272) );
  INV_X1 U14881 ( .A(n13272), .ZN(n13135) );
  INV_X1 U14882 ( .A(n15087), .ZN(n13122) );
  OR2_X1 U14883 ( .A1(n13191), .A2(n13122), .ZN(n13123) );
  NAND2_X1 U14884 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  OAI211_X1 U14885 ( .C1(n13125), .C2(n13237), .A(n13231), .B(n15446), .ZN(
        n13128) );
  OR2_X1 U14886 ( .A1(n13352), .A2(n15162), .ZN(n13127) );
  NAND2_X1 U14887 ( .A1(n15087), .A2(n15225), .ZN(n13126) );
  AND2_X1 U14888 ( .A1(n13127), .A2(n13126), .ZN(n13182) );
  NAND2_X1 U14889 ( .A1(n13128), .A2(n13182), .ZN(n13270) );
  NAND2_X1 U14890 ( .A1(n13270), .A2(n15429), .ZN(n13134) );
  AOI211_X1 U14891 ( .C1(n13274), .C2(n7667), .A(n7418), .B(n13234), .ZN(
        n13271) );
  NOR2_X1 U14892 ( .A1(n13240), .A2(n15456), .ZN(n13132) );
  OAI22_X1 U14893 ( .A1(n15429), .A2(n13130), .B1(n13180), .B2(n15427), .ZN(
        n13131) );
  AOI211_X1 U14894 ( .C1(n13271), .C2(n15461), .A(n13132), .B(n13131), .ZN(
        n13133) );
  OAI211_X1 U14895 ( .C1(n15435), .C2(n13135), .A(n13134), .B(n13133), .ZN(
        P2_U3252) );
  NAND2_X1 U14896 ( .A1(n13136), .A2(n15747), .ZN(n13137) );
  XNOR2_X1 U14897 ( .A(n13659), .B(n15746), .ZN(n13869) );
  NAND2_X1 U14898 ( .A1(n13198), .A2(n13869), .ZN(n13197) );
  INV_X1 U14899 ( .A(n15746), .ZN(n13221) );
  NAND2_X1 U14900 ( .A1(n13197), .A2(n13139), .ZN(n13141) );
  XNOR2_X1 U14901 ( .A(n16697), .B(n15643), .ZN(n13868) );
  INV_X1 U14902 ( .A(n13868), .ZN(n13140) );
  NAND2_X1 U14903 ( .A1(n13141), .A2(n13140), .ZN(n13418) );
  OAI21_X1 U14904 ( .B1(n13141), .B2(n13140), .A(n13418), .ZN(n16703) );
  OR2_X1 U14905 ( .A1(n13201), .A2(n13659), .ZN(n13203) );
  AND2_X1 U14906 ( .A1(n13203), .A2(n16697), .ZN(n13142) );
  NOR2_X1 U14907 ( .A1(n13422), .A2(n13142), .ZN(n16699) );
  INV_X1 U14908 ( .A(n16697), .ZN(n13488) );
  NAND2_X1 U14909 ( .A1(n15744), .A2(n15956), .ZN(n13144) );
  NAND2_X1 U14910 ( .A1(n15746), .A2(n15955), .ZN(n13143) );
  NAND2_X1 U14911 ( .A1(n13144), .A2(n13143), .ZN(n16695) );
  INV_X1 U14912 ( .A(n16695), .ZN(n13145) );
  OAI22_X1 U14913 ( .A1(n16642), .A2(n13145), .B1(n13484), .B2(n16036), .ZN(
        n13146) );
  AOI21_X1 U14914 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n16642), .A(n13146), 
        .ZN(n13147) );
  OAI21_X1 U14915 ( .B1(n13488), .B2(n16587), .A(n13147), .ZN(n13148) );
  AOI21_X1 U14916 ( .B1(n16699), .B2(n15987), .A(n13148), .ZN(n13153) );
  NAND2_X1 U14917 ( .A1(n13656), .A2(n15747), .ZN(n13150) );
  OR2_X1 U14918 ( .A1(n13659), .A2(n15746), .ZN(n13151) );
  XNOR2_X1 U14919 ( .A(n13414), .B(n13868), .ZN(n16706) );
  NAND2_X1 U14920 ( .A1(n16706), .A2(n15929), .ZN(n13152) );
  OAI211_X1 U14921 ( .C1(n16703), .C2(n15970), .A(n13153), .B(n13152), .ZN(
        P1_U3280) );
  INV_X1 U14922 ( .A(n13378), .ZN(n13165) );
  OAI21_X1 U14923 ( .B1(n13155), .B2(n13158), .A(n13154), .ZN(n13373) );
  XOR2_X1 U14924 ( .A(n13373), .B(n13378), .Z(n13156) );
  NAND2_X1 U14925 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13156), .ZN(n13375) );
  OAI211_X1 U14926 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13156), .A(n15797), 
        .B(n13375), .ZN(n13164) );
  NAND2_X1 U14927 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15715)
         );
  INV_X1 U14928 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13159) );
  OAI21_X1 U14929 ( .B1(n13159), .B2(n13158), .A(n13157), .ZN(n13377) );
  XNOR2_X1 U14930 ( .A(n13377), .B(n13165), .ZN(n13160) );
  NAND2_X1 U14931 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n13160), .ZN(n13379) );
  OAI211_X1 U14932 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13160), .A(n15807), 
        .B(n13379), .ZN(n13161) );
  NAND2_X1 U14933 ( .A1(n15715), .A2(n13161), .ZN(n13162) );
  AOI21_X1 U14934 ( .B1(n16283), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n13162), 
        .ZN(n13163) );
  OAI211_X1 U14935 ( .C1(n15791), .C2(n13165), .A(n13164), .B(n13163), .ZN(
        P1_U3261) );
  OAI222_X1 U14936 ( .A1(n16174), .A2(n13167), .B1(P1_U3086), .B2(n13850), 
        .C1(n16178), .C2(n13166), .ZN(P1_U3335) );
  XNOR2_X1 U14937 ( .A(n13240), .B(n7695), .ZN(n13168) );
  NOR2_X1 U14938 ( .A1(n13284), .A2(n15232), .ZN(n13169) );
  NAND2_X1 U14939 ( .A1(n13168), .A2(n13169), .ZN(n13293) );
  INV_X1 U14940 ( .A(n13168), .ZN(n13285) );
  INV_X1 U14941 ( .A(n13169), .ZN(n13170) );
  NAND2_X1 U14942 ( .A1(n13285), .A2(n13170), .ZN(n13171) );
  NAND2_X1 U14943 ( .A1(n13293), .A2(n13171), .ZN(n13178) );
  INV_X1 U14944 ( .A(n13172), .ZN(n13174) );
  NAND2_X1 U14945 ( .A1(n13174), .A2(n13173), .ZN(n13175) );
  INV_X1 U14946 ( .A(n13295), .ZN(n13287) );
  AOI211_X1 U14947 ( .C1(n13178), .C2(n13177), .A(n15077), .B(n13287), .ZN(
        n13179) );
  INV_X1 U14948 ( .A(n13179), .ZN(n13186) );
  INV_X1 U14949 ( .A(n13180), .ZN(n13184) );
  OAI22_X1 U14950 ( .A1(n15076), .A2(n13182), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13181), .ZN(n13183) );
  AOI21_X1 U14951 ( .B1(n13184), .B2(n15074), .A(n13183), .ZN(n13185) );
  OAI211_X1 U14952 ( .C1(n13240), .C2(n15066), .A(n13186), .B(n13185), .ZN(
        P2_U3206) );
  AOI211_X1 U14953 ( .C1(n16523), .C2(n13189), .A(n13188), .B(n13187), .ZN(
        n13193) );
  AOI22_X1 U14954 ( .A1(n13191), .A2(n15536), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n16525), .ZN(n13190) );
  OAI21_X1 U14955 ( .B1(n13193), .B2(n16525), .A(n13190), .ZN(P2_U3511) );
  AOI22_X1 U14956 ( .A1(n13191), .A2(n15599), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n16527), .ZN(n13192) );
  OAI21_X1 U14957 ( .B1(n13193), .B2(n16527), .A(n13192), .ZN(P2_U3466) );
  INV_X1 U14958 ( .A(n13194), .ZN(n13195) );
  AOI21_X1 U14959 ( .B1(n13869), .B2(n13196), .A(n13195), .ZN(n16683) );
  OAI211_X1 U14960 ( .C1(n13198), .C2(n13869), .A(n13197), .B(n16623), .ZN(
        n13200) );
  AOI22_X1 U14961 ( .A1(n15956), .A2(n15745), .B1(n15747), .B2(n15955), .ZN(
        n13199) );
  OAI211_X1 U14962 ( .C1(n16683), .C2(n16619), .A(n13200), .B(n13199), .ZN(
        n16688) );
  NAND2_X1 U14963 ( .A1(n16688), .A2(n16014), .ZN(n13207) );
  OAI22_X1 U14964 ( .A1(n16014), .A2(n11637), .B1(n13326), .B2(n16036), .ZN(
        n13205) );
  NAND2_X1 U14965 ( .A1(n13201), .A2(n13659), .ZN(n13202) );
  NAND2_X1 U14966 ( .A1(n13203), .A2(n13202), .ZN(n16687) );
  INV_X1 U14967 ( .A(n15987), .ZN(n16475) );
  NOR2_X1 U14968 ( .A1(n16687), .A2(n16475), .ZN(n13204) );
  AOI211_X1 U14969 ( .C1(n16632), .C2(n13659), .A(n13205), .B(n13204), .ZN(
        n13206) );
  OAI211_X1 U14970 ( .C1(n16683), .C2(n16006), .A(n13207), .B(n13206), .ZN(
        P1_U3281) );
  OR2_X1 U14971 ( .A1(n8254), .A2(n13209), .ZN(n14390) );
  XNOR2_X1 U14972 ( .A(n13210), .B(n14390), .ZN(n13283) );
  XNOR2_X1 U14973 ( .A(n13211), .B(n14390), .ZN(n13212) );
  AOI222_X1 U14974 ( .A1(n13212), .A2(n16500), .B1(n14403), .B2(n14779), .C1(
        n14391), .C2(n14777), .ZN(n13279) );
  OAI21_X1 U14975 ( .B1(n14894), .B2(n13283), .A(n13279), .ZN(n13228) );
  INV_X1 U14976 ( .A(n13228), .ZN(n13215) );
  AOI22_X1 U14977 ( .A1(n16734), .A2(n13213), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n16733), .ZN(n13214) );
  OAI21_X1 U14978 ( .B1(n13215), .B2(n16733), .A(n13214), .ZN(P3_U3417) );
  AOI21_X1 U14979 ( .B1(n13217), .B2(n13216), .A(n7632), .ZN(n13225) );
  OAI22_X1 U14980 ( .A1(n16723), .A2(n13219), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13218), .ZN(n13223) );
  OAI22_X1 U14981 ( .A1(n13221), .A2(n15717), .B1(n15716), .B2(n13220), .ZN(
        n13222) );
  AOI211_X1 U14982 ( .C1(n13656), .C2(n16719), .A(n13223), .B(n13222), .ZN(
        n13224) );
  OAI21_X1 U14983 ( .B1(n13225), .B2(n15729), .A(n13224), .ZN(P1_U3236) );
  OAI22_X1 U14984 ( .A1(n14872), .A2(n14397), .B1(n16724), .B2(n13226), .ZN(
        n13227) );
  AOI21_X1 U14985 ( .B1(n13228), .B2(n16724), .A(n13227), .ZN(n13229) );
  INV_X1 U14986 ( .A(n13229), .ZN(P3_U3468) );
  NAND2_X1 U14987 ( .A1(n13240), .A2(n15086), .ZN(n13230) );
  XNOR2_X1 U14988 ( .A(n13347), .B(n13340), .ZN(n13233) );
  OAI22_X1 U14989 ( .A1(n15172), .A2(n15162), .B1(n13284), .B2(n15043), .ZN(
        n13289) );
  AOI21_X1 U14990 ( .B1(n13233), .B2(n15446), .A(n13289), .ZN(n15548) );
  INV_X1 U14991 ( .A(n13234), .ZN(n13235) );
  AOI211_X1 U14992 ( .C1(n15545), .C2(n13235), .A(n7418), .B(n13358), .ZN(
        n15544) );
  AOI22_X1 U14993 ( .A1(n15454), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13288), 
        .B2(n15452), .ZN(n13236) );
  OAI21_X1 U14994 ( .B1(n13348), .B2(n15456), .A(n13236), .ZN(n13244) );
  INV_X1 U14995 ( .A(n13237), .ZN(n13238) );
  OR2_X1 U14996 ( .A1(n13240), .A2(n13284), .ZN(n13241) );
  NAND2_X1 U14997 ( .A1(n13242), .A2(n13241), .ZN(n13341) );
  XNOR2_X1 U14998 ( .A(n13341), .B(n13340), .ZN(n15549) );
  NOR2_X1 U14999 ( .A1(n15549), .A2(n15435), .ZN(n13243) );
  AOI211_X1 U15000 ( .C1(n15544), .C2(n15461), .A(n13244), .B(n13243), .ZN(
        n13245) );
  OAI21_X1 U15001 ( .B1(n15454), .B2(n15548), .A(n13245), .ZN(P2_U3251) );
  XNOR2_X1 U15002 ( .A(n14163), .B(n14402), .ZN(n13248) );
  XNOR2_X1 U15003 ( .A(n13248), .B(n14403), .ZN(n14130) );
  NAND2_X1 U15004 ( .A1(n13246), .A2(n13262), .ZN(n14127) );
  AND2_X1 U15005 ( .A1(n14130), .A2(n14127), .ZN(n13247) );
  INV_X1 U15006 ( .A(n13248), .ZN(n13249) );
  XNOR2_X1 U15007 ( .A(n14163), .B(n13250), .ZN(n13310) );
  XNOR2_X1 U15008 ( .A(n13310), .B(n14133), .ZN(n13308) );
  XNOR2_X1 U15009 ( .A(n13309), .B(n13308), .ZN(n13255) );
  AOI22_X1 U15010 ( .A1(n14218), .A2(n14254), .B1(n7422), .B2(n14403), .ZN(
        n13252) );
  OAI211_X1 U15011 ( .C1(n14282), .C2(n16664), .A(n13252), .B(n13251), .ZN(
        n13253) );
  AOI21_X1 U15012 ( .B1(n13367), .B2(n14287), .A(n13253), .ZN(n13254) );
  OAI21_X1 U15013 ( .B1(n13255), .B2(n14295), .A(n13254), .ZN(P3_U3176) );
  INV_X1 U15014 ( .A(n13703), .ZN(n13258) );
  OAI222_X1 U15015 ( .A1(n13257), .A2(P2_U3088), .B1(n15626), .B2(n13258), 
        .C1(n13256), .C2(n15628), .ZN(P2_U3306) );
  INV_X1 U15016 ( .A(n13849), .ZN(n13586) );
  OAI222_X1 U15017 ( .A1(n16174), .A2(n13704), .B1(n13259), .B2(n13258), .C1(
        n13586), .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U15018 ( .A(n13260), .B(n9085), .ZN(n16648) );
  AOI21_X1 U15019 ( .B1(n13261), .B2(n14396), .A(n14817), .ZN(n13265) );
  OAI22_X1 U15020 ( .A1(n14815), .A2(n16497), .B1(n13262), .B2(n16495), .ZN(
        n13263) );
  AOI21_X1 U15021 ( .B1(n13265), .B2(n13264), .A(n13263), .ZN(n16645) );
  AOI22_X1 U15022 ( .A1(n14821), .A2(n14402), .B1(n16508), .B2(n14134), .ZN(
        n13267) );
  NAND2_X1 U15023 ( .A1(n16517), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n13266) );
  OAI211_X1 U15024 ( .C1(n16645), .C2(n16517), .A(n13267), .B(n13266), .ZN(
        n13268) );
  AOI21_X1 U15025 ( .B1(n14824), .B2(n16648), .A(n13268), .ZN(n13269) );
  INV_X1 U15026 ( .A(n13269), .ZN(P3_U3223) );
  AOI211_X1 U15027 ( .C1(n16523), .C2(n13272), .A(n13271), .B(n13270), .ZN(
        n13276) );
  AOI22_X1 U15028 ( .A1(n13274), .A2(n15536), .B1(P2_REG1_REG_13__SCAN_IN), 
        .B2(n16525), .ZN(n13273) );
  OAI21_X1 U15029 ( .B1(n13276), .B2(n16525), .A(n13273), .ZN(P2_U3512) );
  AOI22_X1 U15030 ( .A1(n13274), .A2(n15599), .B1(P2_REG0_REG_13__SCAN_IN), 
        .B2(n16527), .ZN(n13275) );
  OAI21_X1 U15031 ( .B1(n13276), .B2(n16527), .A(n13275), .ZN(P2_U3469) );
  INV_X1 U15032 ( .A(n13277), .ZN(n13278) );
  OAI22_X1 U15033 ( .A1(n14809), .A2(n14397), .B1(n13278), .B2(n14792), .ZN(
        n13281) );
  NOR2_X1 U15034 ( .A1(n13279), .A2(n16517), .ZN(n13280) );
  AOI211_X1 U15035 ( .C1(n16517), .C2(P3_REG2_REG_9__SCAN_IN), .A(n13281), .B(
        n13280), .ZN(n13282) );
  OAI21_X1 U15036 ( .B1(n14813), .B2(n13283), .A(n13282), .ZN(P3_U3224) );
  NOR3_X1 U15037 ( .A1(n13285), .A2(n13284), .A3(n15067), .ZN(n13286) );
  AOI21_X1 U15038 ( .B1(n13287), .B2(n15070), .A(n13286), .ZN(n13300) );
  XNOR2_X1 U15039 ( .A(n13348), .B(n11679), .ZN(n13394) );
  NOR2_X1 U15040 ( .A1(n13352), .A2(n15232), .ZN(n13392) );
  XNOR2_X1 U15041 ( .A(n13394), .B(n13392), .ZN(n13299) );
  INV_X1 U15042 ( .A(n13288), .ZN(n13292) );
  NAND2_X1 U15043 ( .A1(n15033), .A2(n13289), .ZN(n13290) );
  OAI211_X1 U15044 ( .C1(n15052), .C2(n13292), .A(n13291), .B(n13290), .ZN(
        n13297) );
  AND2_X1 U15045 ( .A1(n13299), .A2(n13293), .ZN(n13294) );
  NOR2_X1 U15046 ( .A1(n13395), .A2(n15077), .ZN(n13296) );
  AOI211_X1 U15047 ( .C1(n15545), .C2(n15080), .A(n13297), .B(n13296), .ZN(
        n13298) );
  OAI21_X1 U15048 ( .B1(n13300), .B2(n13299), .A(n13298), .ZN(P2_U3187) );
  INV_X1 U15049 ( .A(n13301), .ZN(n13302) );
  OAI222_X1 U15050 ( .A1(P3_U3151), .A2(n13304), .B1(n14959), .B2(n13303), 
        .C1(n14968), .C2(n13302), .ZN(P3_U3270) );
  INV_X1 U15051 ( .A(n13305), .ZN(n13306) );
  OAI222_X1 U15052 ( .A1(P3_U3151), .A2(n9393), .B1(n14959), .B2(n13307), .C1(
        n14968), .C2(n13306), .ZN(P3_U3271) );
  INV_X1 U15053 ( .A(n13310), .ZN(n13311) );
  NAND2_X1 U15054 ( .A1(n13311), .A2(n14133), .ZN(n13312) );
  NAND2_X1 U15055 ( .A1(n13313), .A2(n13312), .ZN(n13525) );
  XNOR2_X1 U15056 ( .A(n14163), .B(n16673), .ZN(n13527) );
  XNOR2_X1 U15057 ( .A(n13527), .B(n13526), .ZN(n13314) );
  XNOR2_X1 U15058 ( .A(n13525), .B(n13314), .ZN(n13321) );
  AOI21_X1 U15059 ( .B1(n14218), .B2(n14416), .A(n13315), .ZN(n13319) );
  NAND2_X1 U15060 ( .A1(n14287), .A2(n14820), .ZN(n13318) );
  NAND2_X1 U15061 ( .A1(n14292), .A2(n16673), .ZN(n13317) );
  NAND2_X1 U15062 ( .A1(n7422), .A2(n14133), .ZN(n13316) );
  NAND4_X1 U15063 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13320) );
  AOI21_X1 U15064 ( .B1(n13321), .B2(n14273), .A(n13320), .ZN(n13322) );
  INV_X1 U15065 ( .A(n13322), .ZN(P3_U3164) );
  INV_X1 U15066 ( .A(n13659), .ZN(n16685) );
  OAI211_X1 U15067 ( .C1(n13325), .C2(n13324), .A(n13323), .B(n16714), .ZN(
        n13334) );
  INV_X1 U15068 ( .A(n13326), .ZN(n13332) );
  INV_X1 U15069 ( .A(n13327), .ZN(n13330) );
  OAI22_X1 U15070 ( .A1(n15643), .A2(n15717), .B1(n15716), .B2(n13328), .ZN(
        n13329) );
  AOI211_X1 U15071 ( .C1(n13332), .C2(n13331), .A(n13330), .B(n13329), .ZN(
        n13333) );
  OAI211_X1 U15072 ( .C1(n16685), .C2(n15712), .A(n13334), .B(n13333), .ZN(
        P1_U3224) );
  NAND2_X1 U15073 ( .A1(n13729), .A2(n13335), .ZN(n13336) );
  OAI211_X1 U15074 ( .C1(n13730), .C2(n16174), .A(n13336), .B(n13908), .ZN(
        P1_U3332) );
  NAND2_X1 U15075 ( .A1(n13729), .A2(n15617), .ZN(n13338) );
  OAI211_X1 U15076 ( .C1(n13339), .C2(n15628), .A(n13338), .B(n13337), .ZN(
        P2_U3304) );
  NAND2_X1 U15077 ( .A1(n13341), .A2(n13340), .ZN(n13343) );
  OR2_X1 U15078 ( .A1(n13348), .A2(n13352), .ZN(n13342) );
  INV_X1 U15079 ( .A(n13350), .ZN(n15194) );
  NAND2_X1 U15080 ( .A1(n13344), .A2(n15194), .ZN(n13345) );
  NAND2_X1 U15081 ( .A1(n15174), .A2(n13345), .ZN(n13489) );
  INV_X1 U15082 ( .A(n13489), .ZN(n13364) );
  OR2_X1 U15083 ( .A1(n13348), .A2(n15085), .ZN(n13346) );
  NAND2_X1 U15084 ( .A1(n13348), .A2(n15085), .ZN(n13349) );
  XNOR2_X1 U15085 ( .A(n15195), .B(n13350), .ZN(n13351) );
  NAND2_X1 U15086 ( .A1(n13351), .A2(n15446), .ZN(n13356) );
  INV_X1 U15087 ( .A(n15443), .ZN(n15394) );
  NAND2_X1 U15088 ( .A1(n15175), .A2(n15073), .ZN(n13354) );
  OR2_X1 U15089 ( .A1(n13352), .A2(n15043), .ZN(n13353) );
  NAND2_X1 U15090 ( .A1(n13354), .A2(n13353), .ZN(n13456) );
  AOI21_X1 U15091 ( .B1(n13489), .B2(n15394), .A(n13456), .ZN(n13355) );
  NAND2_X1 U15092 ( .A1(n13356), .A2(n13355), .ZN(n13493) );
  NAND2_X1 U15093 ( .A1(n13493), .A2(n15429), .ZN(n13363) );
  OAI22_X1 U15094 ( .A1(n15429), .A2(n13357), .B1(n13458), .B2(n15427), .ZN(
        n13361) );
  OAI21_X1 U15095 ( .B1(n13358), .B2(n15197), .A(n15232), .ZN(n13359) );
  OR2_X1 U15096 ( .A1(n15448), .A2(n13359), .ZN(n13490) );
  NOR2_X1 U15097 ( .A1(n13490), .A2(n15318), .ZN(n13360) );
  AOI211_X1 U15098 ( .C1(n15316), .C2(n13463), .A(n13361), .B(n13360), .ZN(
        n13362) );
  OAI211_X1 U15099 ( .C1(n13364), .C2(n15458), .A(n13363), .B(n13362), .ZN(
        P2_U3250) );
  XNOR2_X1 U15100 ( .A(n13365), .B(n14404), .ZN(n13366) );
  AOI222_X1 U15101 ( .A1(n14403), .A2(n14777), .B1(n16500), .B2(n13366), .C1(
        n14254), .C2(n14779), .ZN(n16662) );
  INV_X1 U15102 ( .A(n13367), .ZN(n13368) );
  OAI22_X1 U15103 ( .A1(n14809), .A2(n16664), .B1(n13368), .B2(n14792), .ZN(
        n13369) );
  AOI21_X1 U15104 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n16517), .A(n13369), 
        .ZN(n13372) );
  XNOR2_X1 U15105 ( .A(n13370), .B(n14404), .ZN(n16667) );
  NAND2_X1 U15106 ( .A1(n16667), .A2(n14824), .ZN(n13371) );
  OAI211_X1 U15107 ( .C1(n16662), .C2(n16517), .A(n13372), .B(n13371), .ZN(
        P3_U3222) );
  NAND2_X1 U15108 ( .A1(n13378), .A2(n13373), .ZN(n13374) );
  NAND2_X1 U15109 ( .A1(n13375), .A2(n13374), .ZN(n13376) );
  XOR2_X1 U15110 ( .A(n13376), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13383) );
  NAND2_X1 U15111 ( .A1(n13378), .A2(n13377), .ZN(n13380) );
  NAND2_X1 U15112 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  XNOR2_X1 U15113 ( .A(n13382), .B(n13381), .ZN(n13384) );
  AOI22_X1 U15114 ( .A1(n13383), .A2(n15797), .B1(n15807), .B2(n13384), .ZN(
        n13389) );
  INV_X1 U15115 ( .A(n13383), .ZN(n13386) );
  NOR2_X1 U15116 ( .A1(n13384), .A2(n16297), .ZN(n13385) );
  AOI211_X1 U15117 ( .C1(n13387), .C2(n13386), .A(n16294), .B(n13385), .ZN(
        n13388) );
  MUX2_X1 U15118 ( .A(n13389), .B(n13388), .S(n10650), .Z(n13390) );
  NAND2_X1 U15119 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15656)
         );
  OAI211_X1 U15120 ( .C1(n13391), .C2(n16301), .A(n13390), .B(n15656), .ZN(
        P1_U3262) );
  INV_X1 U15121 ( .A(n13392), .ZN(n13393) );
  XNOR2_X1 U15122 ( .A(n15197), .B(n7695), .ZN(n13396) );
  NOR2_X1 U15123 ( .A1(n15172), .A2(n15232), .ZN(n13397) );
  NAND2_X1 U15124 ( .A1(n13396), .A2(n13397), .ZN(n13402) );
  INV_X1 U15125 ( .A(n13396), .ZN(n13400) );
  INV_X1 U15126 ( .A(n13397), .ZN(n13398) );
  NAND2_X1 U15127 ( .A1(n13400), .A2(n13398), .ZN(n13399) );
  NAND2_X1 U15128 ( .A1(n13402), .A2(n13399), .ZN(n13459) );
  NOR3_X1 U15129 ( .A1(n13400), .A2(n15172), .A3(n15067), .ZN(n13401) );
  AOI21_X1 U15130 ( .B1(n7590), .B2(n15070), .A(n13401), .ZN(n13412) );
  XNOR2_X1 U15131 ( .A(n15539), .B(n11679), .ZN(n13474) );
  NAND2_X1 U15132 ( .A1(n15175), .A2(n7418), .ZN(n13465) );
  XNOR2_X1 U15133 ( .A(n13474), .B(n13465), .ZN(n13411) );
  AND2_X1 U15134 ( .A1(n13411), .A2(n13402), .ZN(n13403) );
  INV_X1 U15135 ( .A(n13468), .ZN(n13477) );
  NAND2_X1 U15136 ( .A1(n15177), .A2(n15073), .ZN(n13405) );
  INV_X1 U15137 ( .A(n15172), .ZN(n15196) );
  NAND2_X1 U15138 ( .A1(n15196), .A2(n15225), .ZN(n13404) );
  NAND2_X1 U15139 ( .A1(n13405), .A2(n13404), .ZN(n15445) );
  NOR2_X1 U15140 ( .A1(n13406), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16242) );
  AOI21_X1 U15141 ( .B1(n15033), .B2(n15445), .A(n16242), .ZN(n13408) );
  NAND2_X1 U15142 ( .A1(n15074), .A2(n15453), .ZN(n13407) );
  OAI211_X1 U15143 ( .C1(n15457), .C2(n15066), .A(n13408), .B(n13407), .ZN(
        n13409) );
  AOI21_X1 U15144 ( .B1(n13477), .B2(n15070), .A(n13409), .ZN(n13410) );
  OAI21_X1 U15145 ( .B1(n13412), .B2(n13411), .A(n13410), .ZN(P2_U3198) );
  NOR2_X1 U15146 ( .A1(n16697), .A2(n15745), .ZN(n13413) );
  XNOR2_X1 U15147 ( .A(n16137), .B(n15744), .ZN(n13870) );
  OR2_X1 U15148 ( .A1(n13415), .A2(n13420), .ZN(n13416) );
  NAND2_X1 U15149 ( .A1(n13500), .A2(n13416), .ZN(n16141) );
  INV_X1 U15150 ( .A(n15743), .ZN(n16030) );
  AOI21_X1 U15151 ( .B1(n13420), .B2(n13419), .A(n13504), .ZN(n13421) );
  OAI222_X1 U15152 ( .A1(n16031), .A2(n15643), .B1(n16029), .B2(n16030), .C1(
        n16702), .C2(n13421), .ZN(n16136) );
  NAND2_X1 U15153 ( .A1(n16136), .A2(n16014), .ZN(n13429) );
  INV_X1 U15154 ( .A(n13422), .ZN(n13424) );
  INV_X1 U15155 ( .A(n16137), .ZN(n13425) );
  INV_X1 U15156 ( .A(n13508), .ZN(n13423) );
  AOI21_X1 U15157 ( .B1(n16137), .B2(n13424), .A(n13423), .ZN(n16138) );
  NOR2_X1 U15158 ( .A1(n13425), .A2(n16587), .ZN(n13427) );
  OAI22_X1 U15159 ( .A1(n16014), .A2(n11876), .B1(n15642), .B2(n16036), .ZN(
        n13426) );
  AOI211_X1 U15160 ( .C1(n16138), .C2(n15987), .A(n13427), .B(n13426), .ZN(
        n13428) );
  OAI211_X1 U15161 ( .C1(n16141), .C2(n16040), .A(n13429), .B(n13428), .ZN(
        P1_U3279) );
  INV_X1 U15162 ( .A(n13430), .ZN(n13433) );
  INV_X1 U15163 ( .A(n13431), .ZN(n13432) );
  OAI222_X1 U15164 ( .A1(n15628), .A2(n13434), .B1(n15626), .B2(n13433), .C1(
        P2_U3088), .C2(n13432), .ZN(P2_U3305) );
  NOR2_X1 U15165 ( .A1(n13494), .A2(n13437), .ZN(n15133) );
  AOI211_X1 U15166 ( .C1(n13437), .C2(n13494), .A(n15133), .B(n16264), .ZN(
        n13446) );
  NOR2_X1 U15167 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13438), .ZN(n13439) );
  AOI21_X1 U15168 ( .B1(n16270), .B2(n15117), .A(n13439), .ZN(n13444) );
  NOR2_X1 U15169 ( .A1(n13441), .A2(n13440), .ZN(n15116) );
  XNOR2_X1 U15170 ( .A(n15131), .B(n15116), .ZN(n13442) );
  NAND2_X1 U15171 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13442), .ZN(n15118) );
  OAI211_X1 U15172 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n13442), .A(n16257), 
        .B(n15118), .ZN(n13443) );
  OAI211_X1 U15173 ( .C1(n16278), .C2(n8177), .A(n13444), .B(n13443), .ZN(
        n13445) );
  OR2_X1 U15174 ( .A1(n13446), .A2(n13445), .ZN(P2_U3229) );
  AOI21_X1 U15175 ( .B1(n13447), .B2(n14483), .A(n14817), .ZN(n13450) );
  OAI22_X1 U15176 ( .A1(n13526), .A2(n16495), .B1(n14256), .B2(n16497), .ZN(
        n13448) );
  AOI21_X1 U15177 ( .B1(n13450), .B2(n13449), .A(n13448), .ZN(n14897) );
  INV_X1 U15178 ( .A(n14898), .ZN(n14258) );
  INV_X1 U15179 ( .A(n14259), .ZN(n13451) );
  OAI22_X1 U15180 ( .A1(n14819), .A2(n14522), .B1(n13451), .B2(n14792), .ZN(
        n13452) );
  AOI21_X1 U15181 ( .B1(n14258), .B2(n14821), .A(n13452), .ZN(n13455) );
  XNOR2_X1 U15182 ( .A(n13453), .B(n14483), .ZN(n14895) );
  NAND2_X1 U15183 ( .A1(n14895), .A2(n14824), .ZN(n13454) );
  OAI211_X1 U15184 ( .C1(n14897), .C2(n16517), .A(n13455), .B(n13454), .ZN(
        P3_U3220) );
  AOI22_X1 U15185 ( .A1(n15033), .A2(n13456), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13457) );
  OAI21_X1 U15186 ( .B1(n15052), .B2(n13458), .A(n13457), .ZN(n13462) );
  AOI211_X1 U15187 ( .C1(n13460), .C2(n13459), .A(n15077), .B(n7590), .ZN(
        n13461) );
  AOI211_X1 U15188 ( .C1(n13463), .C2(n15080), .A(n13462), .B(n13461), .ZN(
        n13464) );
  INV_X1 U15189 ( .A(n13464), .ZN(P2_U3213) );
  INV_X1 U15190 ( .A(n13474), .ZN(n13466) );
  NAND2_X1 U15191 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  XNOR2_X1 U15192 ( .A(n15598), .B(n11679), .ZN(n14067) );
  NAND2_X1 U15193 ( .A1(n15177), .A2(n7418), .ZN(n14068) );
  XNOR2_X1 U15194 ( .A(n14067), .B(n14068), .ZN(n13475) );
  OR2_X1 U15195 ( .A1(n15203), .A2(n15162), .ZN(n13471) );
  NAND2_X1 U15196 ( .A1(n15175), .A2(n15225), .ZN(n13470) );
  AND2_X1 U15197 ( .A1(n13471), .A2(n13470), .ZN(n15422) );
  INV_X1 U15198 ( .A(n15422), .ZN(n13472) );
  AOI22_X1 U15199 ( .A1(n13472), .A2(n15033), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13473) );
  OAI21_X1 U15200 ( .B1(n15428), .B2(n15052), .A(n13473), .ZN(n13479) );
  INV_X1 U15201 ( .A(n15067), .ZN(n15050) );
  AOI22_X1 U15202 ( .A1(n13474), .A2(n15070), .B1(n15050), .B2(n15175), .ZN(
        n13476) );
  NOR3_X1 U15203 ( .A1(n13477), .A2(n13476), .A3(n13475), .ZN(n13478) );
  AOI211_X1 U15204 ( .C1(n15598), .C2(n15080), .A(n13479), .B(n13478), .ZN(
        n13480) );
  OAI21_X1 U15205 ( .B1(n15077), .B2(n14071), .A(n13480), .ZN(P2_U3200) );
  OAI211_X1 U15206 ( .C1(n13483), .C2(n13482), .A(n13481), .B(n16714), .ZN(
        n13487) );
  AND2_X1 U15207 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n15802) );
  NOR2_X1 U15208 ( .A1(n16723), .A2(n13484), .ZN(n13485) );
  AOI211_X1 U15209 ( .C1(n16716), .C2(n16695), .A(n15802), .B(n13485), .ZN(
        n13486) );
  OAI211_X1 U15210 ( .C1(n13488), .C2(n15712), .A(n13487), .B(n13486), .ZN(
        P1_U3234) );
  NAND2_X1 U15211 ( .A1(n13489), .A2(n11714), .ZN(n13491) );
  NAND2_X1 U15212 ( .A1(n13491), .A2(n13490), .ZN(n13492) );
  NOR2_X1 U15213 ( .A1(n13493), .A2(n13492), .ZN(n13496) );
  MUX2_X1 U15214 ( .A(n13494), .B(n13496), .S(n16526), .Z(n13495) );
  OAI21_X1 U15215 ( .B1(n15197), .B2(n15530), .A(n13495), .ZN(P2_U3514) );
  MUX2_X1 U15216 ( .A(n13497), .B(n13496), .S(n16529), .Z(n13498) );
  OAI21_X1 U15217 ( .B1(n15197), .B2(n15594), .A(n13498), .ZN(P2_U3475) );
  XNOR2_X1 U15218 ( .A(n16718), .B(n15743), .ZN(n13872) );
  NAND2_X1 U15219 ( .A1(n16137), .A2(n15744), .ZN(n13499) );
  INV_X1 U15220 ( .A(n14041), .ZN(n13502) );
  AOI21_X1 U15221 ( .B1(n13872), .B2(n13503), .A(n13502), .ZN(n16135) );
  INV_X1 U15222 ( .A(n15744), .ZN(n13505) );
  AOI21_X1 U15223 ( .B1(n7609), .B2(n13501), .A(n16702), .ZN(n13506) );
  INV_X1 U15224 ( .A(n15742), .ZN(n14042) );
  OAI22_X1 U15225 ( .A1(n14042), .A2(n16029), .B1(n13505), .B2(n16031), .ZN(
        n16717) );
  AOI21_X1 U15226 ( .B1(n13506), .B2(n14024), .A(n16717), .ZN(n16134) );
  OAI21_X1 U15227 ( .B1(n16722), .B2(n16036), .A(n16134), .ZN(n13507) );
  NAND2_X1 U15228 ( .A1(n13507), .A2(n16014), .ZN(n13512) );
  AOI211_X1 U15229 ( .C1(n16718), .C2(n13508), .A(n16686), .B(n7588), .ZN(
        n16132) );
  OAI22_X1 U15230 ( .A1(n8188), .A2(n16587), .B1(n16014), .B2(n13509), .ZN(
        n13510) );
  AOI21_X1 U15231 ( .B1(n16132), .B2(n16636), .A(n13510), .ZN(n13511) );
  OAI211_X1 U15232 ( .C1(n16135), .C2(n16040), .A(n13512), .B(n13511), .ZN(
        P1_U3278) );
  INV_X1 U15233 ( .A(n13749), .ZN(n13515) );
  OAI222_X1 U15234 ( .A1(n15628), .A2(n13514), .B1(n15626), .B2(n13515), .C1(
        P2_U3088), .C2(n13513), .ZN(P2_U3303) );
  OAI222_X1 U15235 ( .A1(n13516), .A2(P1_U3086), .B1(n16174), .B2(n13750), 
        .C1(n13515), .C2(n16178), .ZN(P1_U3331) );
  XNOR2_X1 U15236 ( .A(n13517), .B(n14484), .ZN(n14893) );
  OAI211_X1 U15237 ( .C1(n13519), .C2(n14484), .A(n13518), .B(n16500), .ZN(
        n13521) );
  AOI22_X1 U15238 ( .A1(n14777), .A2(n14416), .B1(n14205), .B2(n14779), .ZN(
        n13520) );
  NAND2_X1 U15239 ( .A1(n13521), .A2(n13520), .ZN(n14890) );
  AOI22_X1 U15240 ( .A1(n16517), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n16508), 
        .B2(n13536), .ZN(n13522) );
  OAI21_X1 U15241 ( .B1(n14889), .B2(n14809), .A(n13522), .ZN(n13523) );
  AOI21_X1 U15242 ( .B1(n14890), .B2(n14819), .A(n13523), .ZN(n13524) );
  OAI21_X1 U15243 ( .B1(n14813), .B2(n14893), .A(n13524), .ZN(P3_U3219) );
  INV_X1 U15244 ( .A(n13525), .ZN(n13528) );
  XNOR2_X1 U15245 ( .A(n14898), .B(n14163), .ZN(n13529) );
  XNOR2_X1 U15246 ( .A(n13529), .B(n14816), .ZN(n14252) );
  NAND2_X1 U15247 ( .A1(n14253), .A2(n14252), .ZN(n14251) );
  NAND2_X1 U15248 ( .A1(n13529), .A2(n14416), .ZN(n13530) );
  XNOR2_X1 U15249 ( .A(n14889), .B(n14163), .ZN(n13549) );
  XNOR2_X1 U15250 ( .A(n13549), .B(n14256), .ZN(n13531) );
  OAI211_X1 U15251 ( .C1(n13532), .C2(n13531), .A(n13551), .B(n14273), .ZN(
        n13538) );
  NAND2_X1 U15252 ( .A1(n7422), .A2(n14416), .ZN(n13534) );
  OR2_X1 U15253 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13533), .ZN(n14539) );
  OAI211_X1 U15254 ( .C1(n14290), .C2(n14805), .A(n13534), .B(n14539), .ZN(
        n13535) );
  AOI21_X1 U15255 ( .B1(n13536), .B2(n14287), .A(n13535), .ZN(n13537) );
  OAI211_X1 U15256 ( .C1(n14282), .C2(n14889), .A(n13538), .B(n13537), .ZN(
        P3_U3155) );
  XNOR2_X1 U15257 ( .A(n13539), .B(n13542), .ZN(n14888) );
  OAI211_X1 U15258 ( .C1(n13542), .C2(n13541), .A(n13540), .B(n16500), .ZN(
        n13544) );
  AOI22_X1 U15259 ( .A1(n14777), .A2(n13557), .B1(n14227), .B2(n14779), .ZN(
        n13543) );
  NAND2_X1 U15260 ( .A1(n13544), .A2(n13543), .ZN(n14885) );
  INV_X1 U15261 ( .A(n14886), .ZN(n13546) );
  AOI22_X1 U15262 ( .A1(n16517), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n16508), 
        .B2(n13556), .ZN(n13545) );
  OAI21_X1 U15263 ( .B1(n13546), .B2(n14809), .A(n13545), .ZN(n13547) );
  AOI21_X1 U15264 ( .B1(n14885), .B2(n14819), .A(n13547), .ZN(n13548) );
  OAI21_X1 U15265 ( .B1(n14888), .B2(n14813), .A(n13548), .ZN(P3_U3218) );
  NAND2_X1 U15266 ( .A1(n13549), .A2(n13557), .ZN(n13550) );
  XNOR2_X1 U15267 ( .A(n14886), .B(n14163), .ZN(n13553) );
  INV_X1 U15268 ( .A(n13553), .ZN(n13552) );
  NAND2_X1 U15269 ( .A1(n13552), .A2(n14205), .ZN(n13922) );
  NAND2_X1 U15270 ( .A1(n13553), .A2(n14805), .ZN(n13920) );
  NAND2_X1 U15271 ( .A1(n13922), .A2(n13920), .ZN(n13554) );
  XNOR2_X1 U15272 ( .A(n13921), .B(n13554), .ZN(n13563) );
  NAND2_X1 U15273 ( .A1(n14886), .A2(n14292), .ZN(n13561) );
  AOI21_X1 U15274 ( .B1(n14218), .B2(n14227), .A(n13555), .ZN(n13560) );
  NAND2_X1 U15275 ( .A1(n14287), .A2(n13556), .ZN(n13559) );
  NAND2_X1 U15276 ( .A1(n7422), .A2(n13557), .ZN(n13558) );
  NAND4_X1 U15277 ( .A1(n13561), .A2(n13560), .A3(n13559), .A4(n13558), .ZN(
        n13562) );
  AOI21_X1 U15278 ( .B1(n13563), .B2(n14273), .A(n13562), .ZN(n13564) );
  INV_X1 U15279 ( .A(n13564), .ZN(P3_U3181) );
  INV_X1 U15280 ( .A(n13567), .ZN(n15611) );
  OAI222_X1 U15281 ( .A1(n16174), .A2(n14300), .B1(P1_U3086), .B2(n13565), 
        .C1(n16178), .C2(n15611), .ZN(P1_U3326) );
  INV_X1 U15282 ( .A(n15613), .ZN(n13566) );
  OAI222_X1 U15283 ( .A1(n16174), .A2(n13802), .B1(n16178), .B2(n13566), .C1(
        n10784), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U15284 ( .A1(n13567), .A2(n13838), .ZN(n13569) );
  OR2_X1 U15285 ( .A1(n10937), .A2(n14300), .ZN(n13568) );
  NAND2_X1 U15286 ( .A1(n13829), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n13576) );
  INV_X1 U15287 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n13570) );
  OR2_X1 U15288 ( .A1(n10679), .A2(n13570), .ZN(n13575) );
  INV_X1 U15289 ( .A(n13571), .ZN(n13714) );
  NAND2_X1 U15290 ( .A1(n13714), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n13713) );
  NAND2_X1 U15291 ( .A1(n13734), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U15292 ( .A1(n13792), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n13791) );
  INV_X1 U15293 ( .A(n13791), .ZN(n13808) );
  NAND2_X1 U15294 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n13808), .ZN(n14034) );
  OR2_X1 U15295 ( .A1(n10700), .A2(n14034), .ZN(n13574) );
  INV_X1 U15296 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n13572) );
  OR2_X1 U15297 ( .A1(n13810), .A2(n13572), .ZN(n13573) );
  NAND2_X1 U15298 ( .A1(n16033), .A2(n13839), .ZN(n13577) );
  NAND2_X1 U15299 ( .A1(n13578), .A2(n13577), .ZN(n13585) );
  MUX2_X1 U15300 ( .A(n13849), .B(n13850), .S(n13585), .Z(n13579) );
  MUX2_X1 U15301 ( .A(n16048), .B(n15827), .S(n13771), .Z(n13821) );
  INV_X1 U15302 ( .A(n13821), .ZN(n13825) );
  AOI21_X1 U15303 ( .B1(n13581), .B2(n13836), .A(n13580), .ZN(n13605) );
  AOI21_X1 U15304 ( .B1(n15756), .B2(n13771), .A(n8105), .ZN(n13604) );
  NAND2_X1 U15305 ( .A1(n13584), .A2(n13583), .ZN(n13592) );
  MUX2_X1 U15306 ( .A(n13828), .B(n13586), .S(n13585), .Z(n13588) );
  NAND2_X1 U15307 ( .A1(n16474), .A2(n13588), .ZN(n13591) );
  AND2_X1 U15308 ( .A1(n16474), .A2(n13587), .ZN(n13589) );
  OAI21_X1 U15309 ( .B1(n13589), .B2(n13588), .A(n8099), .ZN(n13590) );
  OAI211_X1 U15310 ( .C1(n8099), .C2(n13592), .A(n13591), .B(n13590), .ZN(
        n13598) );
  INV_X1 U15311 ( .A(n13598), .ZN(n13595) );
  NAND3_X1 U15312 ( .A1(n13595), .A2(n13594), .A3(n13855), .ZN(n13603) );
  NAND2_X1 U15313 ( .A1(n13598), .A2(n13597), .ZN(n13601) );
  MUX2_X1 U15314 ( .A(n15757), .B(n13599), .S(n13836), .Z(n13600) );
  NAND3_X1 U15315 ( .A1(n13601), .A2(n13855), .A3(n13600), .ZN(n13602) );
  OAI211_X1 U15316 ( .C1(n13605), .C2(n13604), .A(n13603), .B(n13602), .ZN(
        n13606) );
  NAND3_X1 U15317 ( .A1(n13606), .A2(n13856), .A3(n13616), .ZN(n13618) );
  NAND2_X1 U15318 ( .A1(n13607), .A2(n13836), .ZN(n13610) );
  NAND3_X1 U15319 ( .A1(n15755), .A2(n13771), .A3(n13608), .ZN(n13609) );
  OAI21_X1 U15320 ( .B1(n15755), .B2(n13610), .A(n13609), .ZN(n13615) );
  OAI21_X1 U15321 ( .B1(n15754), .B2(n13771), .A(n13611), .ZN(n13614) );
  NAND2_X1 U15322 ( .A1(n15754), .A2(n13771), .ZN(n13612) );
  NAND2_X1 U15323 ( .A1(n13612), .A2(n16546), .ZN(n13613) );
  AOI22_X1 U15324 ( .A1(n13616), .A2(n13615), .B1(n13614), .B2(n13613), .ZN(
        n13617) );
  NAND2_X1 U15325 ( .A1(n13618), .A2(n13617), .ZN(n13622) );
  MUX2_X1 U15326 ( .A(n13619), .B(n15753), .S(n13771), .Z(n13623) );
  NAND2_X1 U15327 ( .A1(n13622), .A2(n13623), .ZN(n13621) );
  MUX2_X1 U15328 ( .A(n13619), .B(n15753), .S(n7421), .Z(n13620) );
  NAND2_X1 U15329 ( .A1(n13621), .A2(n13620), .ZN(n13627) );
  INV_X1 U15330 ( .A(n13622), .ZN(n13625) );
  INV_X1 U15331 ( .A(n13623), .ZN(n13624) );
  NAND2_X1 U15332 ( .A1(n13625), .A2(n13624), .ZN(n13626) );
  MUX2_X1 U15333 ( .A(n13628), .B(n15752), .S(n7421), .Z(n13631) );
  MUX2_X1 U15334 ( .A(n15752), .B(n13628), .S(n7421), .Z(n13629) );
  INV_X1 U15335 ( .A(n13631), .ZN(n13632) );
  MUX2_X1 U15336 ( .A(n13633), .B(n15751), .S(n13771), .Z(n13635) );
  MUX2_X1 U15337 ( .A(n13633), .B(n15751), .S(n7421), .Z(n13634) );
  INV_X1 U15338 ( .A(n13635), .ZN(n13636) );
  MUX2_X1 U15339 ( .A(n15750), .B(n13637), .S(n13771), .Z(n13641) );
  NAND2_X1 U15340 ( .A1(n13640), .A2(n13641), .ZN(n13639) );
  MUX2_X1 U15341 ( .A(n15750), .B(n13637), .S(n7421), .Z(n13638) );
  NAND2_X1 U15342 ( .A1(n13639), .A2(n13638), .ZN(n13645) );
  INV_X1 U15343 ( .A(n13640), .ZN(n13643) );
  INV_X1 U15344 ( .A(n13641), .ZN(n13642) );
  NAND2_X1 U15345 ( .A1(n13643), .A2(n13642), .ZN(n13644) );
  MUX2_X1 U15346 ( .A(n15749), .B(n16633), .S(n7421), .Z(n13648) );
  MUX2_X1 U15347 ( .A(n15749), .B(n16633), .S(n13771), .Z(n13646) );
  MUX2_X1 U15348 ( .A(n15748), .B(n13649), .S(n13771), .Z(n13652) );
  MUX2_X1 U15349 ( .A(n15748), .B(n13649), .S(n7421), .Z(n13650) );
  NAND2_X1 U15350 ( .A1(n13651), .A2(n13650), .ZN(n13655) );
  INV_X1 U15351 ( .A(n13652), .ZN(n13653) );
  MUX2_X1 U15352 ( .A(n15747), .B(n13656), .S(n7421), .Z(n13658) );
  MUX2_X1 U15353 ( .A(n15747), .B(n13656), .S(n13771), .Z(n13657) );
  MUX2_X1 U15354 ( .A(n15746), .B(n13659), .S(n13771), .Z(n13662) );
  MUX2_X1 U15355 ( .A(n15746), .B(n13659), .S(n7421), .Z(n13660) );
  INV_X1 U15356 ( .A(n13662), .ZN(n13663) );
  MUX2_X1 U15357 ( .A(n15745), .B(n16697), .S(n7421), .Z(n13667) );
  MUX2_X1 U15358 ( .A(n16697), .B(n15745), .S(n7421), .Z(n13664) );
  NAND2_X1 U15359 ( .A1(n13665), .A2(n13664), .ZN(n13671) );
  INV_X1 U15360 ( .A(n13666), .ZN(n13669) );
  INV_X1 U15361 ( .A(n13667), .ZN(n13668) );
  NAND2_X1 U15362 ( .A1(n13669), .A2(n13668), .ZN(n13670) );
  MUX2_X1 U15363 ( .A(n15744), .B(n16137), .S(n13771), .Z(n13673) );
  MUX2_X1 U15364 ( .A(n15744), .B(n16137), .S(n7421), .Z(n13672) );
  MUX2_X1 U15365 ( .A(n15743), .B(n16718), .S(n7421), .Z(n13676) );
  MUX2_X1 U15366 ( .A(n15743), .B(n16718), .S(n13771), .Z(n13675) );
  INV_X1 U15367 ( .A(n13676), .ZN(n13677) );
  MUX2_X1 U15368 ( .A(n15742), .B(n16129), .S(n13771), .Z(n13680) );
  MUX2_X1 U15369 ( .A(n16129), .B(n15742), .S(n13771), .Z(n13678) );
  MUX2_X1 U15370 ( .A(n15741), .B(n16123), .S(n7421), .Z(n13684) );
  NAND2_X1 U15371 ( .A1(n13683), .A2(n13684), .ZN(n13682) );
  MUX2_X1 U15372 ( .A(n15741), .B(n16123), .S(n13771), .Z(n13681) );
  NAND2_X1 U15373 ( .A1(n13682), .A2(n13681), .ZN(n13688) );
  INV_X1 U15374 ( .A(n13684), .ZN(n13685) );
  NAND2_X1 U15375 ( .A1(n13686), .A2(n13685), .ZN(n13687) );
  MUX2_X1 U15376 ( .A(n16118), .B(n15740), .S(n7421), .Z(n13690) );
  MUX2_X1 U15377 ( .A(n16118), .B(n15740), .S(n13771), .Z(n13689) );
  MUX2_X1 U15378 ( .A(n15954), .B(n16111), .S(n7421), .Z(n13695) );
  NAND2_X1 U15379 ( .A1(n13694), .A2(n13695), .ZN(n13693) );
  MUX2_X1 U15380 ( .A(n16111), .B(n15954), .S(n7421), .Z(n13692) );
  NAND2_X1 U15381 ( .A1(n13693), .A2(n13692), .ZN(n13699) );
  INV_X1 U15382 ( .A(n13695), .ZN(n13696) );
  NAND2_X1 U15383 ( .A1(n13697), .A2(n13696), .ZN(n13698) );
  MUX2_X1 U15384 ( .A(n15739), .B(n15958), .S(n13771), .Z(n13701) );
  MUX2_X1 U15385 ( .A(n15739), .B(n15958), .S(n7421), .Z(n13700) );
  INV_X1 U15386 ( .A(n13701), .ZN(n13702) );
  NAND2_X1 U15387 ( .A1(n13703), .A2(n13838), .ZN(n13706) );
  OR2_X1 U15388 ( .A1(n10937), .A2(n13704), .ZN(n13705) );
  MUX2_X1 U15389 ( .A(n15957), .B(n15937), .S(n7421), .Z(n13708) );
  MUX2_X1 U15390 ( .A(n15937), .B(n15957), .S(n7421), .Z(n13707) );
  INV_X1 U15391 ( .A(n13708), .ZN(n13709) );
  XNOR2_X1 U15392 ( .A(n13711), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n16181) );
  NAND2_X1 U15393 ( .A1(n13805), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n13719) );
  INV_X1 U15394 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15923) );
  OR2_X1 U15395 ( .A1(n13807), .A2(n15923), .ZN(n13718) );
  OAI21_X1 U15396 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n13714), .A(n13713), 
        .ZN(n15922) );
  OR2_X1 U15397 ( .A1(n10700), .A2(n15922), .ZN(n13717) );
  INV_X1 U15398 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n13715) );
  OR2_X1 U15399 ( .A1(n13810), .A2(n13715), .ZN(n13716) );
  MUX2_X1 U15400 ( .A(n15921), .B(n15665), .S(n7421), .Z(n13725) );
  INV_X1 U15401 ( .A(n13725), .ZN(n13720) );
  NAND2_X1 U15402 ( .A1(n13724), .A2(n13720), .ZN(n13723) );
  MUX2_X1 U15403 ( .A(n15665), .B(n15921), .S(n7421), .Z(n13721) );
  INV_X1 U15404 ( .A(n13721), .ZN(n13722) );
  NAND2_X1 U15405 ( .A1(n13723), .A2(n13722), .ZN(n13728) );
  INV_X1 U15406 ( .A(n13724), .ZN(n13726) );
  NAND2_X1 U15407 ( .A1(n13726), .A2(n13725), .ZN(n13727) );
  NAND2_X1 U15408 ( .A1(n13729), .A2(n13838), .ZN(n13732) );
  OR2_X1 U15409 ( .A1(n10937), .A2(n13730), .ZN(n13731) );
  NAND2_X1 U15410 ( .A1(n13805), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n13739) );
  INV_X1 U15411 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15907) );
  OR2_X1 U15412 ( .A1(n13807), .A2(n15907), .ZN(n13738) );
  OAI21_X1 U15413 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n13734), .A(n13733), 
        .ZN(n15906) );
  OR2_X1 U15414 ( .A1(n10700), .A2(n15906), .ZN(n13737) );
  INV_X1 U15415 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n13735) );
  OR2_X1 U15416 ( .A1(n13810), .A2(n13735), .ZN(n13736) );
  NAND4_X1 U15417 ( .A1(n13739), .A2(n13738), .A3(n13737), .A4(n13736), .ZN(
        n15917) );
  MUX2_X1 U15418 ( .A(n16088), .B(n15917), .S(n13771), .Z(n13741) );
  MUX2_X1 U15419 ( .A(n16088), .B(n15917), .S(n13836), .Z(n13740) );
  NAND2_X1 U15420 ( .A1(n13805), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n13748) );
  INV_X1 U15421 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15891) );
  OR2_X1 U15422 ( .A1(n13807), .A2(n15891), .ZN(n13747) );
  INV_X1 U15423 ( .A(n13742), .ZN(n13762) );
  OAI21_X1 U15424 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n13743), .A(n13762), 
        .ZN(n15890) );
  OR2_X1 U15425 ( .A1(n10700), .A2(n15890), .ZN(n13746) );
  INV_X1 U15426 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n13744) );
  OR2_X1 U15427 ( .A1(n13810), .A2(n13744), .ZN(n13745) );
  NAND4_X1 U15428 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n15737) );
  NAND2_X1 U15429 ( .A1(n13749), .A2(n13838), .ZN(n13752) );
  OR2_X1 U15430 ( .A1(n10937), .A2(n13750), .ZN(n13751) );
  MUX2_X1 U15431 ( .A(n15737), .B(n16082), .S(n13771), .Z(n13756) );
  NAND2_X1 U15432 ( .A1(n13755), .A2(n13756), .ZN(n13754) );
  MUX2_X1 U15433 ( .A(n15737), .B(n16082), .S(n13836), .Z(n13753) );
  INV_X1 U15434 ( .A(n13755), .ZN(n13758) );
  INV_X1 U15435 ( .A(n13756), .ZN(n13757) );
  NAND2_X1 U15436 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  NAND2_X1 U15437 ( .A1(n13805), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n13768) );
  INV_X1 U15438 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15879) );
  OR2_X1 U15439 ( .A1(n13807), .A2(n15879), .ZN(n13767) );
  INV_X1 U15440 ( .A(n13760), .ZN(n13779) );
  INV_X1 U15441 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13761) );
  NAND2_X1 U15442 ( .A1(n13762), .A2(n13761), .ZN(n13763) );
  NAND2_X1 U15443 ( .A1(n13779), .A2(n13763), .ZN(n15878) );
  OR2_X1 U15444 ( .A1(n10700), .A2(n15878), .ZN(n13766) );
  INV_X1 U15445 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n13764) );
  OR2_X1 U15446 ( .A1(n13810), .A2(n13764), .ZN(n13765) );
  NAND4_X1 U15447 ( .A1(n13768), .A2(n13767), .A3(n13766), .A4(n13765), .ZN(
        n15736) );
  NAND2_X1 U15448 ( .A1(n15624), .A2(n13838), .ZN(n13770) );
  OR2_X1 U15449 ( .A1(n10937), .A2(n16179), .ZN(n13769) );
  MUX2_X1 U15450 ( .A(n15736), .B(n16074), .S(n13836), .Z(n13773) );
  MUX2_X1 U15451 ( .A(n15736), .B(n16074), .S(n13771), .Z(n13772) );
  INV_X1 U15452 ( .A(n13773), .ZN(n13774) );
  NAND2_X1 U15453 ( .A1(n15621), .A2(n13838), .ZN(n13776) );
  OR2_X1 U15454 ( .A1(n10937), .A2(n8126), .ZN(n13775) );
  NAND2_X1 U15455 ( .A1(n13805), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n13786) );
  INV_X1 U15456 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13777) );
  OR2_X1 U15457 ( .A1(n13807), .A2(n13777), .ZN(n13785) );
  INV_X1 U15458 ( .A(n13792), .ZN(n13781) );
  INV_X1 U15459 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U15460 ( .A1(n13779), .A2(n13778), .ZN(n13780) );
  NAND2_X1 U15461 ( .A1(n13781), .A2(n13780), .ZN(n15860) );
  INV_X1 U15462 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n13782) );
  OR2_X1 U15463 ( .A1(n13810), .A2(n13782), .ZN(n13783) );
  NAND4_X1 U15464 ( .A1(n13786), .A2(n13785), .A3(n13784), .A4(n13783), .ZN(
        n15735) );
  MUX2_X1 U15465 ( .A(n16069), .B(n15735), .S(n13836), .Z(n13788) );
  MUX2_X1 U15466 ( .A(n15735), .B(n16069), .S(n13836), .Z(n13787) );
  INV_X1 U15467 ( .A(n13788), .ZN(n13789) );
  NAND2_X1 U15468 ( .A1(n13805), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n13797) );
  INV_X1 U15469 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13790) );
  OR2_X1 U15470 ( .A1(n13807), .A2(n13790), .ZN(n13796) );
  OAI21_X1 U15471 ( .B1(n13792), .B2(P1_REG3_REG_27__SCAN_IN), .A(n13791), 
        .ZN(n15849) );
  OR2_X1 U15472 ( .A1(n10700), .A2(n15849), .ZN(n13795) );
  INV_X1 U15473 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13793) );
  OR2_X1 U15474 ( .A1(n13810), .A2(n13793), .ZN(n13794) );
  NAND4_X1 U15475 ( .A1(n13797), .A2(n13796), .A3(n13795), .A4(n13794), .ZN(
        n15734) );
  NAND2_X1 U15476 ( .A1(n16169), .A2(n13838), .ZN(n13799) );
  OR2_X1 U15477 ( .A1(n10937), .A2(n16172), .ZN(n13798) );
  MUX2_X1 U15478 ( .A(n15734), .B(n16062), .S(n13836), .Z(n13801) );
  MUX2_X1 U15479 ( .A(n15734), .B(n16062), .S(n13771), .Z(n13800) );
  NAND2_X1 U15480 ( .A1(n15613), .A2(n13838), .ZN(n13804) );
  OR2_X1 U15481 ( .A1(n10937), .A2(n13802), .ZN(n13803) );
  NAND2_X1 U15482 ( .A1(n13805), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n13814) );
  INV_X1 U15483 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13806) );
  OR2_X1 U15484 ( .A1(n13807), .A2(n13806), .ZN(n13813) );
  OAI21_X1 U15485 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n13808), .A(n14034), 
        .ZN(n15835) );
  OR2_X1 U15486 ( .A1(n10700), .A2(n15835), .ZN(n13812) );
  INV_X1 U15487 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n13809) );
  OR2_X1 U15488 ( .A1(n13810), .A2(n13809), .ZN(n13811) );
  NAND4_X1 U15489 ( .A1(n13814), .A2(n13813), .A3(n13812), .A4(n13811), .ZN(
        n15733) );
  MUX2_X1 U15490 ( .A(n16054), .B(n15733), .S(n13836), .Z(n13815) );
  NAND2_X1 U15491 ( .A1(n13816), .A2(n13815), .ZN(n13819) );
  MUX2_X1 U15492 ( .A(n16054), .B(n15733), .S(n13771), .Z(n13818) );
  AOI21_X1 U15493 ( .B1(n13819), .B2(n13818), .A(n13817), .ZN(n13822) );
  INV_X1 U15494 ( .A(n13822), .ZN(n13824) );
  MUX2_X1 U15495 ( .A(n14031), .B(n15732), .S(n13836), .Z(n13820) );
  NAND2_X1 U15496 ( .A1(n13919), .A2(n13838), .ZN(n13827) );
  INV_X1 U15497 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14297) );
  OR2_X1 U15498 ( .A1(n10937), .A2(n14297), .ZN(n13826) );
  NAND2_X1 U15499 ( .A1(n13827), .A2(n13826), .ZN(n13852) );
  INV_X1 U15500 ( .A(n13828), .ZN(n13834) );
  INV_X1 U15501 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13833) );
  NAND2_X1 U15502 ( .A1(n13829), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U15503 ( .A1(n13830), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n13831) );
  OAI211_X1 U15504 ( .C1(n10679), .C2(n13833), .A(n13832), .B(n13831), .ZN(
        n15731) );
  OAI21_X1 U15505 ( .B1(n15815), .B2(n13834), .A(n15731), .ZN(n13835) );
  MUX2_X1 U15506 ( .A(n16045), .B(n13835), .S(n13836), .Z(n13901) );
  OAI21_X1 U15507 ( .B1(n15815), .B2(n13586), .A(n15731), .ZN(n13837) );
  MUX2_X1 U15508 ( .A(n13837), .B(n16045), .S(n13836), .Z(n13897) );
  INV_X1 U15509 ( .A(n13897), .ZN(n13900) );
  INV_X1 U15510 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16163) );
  XNOR2_X1 U15511 ( .A(n13845), .B(n15815), .ZN(n13909) );
  NAND2_X1 U15512 ( .A1(n13850), .A2(n13839), .ZN(n13841) );
  NAND2_X1 U15513 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  AND2_X1 U15514 ( .A1(n13843), .A2(n13842), .ZN(n13848) );
  INV_X1 U15515 ( .A(n13848), .ZN(n13891) );
  NOR2_X1 U15516 ( .A1(n13891), .A2(n13908), .ZN(n13899) );
  OAI211_X1 U15517 ( .C1(n13901), .C2(n13900), .A(n13909), .B(n13899), .ZN(
        n13913) );
  INV_X1 U15518 ( .A(n15815), .ZN(n13844) );
  NAND2_X1 U15519 ( .A1(n13845), .A2(n13844), .ZN(n13847) );
  NAND2_X1 U15520 ( .A1(n16042), .A2(n15815), .ZN(n13846) );
  MUX2_X1 U15521 ( .A(n13847), .B(n13846), .S(n7421), .Z(n13896) );
  XNOR2_X1 U15522 ( .A(n13896), .B(n13848), .ZN(n13851) );
  OR2_X1 U15523 ( .A1(n13850), .A2(n13849), .ZN(n13890) );
  NAND2_X1 U15524 ( .A1(n13851), .A2(n13890), .ZN(n13888) );
  XNOR2_X1 U15525 ( .A(n13852), .B(n15731), .ZN(n13882) );
  INV_X1 U15526 ( .A(n15733), .ZN(n14051) );
  XNOR2_X1 U15527 ( .A(n16054), .B(n14051), .ZN(n15832) );
  XNOR2_X1 U15528 ( .A(n16069), .B(n15735), .ZN(n15856) );
  INV_X1 U15529 ( .A(n15737), .ZN(n15674) );
  OR2_X1 U15530 ( .A1(n16082), .A2(n15674), .ZN(n14027) );
  NAND2_X1 U15531 ( .A1(n16082), .A2(n15674), .ZN(n13853) );
  NAND2_X1 U15532 ( .A1(n14027), .A2(n13853), .ZN(n15895) );
  XNOR2_X1 U15533 ( .A(n15921), .B(n15738), .ZN(n15927) );
  XNOR2_X1 U15534 ( .A(n16088), .B(n15917), .ZN(n15912) );
  XNOR2_X1 U15535 ( .A(n15958), .B(n15976), .ZN(n14025) );
  XNOR2_X1 U15536 ( .A(n16111), .B(n15954), .ZN(n14048) );
  XNOR2_X1 U15537 ( .A(n16129), .B(n14042), .ZN(n16026) );
  NOR3_X1 U15538 ( .A1(n13859), .A2(n13858), .A3(n13857), .ZN(n13861) );
  NAND3_X1 U15539 ( .A1(n16574), .A2(n13861), .A3(n13860), .ZN(n13862) );
  NOR2_X1 U15540 ( .A1(n13863), .A2(n13862), .ZN(n13865) );
  NAND4_X1 U15541 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n16618), .ZN(
        n13867) );
  NOR2_X1 U15542 ( .A1(n13868), .A2(n13867), .ZN(n13871) );
  NAND4_X1 U15543 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13873) );
  NOR2_X1 U15544 ( .A1(n16026), .A2(n13873), .ZN(n13874) );
  XNOR2_X1 U15545 ( .A(n16118), .B(n15740), .ZN(n15991) );
  XNOR2_X1 U15546 ( .A(n16123), .B(n15741), .ZN(n16015) );
  NAND4_X1 U15547 ( .A1(n14048), .A2(n13874), .A3(n15991), .A4(n16015), .ZN(
        n13875) );
  NOR2_X1 U15548 ( .A1(n14025), .A2(n13875), .ZN(n13876) );
  XNOR2_X1 U15549 ( .A(n15937), .B(n15957), .ZN(n15934) );
  NAND3_X1 U15550 ( .A1(n15912), .A2(n13876), .A3(n15934), .ZN(n13877) );
  NOR3_X1 U15551 ( .A1(n15895), .A2(n15927), .A3(n13877), .ZN(n13879) );
  NAND2_X1 U15552 ( .A1(n16074), .A2(n15736), .ZN(n14049) );
  OR2_X1 U15553 ( .A1(n16074), .A2(n15736), .ZN(n13878) );
  NAND2_X1 U15554 ( .A1(n14049), .A2(n13878), .ZN(n15873) );
  NAND3_X1 U15555 ( .A1(n15856), .A2(n13879), .A3(n15873), .ZN(n13880) );
  NOR2_X1 U15556 ( .A1(n15832), .A2(n13880), .ZN(n13881) );
  XNOR2_X1 U15557 ( .A(n14031), .B(n15732), .ZN(n14052) );
  XNOR2_X1 U15558 ( .A(n16062), .B(n15734), .ZN(n15846) );
  AND4_X1 U15559 ( .A1(n13882), .A2(n13881), .A3(n14052), .A4(n15846), .ZN(
        n13883) );
  NAND2_X1 U15560 ( .A1(n13909), .A2(n13883), .ZN(n13884) );
  XNOR2_X1 U15561 ( .A(n13884), .B(n16033), .ZN(n13886) );
  INV_X1 U15562 ( .A(n13890), .ZN(n13885) );
  NAND2_X1 U15563 ( .A1(n13886), .A2(n13885), .ZN(n13887) );
  NAND2_X1 U15564 ( .A1(n13897), .A2(n13889), .ZN(n13894) );
  INV_X1 U15565 ( .A(n13896), .ZN(n13893) );
  AND2_X1 U15566 ( .A1(n13891), .A2(n13890), .ZN(n13910) );
  INV_X1 U15567 ( .A(n13910), .ZN(n13892) );
  OR3_X1 U15568 ( .A1(n13901), .A2(n13908), .A3(n13892), .ZN(n13895) );
  OAI22_X1 U15569 ( .A1(n13907), .A2(n13894), .B1(n13893), .B2(n13895), .ZN(
        n13912) );
  INV_X1 U15570 ( .A(n13895), .ZN(n13898) );
  NAND3_X1 U15571 ( .A1(n13898), .A2(n13897), .A3(n13896), .ZN(n13906) );
  NAND4_X1 U15572 ( .A1(n13909), .A2(n13901), .A3(n13900), .A4(n13899), .ZN(
        n13905) );
  INV_X1 U15573 ( .A(n16170), .ZN(n16280) );
  NAND3_X1 U15574 ( .A1(n13902), .A2(n16280), .A3(n15955), .ZN(n13903) );
  OAI211_X1 U15575 ( .C1(n16180), .C2(n13908), .A(n13903), .B(P1_B_REG_SCAN_IN), .ZN(n13904) );
  NAND3_X1 U15576 ( .A1(n13906), .A2(n13905), .A3(n13904), .ZN(n13911) );
  INV_X1 U15577 ( .A(n13915), .ZN(n13917) );
  OAI222_X1 U15578 ( .A1(n14968), .A2(n13917), .B1(n14959), .B2(n13916), .C1(
        P3_U3151), .C2(n14510), .ZN(P3_U3267) );
  INV_X1 U15579 ( .A(n13919), .ZN(n14056) );
  INV_X1 U15580 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14302) );
  OAI222_X1 U15581 ( .A1(P2_U3088), .A2(n13918), .B1(n15626), .B2(n14056), 
        .C1(n14302), .C2(n15628), .ZN(P2_U3297) );
  INV_X1 U15582 ( .A(n14720), .ZN(n14689) );
  XNOR2_X1 U15583 ( .A(n14323), .B(n13935), .ZN(n13941) );
  INV_X1 U15584 ( .A(n13941), .ZN(n14119) );
  XNOR2_X1 U15585 ( .A(n14882), .B(n14163), .ZN(n13923) );
  XNOR2_X1 U15586 ( .A(n13923), .B(n14227), .ZN(n14203) );
  INV_X1 U15587 ( .A(n13923), .ZN(n13924) );
  NAND2_X1 U15588 ( .A1(n13924), .A2(n14227), .ZN(n13925) );
  XNOR2_X1 U15589 ( .A(n14796), .B(n14163), .ZN(n13926) );
  XNOR2_X1 U15590 ( .A(n13926), .B(n14778), .ZN(n14225) );
  INV_X1 U15591 ( .A(n13926), .ZN(n13927) );
  NAND2_X1 U15592 ( .A1(n13927), .A2(n14778), .ZN(n13928) );
  XNOR2_X1 U15593 ( .A(n14873), .B(n12268), .ZN(n13929) );
  XNOR2_X1 U15594 ( .A(n13929), .B(n14156), .ZN(n14275) );
  INV_X1 U15595 ( .A(n13929), .ZN(n13930) );
  NAND2_X1 U15596 ( .A1(n13930), .A2(n14156), .ZN(n13931) );
  XNOR2_X1 U15597 ( .A(n14160), .B(n14163), .ZN(n13932) );
  XNOR2_X1 U15598 ( .A(n13932), .B(n14750), .ZN(n14154) );
  NAND2_X1 U15599 ( .A1(n13932), .A2(n14750), .ZN(n13933) );
  XNOR2_X1 U15600 ( .A(n14934), .B(n14163), .ZN(n13934) );
  XNOR2_X1 U15601 ( .A(n13934), .B(n14187), .ZN(n14243) );
  INV_X1 U15602 ( .A(n12268), .ZN(n13935) );
  XNOR2_X1 U15603 ( .A(n14191), .B(n13935), .ZN(n13936) );
  AND2_X1 U15604 ( .A1(n13936), .A2(n14719), .ZN(n14183) );
  INV_X1 U15605 ( .A(n13936), .ZN(n13937) );
  NAND2_X1 U15606 ( .A1(n13937), .A2(n14751), .ZN(n14182) );
  XNOR2_X1 U15607 ( .A(n14854), .B(n14163), .ZN(n13938) );
  XNOR2_X1 U15608 ( .A(n14918), .B(n14163), .ZN(n13943) );
  NOR2_X1 U15609 ( .A1(n13943), .A2(n14673), .ZN(n13945) );
  AOI21_X1 U15610 ( .B1(n14673), .B2(n13943), .A(n13945), .ZN(n14234) );
  INV_X1 U15611 ( .A(n13945), .ZN(n14195) );
  XNOR2_X1 U15612 ( .A(n14681), .B(n12268), .ZN(n13946) );
  NAND2_X1 U15613 ( .A1(n13946), .A2(n14690), .ZN(n13949) );
  INV_X1 U15614 ( .A(n13946), .ZN(n13947) );
  NAND2_X1 U15615 ( .A1(n13947), .A2(n14325), .ZN(n13948) );
  NAND2_X1 U15616 ( .A1(n13949), .A2(n13948), .ZN(n14194) );
  INV_X1 U15617 ( .A(n13949), .ZN(n13950) );
  NOR2_X1 U15618 ( .A1(n14197), .A2(n13950), .ZN(n14286) );
  XNOR2_X1 U15619 ( .A(n14293), .B(n14163), .ZN(n13951) );
  NAND2_X1 U15620 ( .A1(n13951), .A2(n14646), .ZN(n13952) );
  OAI21_X1 U15621 ( .B1(n13951), .B2(n14646), .A(n13952), .ZN(n14285) );
  INV_X1 U15622 ( .A(n13952), .ZN(n13953) );
  XNOR2_X1 U15623 ( .A(n14655), .B(n14163), .ZN(n14176) );
  NAND2_X1 U15624 ( .A1(n14176), .A2(n14661), .ZN(n14164) );
  OAI21_X1 U15625 ( .B1(n14176), .B2(n14661), .A(n14164), .ZN(n13954) );
  AOI22_X1 U15626 ( .A1(n14674), .A2(n7422), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13956) );
  NAND2_X1 U15627 ( .A1(n14654), .A2(n14287), .ZN(n13955) );
  OAI211_X1 U15628 ( .C1(n14647), .C2(n14290), .A(n13956), .B(n13955), .ZN(
        n13957) );
  AOI21_X1 U15629 ( .B1(n14655), .B2(n14292), .A(n13957), .ZN(n13958) );
  OAI21_X1 U15630 ( .B1(n13959), .B2(n14295), .A(n13958), .ZN(P3_U3154) );
  INV_X1 U15631 ( .A(n13960), .ZN(n13961) );
  AOI22_X1 U15632 ( .A1(n15937), .A2(n8750), .B1(n14013), .B2(n15957), .ZN(
        n13963) );
  XNOR2_X1 U15633 ( .A(n13963), .B(n13999), .ZN(n13965) );
  AOI22_X1 U15634 ( .A1(n15937), .A2(n14013), .B1(n14001), .B2(n15957), .ZN(
        n13964) );
  XNOR2_X1 U15635 ( .A(n13965), .B(n13964), .ZN(n15664) );
  NAND2_X1 U15636 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  OAI22_X1 U15637 ( .A1(n15921), .A2(n13968), .B1(n15665), .B2(n13967), .ZN(
        n13972) );
  OAI22_X1 U15638 ( .A1(n15921), .A2(n13969), .B1(n15665), .B2(n13968), .ZN(
        n13970) );
  XNOR2_X1 U15639 ( .A(n13970), .B(n13999), .ZN(n13971) );
  XOR2_X1 U15640 ( .A(n13972), .B(n13971), .Z(n15705) );
  INV_X1 U15641 ( .A(n13971), .ZN(n13974) );
  INV_X1 U15642 ( .A(n13972), .ZN(n13973) );
  NAND2_X1 U15643 ( .A1(n13974), .A2(n13973), .ZN(n13975) );
  NAND2_X1 U15644 ( .A1(n16088), .A2(n8750), .ZN(n13977) );
  NAND2_X1 U15645 ( .A1(n15917), .A2(n14013), .ZN(n13976) );
  NAND2_X1 U15646 ( .A1(n13977), .A2(n13976), .ZN(n13978) );
  XNOR2_X1 U15647 ( .A(n13978), .B(n13999), .ZN(n13979) );
  AOI22_X1 U15648 ( .A1(n16088), .A2(n14013), .B1(n14001), .B2(n15917), .ZN(
        n13980) );
  XNOR2_X1 U15649 ( .A(n13979), .B(n13980), .ZN(n15649) );
  INV_X1 U15650 ( .A(n13979), .ZN(n13981) );
  NAND2_X1 U15651 ( .A1(n16082), .A2(n8750), .ZN(n13983) );
  NAND2_X1 U15652 ( .A1(n15737), .A2(n14005), .ZN(n13982) );
  NAND2_X1 U15653 ( .A1(n13983), .A2(n13982), .ZN(n13984) );
  XNOR2_X1 U15654 ( .A(n13984), .B(n13999), .ZN(n13985) );
  AOI22_X1 U15655 ( .A1(n16082), .A2(n14013), .B1(n14012), .B2(n15737), .ZN(
        n13986) );
  XNOR2_X1 U15656 ( .A(n13985), .B(n13986), .ZN(n15697) );
  INV_X1 U15657 ( .A(n13985), .ZN(n13987) );
  NAND2_X1 U15658 ( .A1(n13987), .A2(n13986), .ZN(n13988) );
  NAND2_X1 U15659 ( .A1(n16074), .A2(n8750), .ZN(n13991) );
  NAND2_X1 U15660 ( .A1(n15736), .A2(n14013), .ZN(n13990) );
  NAND2_X1 U15661 ( .A1(n13991), .A2(n13990), .ZN(n13992) );
  XNOR2_X1 U15662 ( .A(n13992), .B(n13999), .ZN(n13993) );
  AOI22_X1 U15663 ( .A1(n16074), .A2(n14013), .B1(n14001), .B2(n15736), .ZN(
        n13994) );
  XNOR2_X1 U15664 ( .A(n13993), .B(n13994), .ZN(n15673) );
  INV_X1 U15665 ( .A(n13993), .ZN(n13995) );
  NAND2_X1 U15666 ( .A1(n13995), .A2(n13994), .ZN(n13996) );
  NAND2_X1 U15667 ( .A1(n16069), .A2(n8750), .ZN(n13998) );
  NAND2_X1 U15668 ( .A1(n15735), .A2(n14005), .ZN(n13997) );
  NAND2_X1 U15669 ( .A1(n13998), .A2(n13997), .ZN(n14000) );
  XNOR2_X1 U15670 ( .A(n14000), .B(n13999), .ZN(n14002) );
  AOI22_X1 U15671 ( .A1(n16069), .A2(n14005), .B1(n14001), .B2(n15735), .ZN(
        n14003) );
  XNOR2_X1 U15672 ( .A(n14002), .B(n14003), .ZN(n15723) );
  INV_X1 U15673 ( .A(n14002), .ZN(n14004) );
  NAND2_X1 U15674 ( .A1(n16062), .A2(n8750), .ZN(n14007) );
  NAND2_X1 U15675 ( .A1(n15734), .A2(n14005), .ZN(n14006) );
  NAND2_X1 U15676 ( .A1(n14007), .A2(n14006), .ZN(n14008) );
  XNOR2_X1 U15677 ( .A(n14008), .B(n13999), .ZN(n14009) );
  AOI22_X1 U15678 ( .A1(n16062), .A2(n14013), .B1(n14012), .B2(n15734), .ZN(
        n14010) );
  XNOR2_X1 U15679 ( .A(n14009), .B(n14010), .ZN(n15631) );
  INV_X1 U15680 ( .A(n14009), .ZN(n14011) );
  AOI22_X1 U15681 ( .A1(n16054), .A2(n14013), .B1(n14012), .B2(n15733), .ZN(
        n14016) );
  AOI22_X1 U15682 ( .A1(n16054), .A2(n8750), .B1(n14013), .B2(n15733), .ZN(
        n14014) );
  XNOR2_X1 U15683 ( .A(n14014), .B(n13999), .ZN(n14015) );
  XOR2_X1 U15684 ( .A(n14016), .B(n14015), .Z(n14017) );
  INV_X1 U15685 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14018) );
  OAI22_X1 U15686 ( .A1(n16723), .A2(n15835), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14018), .ZN(n14020) );
  INV_X1 U15687 ( .A(n15734), .ZN(n15828) );
  OAI22_X1 U15688 ( .A1(n15827), .A2(n15717), .B1(n15716), .B2(n15828), .ZN(
        n14019) );
  AOI211_X1 U15689 ( .C1(n16054), .C2(n16719), .A(n14020), .B(n14019), .ZN(
        n14021) );
  OAI21_X1 U15690 ( .B1(n14022), .B2(n15729), .A(n14021), .ZN(P1_U3220) );
  INV_X1 U15691 ( .A(n16074), .ZN(n15871) );
  INV_X1 U15692 ( .A(n15740), .ZN(n15977) );
  INV_X1 U15693 ( .A(n16129), .ZN(n14043) );
  INV_X1 U15694 ( .A(n15741), .ZN(n16028) );
  INV_X1 U15695 ( .A(n15927), .ZN(n15916) );
  INV_X1 U15696 ( .A(n16088), .ZN(n15905) );
  INV_X1 U15697 ( .A(n15895), .ZN(n14026) );
  OAI21_X1 U15698 ( .B1(n15871), .B2(n15736), .A(n15872), .ZN(n15857) );
  INV_X1 U15699 ( .A(n15735), .ZN(n15675) );
  NAND2_X1 U15700 ( .A1(n16069), .A2(n15675), .ZN(n14028) );
  NOR2_X1 U15701 ( .A1(n15839), .A2(n15733), .ZN(n14029) );
  OAI22_X1 U15702 ( .A1(n15826), .A2(n14029), .B1(n14051), .B2(n16054), .ZN(
        n14030) );
  INV_X1 U15703 ( .A(n16111), .ZN(n15985) );
  INV_X1 U15704 ( .A(n16082), .ZN(n15889) );
  AOI211_X1 U15705 ( .C1(n14031), .C2(n15834), .A(n16686), .B(n15820), .ZN(
        n16050) );
  INV_X1 U15706 ( .A(P1_B_REG_SCAN_IN), .ZN(n14032) );
  NOR2_X1 U15707 ( .A1(n16170), .A2(n14032), .ZN(n14033) );
  NOR2_X1 U15708 ( .A1(n16029), .A2(n14033), .ZN(n15814) );
  NAND2_X1 U15709 ( .A1(n15731), .A2(n15814), .ZN(n16046) );
  OAI22_X1 U15710 ( .A1(n14035), .A2(n16046), .B1(n14034), .B2(n16036), .ZN(
        n14037) );
  NAND2_X1 U15711 ( .A1(n15733), .A2(n15955), .ZN(n16047) );
  NOR2_X1 U15712 ( .A1(n16642), .A2(n16047), .ZN(n14036) );
  AOI211_X1 U15713 ( .C1(n16642), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14037), 
        .B(n14036), .ZN(n14038) );
  OAI21_X1 U15714 ( .B1(n16048), .B2(n16587), .A(n14038), .ZN(n14039) );
  AOI21_X1 U15715 ( .B1(n16050), .B2(n16636), .A(n14039), .ZN(n14055) );
  OR2_X1 U15716 ( .A1(n16718), .A2(n15743), .ZN(n14040) );
  NAND2_X1 U15717 ( .A1(n14043), .A2(n14042), .ZN(n14044) );
  INV_X1 U15718 ( .A(n16118), .ZN(n15999) );
  NAND2_X1 U15719 ( .A1(n15999), .A2(n15977), .ZN(n14045) );
  NAND2_X1 U15720 ( .A1(n16118), .A2(n15740), .ZN(n14046) );
  OR2_X2 U15721 ( .A1(n15964), .A2(n15963), .ZN(n15966) );
  INV_X1 U15722 ( .A(n14049), .ZN(n14050) );
  INV_X1 U15723 ( .A(n16069), .ZN(n15865) );
  XNOR2_X1 U15724 ( .A(n14053), .B(n14052), .ZN(n16051) );
  NAND2_X1 U15725 ( .A1(n16051), .A2(n15929), .ZN(n14054) );
  OAI211_X1 U15726 ( .C1(n16053), .C2(n15970), .A(n14055), .B(n14054), .ZN(
        P1_U3356) );
  OAI222_X1 U15727 ( .A1(n16174), .A2(n14297), .B1(P1_U3086), .B2(n14057), 
        .C1(n16178), .C2(n14056), .ZN(P1_U3325) );
  AOI22_X1 U15728 ( .A1(n15033), .A2(n14059), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14058), .ZN(n14065) );
  OAI21_X1 U15729 ( .B1(n14062), .B2(n14061), .A(n14060), .ZN(n14063) );
  NAND2_X1 U15730 ( .A1(n15070), .A2(n14063), .ZN(n14064) );
  OAI211_X1 U15731 ( .C1(n14066), .C2(n15066), .A(n14065), .B(n14064), .ZN(
        P2_U3194) );
  NOR2_X1 U15732 ( .A1(n15192), .A2(n15232), .ZN(n14106) );
  XNOR2_X1 U15733 ( .A(n15284), .B(n11679), .ZN(n14104) );
  NAND2_X1 U15734 ( .A1(n15212), .A2(n7418), .ZN(n14088) );
  INV_X1 U15735 ( .A(n14088), .ZN(n14092) );
  XNOR2_X1 U15736 ( .A(n15360), .B(n11679), .ZN(n14089) );
  INV_X1 U15737 ( .A(n14089), .ZN(n14091) );
  INV_X1 U15738 ( .A(n14067), .ZN(n14069) );
  NAND2_X1 U15739 ( .A1(n14069), .A2(n14068), .ZN(n14070) );
  XNOR2_X1 U15740 ( .A(n15595), .B(n7695), .ZN(n14072) );
  NOR2_X1 U15741 ( .A1(n15203), .A2(n15232), .ZN(n14073) );
  NAND2_X1 U15742 ( .A1(n14072), .A2(n14073), .ZN(n14076) );
  INV_X1 U15743 ( .A(n14072), .ZN(n14986) );
  INV_X1 U15744 ( .A(n14073), .ZN(n14074) );
  NAND2_X1 U15745 ( .A1(n14986), .A2(n14074), .ZN(n14075) );
  XNOR2_X1 U15746 ( .A(n15590), .B(n7695), .ZN(n14077) );
  NOR2_X1 U15747 ( .A1(n15181), .A2(n15232), .ZN(n14078) );
  NAND2_X1 U15748 ( .A1(n14077), .A2(n14078), .ZN(n14082) );
  INV_X1 U15749 ( .A(n14077), .ZN(n15039) );
  INV_X1 U15750 ( .A(n14078), .ZN(n14079) );
  NAND2_X1 U15751 ( .A1(n15039), .A2(n14079), .ZN(n14080) );
  AND2_X1 U15752 ( .A1(n14082), .A2(n14080), .ZN(n14984) );
  NAND2_X1 U15753 ( .A1(n15037), .A2(n14082), .ZN(n14087) );
  XNOR2_X1 U15754 ( .A(n15585), .B(n7695), .ZN(n14083) );
  NOR2_X1 U15755 ( .A1(n15183), .A2(n15232), .ZN(n14084) );
  NAND2_X1 U15756 ( .A1(n14083), .A2(n14084), .ZN(n14090) );
  INV_X1 U15757 ( .A(n14083), .ZN(n14992) );
  INV_X1 U15758 ( .A(n14084), .ZN(n14085) );
  NAND2_X1 U15759 ( .A1(n14992), .A2(n14085), .ZN(n14086) );
  AND2_X1 U15760 ( .A1(n14090), .A2(n14086), .ZN(n15036) );
  XNOR2_X1 U15761 ( .A(n14089), .B(n14088), .ZN(n14993) );
  XNOR2_X1 U15762 ( .A(n15342), .B(n11679), .ZN(n14093) );
  INV_X1 U15763 ( .A(n14093), .ZN(n14094) );
  XNOR2_X1 U15764 ( .A(n15496), .B(n11679), .ZN(n15003) );
  AND2_X1 U15765 ( .A1(n15191), .A2(n7418), .ZN(n14097) );
  NAND2_X1 U15766 ( .A1(n15003), .A2(n14097), .ZN(n14098) );
  OAI21_X1 U15767 ( .B1(n15003), .B2(n14097), .A(n14098), .ZN(n15027) );
  INV_X1 U15768 ( .A(n14098), .ZN(n14103) );
  XNOR2_X1 U15769 ( .A(n15299), .B(n11679), .ZN(n14099) );
  AND2_X1 U15770 ( .A1(n15084), .A2(n7418), .ZN(n14100) );
  NAND2_X1 U15771 ( .A1(n14099), .A2(n14100), .ZN(n14105) );
  INV_X1 U15772 ( .A(n14099), .ZN(n15068) );
  INV_X1 U15773 ( .A(n14100), .ZN(n14101) );
  NAND2_X1 U15774 ( .A1(n15068), .A2(n14101), .ZN(n14102) );
  AND2_X1 U15775 ( .A1(n14105), .A2(n14102), .ZN(n15005) );
  XNOR2_X1 U15776 ( .A(n14104), .B(n14106), .ZN(n15081) );
  XNOR2_X1 U15777 ( .A(n15478), .B(n11679), .ZN(n14108) );
  AND2_X1 U15778 ( .A1(n15193), .A2(n7418), .ZN(n14107) );
  NAND2_X1 U15779 ( .A1(n14108), .A2(n14107), .ZN(n14111) );
  OAI21_X1 U15780 ( .B1(n14108), .B2(n14107), .A(n14111), .ZN(n14973) );
  NOR2_X1 U15781 ( .A1(n15220), .A2(n15067), .ZN(n14109) );
  AOI22_X1 U15782 ( .A1(n14972), .A2(n15070), .B1(n14109), .B2(n14108), .ZN(
        n14118) );
  MUX2_X1 U15783 ( .A(n15241), .B(n15474), .S(n15232), .Z(n14110) );
  INV_X1 U15784 ( .A(n14111), .ZN(n14112) );
  NAND2_X1 U15785 ( .A1(n7430), .A2(n8828), .ZN(n14117) );
  AOI22_X1 U15786 ( .A1(n15083), .A2(n15073), .B1(n15225), .B2(n15193), .ZN(
        n15253) );
  INV_X1 U15787 ( .A(n15255), .ZN(n14113) );
  AOI22_X1 U15788 ( .A1(n14113), .A2(n15074), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14114) );
  OAI21_X1 U15789 ( .B1(n15253), .B2(n15076), .A(n14114), .ZN(n14115) );
  OAI21_X1 U15790 ( .B1(n14118), .B2(n7430), .A(n7498), .ZN(P2_U3192) );
  OAI21_X1 U15791 ( .B1(n14120), .B2(n14119), .A(n14232), .ZN(n14121) );
  NOR2_X1 U15792 ( .A1(n14121), .A2(n14720), .ZN(n14235) );
  AOI21_X1 U15793 ( .B1(n14720), .B2(n14121), .A(n14235), .ZN(n14126) );
  AOI22_X1 U15794 ( .A1(n7422), .A2(n14267), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14123) );
  NAND2_X1 U15795 ( .A1(n14287), .A2(n14707), .ZN(n14122) );
  OAI211_X1 U15796 ( .C1(n14702), .C2(n14290), .A(n14123), .B(n14122), .ZN(
        n14124) );
  AOI21_X1 U15797 ( .B1(n14323), .B2(n14292), .A(n14124), .ZN(n14125) );
  OAI21_X1 U15798 ( .B1(n14126), .B2(n14295), .A(n14125), .ZN(P3_U3156) );
  AND2_X1 U15799 ( .A1(n14128), .A2(n14127), .ZN(n14131) );
  OAI211_X1 U15800 ( .C1(n14131), .C2(n14130), .A(n14273), .B(n14129), .ZN(
        n14138) );
  AOI21_X1 U15801 ( .B1(n14292), .B2(n14402), .A(n14132), .ZN(n14137) );
  AOI22_X1 U15802 ( .A1(n14218), .A2(n14133), .B1(n7422), .B2(n14398), .ZN(
        n14136) );
  NAND2_X1 U15803 ( .A1(n14287), .A2(n14134), .ZN(n14135) );
  NAND4_X1 U15804 ( .A1(n14138), .A2(n14137), .A3(n14136), .A4(n14135), .ZN(
        P3_U3157) );
  AND2_X1 U15805 ( .A1(n14140), .A2(n14139), .ZN(n14143) );
  OAI211_X1 U15806 ( .C1(n14143), .C2(n14142), .A(n14273), .B(n14141), .ZN(
        n14150) );
  AOI21_X1 U15807 ( .B1(n14292), .B2(n14145), .A(n14144), .ZN(n14149) );
  AOI22_X1 U15808 ( .A1(n14218), .A2(n14216), .B1(n7422), .B2(n14366), .ZN(
        n14148) );
  NAND2_X1 U15809 ( .A1(n14287), .A2(n14146), .ZN(n14147) );
  NAND4_X1 U15810 ( .A1(n14150), .A2(n14149), .A3(n14148), .A4(n14147), .ZN(
        P3_U3158) );
  INV_X1 U15811 ( .A(n14151), .ZN(n14152) );
  AOI21_X1 U15812 ( .B1(n14154), .B2(n14153), .A(n14152), .ZN(n14162) );
  NOR2_X1 U15813 ( .A1(n14155), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14608) );
  AOI21_X1 U15814 ( .B1(n7422), .B2(n14156), .A(n14608), .ZN(n14158) );
  NAND2_X1 U15815 ( .A1(n14287), .A2(n14766), .ZN(n14157) );
  OAI211_X1 U15816 ( .C1(n14763), .C2(n14290), .A(n14158), .B(n14157), .ZN(
        n14159) );
  AOI21_X1 U15817 ( .B1(n14160), .B2(n14292), .A(n14159), .ZN(n14161) );
  OAI21_X1 U15818 ( .B1(n14162), .B2(n14295), .A(n14161), .ZN(P3_U3159) );
  XNOR2_X1 U15819 ( .A(n14634), .B(n14163), .ZN(n14174) );
  NAND3_X1 U15820 ( .A1(n14174), .A2(n14164), .A3(n14273), .ZN(n14165) );
  INV_X1 U15821 ( .A(n14633), .ZN(n14172) );
  INV_X1 U15822 ( .A(n14287), .ZN(n14171) );
  OAI22_X1 U15823 ( .A1(n14661), .A2(n14167), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14166), .ZN(n14168) );
  AOI21_X1 U15824 ( .B1(n14169), .B2(n14218), .A(n14168), .ZN(n14170) );
  OAI21_X1 U15825 ( .B1(n14172), .B2(n14171), .A(n14170), .ZN(n14173) );
  AOI21_X1 U15826 ( .B1(n14638), .B2(n14292), .A(n14173), .ZN(n14180) );
  INV_X1 U15827 ( .A(n14174), .ZN(n14177) );
  NAND3_X1 U15828 ( .A1(n14175), .A2(n14273), .A3(n14177), .ZN(n14179) );
  NAND4_X1 U15829 ( .A1(n14177), .A2(n14273), .A3(n14661), .A4(n14176), .ZN(
        n14178) );
  NAND4_X1 U15830 ( .A1(n14181), .A2(n14180), .A3(n14179), .A4(n14178), .ZN(
        P3_U3160) );
  INV_X1 U15831 ( .A(n14182), .ZN(n14184) );
  NOR2_X1 U15832 ( .A1(n14184), .A2(n14183), .ZN(n14185) );
  XNOR2_X1 U15833 ( .A(n14186), .B(n14185), .ZN(n14193) );
  AOI22_X1 U15834 ( .A1(n7422), .A2(n14187), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14189) );
  NAND2_X1 U15835 ( .A1(n14287), .A2(n14741), .ZN(n14188) );
  OAI211_X1 U15836 ( .C1(n14737), .C2(n14290), .A(n14189), .B(n14188), .ZN(
        n14190) );
  AOI21_X1 U15837 ( .B1(n14191), .B2(n14292), .A(n14190), .ZN(n14192) );
  OAI21_X1 U15838 ( .B1(n14193), .B2(n14295), .A(n14192), .ZN(P3_U3163) );
  AND3_X1 U15839 ( .A1(n14236), .A2(n14195), .A3(n14194), .ZN(n14196) );
  OAI21_X1 U15840 ( .B1(n14197), .B2(n14196), .A(n14273), .ZN(n14201) );
  AOI22_X1 U15841 ( .A1(n14673), .A2(n7422), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14198) );
  OAI21_X1 U15842 ( .B1(n14646), .B2(n14290), .A(n14198), .ZN(n14199) );
  AOI21_X1 U15843 ( .B1(n14677), .B2(n14287), .A(n14199), .ZN(n14200) );
  OAI211_X1 U15844 ( .C1(n14914), .C2(n14282), .A(n14201), .B(n14200), .ZN(
        P3_U3165) );
  INV_X1 U15845 ( .A(n14882), .ZN(n14810) );
  OAI211_X1 U15846 ( .C1(n14204), .C2(n14203), .A(n14202), .B(n14273), .ZN(
        n14209) );
  NAND2_X1 U15847 ( .A1(n7422), .A2(n14205), .ZN(n14206) );
  NAND2_X1 U15848 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14558)
         );
  OAI211_X1 U15849 ( .C1(n14290), .C2(n14806), .A(n14206), .B(n14558), .ZN(
        n14207) );
  AOI21_X1 U15850 ( .B1(n14807), .B2(n14287), .A(n14207), .ZN(n14208) );
  OAI211_X1 U15851 ( .C1(n14810), .C2(n14282), .A(n14209), .B(n14208), .ZN(
        P3_U3166) );
  OAI21_X1 U15852 ( .B1(n14212), .B2(n14211), .A(n14210), .ZN(n14213) );
  NAND2_X1 U15853 ( .A1(n14213), .A2(n14273), .ZN(n14223) );
  AOI21_X1 U15854 ( .B1(n14292), .B2(n14215), .A(n14214), .ZN(n14222) );
  AOI22_X1 U15855 ( .A1(n14218), .A2(n14217), .B1(n7422), .B2(n14216), .ZN(
        n14221) );
  NAND2_X1 U15856 ( .A1(n14287), .A2(n14219), .ZN(n14220) );
  NAND4_X1 U15857 ( .A1(n14223), .A2(n14222), .A3(n14221), .A4(n14220), .ZN(
        P3_U3167) );
  INV_X1 U15858 ( .A(n14796), .ZN(n14880) );
  OAI211_X1 U15859 ( .C1(n14226), .C2(n14225), .A(n14224), .B(n14273), .ZN(
        n14231) );
  NAND2_X1 U15860 ( .A1(n7422), .A2(n14227), .ZN(n14228) );
  NAND2_X1 U15861 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14571)
         );
  OAI211_X1 U15862 ( .C1(n14290), .C2(n14786), .A(n14228), .B(n14571), .ZN(
        n14229) );
  AOI21_X1 U15863 ( .B1(n14791), .B2(n14287), .A(n14229), .ZN(n14230) );
  OAI211_X1 U15864 ( .C1(n14880), .C2(n14282), .A(n14231), .B(n14230), .ZN(
        P3_U3168) );
  INV_X1 U15865 ( .A(n14232), .ZN(n14233) );
  NOR3_X1 U15866 ( .A1(n14235), .A2(n14234), .A3(n14233), .ZN(n14238) );
  INV_X1 U15867 ( .A(n14236), .ZN(n14237) );
  OAI21_X1 U15868 ( .B1(n14238), .B2(n14237), .A(n14273), .ZN(n14242) );
  AOI22_X1 U15869 ( .A1(n7422), .A2(n14720), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14239) );
  OAI21_X1 U15870 ( .B1(n14690), .B2(n14290), .A(n14239), .ZN(n14240) );
  AOI21_X1 U15871 ( .B1(n14695), .B2(n14287), .A(n14240), .ZN(n14241) );
  AOI21_X1 U15872 ( .B1(n14244), .B2(n14243), .A(n14295), .ZN(n14246) );
  NAND2_X1 U15873 ( .A1(n14246), .A2(n14245), .ZN(n14250) );
  AOI22_X1 U15874 ( .A1(n7422), .A2(n14780), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14247) );
  OAI21_X1 U15875 ( .B1(n14751), .B2(n14290), .A(n14247), .ZN(n14248) );
  AOI21_X1 U15876 ( .B1(n14755), .B2(n14287), .A(n14248), .ZN(n14249) );
  OAI211_X1 U15877 ( .C1(n14934), .C2(n14282), .A(n14250), .B(n14249), .ZN(
        P3_U3173) );
  OAI211_X1 U15878 ( .C1(n14253), .C2(n14252), .A(n14251), .B(n14273), .ZN(
        n14263) );
  NAND2_X1 U15879 ( .A1(n7422), .A2(n14254), .ZN(n14255) );
  OR2_X1 U15880 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9126), .ZN(n14520) );
  OAI211_X1 U15881 ( .C1(n14290), .C2(n14256), .A(n14255), .B(n14520), .ZN(
        n14257) );
  INV_X1 U15882 ( .A(n14257), .ZN(n14262) );
  NAND2_X1 U15883 ( .A1(n14258), .A2(n14292), .ZN(n14261) );
  NAND2_X1 U15884 ( .A1(n14287), .A2(n14259), .ZN(n14260) );
  NAND4_X1 U15885 ( .A1(n14263), .A2(n14262), .A3(n14261), .A4(n14260), .ZN(
        P3_U3174) );
  INV_X1 U15886 ( .A(n14264), .ZN(n14265) );
  AOI21_X1 U15887 ( .B1(n14267), .B2(n14266), .A(n14265), .ZN(n14272) );
  AOI22_X1 U15888 ( .A1(n7422), .A2(n14719), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14269) );
  NAND2_X1 U15889 ( .A1(n14287), .A2(n14723), .ZN(n14268) );
  OAI211_X1 U15890 ( .C1(n14689), .C2(n14290), .A(n14269), .B(n14268), .ZN(
        n14270) );
  AOI21_X1 U15891 ( .B1(n14854), .B2(n14292), .A(n14270), .ZN(n14271) );
  OAI21_X1 U15892 ( .B1(n14272), .B2(n14295), .A(n14271), .ZN(P3_U3175) );
  INV_X1 U15893 ( .A(n14873), .ZN(n14283) );
  OAI211_X1 U15894 ( .C1(n14276), .C2(n14275), .A(n14274), .B(n14273), .ZN(
        n14281) );
  NAND2_X1 U15895 ( .A1(n7422), .A2(n14778), .ZN(n14278) );
  OAI211_X1 U15896 ( .C1(n14290), .C2(n14750), .A(n14278), .B(n14277), .ZN(
        n14279) );
  AOI21_X1 U15897 ( .B1(n14772), .B2(n14287), .A(n14279), .ZN(n14280) );
  OAI211_X1 U15898 ( .C1(n14283), .C2(n14282), .A(n14281), .B(n14280), .ZN(
        P3_U3178) );
  AOI21_X1 U15899 ( .B1(n14286), .B2(n14285), .A(n14284), .ZN(n14296) );
  AOI22_X1 U15900 ( .A1(n14325), .A2(n7422), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14289) );
  NAND2_X1 U15901 ( .A1(n14665), .A2(n14287), .ZN(n14288) );
  OAI211_X1 U15902 ( .C1(n14661), .C2(n14290), .A(n14289), .B(n14288), .ZN(
        n14291) );
  AOI21_X1 U15903 ( .B1(n14293), .B2(n14292), .A(n14291), .ZN(n14294) );
  OAI21_X1 U15904 ( .B1(n14296), .B2(n14295), .A(n14294), .ZN(P3_U3180) );
  OAI22_X1 U15905 ( .A1(n14297), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n14302), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U15906 ( .A1(n14300), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n14299), 
        .B2(n14298), .ZN(n14310) );
  OR2_X1 U15907 ( .A1(n14309), .A2(n14310), .ZN(n14301) );
  OAI21_X1 U15908 ( .B1(n14302), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n14301), 
        .ZN(n14305) );
  AOI22_X1 U15909 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n14303), .B2(n16163), .ZN(n14304) );
  XNOR2_X1 U15910 ( .A(n14305), .B(n14304), .ZN(n14949) );
  NAND2_X1 U15911 ( .A1(n14949), .A2(n8963), .ZN(n14308) );
  INV_X1 U15912 ( .A(SI_31_), .ZN(n14306) );
  OR2_X1 U15913 ( .A1(n9078), .A2(n14306), .ZN(n14307) );
  NAND2_X1 U15914 ( .A1(n14617), .A2(n14313), .ZN(n14498) );
  XNOR2_X1 U15915 ( .A(n14310), .B(n14309), .ZN(n14956) );
  OR2_X1 U15916 ( .A1(n9078), .A2(n14955), .ZN(n14311) );
  NAND2_X1 U15917 ( .A1(n16726), .A2(n14317), .ZN(n14457) );
  INV_X1 U15918 ( .A(n14313), .ZN(n14614) );
  NAND2_X1 U15919 ( .A1(n16726), .A2(n14614), .ZN(n14314) );
  NAND4_X1 U15920 ( .A1(n14498), .A2(n14454), .A3(n14457), .A4(n14314), .ZN(
        n14315) );
  AOI21_X1 U15921 ( .B1(n14316), .B2(n14452), .A(n14315), .ZN(n14321) );
  OR2_X1 U15922 ( .A1(n16726), .A2(n14317), .ZN(n14456) );
  INV_X1 U15923 ( .A(n14456), .ZN(n14318) );
  AND2_X1 U15924 ( .A1(n16735), .A2(n14614), .ZN(n14464) );
  INV_X1 U15925 ( .A(n14322), .ZN(n14509) );
  OAI21_X1 U15926 ( .B1(n14914), .B2(n14325), .A(n14324), .ZN(n14327) );
  AND2_X1 U15927 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  NAND2_X1 U15928 ( .A1(n14329), .A2(n14328), .ZN(n14331) );
  NAND2_X1 U15929 ( .A1(n14331), .A2(n14330), .ZN(n14334) );
  AOI21_X1 U15930 ( .B1(n14336), .B2(n14332), .A(n14334), .ZN(n14333) );
  INV_X1 U15931 ( .A(n14334), .ZN(n14338) );
  NAND2_X1 U15932 ( .A1(n14336), .A2(n14335), .ZN(n14337) );
  AOI22_X1 U15933 ( .A1(n14492), .A2(n7591), .B1(n14338), .B2(n14337), .ZN(
        n14339) );
  MUX2_X1 U15934 ( .A(n14341), .B(n14340), .S(n14455), .Z(n14443) );
  INV_X1 U15935 ( .A(n14342), .ZN(n14467) );
  OR2_X1 U15936 ( .A1(n14776), .A2(n8237), .ZN(n14488) );
  OR2_X1 U15937 ( .A1(n14488), .A2(n14343), .ZN(n14345) );
  NAND2_X1 U15938 ( .A1(n14347), .A2(n7600), .ZN(n14344) );
  NAND4_X1 U15939 ( .A1(n14467), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14352) );
  NAND3_X1 U15940 ( .A1(n14346), .A2(n14880), .A3(n14778), .ZN(n14348) );
  AND2_X1 U15941 ( .A1(n14348), .A2(n14347), .ZN(n14349) );
  OAI211_X1 U15942 ( .C1(n14350), .C2(n14488), .A(n14466), .B(n14349), .ZN(
        n14351) );
  MUX2_X1 U15943 ( .A(n14352), .B(n14351), .S(n14455), .Z(n14433) );
  NAND2_X1 U15944 ( .A1(n14404), .A2(n7598), .ZN(n14354) );
  NAND3_X1 U15945 ( .A1(n14354), .A2(n14411), .A3(n14353), .ZN(n14408) );
  AND2_X1 U15946 ( .A1(n14356), .A2(n14355), .ZN(n14361) );
  NAND2_X1 U15947 ( .A1(n14361), .A2(n14357), .ZN(n14358) );
  OAI21_X1 U15948 ( .B1(n14358), .B2(n16494), .A(n14373), .ZN(n14359) );
  NOR2_X1 U15949 ( .A1(n14360), .A2(n14359), .ZN(n14365) );
  INV_X1 U15950 ( .A(n16494), .ZN(n16489) );
  INV_X1 U15951 ( .A(n14361), .ZN(n14362) );
  NAND3_X1 U15952 ( .A1(n16489), .A2(n14363), .A3(n14362), .ZN(n14364) );
  MUX2_X1 U15953 ( .A(n14365), .B(n14364), .S(n14455), .Z(n14371) );
  INV_X1 U15954 ( .A(n14368), .ZN(n14370) );
  NAND2_X1 U15955 ( .A1(n14366), .A2(n16491), .ZN(n14367) );
  AND2_X1 U15956 ( .A1(n14368), .A2(n14367), .ZN(n14369) );
  OAI22_X1 U15957 ( .A1(n14371), .A2(n14370), .B1(n14369), .B2(n14451), .ZN(
        n14372) );
  OAI211_X1 U15958 ( .C1(n14373), .C2(n14451), .A(n14372), .B(n14470), .ZN(
        n14377) );
  MUX2_X1 U15959 ( .A(n14375), .B(n14374), .S(n14455), .Z(n14376) );
  NAND3_X1 U15960 ( .A1(n14377), .A2(n14473), .A3(n14376), .ZN(n14381) );
  MUX2_X1 U15961 ( .A(n14379), .B(n14378), .S(n14451), .Z(n14380) );
  NAND3_X1 U15962 ( .A1(n14381), .A2(n14474), .A3(n14380), .ZN(n14385) );
  MUX2_X1 U15963 ( .A(n14383), .B(n14382), .S(n14455), .Z(n14384) );
  NAND3_X1 U15964 ( .A1(n14385), .A2(n14475), .A3(n14384), .ZN(n14389) );
  MUX2_X1 U15965 ( .A(n14387), .B(n14386), .S(n14451), .Z(n14388) );
  NAND3_X1 U15966 ( .A1(n14389), .A2(n14479), .A3(n14388), .ZN(n14395) );
  INV_X1 U15967 ( .A(n14390), .ZN(n14471) );
  NAND2_X1 U15968 ( .A1(n14391), .A2(n16595), .ZN(n14392) );
  MUX2_X1 U15969 ( .A(n14393), .B(n14392), .S(n14455), .Z(n14394) );
  NAND3_X1 U15970 ( .A1(n14395), .A2(n14471), .A3(n14394), .ZN(n14401) );
  NAND2_X1 U15971 ( .A1(n14404), .A2(n14396), .ZN(n14478) );
  NOR3_X1 U15972 ( .A1(n14398), .A2(n14397), .A3(n14451), .ZN(n14399) );
  NOR2_X1 U15973 ( .A1(n14478), .A2(n14399), .ZN(n14400) );
  NAND2_X1 U15974 ( .A1(n14401), .A2(n14400), .ZN(n14409) );
  INV_X1 U15975 ( .A(n14402), .ZN(n16646) );
  NAND3_X1 U15976 ( .A1(n14404), .A2(n14403), .A3(n16646), .ZN(n14405) );
  NAND4_X1 U15977 ( .A1(n14409), .A2(n14406), .A3(n14410), .A4(n14405), .ZN(
        n14407) );
  MUX2_X1 U15978 ( .A(n14408), .B(n14407), .S(n14455), .Z(n14414) );
  NOR2_X1 U15979 ( .A1(n14409), .A2(n8254), .ZN(n14413) );
  MUX2_X1 U15980 ( .A(n14411), .B(n14410), .S(n14451), .Z(n14412) );
  OAI21_X1 U15981 ( .B1(n14414), .B2(n14413), .A(n14412), .ZN(n14415) );
  NAND2_X1 U15982 ( .A1(n14415), .A2(n14483), .ZN(n14421) );
  NAND2_X1 U15983 ( .A1(n14898), .A2(n14416), .ZN(n14417) );
  MUX2_X1 U15984 ( .A(n14418), .B(n14417), .S(n14451), .Z(n14419) );
  NAND3_X1 U15985 ( .A1(n14421), .A2(n14420), .A3(n14419), .ZN(n14425) );
  MUX2_X1 U15986 ( .A(n14423), .B(n14422), .S(n14455), .Z(n14424) );
  NAND3_X1 U15987 ( .A1(n14425), .A2(n8370), .A3(n14424), .ZN(n14430) );
  INV_X1 U15988 ( .A(n14488), .ZN(n14429) );
  OR2_X1 U15989 ( .A1(n14886), .A2(n14805), .ZN(n14427) );
  MUX2_X1 U15990 ( .A(n14427), .B(n14426), .S(n14455), .Z(n14428) );
  AND4_X1 U15991 ( .A1(n14430), .A2(n14429), .A3(n14803), .A4(n14428), .ZN(
        n14432) );
  MUX2_X1 U15992 ( .A(n14466), .B(n14467), .S(n14455), .Z(n14431) );
  OAI211_X1 U15993 ( .C1(n14433), .C2(n14432), .A(n9365), .B(n14431), .ZN(
        n14437) );
  MUX2_X1 U15994 ( .A(n14435), .B(n14434), .S(n14451), .Z(n14436) );
  NAND3_X1 U15995 ( .A1(n14437), .A2(n14436), .A3(n14733), .ZN(n14441) );
  MUX2_X1 U15996 ( .A(n14439), .B(n14438), .S(n14455), .Z(n14440) );
  NAND3_X1 U15997 ( .A1(n14493), .A2(n14441), .A3(n14440), .ZN(n14442) );
  NAND4_X1 U15998 ( .A1(n14492), .A2(n14700), .A3(n14443), .A4(n14442), .ZN(
        n14444) );
  INV_X1 U15999 ( .A(n14445), .ZN(n14447) );
  MUX2_X1 U16000 ( .A(n14447), .B(n14446), .S(n14455), .Z(n14448) );
  NOR2_X1 U16001 ( .A1(n14495), .A2(n14448), .ZN(n14449) );
  NAND2_X1 U16002 ( .A1(n14456), .A2(n14457), .ZN(n14496) );
  AOI21_X1 U16003 ( .B1(n14450), .B2(n14449), .A(n14496), .ZN(n14453) );
  NAND3_X1 U16004 ( .A1(n14453), .A2(n14452), .A3(n14451), .ZN(n14463) );
  INV_X1 U16005 ( .A(n14453), .ZN(n14461) );
  INV_X1 U16006 ( .A(n14454), .ZN(n14460) );
  NAND2_X1 U16007 ( .A1(n14456), .A2(n14455), .ZN(n14458) );
  NAND2_X1 U16008 ( .A1(n14458), .A2(n14457), .ZN(n14459) );
  OAI21_X1 U16009 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(n14462) );
  NAND3_X1 U16010 ( .A1(n14463), .A2(n14498), .A3(n14462), .ZN(n14465) );
  INV_X1 U16011 ( .A(n14464), .ZN(n14497) );
  NAND2_X1 U16012 ( .A1(n14465), .A2(n14497), .ZN(n14506) );
  NAND2_X1 U16013 ( .A1(n14467), .A2(n14466), .ZN(n14765) );
  INV_X1 U16014 ( .A(n12707), .ZN(n14469) );
  NAND4_X1 U16015 ( .A1(n14471), .A2(n14470), .A3(n14469), .A4(n14468), .ZN(
        n14477) );
  NAND4_X1 U16016 ( .A1(n14475), .A2(n14474), .A3(n14473), .A4(n14472), .ZN(
        n14476) );
  NOR2_X1 U16017 ( .A1(n14477), .A2(n14476), .ZN(n14482) );
  INV_X1 U16018 ( .A(n14478), .ZN(n14481) );
  AND2_X1 U16019 ( .A1(n16489), .A2(n14479), .ZN(n14480) );
  NAND4_X1 U16020 ( .A1(n14482), .A2(n14822), .A3(n14481), .A4(n14480), .ZN(
        n14485) );
  NOR3_X1 U16021 ( .A1(n14485), .A2(n14484), .A3(n9133), .ZN(n14486) );
  NAND3_X1 U16022 ( .A1(n14803), .A2(n14486), .A3(n8370), .ZN(n14487) );
  OR2_X1 U16023 ( .A1(n14488), .A2(n14487), .ZN(n14489) );
  NOR2_X1 U16024 ( .A1(n14765), .A2(n14489), .ZN(n14490) );
  AND3_X1 U16025 ( .A1(n9365), .A2(n14733), .A3(n14490), .ZN(n14491) );
  NAND4_X1 U16026 ( .A1(n14700), .A2(n14493), .A3(n14492), .A4(n14491), .ZN(
        n14494) );
  NAND3_X1 U16027 ( .A1(n14499), .A2(n14498), .A3(n14497), .ZN(n14501) );
  XNOR2_X1 U16028 ( .A(n14501), .B(n14500), .ZN(n14502) );
  AOI22_X1 U16029 ( .A1(n14506), .A2(n14504), .B1(n14503), .B2(n14502), .ZN(
        n14505) );
  OAI21_X1 U16030 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n14508) );
  NOR3_X1 U16031 ( .A1(n14511), .A2(n14594), .A3(n14510), .ZN(n14514) );
  OAI21_X1 U16032 ( .B1(n14515), .B2(n14512), .A(P3_B_REG_SCAN_IN), .ZN(n14513) );
  OAI21_X1 U16033 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(n14519) );
  NAND2_X1 U16034 ( .A1(n14519), .A2(n14604), .ZN(n14530) );
  OAI21_X1 U16035 ( .B1(n7608), .B2(P3_REG1_REG_13__SCAN_IN), .A(n7455), .ZN(
        n14527) );
  INV_X1 U16036 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n16410) );
  OAI21_X1 U16037 ( .B1(n14572), .B2(n16410), .A(n14520), .ZN(n14526) );
  AOI21_X1 U16038 ( .B1(n14523), .B2(n14522), .A(n14521), .ZN(n14524) );
  NOR2_X1 U16039 ( .A1(n14541), .A2(n14524), .ZN(n14525) );
  AOI211_X1 U16040 ( .C1(n14528), .C2(n14527), .A(n14526), .B(n14525), .ZN(
        n14529) );
  OAI211_X1 U16041 ( .C1(n14606), .C2(n14531), .A(n14530), .B(n14529), .ZN(
        P3_U3195) );
  AOI21_X1 U16042 ( .B1(n14534), .B2(n14533), .A(n14532), .ZN(n14549) );
  AOI21_X1 U16043 ( .B1(n14537), .B2(n14536), .A(n14535), .ZN(n14540) );
  INV_X1 U16044 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n16414) );
  OR2_X1 U16045 ( .A1(n14572), .A2(n16414), .ZN(n14538) );
  OAI211_X1 U16046 ( .C1(n14541), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        n14546) );
  AOI211_X1 U16047 ( .C1(n14544), .C2(n14543), .A(n14574), .B(n14542), .ZN(
        n14545) );
  AOI211_X1 U16048 ( .C1(n14580), .C2(n14547), .A(n14546), .B(n14545), .ZN(
        n14548) );
  OAI21_X1 U16049 ( .B1(n14549), .B2(n14611), .A(n14548), .ZN(P3_U3196) );
  AOI21_X1 U16050 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14567) );
  INV_X1 U16051 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14560) );
  AND2_X1 U16052 ( .A1(n14555), .A2(n14554), .ZN(n14556) );
  OAI21_X1 U16053 ( .B1(n14557), .B2(n14556), .A(n14603), .ZN(n14559) );
  OAI211_X1 U16054 ( .C1(n14560), .C2(n14572), .A(n14559), .B(n14558), .ZN(
        n14565) );
  AOI211_X1 U16055 ( .C1(n14563), .C2(n14562), .A(n14574), .B(n14561), .ZN(
        n14564) );
  AOI211_X1 U16056 ( .C1(n14580), .C2(n7899), .A(n14565), .B(n14564), .ZN(
        n14566) );
  OAI21_X1 U16057 ( .B1(n14567), .B2(n14611), .A(n14566), .ZN(P3_U3198) );
  AOI21_X1 U16058 ( .B1(n14570), .B2(n14569), .A(n14568), .ZN(n14586) );
  INV_X1 U16059 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n16449) );
  OAI21_X1 U16060 ( .B1(n14572), .B2(n16449), .A(n14571), .ZN(n14578) );
  AOI211_X1 U16061 ( .C1(n14576), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14577) );
  AOI211_X1 U16062 ( .C1(n14580), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        n14585) );
  INV_X1 U16063 ( .A(n14581), .ZN(n14582) );
  NOR2_X1 U16064 ( .A1(n14582), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n14583) );
  OAI21_X1 U16065 ( .B1(n14583), .B2(n8331), .A(n14603), .ZN(n14584) );
  OAI211_X1 U16066 ( .C1(n14586), .C2(n14611), .A(n14585), .B(n14584), .ZN(
        P3_U3199) );
  XNOR2_X1 U16067 ( .A(n14605), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n14595) );
  XNOR2_X1 U16068 ( .A(n14589), .B(n14595), .ZN(n14612) );
  INV_X1 U16069 ( .A(n14590), .ZN(n14592) );
  XNOR2_X1 U16070 ( .A(n14605), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n14600) );
  MUX2_X1 U16071 ( .A(n14595), .B(n14600), .S(n14594), .Z(n14596) );
  INV_X1 U16072 ( .A(n14597), .ZN(n14598) );
  NOR2_X1 U16073 ( .A1(n14599), .A2(n14598), .ZN(n14601) );
  XNOR2_X1 U16074 ( .A(n14601), .B(n14600), .ZN(n14602) );
  NOR2_X1 U16075 ( .A1(n14606), .A2(n14605), .ZN(n14607) );
  AOI211_X1 U16076 ( .C1(P3_ADDR_REG_19__SCAN_IN), .C2(n14609), .A(n14608), 
        .B(n14607), .ZN(n14610) );
  NOR2_X1 U16077 ( .A1(n14614), .A2(n14613), .ZN(n16728) );
  OAI21_X1 U16078 ( .B1(n14615), .B2(n14792), .A(n14819), .ZN(n14622) );
  NOR2_X1 U16079 ( .A1(n16728), .A2(n14622), .ZN(n14619) );
  NOR2_X1 U16080 ( .A1(n14819), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n14616) );
  OAI22_X1 U16081 ( .A1(n14617), .A2(n14809), .B1(n14619), .B2(n14616), .ZN(
        P3_U3202) );
  INV_X1 U16082 ( .A(n16726), .ZN(n14620) );
  NOR2_X1 U16083 ( .A1(n14819), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n14618) );
  OAI22_X1 U16084 ( .A1(n14620), .A2(n14809), .B1(n14619), .B2(n14618), .ZN(
        P3_U3203) );
  INV_X1 U16085 ( .A(n14621), .ZN(n14623) );
  OAI22_X1 U16086 ( .A1(n14623), .A2(n14622), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14819), .ZN(n14626) );
  NAND2_X1 U16087 ( .A1(n14624), .A2(n14821), .ZN(n14625) );
  OAI211_X1 U16088 ( .C1(n14627), .C2(n14813), .A(n14626), .B(n14625), .ZN(
        P3_U3204) );
  OAI211_X1 U16089 ( .C1(n14629), .C2(n14634), .A(n14628), .B(n16500), .ZN(
        n14631) );
  OR2_X1 U16090 ( .A1(n14661), .A2(n16495), .ZN(n14630) );
  OAI211_X1 U16091 ( .C1(n14632), .C2(n16497), .A(n14631), .B(n14630), .ZN(
        n14829) );
  NAND2_X1 U16092 ( .A1(n14829), .A2(n14819), .ZN(n14642) );
  AOI22_X1 U16093 ( .A1(n14633), .A2(n16508), .B1(n16517), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n14641) );
  AND2_X1 U16094 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  NAND2_X1 U16095 ( .A1(n14830), .A2(n14824), .ZN(n14640) );
  NAND2_X1 U16096 ( .A1(n14638), .A2(n14821), .ZN(n14639) );
  NAND4_X1 U16097 ( .A1(n14642), .A2(n14641), .A3(n14640), .A4(n14639), .ZN(
        P3_U3205) );
  AOI21_X1 U16098 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n14653) );
  OAI22_X1 U16099 ( .A1(n14647), .A2(n16497), .B1(n14646), .B2(n16495), .ZN(
        n14648) );
  INV_X1 U16100 ( .A(n14648), .ZN(n14652) );
  NAND2_X1 U16101 ( .A1(n8261), .A2(n7777), .ZN(n14649) );
  NAND2_X1 U16102 ( .A1(n14650), .A2(n14649), .ZN(n14833) );
  NAND2_X1 U16103 ( .A1(n14833), .A2(n16678), .ZN(n14651) );
  NAND2_X1 U16104 ( .A1(n14832), .A2(n14819), .ZN(n14659) );
  AOI22_X1 U16105 ( .A1(n14654), .A2(n16508), .B1(n16517), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n14658) );
  NAND2_X1 U16106 ( .A1(n14833), .A2(n14758), .ZN(n14657) );
  NAND2_X1 U16107 ( .A1(n14655), .A2(n14821), .ZN(n14656) );
  NAND4_X1 U16108 ( .A1(n14659), .A2(n14658), .A3(n14657), .A4(n14656), .ZN(
        P3_U3206) );
  XOR2_X1 U16109 ( .A(n14664), .B(n14660), .Z(n14662) );
  OAI222_X1 U16110 ( .A1(n14662), .A2(n14817), .B1(n16497), .B2(n14661), .C1(
        n16495), .C2(n14690), .ZN(n14836) );
  INV_X1 U16111 ( .A(n14836), .ZN(n14669) );
  XOR2_X1 U16112 ( .A(n14664), .B(n14663), .Z(n14837) );
  AOI22_X1 U16113 ( .A1(n16508), .A2(n14665), .B1(n16517), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n14666) );
  OAI21_X1 U16114 ( .B1(n14910), .B2(n14809), .A(n14666), .ZN(n14667) );
  AOI21_X1 U16115 ( .B1(n14837), .B2(n14824), .A(n14667), .ZN(n14668) );
  OAI21_X1 U16116 ( .B1(n14669), .B2(n16517), .A(n14668), .ZN(P3_U3207) );
  NAND2_X1 U16117 ( .A1(n14670), .A2(n14682), .ZN(n14671) );
  NAND3_X1 U16118 ( .A1(n14672), .A2(n16500), .A3(n14671), .ZN(n14676) );
  AOI22_X1 U16119 ( .A1(n14779), .A2(n14674), .B1(n14673), .B2(n14777), .ZN(
        n14675) );
  INV_X1 U16120 ( .A(n14677), .ZN(n14679) );
  INV_X1 U16121 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n14678) );
  OAI22_X1 U16122 ( .A1(n14679), .A2(n14792), .B1(n14678), .B2(n14819), .ZN(
        n14680) );
  AOI21_X1 U16123 ( .B1(n14681), .B2(n14821), .A(n14680), .ZN(n14685) );
  XNOR2_X1 U16124 ( .A(n14683), .B(n8344), .ZN(n14840) );
  NAND2_X1 U16125 ( .A1(n14840), .A2(n14824), .ZN(n14684) );
  OAI211_X1 U16126 ( .C1(n14842), .C2(n16517), .A(n14685), .B(n14684), .ZN(
        P3_U3208) );
  XNOR2_X1 U16127 ( .A(n14686), .B(n14687), .ZN(n14694) );
  XNOR2_X1 U16128 ( .A(n14688), .B(n14687), .ZN(n14692) );
  OAI22_X1 U16129 ( .A1(n14690), .A2(n16497), .B1(n14689), .B2(n16495), .ZN(
        n14691) );
  AOI21_X1 U16130 ( .B1(n14692), .B2(n16500), .A(n14691), .ZN(n14693) );
  OAI21_X1 U16131 ( .B1(n16503), .B2(n14694), .A(n14693), .ZN(n14845) );
  INV_X1 U16132 ( .A(n14845), .ZN(n14699) );
  INV_X1 U16133 ( .A(n14694), .ZN(n14846) );
  AOI22_X1 U16134 ( .A1(n16517), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n16508), 
        .B2(n14695), .ZN(n14696) );
  OAI21_X1 U16135 ( .B1(n14918), .B2(n14809), .A(n14696), .ZN(n14697) );
  AOI21_X1 U16136 ( .B1(n14846), .B2(n14758), .A(n14697), .ZN(n14698) );
  OAI21_X1 U16137 ( .B1(n14699), .B2(n16517), .A(n14698), .ZN(P3_U3209) );
  XNOR2_X1 U16138 ( .A(n14701), .B(n14700), .ZN(n14704) );
  OAI22_X1 U16139 ( .A1(n14702), .A2(n16497), .B1(n14737), .B2(n16495), .ZN(
        n14703) );
  AOI21_X1 U16140 ( .B1(n14704), .B2(n16500), .A(n14703), .ZN(n14851) );
  XNOR2_X1 U16141 ( .A(n14706), .B(n14705), .ZN(n14849) );
  AOI22_X1 U16142 ( .A1(n16517), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n16508), 
        .B2(n14707), .ZN(n14708) );
  OAI21_X1 U16143 ( .B1(n14922), .B2(n14809), .A(n14708), .ZN(n14709) );
  AOI21_X1 U16144 ( .B1(n14849), .B2(n14824), .A(n14709), .ZN(n14710) );
  OAI21_X1 U16145 ( .B1(n14851), .B2(n16517), .A(n14710), .ZN(P3_U3210) );
  NAND2_X1 U16146 ( .A1(n14711), .A2(n14716), .ZN(n14712) );
  NAND2_X1 U16147 ( .A1(n14713), .A2(n14712), .ZN(n14855) );
  INV_X1 U16148 ( .A(n14758), .ZN(n14729) );
  NAND2_X1 U16149 ( .A1(n14715), .A2(n14714), .ZN(n14717) );
  XNOR2_X1 U16150 ( .A(n14717), .B(n14716), .ZN(n14718) );
  NAND2_X1 U16151 ( .A1(n14718), .A2(n16500), .ZN(n14722) );
  AOI22_X1 U16152 ( .A1(n14720), .A2(n14779), .B1(n14777), .B2(n14719), .ZN(
        n14721) );
  OAI211_X1 U16153 ( .C1(n16503), .C2(n14855), .A(n14722), .B(n14721), .ZN(
        n14856) );
  NAND2_X1 U16154 ( .A1(n14856), .A2(n14819), .ZN(n14728) );
  INV_X1 U16155 ( .A(n14723), .ZN(n14724) );
  OAI22_X1 U16156 ( .A1(n14819), .A2(n14725), .B1(n14724), .B2(n14792), .ZN(
        n14726) );
  AOI21_X1 U16157 ( .B1(n14854), .B2(n14821), .A(n14726), .ZN(n14727) );
  OAI211_X1 U16158 ( .C1(n14855), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        P3_U3211) );
  NAND2_X1 U16159 ( .A1(n14731), .A2(n14730), .ZN(n14732) );
  XOR2_X1 U16160 ( .A(n14733), .B(n14732), .Z(n14740) );
  OR2_X1 U16161 ( .A1(n14734), .A2(n14733), .ZN(n14735) );
  NAND2_X1 U16162 ( .A1(n14736), .A2(n14735), .ZN(n14861) );
  OAI22_X1 U16163 ( .A1(n14737), .A2(n16497), .B1(n14763), .B2(n16495), .ZN(
        n14738) );
  AOI21_X1 U16164 ( .B1(n14861), .B2(n16678), .A(n14738), .ZN(n14739) );
  OAI21_X1 U16165 ( .B1(n14740), .B2(n14817), .A(n14739), .ZN(n14860) );
  INV_X1 U16166 ( .A(n14860), .ZN(n14745) );
  AOI22_X1 U16167 ( .A1(n16517), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n16508), 
        .B2(n14741), .ZN(n14742) );
  OAI21_X1 U16168 ( .B1(n14930), .B2(n14809), .A(n14742), .ZN(n14743) );
  AOI21_X1 U16169 ( .B1(n14861), .B2(n14758), .A(n14743), .ZN(n14744) );
  OAI21_X1 U16170 ( .B1(n14745), .B2(n16517), .A(n14744), .ZN(P3_U3212) );
  XNOR2_X1 U16171 ( .A(n14747), .B(n14746), .ZN(n14754) );
  OAI21_X1 U16172 ( .B1(n14749), .B2(n9365), .A(n14748), .ZN(n14865) );
  OAI22_X1 U16173 ( .A1(n14751), .A2(n16497), .B1(n14750), .B2(n16495), .ZN(
        n14752) );
  AOI21_X1 U16174 ( .B1(n14865), .B2(n16678), .A(n14752), .ZN(n14753) );
  OAI21_X1 U16175 ( .B1(n14754), .B2(n14817), .A(n14753), .ZN(n14864) );
  INV_X1 U16176 ( .A(n14864), .ZN(n14760) );
  AOI22_X1 U16177 ( .A1(n16517), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n16508), 
        .B2(n14755), .ZN(n14756) );
  OAI21_X1 U16178 ( .B1(n14934), .B2(n14809), .A(n14756), .ZN(n14757) );
  AOI21_X1 U16179 ( .B1(n14865), .B2(n14758), .A(n14757), .ZN(n14759) );
  OAI21_X1 U16180 ( .B1(n14760), .B2(n16517), .A(n14759), .ZN(P3_U3213) );
  XOR2_X1 U16181 ( .A(n14765), .B(n14761), .Z(n14762) );
  OAI222_X1 U16182 ( .A1(n16497), .A2(n14763), .B1(n16495), .B2(n14786), .C1(
        n14762), .C2(n14817), .ZN(n14868) );
  INV_X1 U16183 ( .A(n14868), .ZN(n14770) );
  XOR2_X1 U16184 ( .A(n14765), .B(n14764), .Z(n14869) );
  AOI22_X1 U16185 ( .A1(n16517), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n16508), 
        .B2(n14766), .ZN(n14767) );
  OAI21_X1 U16186 ( .B1(n14939), .B2(n14809), .A(n14767), .ZN(n14768) );
  AOI21_X1 U16187 ( .B1(n14869), .B2(n14824), .A(n14768), .ZN(n14769) );
  OAI21_X1 U16188 ( .B1(n14770), .B2(n16517), .A(n14769), .ZN(P3_U3214) );
  XNOR2_X1 U16189 ( .A(n14771), .B(n14776), .ZN(n14876) );
  INV_X1 U16190 ( .A(n14772), .ZN(n14773) );
  OAI22_X1 U16191 ( .A1(n14819), .A2(n14774), .B1(n14773), .B2(n14792), .ZN(
        n14783) );
  OAI21_X1 U16192 ( .B1(n7566), .B2(n14776), .A(n14775), .ZN(n14781) );
  AOI222_X1 U16193 ( .A1(n14781), .A2(n16500), .B1(n14780), .B2(n14779), .C1(
        n14778), .C2(n14777), .ZN(n14875) );
  NOR2_X1 U16194 ( .A1(n14875), .A2(n16517), .ZN(n14782) );
  AOI211_X1 U16195 ( .C1(n14821), .C2(n14873), .A(n14783), .B(n14782), .ZN(
        n14784) );
  OAI21_X1 U16196 ( .B1(n14813), .B2(n14876), .A(n14784), .ZN(P3_U3215) );
  AOI21_X1 U16197 ( .B1(n14785), .B2(n14797), .A(n14817), .ZN(n14790) );
  OAI22_X1 U16198 ( .A1(n14787), .A2(n16495), .B1(n14786), .B2(n16497), .ZN(
        n14788) );
  AOI21_X1 U16199 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14879) );
  INV_X1 U16200 ( .A(n14791), .ZN(n14793) );
  OAI22_X1 U16201 ( .A1(n14819), .A2(n14794), .B1(n14793), .B2(n14792), .ZN(
        n14795) );
  AOI21_X1 U16202 ( .B1(n14796), .B2(n14821), .A(n14795), .ZN(n14800) );
  XNOR2_X1 U16203 ( .A(n14798), .B(n14797), .ZN(n14877) );
  NAND2_X1 U16204 ( .A1(n14877), .A2(n14824), .ZN(n14799) );
  OAI211_X1 U16205 ( .C1(n14879), .C2(n16517), .A(n14800), .B(n14799), .ZN(
        P3_U3216) );
  XOR2_X1 U16206 ( .A(n14801), .B(n14803), .Z(n14884) );
  AOI21_X1 U16207 ( .B1(n14803), .B2(n14802), .A(n7610), .ZN(n14804) );
  OAI222_X1 U16208 ( .A1(n16497), .A2(n14806), .B1(n16495), .B2(n14805), .C1(
        n14804), .C2(n14817), .ZN(n14881) );
  AOI22_X1 U16209 ( .A1(n16517), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n16508), 
        .B2(n14807), .ZN(n14808) );
  OAI21_X1 U16210 ( .B1(n14810), .B2(n14809), .A(n14808), .ZN(n14811) );
  AOI21_X1 U16211 ( .B1(n14881), .B2(n14819), .A(n14811), .ZN(n14812) );
  OAI21_X1 U16212 ( .B1(n14813), .B2(n14884), .A(n14812), .ZN(P3_U3217) );
  XOR2_X1 U16213 ( .A(n14822), .B(n14814), .Z(n14818) );
  OAI222_X1 U16214 ( .A1(n14818), .A2(n14817), .B1(n16497), .B2(n14816), .C1(
        n16495), .C2(n14815), .ZN(n16671) );
  NAND2_X1 U16215 ( .A1(n16671), .A2(n14819), .ZN(n14828) );
  AOI22_X1 U16216 ( .A1(n14821), .A2(n16673), .B1(n16508), .B2(n14820), .ZN(
        n14827) );
  XOR2_X1 U16217 ( .A(n14823), .B(n14822), .Z(n16675) );
  INV_X1 U16218 ( .A(n16675), .ZN(n16679) );
  NAND2_X1 U16219 ( .A1(n16679), .A2(n14824), .ZN(n14826) );
  NAND2_X1 U16220 ( .A1(n16517), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n14825) );
  NAND4_X1 U16221 ( .A1(n14828), .A2(n14827), .A3(n14826), .A4(n14825), .ZN(
        P3_U3221) );
  MUX2_X1 U16222 ( .A(n14834), .B(n14903), .S(n16724), .Z(n14835) );
  INV_X1 U16223 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14838) );
  AOI21_X1 U16224 ( .B1(n16666), .B2(n14837), .A(n14836), .ZN(n14907) );
  MUX2_X1 U16225 ( .A(n14838), .B(n14907), .S(n16724), .Z(n14839) );
  OAI21_X1 U16226 ( .B1(n14910), .B2(n14872), .A(n14839), .ZN(P3_U3485) );
  NAND2_X1 U16227 ( .A1(n14840), .A2(n16666), .ZN(n14841) );
  NAND2_X1 U16228 ( .A1(n14842), .A2(n14841), .ZN(n14911) );
  MUX2_X1 U16229 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n14911), .S(n16724), .Z(
        n14843) );
  INV_X1 U16230 ( .A(n14843), .ZN(n14844) );
  OAI21_X1 U16231 ( .B1(n14914), .B2(n14872), .A(n14844), .ZN(P3_U3484) );
  AOI21_X1 U16232 ( .B1(n16643), .B2(n14846), .A(n14845), .ZN(n14915) );
  MUX2_X1 U16233 ( .A(n14847), .B(n14915), .S(n16724), .Z(n14848) );
  OAI21_X1 U16234 ( .B1(n14872), .B2(n14918), .A(n14848), .ZN(P3_U3483) );
  NAND2_X1 U16235 ( .A1(n14849), .A2(n16666), .ZN(n14850) );
  NAND2_X1 U16236 ( .A1(n14851), .A2(n14850), .ZN(n14919) );
  MUX2_X1 U16237 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n14919), .S(n16724), .Z(
        n14852) );
  INV_X1 U16238 ( .A(n14852), .ZN(n14853) );
  OAI21_X1 U16239 ( .B1(n14922), .B2(n14872), .A(n14853), .ZN(P3_U3482) );
  INV_X1 U16240 ( .A(n14854), .ZN(n14926) );
  INV_X1 U16241 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n14858) );
  INV_X1 U16242 ( .A(n14855), .ZN(n14857) );
  AOI21_X1 U16243 ( .B1(n16643), .B2(n14857), .A(n14856), .ZN(n14923) );
  MUX2_X1 U16244 ( .A(n14858), .B(n14923), .S(n16724), .Z(n14859) );
  OAI21_X1 U16245 ( .B1(n14926), .B2(n14872), .A(n14859), .ZN(P3_U3481) );
  INV_X1 U16246 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14862) );
  AOI21_X1 U16247 ( .B1(n16643), .B2(n14861), .A(n14860), .ZN(n14927) );
  MUX2_X1 U16248 ( .A(n14862), .B(n14927), .S(n16724), .Z(n14863) );
  OAI21_X1 U16249 ( .B1(n14930), .B2(n14872), .A(n14863), .ZN(P3_U3480) );
  INV_X1 U16250 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n14866) );
  AOI21_X1 U16251 ( .B1(n16643), .B2(n14865), .A(n14864), .ZN(n14931) );
  MUX2_X1 U16252 ( .A(n14866), .B(n14931), .S(n16724), .Z(n14867) );
  OAI21_X1 U16253 ( .B1(n14934), .B2(n14872), .A(n14867), .ZN(P3_U3479) );
  INV_X1 U16254 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14870) );
  AOI21_X1 U16255 ( .B1(n14869), .B2(n16666), .A(n14868), .ZN(n14935) );
  MUX2_X1 U16256 ( .A(n14870), .B(n14935), .S(n16724), .Z(n14871) );
  OAI21_X1 U16257 ( .B1(n14939), .B2(n14872), .A(n14871), .ZN(P3_U3478) );
  NAND2_X1 U16258 ( .A1(n14873), .A2(n16672), .ZN(n14874) );
  OAI211_X1 U16259 ( .C1(n14894), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        n14940) );
  MUX2_X1 U16260 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n14940), .S(n16724), .Z(
        P3_U3477) );
  NAND2_X1 U16261 ( .A1(n14877), .A2(n16666), .ZN(n14878) );
  OAI211_X1 U16262 ( .C1(n14880), .C2(n16663), .A(n14879), .B(n14878), .ZN(
        n14941) );
  MUX2_X1 U16263 ( .A(n14941), .B(P3_REG1_REG_17__SCAN_IN), .S(n7821), .Z(
        P3_U3476) );
  AOI21_X1 U16264 ( .B1(n16672), .B2(n14882), .A(n14881), .ZN(n14883) );
  OAI21_X1 U16265 ( .B1(n14894), .B2(n14884), .A(n14883), .ZN(n14942) );
  MUX2_X1 U16266 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n14942), .S(n16724), .Z(
        P3_U3475) );
  AOI21_X1 U16267 ( .B1(n16672), .B2(n14886), .A(n14885), .ZN(n14887) );
  OAI21_X1 U16268 ( .B1(n14894), .B2(n14888), .A(n14887), .ZN(n14943) );
  MUX2_X1 U16269 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n14943), .S(n16724), .Z(
        P3_U3474) );
  INV_X1 U16270 ( .A(n14889), .ZN(n14891) );
  AOI21_X1 U16271 ( .B1(n14891), .B2(n16672), .A(n14890), .ZN(n14892) );
  OAI21_X1 U16272 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(n14944) );
  MUX2_X1 U16273 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n14944), .S(n16724), .Z(
        P3_U3473) );
  NAND2_X1 U16274 ( .A1(n14895), .A2(n16666), .ZN(n14896) );
  OAI211_X1 U16275 ( .C1(n16663), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        n14945) );
  MUX2_X1 U16276 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n14945), .S(n16724), .Z(
        P3_U3472) );
  INV_X1 U16277 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n14900) );
  MUX2_X1 U16278 ( .A(n14900), .B(n14899), .S(n16727), .Z(n14901) );
  INV_X1 U16279 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n14904) );
  MUX2_X1 U16280 ( .A(n14904), .B(n14903), .S(n16727), .Z(n14905) );
  INV_X1 U16281 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14908) );
  MUX2_X1 U16282 ( .A(n14908), .B(n14907), .S(n16727), .Z(n14909) );
  OAI21_X1 U16283 ( .B1(n14910), .B2(n14938), .A(n14909), .ZN(P3_U3453) );
  MUX2_X1 U16284 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n14911), .S(n16727), .Z(
        n14912) );
  INV_X1 U16285 ( .A(n14912), .ZN(n14913) );
  OAI21_X1 U16286 ( .B1(n14914), .B2(n14938), .A(n14913), .ZN(P3_U3452) );
  INV_X1 U16287 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14916) );
  MUX2_X1 U16288 ( .A(n14916), .B(n14915), .S(n16727), .Z(n14917) );
  OAI21_X1 U16289 ( .B1(n14938), .B2(n14918), .A(n14917), .ZN(P3_U3451) );
  MUX2_X1 U16290 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n14919), .S(n16727), .Z(
        n14920) );
  INV_X1 U16291 ( .A(n14920), .ZN(n14921) );
  OAI21_X1 U16292 ( .B1(n14922), .B2(n14938), .A(n14921), .ZN(P3_U3450) );
  INV_X1 U16293 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14924) );
  MUX2_X1 U16294 ( .A(n14924), .B(n14923), .S(n16727), .Z(n14925) );
  OAI21_X1 U16295 ( .B1(n14926), .B2(n14938), .A(n14925), .ZN(P3_U3449) );
  INV_X1 U16296 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14928) );
  MUX2_X1 U16297 ( .A(n14928), .B(n14927), .S(n16727), .Z(n14929) );
  OAI21_X1 U16298 ( .B1(n14930), .B2(n14938), .A(n14929), .ZN(P3_U3448) );
  INV_X1 U16299 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14932) );
  MUX2_X1 U16300 ( .A(n14932), .B(n14931), .S(n16727), .Z(n14933) );
  OAI21_X1 U16301 ( .B1(n14934), .B2(n14938), .A(n14933), .ZN(P3_U3447) );
  INV_X1 U16302 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14936) );
  MUX2_X1 U16303 ( .A(n14936), .B(n14935), .S(n16727), .Z(n14937) );
  OAI21_X1 U16304 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(P3_U3446) );
  MUX2_X1 U16305 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n14940), .S(n16727), .Z(
        P3_U3444) );
  MUX2_X1 U16306 ( .A(n14941), .B(P3_REG0_REG_17__SCAN_IN), .S(n16733), .Z(
        P3_U3441) );
  MUX2_X1 U16307 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n14942), .S(n16727), .Z(
        P3_U3438) );
  MUX2_X1 U16308 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n14943), .S(n16727), .Z(
        P3_U3435) );
  MUX2_X1 U16309 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n14944), .S(n16727), .Z(
        P3_U3432) );
  MUX2_X1 U16310 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n14945), .S(n16727), .Z(
        P3_U3429) );
  MUX2_X1 U16311 ( .A(n14946), .B(P3_D_REG_1__SCAN_IN), .S(n14947), .Z(
        P3_U3377) );
  MUX2_X1 U16312 ( .A(n14948), .B(P3_D_REG_0__SCAN_IN), .S(n14947), .Z(
        P3_U3376) );
  INV_X1 U16313 ( .A(n14949), .ZN(n14954) );
  NOR4_X1 U16314 ( .A1(n14950), .A2(P3_IR_REG_30__SCAN_IN), .A3(n9386), .A4(
        P3_U3151), .ZN(n14951) );
  AOI21_X1 U16315 ( .B1(SI_31_), .B2(n14952), .A(n14951), .ZN(n14953) );
  OAI21_X1 U16316 ( .B1(n14954), .B2(n14968), .A(n14953), .ZN(P3_U3264) );
  OAI222_X1 U16317 ( .A1(P3_U3151), .A2(n14957), .B1(n14968), .B2(n14956), 
        .C1(n14955), .C2(n14959), .ZN(P3_U3265) );
  INV_X1 U16318 ( .A(n14958), .ZN(n14961) );
  OAI222_X1 U16319 ( .A1(P3_U3151), .A2(n14962), .B1(n14968), .B2(n14961), 
        .C1(n14960), .C2(n14959), .ZN(P3_U3266) );
  INV_X1 U16320 ( .A(n14963), .ZN(n14965) );
  OAI222_X1 U16321 ( .A1(n14968), .A2(n14965), .B1(n14959), .B2(n14964), .C1(
        P3_U3151), .C2(n10915), .ZN(P3_U3268) );
  INV_X1 U16322 ( .A(n14966), .ZN(n14967) );
  OAI222_X1 U16323 ( .A1(P3_U3151), .A2(n14970), .B1(n14959), .B2(n14969), 
        .C1(n14968), .C2(n14967), .ZN(P3_U3269) );
  AOI22_X1 U16324 ( .A1(n15225), .A2(n15219), .B1(n15226), .B2(n15073), .ZN(
        n15270) );
  NAND2_X1 U16325 ( .A1(n15478), .A2(n15080), .ZN(n14975) );
  AOI22_X1 U16326 ( .A1(n15264), .A2(n15074), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14974) );
  OAI211_X1 U16327 ( .C1(n15270), .C2(n15076), .A(n14975), .B(n14974), .ZN(
        n14976) );
  AOI22_X1 U16328 ( .A1(n14977), .A2(n15070), .B1(n15050), .B2(n15216), .ZN(
        n14982) );
  AND2_X1 U16329 ( .A1(n15215), .A2(n15225), .ZN(n14978) );
  AOI21_X1 U16330 ( .B1(n15191), .B2(n15073), .A(n14978), .ZN(n15325) );
  AOI22_X1 U16331 ( .A1(n15329), .A2(n15074), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14979) );
  OAI21_X1 U16332 ( .B1(n15325), .B2(n15076), .A(n14979), .ZN(n14980) );
  AOI21_X1 U16333 ( .B1(n15503), .B2(n15080), .A(n14980), .ZN(n14981) );
  OAI21_X1 U16334 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(P2_U3188) );
  INV_X1 U16335 ( .A(n14984), .ZN(n14985) );
  AOI21_X1 U16336 ( .B1(n14985), .B2(n15061), .A(n15077), .ZN(n14988) );
  NOR3_X1 U16337 ( .A1(n14986), .A2(n15203), .A3(n15067), .ZN(n14987) );
  OAI21_X1 U16338 ( .B1(n14988), .B2(n14987), .A(n15037), .ZN(n14991) );
  OAI22_X1 U16339 ( .A1(n15183), .A2(n15162), .B1(n15203), .B2(n15043), .ZN(
        n15393) );
  AND2_X1 U16340 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n15147) );
  NOR2_X1 U16341 ( .A1(n15052), .A2(n15387), .ZN(n14989) );
  AOI211_X1 U16342 ( .C1(n15033), .C2(n15393), .A(n15147), .B(n14989), .ZN(
        n14990) );
  OAI211_X1 U16343 ( .C1(n15590), .C2(n15066), .A(n14991), .B(n14990), .ZN(
        P2_U3191) );
  NOR3_X1 U16344 ( .A1(n14992), .A2(n15183), .A3(n15067), .ZN(n14997) );
  AOI21_X1 U16345 ( .B1(n14993), .B2(n15040), .A(n15077), .ZN(n14996) );
  INV_X1 U16346 ( .A(n14994), .ZN(n14995) );
  OAI21_X1 U16347 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(n15002) );
  INV_X1 U16348 ( .A(n14998), .ZN(n15358) );
  AOI22_X1 U16349 ( .A1(n15215), .A2(n15073), .B1(n15225), .B2(n15210), .ZN(
        n15364) );
  OAI22_X1 U16350 ( .A1(n15364), .A2(n15076), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14999), .ZN(n15000) );
  AOI21_X1 U16351 ( .B1(n15358), .B2(n15074), .A(n15000), .ZN(n15001) );
  OAI211_X1 U16352 ( .C1(n15360), .C2(n15066), .A(n15002), .B(n15001), .ZN(
        P2_U3195) );
  NAND3_X1 U16353 ( .A1(n15003), .A2(n15050), .A3(n15191), .ZN(n15008) );
  OAI21_X1 U16354 ( .B1(n15004), .B2(n15005), .A(n15070), .ZN(n15007) );
  INV_X1 U16355 ( .A(n15006), .ZN(n15071) );
  AOI21_X1 U16356 ( .B1(n15008), .B2(n15007), .A(n15071), .ZN(n15009) );
  INV_X1 U16357 ( .A(n15009), .ZN(n15014) );
  OAI22_X1 U16358 ( .A1(n15192), .A2(n15162), .B1(n15010), .B2(n15043), .ZN(
        n15291) );
  OAI22_X1 U16359 ( .A1(n15297), .A2(n15052), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15011), .ZN(n15012) );
  AOI21_X1 U16360 ( .B1(n15291), .B2(n15033), .A(n15012), .ZN(n15013) );
  OAI211_X1 U16361 ( .C1(n15568), .C2(n15066), .A(n15014), .B(n15013), .ZN(
        P2_U3197) );
  OAI21_X1 U16362 ( .B1(n15017), .B2(n15016), .A(n15015), .ZN(n15018) );
  NAND2_X1 U16363 ( .A1(n15018), .A2(n15070), .ZN(n15026) );
  AOI21_X1 U16364 ( .B1(n15033), .B2(n15020), .A(n15019), .ZN(n15025) );
  NAND2_X1 U16365 ( .A1(n15074), .A2(n15021), .ZN(n15024) );
  NAND2_X1 U16366 ( .A1(n15080), .A2(n15022), .ZN(n15023) );
  NAND4_X1 U16367 ( .A1(n15026), .A2(n15025), .A3(n15024), .A4(n15023), .ZN(
        P2_U3199) );
  AOI211_X1 U16368 ( .C1(n7494), .C2(n15027), .A(n15077), .B(n15004), .ZN(
        n15028) );
  INV_X1 U16369 ( .A(n15028), .ZN(n15035) );
  NAND2_X1 U16370 ( .A1(n15084), .A2(n15073), .ZN(n15030) );
  NAND2_X1 U16371 ( .A1(n15216), .A2(n15225), .ZN(n15029) );
  NAND2_X1 U16372 ( .A1(n15030), .A2(n15029), .ZN(n15310) );
  OAI22_X1 U16373 ( .A1(n15314), .A2(n15052), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15031), .ZN(n15032) );
  AOI21_X1 U16374 ( .B1(n15310), .B2(n15033), .A(n15032), .ZN(n15034) );
  OAI211_X1 U16375 ( .C1(n15572), .C2(n15066), .A(n15035), .B(n15034), .ZN(
        P2_U3201) );
  INV_X1 U16376 ( .A(n15036), .ZN(n15038) );
  AOI21_X1 U16377 ( .B1(n15038), .B2(n15037), .A(n15077), .ZN(n15042) );
  NOR3_X1 U16378 ( .A1(n15039), .A2(n15181), .A3(n15067), .ZN(n15041) );
  OAI21_X1 U16379 ( .B1(n15042), .B2(n15041), .A(n15040), .ZN(n15048) );
  OAI22_X1 U16380 ( .A1(n15184), .A2(n15162), .B1(n15181), .B2(n15043), .ZN(
        n15369) );
  INV_X1 U16381 ( .A(n15369), .ZN(n15045) );
  OAI22_X1 U16382 ( .A1(n15045), .A2(n15076), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15044), .ZN(n15046) );
  AOI21_X1 U16383 ( .B1(n15373), .B2(n15074), .A(n15046), .ZN(n15047) );
  OAI211_X1 U16384 ( .C1(n15585), .C2(n15066), .A(n15048), .B(n15047), .ZN(
        P2_U3205) );
  INV_X1 U16385 ( .A(n15049), .ZN(n15058) );
  AOI22_X1 U16386 ( .A1(n15051), .A2(n15070), .B1(n15050), .B2(n15215), .ZN(
        n15057) );
  NOR2_X1 U16387 ( .A1(n15052), .A2(n15343), .ZN(n15055) );
  AOI22_X1 U16388 ( .A1(n15216), .A2(n15073), .B1(n15225), .B2(n15212), .ZN(
        n15349) );
  OAI22_X1 U16389 ( .A1(n15349), .A2(n15076), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15053), .ZN(n15054) );
  AOI211_X1 U16390 ( .C1(n15342), .C2(n15080), .A(n15055), .B(n15054), .ZN(
        n15056) );
  OAI21_X1 U16391 ( .B1(n15058), .B2(n15057), .A(n15056), .ZN(P2_U3207) );
  AOI21_X1 U16392 ( .B1(n15060), .B2(n15059), .A(n15077), .ZN(n15062) );
  NAND2_X1 U16393 ( .A1(n15062), .A2(n15061), .ZN(n15065) );
  AOI22_X1 U16394 ( .A1(n15208), .A2(n15073), .B1(n15225), .B2(n15177), .ZN(
        n15405) );
  OAI22_X1 U16395 ( .A1(n15405), .A2(n15076), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15127), .ZN(n15063) );
  AOI21_X1 U16396 ( .B1(n15410), .B2(n15074), .A(n15063), .ZN(n15064) );
  OAI211_X1 U16397 ( .C1(n15595), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        P2_U3210) );
  INV_X1 U16398 ( .A(n15084), .ZN(n15218) );
  NOR3_X1 U16399 ( .A1(n15068), .A2(n15218), .A3(n15067), .ZN(n15069) );
  AOI21_X1 U16400 ( .B1(n15071), .B2(n15070), .A(n15069), .ZN(n15082) );
  AND2_X1 U16401 ( .A1(n15084), .A2(n15225), .ZN(n15072) );
  AOI21_X1 U16402 ( .B1(n15193), .B2(n15073), .A(n15072), .ZN(n15277) );
  AOI22_X1 U16403 ( .A1(n15281), .A2(n15074), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n15075) );
  OAI21_X1 U16404 ( .B1(n15277), .B2(n15076), .A(n15075), .ZN(n15079) );
  MUX2_X1 U16405 ( .A(n15163), .B(P2_DATAO_REG_31__SCAN_IN), .S(n15098), .Z(
        P2_U3562) );
  MUX2_X1 U16406 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n15228), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U16407 ( .A(n15083), .B(P2_DATAO_REG_29__SCAN_IN), .S(n15098), .Z(
        P2_U3560) );
  MUX2_X1 U16408 ( .A(n15226), .B(P2_DATAO_REG_28__SCAN_IN), .S(n15098), .Z(
        P2_U3559) );
  MUX2_X1 U16409 ( .A(n15193), .B(P2_DATAO_REG_27__SCAN_IN), .S(n15098), .Z(
        P2_U3558) );
  MUX2_X1 U16410 ( .A(n15084), .B(P2_DATAO_REG_25__SCAN_IN), .S(n15098), .Z(
        P2_U3556) );
  MUX2_X1 U16411 ( .A(n15216), .B(P2_DATAO_REG_23__SCAN_IN), .S(n15098), .Z(
        P2_U3554) );
  MUX2_X1 U16412 ( .A(n15212), .B(P2_DATAO_REG_21__SCAN_IN), .S(n15098), .Z(
        P2_U3552) );
  MUX2_X1 U16413 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n15210), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U16414 ( .A(n15208), .B(P2_DATAO_REG_19__SCAN_IN), .S(n15098), .Z(
        P2_U3550) );
  MUX2_X1 U16415 ( .A(n15205), .B(P2_DATAO_REG_18__SCAN_IN), .S(n15098), .Z(
        P2_U3549) );
  MUX2_X1 U16416 ( .A(n15177), .B(P2_DATAO_REG_17__SCAN_IN), .S(n15098), .Z(
        P2_U3548) );
  MUX2_X1 U16417 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n15175), .S(P2_U3947), .Z(
        P2_U3547) );
  MUX2_X1 U16418 ( .A(n15196), .B(P2_DATAO_REG_15__SCAN_IN), .S(n15098), .Z(
        P2_U3546) );
  MUX2_X1 U16419 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n15085), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U16420 ( .A(n15086), .B(P2_DATAO_REG_13__SCAN_IN), .S(n15098), .Z(
        P2_U3544) );
  MUX2_X1 U16421 ( .A(n15087), .B(P2_DATAO_REG_12__SCAN_IN), .S(n15098), .Z(
        P2_U3543) );
  MUX2_X1 U16422 ( .A(n15088), .B(P2_DATAO_REG_11__SCAN_IN), .S(n15098), .Z(
        P2_U3542) );
  MUX2_X1 U16423 ( .A(n15089), .B(P2_DATAO_REG_10__SCAN_IN), .S(n15098), .Z(
        P2_U3541) );
  MUX2_X1 U16424 ( .A(n15090), .B(P2_DATAO_REG_9__SCAN_IN), .S(n15098), .Z(
        P2_U3540) );
  MUX2_X1 U16425 ( .A(n15091), .B(P2_DATAO_REG_8__SCAN_IN), .S(n15098), .Z(
        P2_U3539) );
  MUX2_X1 U16426 ( .A(n15092), .B(P2_DATAO_REG_7__SCAN_IN), .S(n15098), .Z(
        P2_U3538) );
  MUX2_X1 U16427 ( .A(n15093), .B(P2_DATAO_REG_6__SCAN_IN), .S(n15098), .Z(
        P2_U3537) );
  MUX2_X1 U16428 ( .A(n15094), .B(P2_DATAO_REG_5__SCAN_IN), .S(n15098), .Z(
        P2_U3536) );
  MUX2_X1 U16429 ( .A(n15095), .B(P2_DATAO_REG_4__SCAN_IN), .S(n15098), .Z(
        P2_U3535) );
  MUX2_X1 U16430 ( .A(n15096), .B(P2_DATAO_REG_3__SCAN_IN), .S(n15098), .Z(
        P2_U3534) );
  MUX2_X1 U16431 ( .A(n15097), .B(P2_DATAO_REG_2__SCAN_IN), .S(n15098), .Z(
        P2_U3533) );
  MUX2_X1 U16432 ( .A(n9875), .B(P2_DATAO_REG_1__SCAN_IN), .S(n15098), .Z(
        P2_U3532) );
  MUX2_X1 U16433 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n15099), .S(P2_U3947), .Z(
        P2_U3531) );
  INV_X1 U16434 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n16305) );
  OR2_X1 U16435 ( .A1(n16305), .A2(n16278), .ZN(n15112) );
  AOI22_X1 U16436 ( .A1(n16270), .A2(n15100), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(P2_U3088), .ZN(n15111) );
  INV_X1 U16437 ( .A(n15101), .ZN(n15105) );
  OAI21_X1 U16438 ( .B1(n11525), .B2(n15103), .A(n15102), .ZN(n15104) );
  NAND3_X1 U16439 ( .A1(n16257), .A2(n15105), .A3(n15104), .ZN(n15110) );
  OAI211_X1 U16440 ( .C1(n15108), .C2(n15107), .A(n16230), .B(n15106), .ZN(
        n15109) );
  NAND4_X1 U16441 ( .A1(n15112), .A2(n15111), .A3(n15110), .A4(n15109), .ZN(
        P2_U3215) );
  INV_X1 U16442 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16443 ( .A1(n15122), .A2(n15121), .ZN(n15113) );
  AOI21_X1 U16444 ( .B1(n15121), .B2(n15122), .A(n15113), .ZN(n16259) );
  NOR2_X1 U16445 ( .A1(n15120), .A2(n15114), .ZN(n15115) );
  AOI21_X1 U16446 ( .B1(n15114), .B2(n15120), .A(n15115), .ZN(n16245) );
  NAND2_X1 U16447 ( .A1(n15117), .A2(n15116), .ZN(n15119) );
  NAND2_X1 U16448 ( .A1(n15119), .A2(n15118), .ZN(n16246) );
  NAND2_X1 U16449 ( .A1(n16245), .A2(n16246), .ZN(n16244) );
  OAI21_X1 U16450 ( .B1(n15120), .B2(n15114), .A(n16244), .ZN(n16258) );
  NAND2_X1 U16451 ( .A1(n16259), .A2(n16258), .ZN(n16256) );
  OAI21_X1 U16452 ( .B1(n15122), .B2(n15121), .A(n16256), .ZN(n15124) );
  INV_X1 U16453 ( .A(n15124), .ZN(n15125) );
  OR2_X1 U16454 ( .A1(n15124), .A2(n15123), .ZN(n15148) );
  OAI21_X1 U16455 ( .B1(n15125), .B2(n15135), .A(n15148), .ZN(n15126) );
  NOR2_X1 U16456 ( .A1(n15126), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n15150) );
  AOI21_X1 U16457 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n15126), .A(n15150), 
        .ZN(n15140) );
  NOR2_X1 U16458 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15127), .ZN(n15130) );
  NOR2_X1 U16459 ( .A1(n15128), .A2(n15135), .ZN(n15129) );
  AOI211_X1 U16460 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n16224), .A(n15130), 
        .B(n15129), .ZN(n15139) );
  NOR2_X1 U16461 ( .A1(n15132), .A2(n15131), .ZN(n15134) );
  XNOR2_X1 U16462 ( .A(n16243), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n16239) );
  NOR2_X1 U16463 ( .A1(n16240), .A2(n16239), .ZN(n16238) );
  XNOR2_X1 U16464 ( .A(n16255), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n16251) );
  AOI21_X1 U16465 ( .B1(n15136), .B2(n15135), .A(n15141), .ZN(n15137) );
  NAND2_X1 U16466 ( .A1(n15137), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n15143) );
  OAI211_X1 U16467 ( .C1(n15137), .C2(P2_REG1_REG_18__SCAN_IN), .A(n15143), 
        .B(n16230), .ZN(n15138) );
  OAI211_X1 U16468 ( .C1(n15140), .C2(n16272), .A(n15139), .B(n15138), .ZN(
        P2_U3232) );
  INV_X1 U16469 ( .A(n15141), .ZN(n15142) );
  NAND2_X1 U16470 ( .A1(n15143), .A2(n15142), .ZN(n15145) );
  INV_X1 U16471 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15523) );
  XNOR2_X1 U16472 ( .A(n10515), .B(n15523), .ZN(n15144) );
  XNOR2_X1 U16473 ( .A(n15145), .B(n15144), .ZN(n15156) );
  AND2_X1 U16474 ( .A1(n16270), .A2(n10515), .ZN(n15146) );
  AOI211_X1 U16475 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n16224), .A(n15147), 
        .B(n15146), .ZN(n15155) );
  INV_X1 U16476 ( .A(n15148), .ZN(n15149) );
  NOR2_X1 U16477 ( .A1(n15150), .A2(n15149), .ZN(n15152) );
  MUX2_X1 U16478 ( .A(n15388), .B(P2_REG2_REG_19__SCAN_IN), .S(n10515), .Z(
        n15151) );
  XNOR2_X1 U16479 ( .A(n15152), .B(n15151), .ZN(n15153) );
  NAND2_X1 U16480 ( .A1(n15153), .A2(n16257), .ZN(n15154) );
  OAI211_X1 U16481 ( .C1(n15156), .C2(n16264), .A(n15155), .B(n15154), .ZN(
        P2_U3233) );
  AND2_X1 U16482 ( .A1(n15595), .A2(n15426), .ZN(n15407) );
  NAND2_X1 U16483 ( .A1(n15284), .A2(n15295), .ZN(n15280) );
  XNOR2_X1 U16484 ( .A(n15166), .B(n15552), .ZN(n15157) );
  NOR2_X1 U16485 ( .A1(n15429), .A2(n15158), .ZN(n15164) );
  INV_X1 U16486 ( .A(P2_B_REG_SCAN_IN), .ZN(n15159) );
  NOR2_X1 U16487 ( .A1(n15160), .A2(n15159), .ZN(n15161) );
  NOR2_X1 U16488 ( .A1(n15162), .A2(n15161), .ZN(n15227) );
  NAND2_X1 U16489 ( .A1(n15163), .A2(n15227), .ZN(n15464) );
  NOR2_X1 U16490 ( .A1(n15454), .A2(n15464), .ZN(n15170) );
  AOI211_X1 U16491 ( .C1(n15552), .C2(n15316), .A(n15164), .B(n15170), .ZN(
        n15165) );
  OAI21_X1 U16492 ( .B1(n15463), .B2(n15318), .A(n15165), .ZN(P2_U3234) );
  AOI21_X1 U16493 ( .B1(n15467), .B2(n15231), .A(n7418), .ZN(n15168) );
  INV_X1 U16494 ( .A(n15166), .ZN(n15167) );
  NAND2_X1 U16495 ( .A1(n15168), .A2(n15167), .ZN(n15465) );
  NOR2_X1 U16496 ( .A1(n15560), .A2(n15456), .ZN(n15169) );
  AOI211_X1 U16497 ( .C1(n15454), .C2(P2_REG2_REG_30__SCAN_IN), .A(n15170), 
        .B(n15169), .ZN(n15171) );
  OAI21_X1 U16498 ( .B1(n15318), .B2(n15465), .A(n15171), .ZN(P2_U3235) );
  INV_X1 U16499 ( .A(n15403), .ZN(n15402) );
  NAND2_X1 U16500 ( .A1(n15197), .A2(n15172), .ZN(n15173) );
  INV_X1 U16501 ( .A(n15437), .ZN(n15439) );
  NAND2_X1 U16502 ( .A1(n15539), .A2(n15175), .ZN(n15176) );
  INV_X1 U16503 ( .A(n15418), .ZN(n15416) );
  OR2_X1 U16504 ( .A1(n15598), .A2(n15177), .ZN(n15178) );
  NAND2_X1 U16505 ( .A1(n15179), .A2(n15178), .ZN(n15401) );
  NAND2_X1 U16506 ( .A1(n15402), .A2(n15401), .ZN(n15400) );
  NAND2_X1 U16507 ( .A1(n15595), .A2(n15203), .ZN(n15180) );
  INV_X1 U16508 ( .A(n15391), .ZN(n15382) );
  NAND2_X1 U16509 ( .A1(n15590), .A2(n15181), .ZN(n15182) );
  NAND2_X1 U16510 ( .A1(n15360), .A2(n15184), .ZN(n15185) );
  NAND2_X1 U16511 ( .A1(n15342), .A2(n15215), .ZN(n15186) );
  NAND2_X1 U16512 ( .A1(n15187), .A2(n15186), .ZN(n15335) );
  NAND2_X1 U16513 ( .A1(n15335), .A2(n15333), .ZN(n15190) );
  OR2_X1 U16514 ( .A1(n15576), .A2(n15188), .ZN(n15189) );
  NAND2_X1 U16515 ( .A1(n15242), .A2(n15241), .ZN(n15240) );
  NAND2_X1 U16516 ( .A1(n15197), .A2(n15196), .ZN(n15198) );
  NAND2_X1 U16517 ( .A1(n15539), .A2(n15200), .ZN(n15201) );
  NAND2_X1 U16518 ( .A1(n15409), .A2(n15203), .ZN(n15204) );
  NAND2_X1 U16519 ( .A1(n15595), .A2(n15205), .ZN(n15206) );
  AND2_X1 U16520 ( .A1(n15590), .A2(n15208), .ZN(n15207) );
  OR2_X1 U16521 ( .A1(n15590), .A2(n15208), .ZN(n15209) );
  NOR2_X1 U16522 ( .A1(n15360), .A2(n15212), .ZN(n15211) );
  NAND2_X1 U16523 ( .A1(n15360), .A2(n15212), .ZN(n15213) );
  INV_X1 U16524 ( .A(n15241), .ZN(n15251) );
  NAND2_X1 U16525 ( .A1(n15252), .A2(n15251), .ZN(n15250) );
  NAND2_X1 U16526 ( .A1(n15250), .A2(n15221), .ZN(n15224) );
  NAND2_X1 U16527 ( .A1(n15226), .A2(n15225), .ZN(n15230) );
  OAI211_X1 U16528 ( .C1(n15470), .C2(n15246), .A(n15232), .B(n15231), .ZN(
        n15469) );
  INV_X1 U16529 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U16530 ( .A1(n15234), .A2(n15427), .B1(n15233), .B2(n15429), .ZN(
        n15235) );
  AOI21_X1 U16531 ( .B1(n15236), .B2(n15316), .A(n15235), .ZN(n15237) );
  OAI21_X1 U16532 ( .B1(n15469), .B2(n15318), .A(n15237), .ZN(n15238) );
  AOI21_X1 U16533 ( .B1(n7448), .B2(n15429), .A(n15238), .ZN(n15239) );
  OAI21_X1 U16534 ( .B1(n8839), .B2(n15435), .A(n15239), .ZN(P2_U3236) );
  OAI21_X1 U16535 ( .B1(n15242), .B2(n15241), .A(n15240), .ZN(n15243) );
  INV_X1 U16536 ( .A(n15243), .ZN(n15475) );
  NAND2_X1 U16537 ( .A1(n15474), .A2(n15263), .ZN(n15244) );
  NAND2_X1 U16538 ( .A1(n15244), .A2(n15232), .ZN(n15245) );
  NOR2_X1 U16539 ( .A1(n15246), .A2(n15245), .ZN(n15473) );
  INV_X1 U16540 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n15247) );
  OAI22_X1 U16541 ( .A1(n15248), .A2(n15456), .B1(n15429), .B2(n15247), .ZN(
        n15249) );
  AOI21_X1 U16542 ( .B1(n15473), .B2(n15461), .A(n15249), .ZN(n15258) );
  OAI211_X1 U16543 ( .C1(n15252), .C2(n15251), .A(n15250), .B(n15446), .ZN(
        n15254) );
  NOR2_X1 U16544 ( .A1(n15255), .A2(n15427), .ZN(n15256) );
  OAI21_X1 U16545 ( .B1(n15472), .B2(n15256), .A(n15429), .ZN(n15257) );
  OAI211_X1 U16546 ( .C1(n15475), .C2(n15435), .A(n15258), .B(n15257), .ZN(
        P2_U3237) );
  AOI21_X1 U16547 ( .B1(n15261), .B2(n15260), .A(n15259), .ZN(n15262) );
  INV_X1 U16548 ( .A(n15262), .ZN(n15480) );
  AOI211_X1 U16549 ( .C1(n15478), .C2(n15280), .A(n7418), .B(n7664), .ZN(
        n15477) );
  INV_X1 U16550 ( .A(n15478), .ZN(n15266) );
  AOI22_X1 U16551 ( .A1(n15264), .A2(n15452), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15454), .ZN(n15265) );
  OAI21_X1 U16552 ( .B1(n15266), .B2(n15456), .A(n15265), .ZN(n15267) );
  AOI21_X1 U16553 ( .B1(n15477), .B2(n15461), .A(n15267), .ZN(n15273) );
  XNOR2_X1 U16554 ( .A(n15269), .B(n15268), .ZN(n15271) );
  OAI21_X1 U16555 ( .B1(n15271), .B2(n11226), .A(n15270), .ZN(n15476) );
  NAND2_X1 U16556 ( .A1(n15476), .A2(n15429), .ZN(n15272) );
  OAI211_X1 U16557 ( .C1(n15480), .C2(n15435), .A(n15273), .B(n15272), .ZN(
        P2_U3238) );
  XNOR2_X1 U16558 ( .A(n15274), .B(n15276), .ZN(n15485) );
  XOR2_X1 U16559 ( .A(n15276), .B(n15275), .Z(n15278) );
  OAI21_X1 U16560 ( .B1(n15278), .B2(n11226), .A(n15277), .ZN(n15481) );
  OR2_X1 U16561 ( .A1(n15284), .A2(n15295), .ZN(n15279) );
  AND3_X1 U16562 ( .A1(n15280), .A2(n15279), .A3(n15232), .ZN(n15482) );
  NAND2_X1 U16563 ( .A1(n15482), .A2(n15461), .ZN(n15283) );
  AOI22_X1 U16564 ( .A1(n15281), .A2(n15452), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15454), .ZN(n15282) );
  OAI211_X1 U16565 ( .C1(n15284), .C2(n15456), .A(n15283), .B(n15282), .ZN(
        n15285) );
  AOI21_X1 U16566 ( .B1(n15481), .B2(n15429), .A(n15285), .ZN(n15286) );
  OAI21_X1 U16567 ( .B1(n15485), .B2(n15435), .A(n15286), .ZN(P2_U3239) );
  INV_X1 U16568 ( .A(n15289), .ZN(n15287) );
  XNOR2_X1 U16569 ( .A(n15288), .B(n15287), .ZN(n15486) );
  INV_X1 U16570 ( .A(n15486), .ZN(n15304) );
  XNOR2_X1 U16571 ( .A(n15290), .B(n15289), .ZN(n15292) );
  AOI21_X1 U16572 ( .B1(n15292), .B2(n15446), .A(n15291), .ZN(n15489) );
  INV_X1 U16573 ( .A(n15489), .ZN(n15302) );
  NAND2_X1 U16574 ( .A1(n15312), .A2(n15299), .ZN(n15293) );
  NAND2_X1 U16575 ( .A1(n15293), .A2(n15232), .ZN(n15294) );
  OR2_X1 U16576 ( .A1(n15295), .A2(n15294), .ZN(n15487) );
  INV_X1 U16577 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n15296) );
  OAI22_X1 U16578 ( .A1(n15297), .A2(n15427), .B1(n15296), .B2(n15429), .ZN(
        n15298) );
  AOI21_X1 U16579 ( .B1(n15299), .B2(n15316), .A(n15298), .ZN(n15300) );
  OAI21_X1 U16580 ( .B1(n15487), .B2(n15318), .A(n15300), .ZN(n15301) );
  AOI21_X1 U16581 ( .B1(n15302), .B2(n15429), .A(n15301), .ZN(n15303) );
  OAI21_X1 U16582 ( .B1(n15304), .B2(n15435), .A(n15303), .ZN(P2_U3240) );
  XNOR2_X1 U16583 ( .A(n15305), .B(n15306), .ZN(n15494) );
  NAND2_X1 U16584 ( .A1(n15307), .A2(n15306), .ZN(n15308) );
  NAND2_X1 U16585 ( .A1(n15309), .A2(n15308), .ZN(n15311) );
  AOI21_X1 U16586 ( .B1(n15311), .B2(n15446), .A(n15310), .ZN(n15493) );
  INV_X1 U16587 ( .A(n15493), .ZN(n15320) );
  OAI211_X1 U16588 ( .C1(n7592), .C2(n15572), .A(n15232), .B(n15312), .ZN(
        n15492) );
  INV_X1 U16589 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n15313) );
  OAI22_X1 U16590 ( .A1(n15314), .A2(n15427), .B1(n15313), .B2(n15429), .ZN(
        n15315) );
  AOI21_X1 U16591 ( .B1(n15496), .B2(n15316), .A(n15315), .ZN(n15317) );
  OAI21_X1 U16592 ( .B1(n15492), .B2(n15318), .A(n15317), .ZN(n15319) );
  AOI21_X1 U16593 ( .B1(n15320), .B2(n15429), .A(n15319), .ZN(n15321) );
  OAI21_X1 U16594 ( .B1(n15435), .B2(n15494), .A(n15321), .ZN(P2_U3241) );
  NAND2_X1 U16595 ( .A1(n15322), .A2(n15333), .ZN(n15323) );
  NAND3_X1 U16596 ( .A1(n15324), .A2(n15446), .A3(n15323), .ZN(n15326) );
  NAND2_X1 U16597 ( .A1(n15340), .A2(n15503), .ZN(n15327) );
  NAND2_X1 U16598 ( .A1(n15327), .A2(n15232), .ZN(n15328) );
  OR2_X1 U16599 ( .A1(n7592), .A2(n15328), .ZN(n15499) );
  INV_X1 U16600 ( .A(n15499), .ZN(n15332) );
  AOI22_X1 U16601 ( .A1(n15329), .A2(n15452), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n15454), .ZN(n15330) );
  OAI21_X1 U16602 ( .B1(n15576), .B2(n15456), .A(n15330), .ZN(n15331) );
  AOI21_X1 U16603 ( .B1(n15332), .B2(n15461), .A(n15331), .ZN(n15338) );
  INV_X1 U16604 ( .A(n15333), .ZN(n15334) );
  XNOR2_X1 U16605 ( .A(n15335), .B(n15334), .ZN(n15498) );
  NAND2_X1 U16606 ( .A1(n15498), .A2(n15336), .ZN(n15337) );
  OAI211_X1 U16607 ( .C1(n15501), .C2(n15454), .A(n15338), .B(n15337), .ZN(
        P2_U3242) );
  XOR2_X1 U16608 ( .A(n15339), .B(n15348), .Z(n15507) );
  INV_X1 U16609 ( .A(n15507), .ZN(n15353) );
  INV_X1 U16610 ( .A(n15340), .ZN(n15341) );
  AOI211_X1 U16611 ( .C1(n15342), .C2(n15355), .A(n7418), .B(n15341), .ZN(
        n15505) );
  INV_X1 U16612 ( .A(n15343), .ZN(n15344) );
  AOI22_X1 U16613 ( .A1(n15344), .A2(n15452), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n15454), .ZN(n15345) );
  OAI21_X1 U16614 ( .B1(n15580), .B2(n15456), .A(n15345), .ZN(n15346) );
  AOI21_X1 U16615 ( .B1(n15505), .B2(n15461), .A(n15346), .ZN(n15352) );
  XNOR2_X1 U16616 ( .A(n15347), .B(n15348), .ZN(n15350) );
  OAI21_X1 U16617 ( .B1(n15350), .B2(n11226), .A(n15349), .ZN(n15506) );
  NAND2_X1 U16618 ( .A1(n15506), .A2(n15429), .ZN(n15351) );
  OAI211_X1 U16619 ( .C1(n15353), .C2(n15435), .A(n15352), .B(n15351), .ZN(
        P2_U3243) );
  XNOR2_X1 U16620 ( .A(n15362), .B(n15354), .ZN(n15513) );
  INV_X1 U16621 ( .A(n15372), .ZN(n15357) );
  INV_X1 U16622 ( .A(n15355), .ZN(n15356) );
  AOI211_X1 U16623 ( .C1(n8227), .C2(n15357), .A(n7418), .B(n15356), .ZN(
        n15510) );
  AOI22_X1 U16624 ( .A1(n15358), .A2(n15452), .B1(n15454), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n15359) );
  OAI21_X1 U16625 ( .B1(n15360), .B2(n15456), .A(n15359), .ZN(n15361) );
  AOI21_X1 U16626 ( .B1(n15510), .B2(n15461), .A(n15361), .ZN(n15367) );
  XNOR2_X1 U16627 ( .A(n15363), .B(n15362), .ZN(n15365) );
  OAI21_X1 U16628 ( .B1(n15365), .B2(n11226), .A(n15364), .ZN(n15511) );
  NAND2_X1 U16629 ( .A1(n15511), .A2(n15429), .ZN(n15366) );
  OAI211_X1 U16630 ( .C1(n15513), .C2(n15435), .A(n15367), .B(n15366), .ZN(
        P2_U3244) );
  XNOR2_X1 U16631 ( .A(n15368), .B(n15375), .ZN(n15370) );
  AOI21_X1 U16632 ( .B1(n15370), .B2(n15446), .A(n15369), .ZN(n15515) );
  OAI21_X1 U16633 ( .B1(n15585), .B2(n15384), .A(n15232), .ZN(n15371) );
  OR2_X1 U16634 ( .A1(n15372), .A2(n15371), .ZN(n15514) );
  INV_X1 U16635 ( .A(n15514), .ZN(n15379) );
  AOI22_X1 U16636 ( .A1(n15454), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n15373), 
        .B2(n15452), .ZN(n15374) );
  OAI21_X1 U16637 ( .B1(n15585), .B2(n15456), .A(n15374), .ZN(n15378) );
  XNOR2_X1 U16638 ( .A(n15376), .B(n15375), .ZN(n15516) );
  NOR2_X1 U16639 ( .A1(n15516), .A2(n15435), .ZN(n15377) );
  AOI211_X1 U16640 ( .C1(n15379), .C2(n15461), .A(n15378), .B(n15377), .ZN(
        n15380) );
  OAI21_X1 U16641 ( .B1(n15454), .B2(n15515), .A(n15380), .ZN(P2_U3245) );
  OAI21_X1 U16642 ( .B1(n15383), .B2(n15382), .A(n15381), .ZN(n15522) );
  INV_X1 U16643 ( .A(n15522), .ZN(n15399) );
  INV_X1 U16644 ( .A(n15407), .ZN(n15385) );
  AOI211_X1 U16645 ( .C1(n15386), .C2(n15385), .A(n7418), .B(n15384), .ZN(
        n15521) );
  NOR2_X1 U16646 ( .A1(n15590), .A2(n15456), .ZN(n15390) );
  OAI22_X1 U16647 ( .A1(n15429), .A2(n15388), .B1(n15387), .B2(n15427), .ZN(
        n15389) );
  AOI211_X1 U16648 ( .C1(n15521), .C2(n15461), .A(n15390), .B(n15389), .ZN(
        n15398) );
  XNOR2_X1 U16649 ( .A(n15392), .B(n15391), .ZN(n15396) );
  AOI21_X1 U16650 ( .B1(n15522), .B2(n15394), .A(n15393), .ZN(n15395) );
  OAI21_X1 U16651 ( .B1(n11226), .B2(n15396), .A(n15395), .ZN(n15520) );
  NAND2_X1 U16652 ( .A1(n15520), .A2(n15429), .ZN(n15397) );
  OAI211_X1 U16653 ( .C1(n15399), .C2(n15458), .A(n15398), .B(n15397), .ZN(
        P2_U3246) );
  OAI21_X1 U16654 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15527) );
  INV_X1 U16655 ( .A(n15527), .ZN(n15415) );
  XNOR2_X1 U16656 ( .A(n15404), .B(n15403), .ZN(n15406) );
  OAI21_X1 U16657 ( .B1(n15406), .B2(n11226), .A(n15405), .ZN(n15525) );
  NAND2_X1 U16658 ( .A1(n15525), .A2(n15429), .ZN(n15414) );
  INV_X1 U16659 ( .A(n15426), .ZN(n15408) );
  AOI211_X1 U16660 ( .C1(n15409), .C2(n15408), .A(n7418), .B(n15407), .ZN(
        n15526) );
  AOI22_X1 U16661 ( .A1(n15454), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n15410), 
        .B2(n15452), .ZN(n15411) );
  OAI21_X1 U16662 ( .B1(n15595), .B2(n15456), .A(n15411), .ZN(n15412) );
  AOI21_X1 U16663 ( .B1(n15526), .B2(n15461), .A(n15412), .ZN(n15413) );
  OAI211_X1 U16664 ( .C1(n15415), .C2(n15435), .A(n15414), .B(n15413), .ZN(
        P2_U3247) );
  XNOR2_X1 U16665 ( .A(n15417), .B(n15416), .ZN(n15531) );
  INV_X1 U16666 ( .A(n15531), .ZN(n15436) );
  NAND2_X1 U16667 ( .A1(n15419), .A2(n15418), .ZN(n15420) );
  NAND3_X1 U16668 ( .A1(n15421), .A2(n15446), .A3(n15420), .ZN(n15423) );
  NAND2_X1 U16669 ( .A1(n15423), .A2(n15422), .ZN(n15534) );
  NAND2_X1 U16670 ( .A1(n15534), .A2(n15429), .ZN(n15434) );
  NAND2_X1 U16671 ( .A1(n15598), .A2(n15449), .ZN(n15424) );
  NAND2_X1 U16672 ( .A1(n15424), .A2(n15232), .ZN(n15425) );
  NOR2_X1 U16673 ( .A1(n15426), .A2(n15425), .ZN(n15532) );
  OAI22_X1 U16674 ( .A1(n15429), .A2(n15121), .B1(n15428), .B2(n15427), .ZN(
        n15432) );
  NOR2_X1 U16675 ( .A1(n15430), .A2(n15456), .ZN(n15431) );
  AOI211_X1 U16676 ( .C1(n15532), .C2(n15461), .A(n15432), .B(n15431), .ZN(
        n15433) );
  OAI211_X1 U16677 ( .C1(n15436), .C2(n15435), .A(n15434), .B(n15433), .ZN(
        P2_U3248) );
  XNOR2_X1 U16678 ( .A(n15438), .B(n15437), .ZN(n15447) );
  NAND2_X1 U16679 ( .A1(n15440), .A2(n15439), .ZN(n15441) );
  NAND2_X1 U16680 ( .A1(n15442), .A2(n15441), .ZN(n15542) );
  NOR2_X1 U16681 ( .A1(n15542), .A2(n15443), .ZN(n15444) );
  AOI211_X1 U16682 ( .C1(n15447), .C2(n15446), .A(n15445), .B(n15444), .ZN(
        n15541) );
  INV_X1 U16683 ( .A(n15448), .ZN(n15451) );
  INV_X1 U16684 ( .A(n15449), .ZN(n15450) );
  AOI211_X1 U16685 ( .C1(n15539), .C2(n15451), .A(n7418), .B(n15450), .ZN(
        n15538) );
  AOI22_X1 U16686 ( .A1(n15454), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n15453), 
        .B2(n15452), .ZN(n15455) );
  OAI21_X1 U16687 ( .B1(n15457), .B2(n15456), .A(n15455), .ZN(n15460) );
  NOR2_X1 U16688 ( .A1(n15542), .A2(n15458), .ZN(n15459) );
  AOI211_X1 U16689 ( .C1(n15538), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15462) );
  OAI21_X1 U16690 ( .B1(n15541), .B2(n15454), .A(n15462), .ZN(P2_U3249) );
  NAND2_X1 U16691 ( .A1(n15465), .A2(n15464), .ZN(n15557) );
  MUX2_X1 U16692 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n15557), .S(n16526), .Z(
        n15466) );
  AOI21_X1 U16693 ( .B1(n15536), .B2(n15467), .A(n15466), .ZN(n15468) );
  INV_X1 U16694 ( .A(n15468), .ZN(P2_U3529) );
  OAI21_X1 U16695 ( .B1(n15550), .B2(n15480), .A(n15479), .ZN(n15563) );
  MUX2_X1 U16696 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n15563), .S(n16526), .Z(
        P2_U3526) );
  AOI211_X1 U16697 ( .C1(n15546), .C2(n15483), .A(n15482), .B(n15481), .ZN(
        n15484) );
  OAI21_X1 U16698 ( .B1(n15550), .B2(n15485), .A(n15484), .ZN(n15564) );
  MUX2_X1 U16699 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n15564), .S(n16526), .Z(
        P2_U3525) );
  NAND2_X1 U16700 ( .A1(n15486), .A2(n16523), .ZN(n15488) );
  AND3_X1 U16701 ( .A1(n15489), .A2(n15488), .A3(n15487), .ZN(n15565) );
  MUX2_X1 U16702 ( .A(n15490), .B(n15565), .S(n16526), .Z(n15491) );
  OAI21_X1 U16703 ( .B1(n15568), .B2(n15530), .A(n15491), .ZN(P2_U3524) );
  OAI211_X1 U16704 ( .C1(n15550), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15569) );
  MUX2_X1 U16705 ( .A(n15569), .B(P2_REG1_REG_24__SCAN_IN), .S(n16525), .Z(
        n15495) );
  AOI21_X1 U16706 ( .B1(n15536), .B2(n15496), .A(n15495), .ZN(n15497) );
  INV_X1 U16707 ( .A(n15497), .ZN(P2_U3523) );
  NAND2_X1 U16708 ( .A1(n15498), .A2(n16523), .ZN(n15500) );
  NAND3_X1 U16709 ( .A1(n15501), .A2(n15500), .A3(n15499), .ZN(n15573) );
  MUX2_X1 U16710 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n15573), .S(n16526), .Z(
        n15502) );
  AOI21_X1 U16711 ( .B1(n15536), .B2(n15503), .A(n15502), .ZN(n15504) );
  INV_X1 U16712 ( .A(n15504), .ZN(P2_U3522) );
  AOI211_X1 U16713 ( .C1(n16523), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        n15577) );
  MUX2_X1 U16714 ( .A(n15508), .B(n15577), .S(n16526), .Z(n15509) );
  OAI21_X1 U16715 ( .B1(n15580), .B2(n15530), .A(n15509), .ZN(P2_U3521) );
  AOI211_X1 U16716 ( .C1(n15546), .C2(n8227), .A(n15511), .B(n15510), .ZN(
        n15512) );
  OAI21_X1 U16717 ( .B1(n15550), .B2(n15513), .A(n15512), .ZN(n15581) );
  MUX2_X1 U16718 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n15581), .S(n16526), .Z(
        P2_U3520) );
  OAI211_X1 U16719 ( .C1(n15550), .C2(n15516), .A(n15515), .B(n15514), .ZN(
        n15582) );
  MUX2_X1 U16720 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n15582), .S(n16526), .Z(
        n15517) );
  AOI21_X1 U16721 ( .B1(n15536), .B2(n15518), .A(n15517), .ZN(n15519) );
  INV_X1 U16722 ( .A(n15519), .ZN(P2_U3519) );
  AOI211_X1 U16723 ( .C1(n11714), .C2(n15522), .A(n15521), .B(n15520), .ZN(
        n15587) );
  MUX2_X1 U16724 ( .A(n15523), .B(n15587), .S(n16526), .Z(n15524) );
  OAI21_X1 U16725 ( .B1(n15590), .B2(n15530), .A(n15524), .ZN(P2_U3518) );
  INV_X1 U16726 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15528) );
  AOI211_X1 U16727 ( .C1(n16523), .C2(n15527), .A(n15526), .B(n15525), .ZN(
        n15591) );
  MUX2_X1 U16728 ( .A(n15528), .B(n15591), .S(n16526), .Z(n15529) );
  OAI21_X1 U16729 ( .B1(n15595), .B2(n15530), .A(n15529), .ZN(P2_U3517) );
  AND2_X1 U16730 ( .A1(n15531), .A2(n16523), .ZN(n15533) );
  MUX2_X1 U16731 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n15596), .S(n16526), .Z(
        n15535) );
  AOI21_X1 U16732 ( .B1(n15536), .B2(n15598), .A(n15535), .ZN(n15537) );
  INV_X1 U16733 ( .A(n15537), .ZN(P2_U3516) );
  AOI21_X1 U16734 ( .B1(n15546), .B2(n15539), .A(n15538), .ZN(n15540) );
  OAI211_X1 U16735 ( .C1(n15543), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        n15601) );
  MUX2_X1 U16736 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n15601), .S(n16526), .Z(
        P2_U3515) );
  AOI21_X1 U16737 ( .B1(n15546), .B2(n15545), .A(n15544), .ZN(n15547) );
  OAI211_X1 U16738 ( .C1(n15550), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        n15602) );
  MUX2_X1 U16739 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n15602), .S(n16526), .Z(
        P2_U3513) );
  MUX2_X1 U16740 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n15551), .S(n16526), .Z(
        P2_U3499) );
  INV_X1 U16741 ( .A(n15552), .ZN(n15556) );
  OAI21_X1 U16742 ( .B1(n15556), .B2(n15594), .A(n15555), .ZN(P2_U3498) );
  MUX2_X1 U16743 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n15557), .S(n16529), .Z(
        n15558) );
  INV_X1 U16744 ( .A(n15558), .ZN(n15559) );
  OAI21_X1 U16745 ( .B1(n15560), .B2(n15594), .A(n15559), .ZN(P2_U3497) );
  MUX2_X1 U16746 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n15562), .S(n15586), .Z(
        P2_U3495) );
  MUX2_X1 U16747 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n15563), .S(n15586), .Z(
        P2_U3494) );
  MUX2_X1 U16748 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n15564), .S(n15586), .Z(
        P2_U3493) );
  INV_X1 U16749 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15566) );
  MUX2_X1 U16750 ( .A(n15566), .B(n15565), .S(n15586), .Z(n15567) );
  OAI21_X1 U16751 ( .B1(n15568), .B2(n15594), .A(n15567), .ZN(P2_U3492) );
  MUX2_X1 U16752 ( .A(n15569), .B(P2_REG0_REG_24__SCAN_IN), .S(n16527), .Z(
        n15570) );
  INV_X1 U16753 ( .A(n15570), .ZN(n15571) );
  OAI21_X1 U16754 ( .B1(n15572), .B2(n15594), .A(n15571), .ZN(P2_U3491) );
  MUX2_X1 U16755 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n15573), .S(n16529), .Z(
        n15574) );
  INV_X1 U16756 ( .A(n15574), .ZN(n15575) );
  OAI21_X1 U16757 ( .B1(n15576), .B2(n15594), .A(n15575), .ZN(P2_U3490) );
  INV_X1 U16758 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n15578) );
  MUX2_X1 U16759 ( .A(n15578), .B(n15577), .S(n16529), .Z(n15579) );
  OAI21_X1 U16760 ( .B1(n15580), .B2(n15594), .A(n15579), .ZN(P2_U3489) );
  MUX2_X1 U16761 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n15581), .S(n16529), .Z(
        P2_U3488) );
  MUX2_X1 U16762 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n15582), .S(n15586), .Z(
        n15583) );
  INV_X1 U16763 ( .A(n15583), .ZN(n15584) );
  OAI21_X1 U16764 ( .B1(n15585), .B2(n15594), .A(n15584), .ZN(P2_U3487) );
  INV_X1 U16765 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15588) );
  MUX2_X1 U16766 ( .A(n15588), .B(n15587), .S(n15586), .Z(n15589) );
  OAI21_X1 U16767 ( .B1(n15590), .B2(n15594), .A(n15589), .ZN(P2_U3486) );
  INV_X1 U16768 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n15592) );
  MUX2_X1 U16769 ( .A(n15592), .B(n15591), .S(n16529), .Z(n15593) );
  OAI21_X1 U16770 ( .B1(n15595), .B2(n15594), .A(n15593), .ZN(P2_U3484) );
  MUX2_X1 U16771 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n15596), .S(n16529), .Z(
        n15597) );
  AOI21_X1 U16772 ( .B1(n15599), .B2(n15598), .A(n15597), .ZN(n15600) );
  INV_X1 U16773 ( .A(n15600), .ZN(P2_U3481) );
  MUX2_X1 U16774 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n15601), .S(n16529), .Z(
        P2_U3478) );
  MUX2_X1 U16775 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n15602), .S(n16529), .Z(
        P2_U3472) );
  INV_X1 U16776 ( .A(n15603), .ZN(n16168) );
  INV_X1 U16777 ( .A(n15604), .ZN(n15606) );
  NOR4_X1 U16778 ( .A1(n15606), .A2(P2_IR_REG_30__SCAN_IN), .A3(n15605), .A4(
        P2_U3088), .ZN(n15607) );
  AOI21_X1 U16779 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n15608), .A(n15607), 
        .ZN(n15609) );
  OAI21_X1 U16780 ( .B1(n16168), .B2(n15626), .A(n15609), .ZN(P2_U3296) );
  OAI222_X1 U16781 ( .A1(P2_U3088), .A2(n15612), .B1(n15626), .B2(n15611), 
        .C1(n15610), .C2(n15628), .ZN(P2_U3298) );
  NAND2_X1 U16782 ( .A1(n15613), .A2(n15617), .ZN(n15615) );
  OAI211_X1 U16783 ( .C1(n15628), .C2(n15616), .A(n15615), .B(n15614), .ZN(
        P2_U3299) );
  NAND2_X1 U16784 ( .A1(n16169), .A2(n15617), .ZN(n15619) );
  OAI211_X1 U16785 ( .C1(n15628), .C2(n15620), .A(n15619), .B(n15618), .ZN(
        P2_U3300) );
  INV_X1 U16786 ( .A(n15621), .ZN(n16173) );
  OAI222_X1 U16787 ( .A1(n15628), .A2(n15623), .B1(n15626), .B2(n16173), .C1(
        P2_U3088), .C2(n15622), .ZN(P2_U3301) );
  INV_X1 U16788 ( .A(n15624), .ZN(n16177) );
  OAI222_X1 U16789 ( .A1(n15628), .A2(n15627), .B1(n15626), .B2(n16177), .C1(
        n15625), .C2(P2_U3088), .ZN(P2_U3302) );
  MUX2_X1 U16790 ( .A(P2_IR_REG_0__SCAN_IN), .B(n15629), .S(P2_U3088), .Z(
        P2_U3327) );
  XOR2_X1 U16791 ( .A(n15631), .B(n15630), .Z(n15637) );
  NAND2_X1 U16792 ( .A1(n15733), .A2(n15956), .ZN(n15633) );
  NAND2_X1 U16793 ( .A1(n15735), .A2(n15955), .ZN(n15632) );
  NAND2_X1 U16794 ( .A1(n15633), .A2(n15632), .ZN(n16061) );
  AOI22_X1 U16795 ( .A1(n16716), .A2(n16061), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15634) );
  OAI21_X1 U16796 ( .B1(n15849), .B2(n16723), .A(n15634), .ZN(n15635) );
  AOI21_X1 U16797 ( .B1(n16062), .B2(n16719), .A(n15635), .ZN(n15636) );
  OAI21_X1 U16798 ( .B1(n15637), .B2(n15729), .A(n15636), .ZN(P1_U3214) );
  AOI21_X1 U16799 ( .B1(n15640), .B2(n15639), .A(n15638), .ZN(n15647) );
  OAI21_X1 U16800 ( .B1(n16723), .B2(n15642), .A(n15641), .ZN(n15645) );
  OAI22_X1 U16801 ( .A1(n16030), .A2(n15717), .B1(n15716), .B2(n15643), .ZN(
        n15644) );
  AOI211_X1 U16802 ( .C1(n16137), .C2(n16719), .A(n15645), .B(n15644), .ZN(
        n15646) );
  OAI21_X1 U16803 ( .B1(n15647), .B2(n15729), .A(n15646), .ZN(P1_U3215) );
  XOR2_X1 U16804 ( .A(n15649), .B(n15648), .Z(n15653) );
  OAI22_X1 U16805 ( .A1(n15674), .A2(n16029), .B1(n15665), .B2(n16031), .ZN(
        n15902) );
  AOI22_X1 U16806 ( .A1(n16716), .A2(n15902), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15650) );
  OAI21_X1 U16807 ( .B1(n15906), .B2(n16723), .A(n15650), .ZN(n15651) );
  AOI21_X1 U16808 ( .B1(n16088), .B2(n16719), .A(n15651), .ZN(n15652) );
  OAI21_X1 U16809 ( .B1(n15653), .B2(n15729), .A(n15652), .ZN(P1_U3216) );
  XOR2_X1 U16810 ( .A(n15655), .B(n15654), .Z(n15660) );
  OAI21_X1 U16811 ( .B1(n15979), .B2(n16723), .A(n15656), .ZN(n15658) );
  OAI22_X1 U16812 ( .A1(n15976), .A2(n15717), .B1(n15977), .B2(n15716), .ZN(
        n15657) );
  AOI211_X1 U16813 ( .C1(n16111), .C2(n16719), .A(n15658), .B(n15657), .ZN(
        n15659) );
  OAI21_X1 U16814 ( .B1(n15660), .B2(n15729), .A(n15659), .ZN(P1_U3219) );
  INV_X1 U16815 ( .A(n15661), .ZN(n15662) );
  AOI21_X1 U16816 ( .B1(n15664), .B2(n15663), .A(n15662), .ZN(n15671) );
  NOR2_X1 U16817 ( .A1(n15665), .A2(n16029), .ZN(n15666) );
  AOI21_X1 U16818 ( .B1(n15739), .B2(n15955), .A(n15666), .ZN(n16097) );
  NOR2_X1 U16819 ( .A1(n16097), .A2(n15691), .ZN(n15669) );
  INV_X1 U16820 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15667) );
  OAI22_X1 U16821 ( .A1(n15942), .A2(n16723), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15667), .ZN(n15668) );
  AOI211_X1 U16822 ( .C1(n15937), .C2(n16719), .A(n15669), .B(n15668), .ZN(
        n15670) );
  OAI21_X1 U16823 ( .B1(n15671), .B2(n15729), .A(n15670), .ZN(P1_U3223) );
  XOR2_X1 U16824 ( .A(n15673), .B(n15672), .Z(n15679) );
  OAI22_X1 U16825 ( .A1(n15675), .A2(n16029), .B1(n15674), .B2(n16031), .ZN(
        n16073) );
  AOI22_X1 U16826 ( .A1(n16073), .A2(n16716), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15676) );
  OAI21_X1 U16827 ( .B1(n15878), .B2(n16723), .A(n15676), .ZN(n15677) );
  AOI21_X1 U16828 ( .B1(n16074), .B2(n16719), .A(n15677), .ZN(n15678) );
  OAI21_X1 U16829 ( .B1(n15679), .B2(n15729), .A(n15678), .ZN(P1_U3225) );
  XOR2_X1 U16830 ( .A(n15680), .B(n15681), .Z(n15686) );
  OAI21_X1 U16831 ( .B1(n16723), .B2(n16035), .A(n15682), .ZN(n15684) );
  OAI22_X1 U16832 ( .A1(n16028), .A2(n15717), .B1(n15716), .B2(n16030), .ZN(
        n15683) );
  AOI211_X1 U16833 ( .C1(n16129), .C2(n16719), .A(n15684), .B(n15683), .ZN(
        n15685) );
  OAI21_X1 U16834 ( .B1(n15686), .B2(n15729), .A(n15685), .ZN(P1_U3226) );
  XOR2_X1 U16835 ( .A(n15688), .B(n15687), .Z(n15695) );
  NOR2_X1 U16836 ( .A1(n16723), .A2(n16013), .ZN(n15693) );
  AND2_X1 U16837 ( .A1(n15742), .A2(n15955), .ZN(n15689) );
  AOI21_X1 U16838 ( .B1(n15740), .B2(n15956), .A(n15689), .ZN(n16008) );
  OAI21_X1 U16839 ( .B1(n16008), .B2(n15691), .A(n15690), .ZN(n15692) );
  AOI211_X1 U16840 ( .C1(n16123), .C2(n16719), .A(n15693), .B(n15692), .ZN(
        n15694) );
  OAI21_X1 U16841 ( .B1(n15695), .B2(n15729), .A(n15694), .ZN(P1_U3228) );
  XOR2_X1 U16842 ( .A(n15697), .B(n15696), .Z(n15702) );
  INV_X1 U16843 ( .A(n15736), .ZN(n15698) );
  INV_X1 U16844 ( .A(n15917), .ZN(n15707) );
  OAI22_X1 U16845 ( .A1(n15698), .A2(n16029), .B1(n15707), .B2(n16031), .ZN(
        n15884) );
  AOI22_X1 U16846 ( .A1(n16716), .A2(n15884), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15699) );
  OAI21_X1 U16847 ( .B1(n15890), .B2(n16723), .A(n15699), .ZN(n15700) );
  AOI21_X1 U16848 ( .B1(n16082), .B2(n16719), .A(n15700), .ZN(n15701) );
  OAI21_X1 U16849 ( .B1(n15702), .B2(n15729), .A(n15701), .ZN(P1_U3229) );
  OAI21_X1 U16850 ( .B1(n15705), .B2(n15704), .A(n15703), .ZN(n15706) );
  NAND2_X1 U16851 ( .A1(n15706), .A2(n16714), .ZN(n15711) );
  NOR2_X1 U16852 ( .A1(n16723), .A2(n15922), .ZN(n15709) );
  OAI22_X1 U16853 ( .A1(n8149), .A2(n15716), .B1(n15707), .B2(n15717), .ZN(
        n15708) );
  AOI211_X1 U16854 ( .C1(P1_REG3_REG_22__SCAN_IN), .C2(P1_U3086), .A(n15709), 
        .B(n15708), .ZN(n15710) );
  OAI211_X1 U16855 ( .C1(n15712), .C2(n15921), .A(n15711), .B(n15710), .ZN(
        P1_U3235) );
  XOR2_X1 U16856 ( .A(n15713), .B(n15714), .Z(n15721) );
  OAI21_X1 U16857 ( .B1(n16723), .B2(n16000), .A(n15715), .ZN(n15719) );
  OAI22_X1 U16858 ( .A1(n15996), .A2(n15717), .B1(n16028), .B2(n15716), .ZN(
        n15718) );
  AOI211_X1 U16859 ( .C1(n16118), .C2(n16719), .A(n15719), .B(n15718), .ZN(
        n15720) );
  OAI21_X1 U16860 ( .B1(n15721), .B2(n15729), .A(n15720), .ZN(P1_U3238) );
  XOR2_X1 U16861 ( .A(n15723), .B(n15722), .Z(n15730) );
  NAND2_X1 U16862 ( .A1(n15736), .A2(n15955), .ZN(n15725) );
  NAND2_X1 U16863 ( .A1(n15734), .A2(n15956), .ZN(n15724) );
  NAND2_X1 U16864 ( .A1(n15725), .A2(n15724), .ZN(n16068) );
  AOI22_X1 U16865 ( .A1(n16716), .A2(n16068), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15726) );
  OAI21_X1 U16866 ( .B1(n15860), .B2(n16723), .A(n15726), .ZN(n15727) );
  AOI21_X1 U16867 ( .B1(n16069), .B2(n16719), .A(n15727), .ZN(n15728) );
  OAI21_X1 U16868 ( .B1(n15730), .B2(n15729), .A(n15728), .ZN(P1_U3240) );
  MUX2_X1 U16869 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15731), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16870 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15732), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16871 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15733), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16872 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15734), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16873 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15735), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16874 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15736), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16875 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15737), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16876 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15917), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16877 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15738), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16878 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15957), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16879 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15739), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16880 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15740), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16881 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15741), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16882 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15742), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16883 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15743), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16884 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15744), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16885 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15745), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16886 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15746), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16887 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15747), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16888 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15748), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16889 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15749), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16890 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15750), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16891 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15751), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16892 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15752), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16893 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15753), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16894 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15754), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16895 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15755), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16896 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n15756), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16897 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15757), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16898 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8099), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI21_X1 U16899 ( .B1(n16280), .B2(n15758), .A(n10784), .ZN(n16279) );
  MUX2_X1 U16900 ( .A(n15760), .B(n15759), .S(n16280), .Z(n15762) );
  NAND2_X1 U16901 ( .A1(n15762), .A2(n15761), .ZN(n15763) );
  OAI211_X1 U16902 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n16279), .A(n15763), .B(
        P1_U4016), .ZN(n15796) );
  AOI22_X1 U16903 ( .A1(n16283), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n15775) );
  XOR2_X1 U16904 ( .A(n15765), .B(n15764), .Z(n15773) );
  OAI21_X1 U16905 ( .B1(n15768), .B2(n15767), .A(n15766), .ZN(n15771) );
  NAND2_X1 U16906 ( .A1(n16294), .A2(n15769), .ZN(n15770) );
  OAI21_X1 U16907 ( .B1(n16297), .B2(n15771), .A(n15770), .ZN(n15772) );
  AOI21_X1 U16908 ( .B1(n15797), .B2(n15773), .A(n15772), .ZN(n15774) );
  NAND3_X1 U16909 ( .A1(n15796), .A2(n15775), .A3(n15774), .ZN(P1_U3245) );
  NAND2_X1 U16910 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n16283), .ZN(n15795) );
  INV_X1 U16911 ( .A(n15776), .ZN(n15781) );
  NOR3_X1 U16912 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n15780) );
  NOR3_X1 U16913 ( .A1(n16291), .A2(n15781), .A3(n15780), .ZN(n15793) );
  MUX2_X1 U16914 ( .A(n11359), .B(P1_REG1_REG_4__SCAN_IN), .S(n15782), .Z(
        n15783) );
  NAND3_X1 U16915 ( .A1(n15785), .A2(n15784), .A3(n15783), .ZN(n15786) );
  NAND3_X1 U16916 ( .A1(n15807), .A2(n15787), .A3(n15786), .ZN(n15789) );
  OAI211_X1 U16917 ( .C1(n15791), .C2(n15790), .A(n15789), .B(n15788), .ZN(
        n15792) );
  NOR2_X1 U16918 ( .A1(n15793), .A2(n15792), .ZN(n15794) );
  NAND3_X1 U16919 ( .A1(n15796), .A2(n15795), .A3(n15794), .ZN(P1_U3247) );
  OAI211_X1 U16920 ( .C1(n15800), .C2(n15799), .A(n15798), .B(n15797), .ZN(
        n15812) );
  INV_X1 U16921 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n16413) );
  NOR2_X1 U16922 ( .A1(n16301), .A2(n16413), .ZN(n15801) );
  AOI211_X1 U16923 ( .C1(n16294), .C2(n15804), .A(n15802), .B(n15801), .ZN(
        n15811) );
  INV_X1 U16924 ( .A(n15803), .ZN(n15809) );
  MUX2_X1 U16925 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15805), .S(n15804), .Z(
        n15808) );
  OAI211_X1 U16926 ( .C1(n15809), .C2(n15808), .A(n15807), .B(n15806), .ZN(
        n15810) );
  NAND3_X1 U16927 ( .A1(n15812), .A2(n15811), .A3(n15810), .ZN(P1_U3256) );
  NAND2_X1 U16928 ( .A1(n16045), .A2(n15820), .ZN(n15819) );
  XNOR2_X1 U16929 ( .A(n15819), .B(n16042), .ZN(n15813) );
  NAND2_X1 U16930 ( .A1(n15813), .A2(n16698), .ZN(n16041) );
  NAND2_X1 U16931 ( .A1(n16642), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n15816) );
  NAND2_X1 U16932 ( .A1(n15815), .A2(n15814), .ZN(n16043) );
  OR2_X1 U16933 ( .A1(n16642), .A2(n16043), .ZN(n15821) );
  OAI211_X1 U16934 ( .C1(n16042), .C2(n16587), .A(n15816), .B(n15821), .ZN(
        n15817) );
  INV_X1 U16935 ( .A(n15817), .ZN(n15818) );
  OAI21_X1 U16936 ( .B1(n16041), .B2(n15825), .A(n15818), .ZN(P1_U3263) );
  OAI211_X1 U16937 ( .C1(n15820), .C2(n16045), .A(n15819), .B(n16698), .ZN(
        n16044) );
  INV_X1 U16938 ( .A(n15821), .ZN(n15823) );
  NOR2_X1 U16939 ( .A1(n16045), .A2(n16587), .ZN(n15822) );
  AOI211_X1 U16940 ( .C1(n16642), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15823), 
        .B(n15822), .ZN(n15824) );
  OAI21_X1 U16941 ( .B1(n15825), .B2(n16044), .A(n15824), .ZN(P1_U3264) );
  XNOR2_X1 U16942 ( .A(n15826), .B(n8057), .ZN(n15830) );
  OAI22_X1 U16943 ( .A1(n15828), .A2(n16031), .B1(n15827), .B2(n16029), .ZN(
        n15829) );
  AOI21_X2 U16944 ( .B1(n15830), .B2(n16623), .A(n15829), .ZN(n16057) );
  OAI21_X1 U16945 ( .B1(n7495), .B2(n15832), .A(n15831), .ZN(n16058) );
  INV_X1 U16946 ( .A(n16058), .ZN(n15841) );
  OR2_X1 U16947 ( .A1(n15839), .A2(n7470), .ZN(n15833) );
  AND2_X1 U16948 ( .A1(n15834), .A2(n15833), .ZN(n16055) );
  NAND2_X1 U16949 ( .A1(n16055), .A2(n15987), .ZN(n15838) );
  INV_X1 U16950 ( .A(n15835), .ZN(n15836) );
  AOI22_X1 U16951 ( .A1(n16642), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n15836), 
        .B2(n16631), .ZN(n15837) );
  OAI211_X1 U16952 ( .C1(n15839), .C2(n16587), .A(n15838), .B(n15837), .ZN(
        n15840) );
  AOI21_X1 U16953 ( .B1(n15841), .B2(n15929), .A(n15840), .ZN(n15842) );
  OAI21_X1 U16954 ( .B1(n16057), .B2(n16642), .A(n15842), .ZN(P1_U3265) );
  AOI21_X1 U16955 ( .B1(n15846), .B2(n15844), .A(n15843), .ZN(n16065) );
  XNOR2_X1 U16956 ( .A(n15845), .B(n15846), .ZN(n16059) );
  NAND2_X1 U16957 ( .A1(n16059), .A2(n15948), .ZN(n15855) );
  NAND2_X1 U16958 ( .A1(n16062), .A2(n15858), .ZN(n15847) );
  NAND2_X1 U16959 ( .A1(n15847), .A2(n16698), .ZN(n15848) );
  NOR2_X1 U16960 ( .A1(n7470), .A2(n15848), .ZN(n16060) );
  INV_X1 U16961 ( .A(n16061), .ZN(n15850) );
  OAI22_X1 U16962 ( .A1(n16642), .A2(n15850), .B1(n15849), .B2(n16036), .ZN(
        n15851) );
  AOI21_X1 U16963 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(n16642), .A(n15851), 
        .ZN(n15852) );
  OAI21_X1 U16964 ( .B1(n8196), .B2(n16587), .A(n15852), .ZN(n15853) );
  AOI21_X1 U16965 ( .B1(n16060), .B2(n16636), .A(n15853), .ZN(n15854) );
  OAI211_X1 U16966 ( .C1(n16065), .C2(n15897), .A(n15855), .B(n15854), .ZN(
        P1_U3266) );
  XNOR2_X1 U16967 ( .A(n7548), .B(n15856), .ZN(n16072) );
  XNOR2_X1 U16968 ( .A(n15857), .B(n15856), .ZN(n16066) );
  AOI21_X1 U16969 ( .B1(n16069), .B2(n15870), .A(n16686), .ZN(n15859) );
  AND2_X1 U16970 ( .A1(n15859), .A2(n15858), .ZN(n16067) );
  NAND2_X1 U16971 ( .A1(n16067), .A2(n16636), .ZN(n15864) );
  INV_X1 U16972 ( .A(n16068), .ZN(n15861) );
  OAI22_X1 U16973 ( .A1(n16642), .A2(n15861), .B1(n15860), .B2(n16036), .ZN(
        n15862) );
  AOI21_X1 U16974 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n16642), .A(n15862), 
        .ZN(n15863) );
  OAI211_X1 U16975 ( .C1(n15865), .C2(n16587), .A(n15864), .B(n15863), .ZN(
        n15866) );
  AOI21_X1 U16976 ( .B1(n16066), .B2(n15948), .A(n15866), .ZN(n15867) );
  OAI21_X1 U16977 ( .B1(n16072), .B2(n16040), .A(n15867), .ZN(P1_U3267) );
  AOI21_X1 U16978 ( .B1(n15873), .B2(n15869), .A(n15868), .ZN(n16075) );
  INV_X1 U16979 ( .A(n16075), .ZN(n15883) );
  OAI211_X1 U16980 ( .C1(n15871), .C2(n15887), .A(n16698), .B(n15870), .ZN(
        n16076) );
  OAI21_X1 U16981 ( .B1(n15874), .B2(n15873), .A(n15872), .ZN(n15875) );
  NAND2_X1 U16982 ( .A1(n15875), .A2(n16623), .ZN(n16079) );
  INV_X1 U16983 ( .A(n16073), .ZN(n15876) );
  OAI211_X1 U16984 ( .C1(n10650), .C2(n16076), .A(n16079), .B(n15876), .ZN(
        n15877) );
  NAND2_X1 U16985 ( .A1(n15877), .A2(n16014), .ZN(n15882) );
  OAI22_X1 U16986 ( .A1(n16014), .A2(n15879), .B1(n15878), .B2(n16036), .ZN(
        n15880) );
  AOI21_X1 U16987 ( .B1(n16074), .B2(n16632), .A(n15880), .ZN(n15881) );
  OAI211_X1 U16988 ( .C1(n15883), .C2(n16040), .A(n15882), .B(n15881), .ZN(
        P1_U3268) );
  AOI21_X1 U16989 ( .B1(n7508), .B2(n15895), .A(n16702), .ZN(n15886) );
  AOI21_X1 U16990 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n16084) );
  INV_X1 U16991 ( .A(n15904), .ZN(n15888) );
  AOI211_X1 U16992 ( .C1(n16082), .C2(n15888), .A(n16686), .B(n15887), .ZN(
        n16081) );
  NOR2_X1 U16993 ( .A1(n15889), .A2(n16587), .ZN(n15893) );
  OAI22_X1 U16994 ( .A1(n16014), .A2(n15891), .B1(n15890), .B2(n16036), .ZN(
        n15892) );
  AOI211_X1 U16995 ( .C1(n16081), .C2(n16636), .A(n15893), .B(n15892), .ZN(
        n15900) );
  OAI21_X1 U16996 ( .B1(n15896), .B2(n15895), .A(n15894), .ZN(n16080) );
  INV_X1 U16997 ( .A(n15897), .ZN(n15898) );
  NAND2_X1 U16998 ( .A1(n16080), .A2(n15898), .ZN(n15899) );
  OAI211_X1 U16999 ( .C1(n16084), .C2(n16642), .A(n15900), .B(n15899), .ZN(
        P1_U3269) );
  XNOR2_X1 U17000 ( .A(n15901), .B(n15912), .ZN(n15903) );
  AOI21_X1 U17001 ( .B1(n15903), .B2(n16623), .A(n15902), .ZN(n16090) );
  AOI211_X1 U17002 ( .C1(n16088), .C2(n15919), .A(n16686), .B(n15904), .ZN(
        n16087) );
  NOR2_X1 U17003 ( .A1(n15905), .A2(n16587), .ZN(n15909) );
  OAI22_X1 U17004 ( .A1(n16014), .A2(n15907), .B1(n15906), .B2(n16036), .ZN(
        n15908) );
  AOI211_X1 U17005 ( .C1(n16087), .C2(n16636), .A(n15909), .B(n15908), .ZN(
        n15914) );
  AOI21_X1 U17006 ( .B1(n15912), .B2(n15911), .A(n15910), .ZN(n16086) );
  NAND2_X1 U17007 ( .A1(n16086), .A2(n15929), .ZN(n15913) );
  OAI211_X1 U17008 ( .C1(n16090), .C2(n16642), .A(n15914), .B(n15913), .ZN(
        P1_U3270) );
  OAI21_X1 U17009 ( .B1(n15916), .B2(n7525), .A(n15915), .ZN(n15918) );
  AOI222_X1 U17010 ( .A1(n16623), .A2(n15918), .B1(n15957), .B2(n15955), .C1(
        n15917), .C2(n15956), .ZN(n16095) );
  INV_X1 U17011 ( .A(n15919), .ZN(n15920) );
  AOI21_X1 U17012 ( .B1(n8191), .B2(n8192), .A(n15920), .ZN(n16093) );
  NOR2_X1 U17013 ( .A1(n15921), .A2(n16587), .ZN(n15925) );
  OAI22_X1 U17014 ( .A1(n16014), .A2(n15923), .B1(n15922), .B2(n16036), .ZN(
        n15924) );
  AOI211_X1 U17015 ( .C1(n16093), .C2(n15987), .A(n15925), .B(n15924), .ZN(
        n15931) );
  OAI21_X1 U17016 ( .B1(n15928), .B2(n15927), .A(n15926), .ZN(n16092) );
  NAND2_X1 U17017 ( .A1(n16092), .A2(n15929), .ZN(n15930) );
  OAI211_X1 U17018 ( .C1(n16095), .C2(n16642), .A(n15931), .B(n15930), .ZN(
        P1_U3271) );
  XOR2_X1 U17019 ( .A(n15932), .B(n15934), .Z(n16102) );
  INV_X1 U17020 ( .A(n15933), .ZN(n15936) );
  AOI21_X1 U17021 ( .B1(n15936), .B2(n8047), .A(n15935), .ZN(n16100) );
  NAND2_X1 U17022 ( .A1(n15937), .A2(n15952), .ZN(n15938) );
  NAND2_X1 U17023 ( .A1(n15938), .A2(n16698), .ZN(n15939) );
  NOR2_X1 U17024 ( .A1(n15940), .A2(n15939), .ZN(n16099) );
  NAND2_X1 U17025 ( .A1(n16099), .A2(n16636), .ZN(n15946) );
  INV_X1 U17026 ( .A(n16097), .ZN(n15944) );
  INV_X1 U17027 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15941) );
  OAI22_X1 U17028 ( .A1(n15942), .A2(n16036), .B1(n15941), .B2(n16014), .ZN(
        n15943) );
  AOI21_X1 U17029 ( .B1(n15944), .B2(n16014), .A(n15943), .ZN(n15945) );
  OAI211_X1 U17030 ( .C1(n8066), .C2(n16587), .A(n15946), .B(n15945), .ZN(
        n15947) );
  AOI21_X1 U17031 ( .B1(n16100), .B2(n15948), .A(n15947), .ZN(n15949) );
  OAI21_X1 U17032 ( .B1(n16102), .B2(n16040), .A(n15949), .ZN(P1_U3272) );
  OAI21_X1 U17033 ( .B1(n15951), .B2(n15963), .A(n15950), .ZN(n16110) );
  INV_X1 U17034 ( .A(n15952), .ZN(n15953) );
  AOI21_X1 U17035 ( .B1(n15958), .B2(n15983), .A(n15953), .ZN(n16108) );
  AOI22_X1 U17036 ( .A1(n15957), .A2(n15956), .B1(n15955), .B2(n15954), .ZN(
        n16103) );
  NAND2_X1 U17037 ( .A1(n15958), .A2(n16632), .ZN(n15962) );
  INV_X1 U17038 ( .A(n15959), .ZN(n15960) );
  AOI22_X1 U17039 ( .A1(n15960), .A2(n16631), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n16642), .ZN(n15961) );
  OAI211_X1 U17040 ( .C1(n16642), .C2(n16103), .A(n15962), .B(n15961), .ZN(
        n15968) );
  NAND2_X1 U17041 ( .A1(n15964), .A2(n15963), .ZN(n15965) );
  NAND2_X1 U17042 ( .A1(n15966), .A2(n15965), .ZN(n16105) );
  NOR2_X1 U17043 ( .A1(n16105), .A2(n16040), .ZN(n15967) );
  AOI211_X1 U17044 ( .C1(n16108), .C2(n15987), .A(n15968), .B(n15967), .ZN(
        n15969) );
  OAI21_X1 U17045 ( .B1(n16110), .B2(n15970), .A(n15969), .ZN(P1_U3273) );
  XNOR2_X1 U17046 ( .A(n15971), .B(n15974), .ZN(n16115) );
  AOI21_X1 U17047 ( .B1(n15974), .B2(n15973), .A(n15972), .ZN(n15975) );
  OAI222_X1 U17048 ( .A1(n16031), .A2(n15977), .B1(n16029), .B2(n15976), .C1(
        n16702), .C2(n15975), .ZN(n15978) );
  INV_X1 U17049 ( .A(n15978), .ZN(n16114) );
  OAI21_X1 U17050 ( .B1(n15979), .B2(n16036), .A(n16114), .ZN(n15980) );
  NAND2_X1 U17051 ( .A1(n15980), .A2(n16014), .ZN(n15989) );
  INV_X1 U17052 ( .A(n15998), .ZN(n15981) );
  NAND2_X1 U17053 ( .A1(n15981), .A2(n16111), .ZN(n15982) );
  AND2_X1 U17054 ( .A1(n15983), .A2(n15982), .ZN(n16112) );
  INV_X1 U17055 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15984) );
  OAI22_X1 U17056 ( .A1(n15985), .A2(n16587), .B1(n16014), .B2(n15984), .ZN(
        n15986) );
  AOI21_X1 U17057 ( .B1(n16112), .B2(n15987), .A(n15986), .ZN(n15988) );
  OAI211_X1 U17058 ( .C1(n16115), .C2(n16040), .A(n15989), .B(n15988), .ZN(
        P1_U3274) );
  XNOR2_X1 U17059 ( .A(n15990), .B(n15991), .ZN(n15995) );
  INV_X1 U17060 ( .A(n15995), .ZN(n16121) );
  OAI211_X1 U17061 ( .C1(n15992), .C2(n15991), .A(n7565), .B(n16623), .ZN(
        n15993) );
  OAI21_X1 U17062 ( .B1(n16028), .B2(n16031), .A(n15993), .ZN(n15994) );
  AOI21_X1 U17063 ( .B1(n16579), .B2(n15995), .A(n15994), .ZN(n16120) );
  INV_X1 U17064 ( .A(n16120), .ZN(n15997) );
  NOR2_X1 U17065 ( .A1(n15996), .A2(n16029), .ZN(n16117) );
  OAI21_X1 U17066 ( .B1(n15997), .B2(n16117), .A(n16014), .ZN(n16005) );
  AOI211_X1 U17067 ( .C1(n16118), .C2(n16007), .A(n16686), .B(n15998), .ZN(
        n16116) );
  NOR2_X1 U17068 ( .A1(n15999), .A2(n16587), .ZN(n16003) );
  OAI22_X1 U17069 ( .A1(n16014), .A2(n16001), .B1(n16000), .B2(n16036), .ZN(
        n16002) );
  AOI211_X1 U17070 ( .C1(n16116), .C2(n16636), .A(n16003), .B(n16002), .ZN(
        n16004) );
  OAI211_X1 U17071 ( .C1(n16121), .C2(n16006), .A(n16005), .B(n16004), .ZN(
        P1_U3275) );
  OAI211_X1 U17072 ( .C1(n8184), .C2(n7599), .A(n16007), .B(n16698), .ZN(
        n16009) );
  NAND2_X1 U17073 ( .A1(n16009), .A2(n16008), .ZN(n16122) );
  XNOR2_X1 U17074 ( .A(n16010), .B(n16015), .ZN(n16011) );
  NAND2_X1 U17075 ( .A1(n16011), .A2(n16623), .ZN(n16125) );
  INV_X1 U17076 ( .A(n16125), .ZN(n16012) );
  AOI21_X1 U17077 ( .B1(n16033), .B2(n16122), .A(n16012), .ZN(n16021) );
  OAI22_X1 U17078 ( .A1(n16014), .A2(n13155), .B1(n16013), .B2(n16036), .ZN(
        n16019) );
  INV_X1 U17079 ( .A(n16015), .ZN(n16017) );
  OAI21_X1 U17080 ( .B1(n7606), .B2(n16017), .A(n16016), .ZN(n16126) );
  NOR2_X1 U17081 ( .A1(n16126), .A2(n16040), .ZN(n16018) );
  AOI211_X1 U17082 ( .C1(n16632), .C2(n16123), .A(n16019), .B(n16018), .ZN(
        n16020) );
  OAI21_X1 U17083 ( .B1(n16021), .B2(n16642), .A(n16020), .ZN(P1_U3276) );
  XOR2_X1 U17084 ( .A(n16022), .B(n16026), .Z(n16131) );
  INV_X1 U17085 ( .A(n16023), .ZN(n16024) );
  AOI21_X1 U17086 ( .B1(n16026), .B2(n16025), .A(n16024), .ZN(n16027) );
  OAI222_X1 U17087 ( .A1(n16031), .A2(n16030), .B1(n16029), .B2(n16028), .C1(
        n16702), .C2(n16027), .ZN(n16127) );
  XNOR2_X1 U17088 ( .A(n16129), .B(n7588), .ZN(n16032) );
  AND2_X1 U17089 ( .A1(n16032), .A2(n16698), .ZN(n16128) );
  NAND2_X1 U17090 ( .A1(n16128), .A2(n16033), .ZN(n16034) );
  OAI21_X1 U17091 ( .B1(n16036), .B2(n16035), .A(n16034), .ZN(n16037) );
  OAI21_X1 U17092 ( .B1(n16127), .B2(n16037), .A(n16014), .ZN(n16039) );
  AOI22_X1 U17093 ( .A1(n16129), .A2(n16632), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n16642), .ZN(n16038) );
  OAI211_X1 U17094 ( .C1(n16131), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P1_U3277) );
  OAI211_X1 U17095 ( .C1(n16042), .C2(n16684), .A(n16041), .B(n16043), .ZN(
        n16144) );
  MUX2_X1 U17096 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n16144), .S(n16708), .Z(
        P1_U3559) );
  OAI211_X1 U17097 ( .C1(n16045), .C2(n16684), .A(n16044), .B(n16043), .ZN(
        n16145) );
  MUX2_X1 U17098 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n16145), .S(n16708), .Z(
        P1_U3558) );
  OAI211_X1 U17099 ( .C1(n16048), .C2(n16684), .A(n16047), .B(n16046), .ZN(
        n16049) );
  NOR2_X1 U17100 ( .A1(n16050), .A2(n16049), .ZN(n16052) );
  MUX2_X1 U17101 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n16146), .S(n16708), .Z(
        P1_U3557) );
  AOI22_X1 U17102 ( .A1(n16055), .A2(n16698), .B1(n16696), .B2(n16054), .ZN(
        n16056) );
  OAI211_X1 U17103 ( .C1(n16142), .C2(n16058), .A(n16057), .B(n16056), .ZN(
        n16147) );
  MUX2_X1 U17104 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n16147), .S(n16708), .Z(
        P1_U3556) );
  NAND2_X1 U17105 ( .A1(n16059), .A2(n16623), .ZN(n16064) );
  AOI211_X1 U17106 ( .C1(n16696), .C2(n16062), .A(n16061), .B(n16060), .ZN(
        n16063) );
  OAI211_X1 U17107 ( .C1(n16142), .C2(n16065), .A(n16064), .B(n16063), .ZN(
        n16148) );
  MUX2_X1 U17108 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n16148), .S(n16708), .Z(
        P1_U3555) );
  NAND2_X1 U17109 ( .A1(n16066), .A2(n16623), .ZN(n16071) );
  AOI211_X1 U17110 ( .C1(n16696), .C2(n16069), .A(n16068), .B(n16067), .ZN(
        n16070) );
  OAI211_X1 U17111 ( .C1(n16142), .C2(n16072), .A(n16071), .B(n16070), .ZN(
        n16149) );
  MUX2_X1 U17112 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n16149), .S(n16708), .Z(
        P1_U3554) );
  AOI21_X1 U17113 ( .B1(n16074), .B2(n16696), .A(n16073), .ZN(n16078) );
  NAND2_X1 U17114 ( .A1(n16075), .A2(n16705), .ZN(n16077) );
  NAND4_X1 U17115 ( .A1(n16079), .A2(n16078), .A3(n16077), .A4(n16076), .ZN(
        n16150) );
  MUX2_X1 U17116 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n16150), .S(n16708), .Z(
        P1_U3553) );
  INV_X1 U17117 ( .A(n16080), .ZN(n16085) );
  AOI21_X1 U17118 ( .B1(n16696), .B2(n16082), .A(n16081), .ZN(n16083) );
  OAI211_X1 U17119 ( .C1(n16142), .C2(n16085), .A(n16084), .B(n16083), .ZN(
        n16151) );
  MUX2_X1 U17120 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n16151), .S(n16708), .Z(
        P1_U3552) );
  INV_X1 U17121 ( .A(n16086), .ZN(n16091) );
  AOI21_X1 U17122 ( .B1(n16696), .B2(n16088), .A(n16087), .ZN(n16089) );
  OAI211_X1 U17123 ( .C1(n16142), .C2(n16091), .A(n16090), .B(n16089), .ZN(
        n16152) );
  MUX2_X1 U17124 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n16152), .S(n16708), .Z(
        P1_U3551) );
  INV_X1 U17125 ( .A(n16092), .ZN(n16096) );
  AOI22_X1 U17126 ( .A1(n16093), .A2(n16698), .B1(n8191), .B2(n16696), .ZN(
        n16094) );
  OAI211_X1 U17127 ( .C1(n16142), .C2(n16096), .A(n16095), .B(n16094), .ZN(
        n16153) );
  MUX2_X1 U17128 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n16153), .S(n16708), .Z(
        P1_U3550) );
  OAI21_X1 U17129 ( .B1(n8066), .B2(n16684), .A(n16097), .ZN(n16098) );
  AOI211_X1 U17130 ( .C1(n16100), .C2(n16623), .A(n16099), .B(n16098), .ZN(
        n16101) );
  OAI21_X1 U17131 ( .B1(n16142), .B2(n16102), .A(n16101), .ZN(n16154) );
  MUX2_X1 U17132 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n16154), .S(n16708), .Z(
        P1_U3549) );
  OAI21_X1 U17133 ( .B1(n16104), .B2(n16684), .A(n16103), .ZN(n16107) );
  NOR2_X1 U17134 ( .A1(n16105), .A2(n16142), .ZN(n16106) );
  AOI211_X1 U17135 ( .C1(n16698), .C2(n16108), .A(n16107), .B(n16106), .ZN(
        n16109) );
  OAI21_X1 U17136 ( .B1(n16110), .B2(n16702), .A(n16109), .ZN(n16155) );
  MUX2_X1 U17137 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n16155), .S(n16708), .Z(
        P1_U3548) );
  AOI22_X1 U17138 ( .A1(n16112), .A2(n16698), .B1(n16696), .B2(n16111), .ZN(
        n16113) );
  OAI211_X1 U17139 ( .C1(n16142), .C2(n16115), .A(n16114), .B(n16113), .ZN(
        n16156) );
  MUX2_X1 U17140 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n16156), .S(n16708), .Z(
        P1_U3547) );
  AOI211_X1 U17141 ( .C1(n16696), .C2(n16118), .A(n16117), .B(n16116), .ZN(
        n16119) );
  OAI211_X1 U17142 ( .C1(n16121), .C2(n16602), .A(n16120), .B(n16119), .ZN(
        n16157) );
  MUX2_X1 U17143 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n16157), .S(n16708), .Z(
        P1_U3546) );
  AOI21_X1 U17144 ( .B1(n16696), .B2(n16123), .A(n16122), .ZN(n16124) );
  OAI211_X1 U17145 ( .C1(n16142), .C2(n16126), .A(n16125), .B(n16124), .ZN(
        n16158) );
  MUX2_X1 U17146 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n16158), .S(n16708), .Z(
        P1_U3545) );
  AOI211_X1 U17147 ( .C1(n16696), .C2(n16129), .A(n16128), .B(n16127), .ZN(
        n16130) );
  OAI21_X1 U17148 ( .B1(n16142), .B2(n16131), .A(n16130), .ZN(n16159) );
  MUX2_X1 U17149 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n16159), .S(n16708), .Z(
        P1_U3544) );
  AOI21_X1 U17150 ( .B1(n16696), .B2(n16718), .A(n16132), .ZN(n16133) );
  OAI211_X1 U17151 ( .C1(n16142), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        n16160) );
  MUX2_X1 U17152 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n16160), .S(n16708), .Z(
        P1_U3543) );
  INV_X1 U17153 ( .A(n16136), .ZN(n16140) );
  AOI22_X1 U17154 ( .A1(n16138), .A2(n16698), .B1(n16696), .B2(n16137), .ZN(
        n16139) );
  OAI211_X1 U17155 ( .C1(n16142), .C2(n16141), .A(n16140), .B(n16139), .ZN(
        n16161) );
  MUX2_X1 U17156 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n16161), .S(n16708), .Z(
        P1_U3542) );
  MUX2_X1 U17157 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n16143), .S(n16708), .Z(
        P1_U3528) );
  MUX2_X1 U17158 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n16144), .S(n16694), .Z(
        P1_U3527) );
  MUX2_X1 U17159 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n16145), .S(n16694), .Z(
        P1_U3526) );
  MUX2_X1 U17160 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n16146), .S(n16694), .Z(
        P1_U3525) );
  MUX2_X1 U17161 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n16147), .S(n16694), .Z(
        P1_U3524) );
  MUX2_X1 U17162 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n16148), .S(n16694), .Z(
        P1_U3523) );
  MUX2_X1 U17163 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n16149), .S(n16694), .Z(
        P1_U3522) );
  MUX2_X1 U17164 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n16150), .S(n16694), .Z(
        P1_U3521) );
  MUX2_X1 U17165 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n16151), .S(n16694), .Z(
        P1_U3520) );
  MUX2_X1 U17166 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n16152), .S(n16694), .Z(
        P1_U3519) );
  MUX2_X1 U17167 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n16153), .S(n16694), .Z(
        P1_U3518) );
  MUX2_X1 U17168 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n16154), .S(n16694), .Z(
        P1_U3517) );
  MUX2_X1 U17169 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n16155), .S(n16694), .Z(
        P1_U3516) );
  MUX2_X1 U17170 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n16156), .S(n16694), .Z(
        P1_U3515) );
  MUX2_X1 U17171 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n16157), .S(n16694), .Z(
        P1_U3513) );
  MUX2_X1 U17172 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n16158), .S(n16694), .Z(
        P1_U3510) );
  MUX2_X1 U17173 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n16159), .S(n16694), .Z(
        P1_U3507) );
  MUX2_X1 U17174 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n16160), .S(n16694), .Z(
        P1_U3504) );
  MUX2_X1 U17175 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n16161), .S(n16694), .Z(
        P1_U3501) );
  INV_X1 U17176 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n16162) );
  NAND3_X1 U17177 ( .A1(n16162), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n16164) );
  OAI22_X1 U17178 ( .A1(n16165), .A2(n16164), .B1(n16163), .B2(n16174), .ZN(
        n16166) );
  INV_X1 U17179 ( .A(n16166), .ZN(n16167) );
  OAI21_X1 U17180 ( .B1(n16168), .B2(n16178), .A(n16167), .ZN(P1_U3324) );
  INV_X1 U17181 ( .A(n16169), .ZN(n16171) );
  OAI222_X1 U17182 ( .A1(n16174), .A2(n16172), .B1(n16178), .B2(n16171), .C1(
        n16170), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U17183 ( .A1(n16175), .A2(P1_U3086), .B1(n16174), .B2(n8126), .C1(
        n16173), .C2(n16178), .ZN(P1_U3329) );
  OAI222_X1 U17184 ( .A1(n16174), .A2(n16179), .B1(n16178), .B2(n16177), .C1(
        n16176), .C2(P1_U3086), .ZN(P1_U3330) );
  MUX2_X1 U17185 ( .A(n16181), .B(n16180), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U17186 ( .A(n16182), .ZN(n16183) );
  MUX2_X1 U17187 ( .A(P1_IR_REG_0__SCAN_IN), .B(n16183), .S(P1_U3086), .Z(
        P1_U3355) );
  INV_X1 U17188 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n16184) );
  NOR2_X1 U17189 ( .A1(n16214), .A2(n16184), .ZN(P1_U3323) );
  INV_X1 U17190 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n16185) );
  NOR2_X1 U17191 ( .A1(n16214), .A2(n16185), .ZN(P1_U3322) );
  INV_X1 U17192 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n16186) );
  NOR2_X1 U17193 ( .A1(n16214), .A2(n16186), .ZN(P1_U3321) );
  INV_X1 U17194 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n16187) );
  NOR2_X1 U17195 ( .A1(n16214), .A2(n16187), .ZN(P1_U3320) );
  INV_X1 U17196 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n16188) );
  NOR2_X1 U17197 ( .A1(n16214), .A2(n16188), .ZN(P1_U3319) );
  INV_X1 U17198 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n16189) );
  NOR2_X1 U17199 ( .A1(n16214), .A2(n16189), .ZN(P1_U3318) );
  INV_X1 U17200 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n16190) );
  NOR2_X1 U17201 ( .A1(n16214), .A2(n16190), .ZN(P1_U3317) );
  INV_X1 U17202 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n16191) );
  NOR2_X1 U17203 ( .A1(n16214), .A2(n16191), .ZN(P1_U3316) );
  INV_X1 U17204 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n16192) );
  NOR2_X1 U17205 ( .A1(n16214), .A2(n16192), .ZN(P1_U3315) );
  INV_X1 U17206 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n16193) );
  NOR2_X1 U17207 ( .A1(n16214), .A2(n16193), .ZN(P1_U3314) );
  INV_X1 U17208 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n16194) );
  NOR2_X1 U17209 ( .A1(n16214), .A2(n16194), .ZN(P1_U3313) );
  INV_X1 U17210 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n16195) );
  NOR2_X1 U17211 ( .A1(n16214), .A2(n16195), .ZN(P1_U3312) );
  INV_X1 U17212 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n16196) );
  NOR2_X1 U17213 ( .A1(n16214), .A2(n16196), .ZN(P1_U3311) );
  INV_X1 U17214 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n16197) );
  NOR2_X1 U17215 ( .A1(n16214), .A2(n16197), .ZN(P1_U3310) );
  INV_X1 U17216 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n16198) );
  NOR2_X1 U17217 ( .A1(n16214), .A2(n16198), .ZN(P1_U3309) );
  INV_X1 U17218 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n16199) );
  NOR2_X1 U17219 ( .A1(n16214), .A2(n16199), .ZN(P1_U3308) );
  INV_X1 U17220 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n16200) );
  NOR2_X1 U17221 ( .A1(n16214), .A2(n16200), .ZN(P1_U3307) );
  INV_X1 U17222 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n16201) );
  NOR2_X1 U17223 ( .A1(n16214), .A2(n16201), .ZN(P1_U3306) );
  INV_X1 U17224 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n16202) );
  NOR2_X1 U17225 ( .A1(n16214), .A2(n16202), .ZN(P1_U3305) );
  INV_X1 U17226 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n16203) );
  NOR2_X1 U17227 ( .A1(n16214), .A2(n16203), .ZN(P1_U3304) );
  INV_X1 U17228 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n16204) );
  NOR2_X1 U17229 ( .A1(n16214), .A2(n16204), .ZN(P1_U3303) );
  INV_X1 U17230 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n16205) );
  NOR2_X1 U17231 ( .A1(n16214), .A2(n16205), .ZN(P1_U3302) );
  INV_X1 U17232 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n16206) );
  NOR2_X1 U17233 ( .A1(n16214), .A2(n16206), .ZN(P1_U3301) );
  INV_X1 U17234 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n16207) );
  NOR2_X1 U17235 ( .A1(n16214), .A2(n16207), .ZN(P1_U3300) );
  INV_X1 U17236 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n16208) );
  NOR2_X1 U17237 ( .A1(n16214), .A2(n16208), .ZN(P1_U3299) );
  INV_X1 U17238 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n16209) );
  NOR2_X1 U17239 ( .A1(n16214), .A2(n16209), .ZN(P1_U3298) );
  NOR2_X1 U17240 ( .A1(n16214), .A2(n16210), .ZN(P1_U3297) );
  NOR2_X1 U17241 ( .A1(n16214), .A2(n16211), .ZN(P1_U3296) );
  NOR2_X1 U17242 ( .A1(n16214), .A2(n16212), .ZN(P1_U3295) );
  NOR2_X1 U17243 ( .A1(n16214), .A2(n16213), .ZN(P1_U3294) );
  INV_X1 U17244 ( .A(n16215), .ZN(n16216) );
  AOI21_X1 U17245 ( .B1(n16217), .B2(n16220), .A(n16216), .ZN(P2_U3417) );
  AND2_X1 U17246 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n16219), .ZN(P2_U3295) );
  AND2_X1 U17247 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n16219), .ZN(P2_U3294) );
  AND2_X1 U17248 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n16219), .ZN(P2_U3293) );
  AND2_X1 U17249 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n16219), .ZN(P2_U3292) );
  AND2_X1 U17250 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n16219), .ZN(P2_U3291) );
  AND2_X1 U17251 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n16219), .ZN(P2_U3290) );
  AND2_X1 U17252 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n16219), .ZN(P2_U3289) );
  AND2_X1 U17253 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n16219), .ZN(P2_U3288) );
  AND2_X1 U17254 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n16219), .ZN(P2_U3287) );
  AND2_X1 U17255 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n16219), .ZN(P2_U3286) );
  AND2_X1 U17256 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n16219), .ZN(P2_U3285) );
  AND2_X1 U17257 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n16219), .ZN(P2_U3284) );
  AND2_X1 U17258 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n16219), .ZN(P2_U3283) );
  AND2_X1 U17259 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n16219), .ZN(P2_U3282) );
  AND2_X1 U17260 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n16219), .ZN(P2_U3281) );
  AND2_X1 U17261 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n16219), .ZN(P2_U3280) );
  AND2_X1 U17262 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n16219), .ZN(P2_U3279) );
  AND2_X1 U17263 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n16219), .ZN(P2_U3278) );
  AND2_X1 U17264 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n16219), .ZN(P2_U3277) );
  AND2_X1 U17265 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n16219), .ZN(P2_U3276) );
  AND2_X1 U17266 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n16219), .ZN(P2_U3275) );
  AND2_X1 U17267 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n16219), .ZN(P2_U3274) );
  AND2_X1 U17268 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n16219), .ZN(P2_U3273) );
  AND2_X1 U17269 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n16219), .ZN(P2_U3272) );
  AND2_X1 U17270 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n16219), .ZN(P2_U3271) );
  AND2_X1 U17271 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n16219), .ZN(P2_U3270) );
  AND2_X1 U17272 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n16219), .ZN(P2_U3269) );
  AND2_X1 U17273 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n16219), .ZN(P2_U3268) );
  AND2_X1 U17274 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n16219), .ZN(P2_U3267) );
  AND2_X1 U17275 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n16219), .ZN(P2_U3266) );
  NOR2_X1 U17276 ( .A1(n16224), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U17277 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n16221) );
  AOI22_X1 U17278 ( .A1(n16223), .A2(n16222), .B1(n16221), .B2(n16220), .ZN(
        P2_U3416) );
  AOI22_X1 U17279 ( .A1(n16224), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n16237) );
  NOR2_X1 U17280 ( .A1(n16226), .A2(n16225), .ZN(n16227) );
  AOI22_X1 U17281 ( .A1(n16230), .A2(n16229), .B1(n16270), .B2(n16228), .ZN(
        n16236) );
  AOI211_X1 U17282 ( .C1(n16233), .C2(n16232), .A(n16231), .B(n16272), .ZN(
        n16234) );
  INV_X1 U17283 ( .A(n16234), .ZN(n16235) );
  NAND3_X1 U17284 ( .A1(n16237), .A2(n16236), .A3(n16235), .ZN(P2_U3216) );
  INV_X1 U17285 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n16441) );
  AOI211_X1 U17286 ( .C1(n16240), .C2(n16239), .A(n16238), .B(n16264), .ZN(
        n16241) );
  AOI211_X1 U17287 ( .C1(n16243), .C2(n16270), .A(n16242), .B(n16241), .ZN(
        n16248) );
  OAI211_X1 U17288 ( .C1(n16246), .C2(n16245), .A(n16257), .B(n16244), .ZN(
        n16247) );
  OAI211_X1 U17289 ( .C1(n16278), .C2(n16441), .A(n16248), .B(n16247), .ZN(
        P2_U3230) );
  INV_X1 U17290 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n16437) );
  AND2_X1 U17291 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n16254) );
  AOI211_X1 U17292 ( .C1(n16252), .C2(n16251), .A(n16250), .B(n16264), .ZN(
        n16253) );
  AOI211_X1 U17293 ( .C1(n16270), .C2(n16255), .A(n16254), .B(n16253), .ZN(
        n16261) );
  OAI211_X1 U17294 ( .C1(n16259), .C2(n16258), .A(n16257), .B(n16256), .ZN(
        n16260) );
  OAI211_X1 U17295 ( .C1(n16278), .C2(n16437), .A(n16261), .B(n16260), .ZN(
        P2_U3231) );
  INV_X1 U17296 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n16386) );
  NOR2_X1 U17297 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n16262), .ZN(n16268) );
  AOI211_X1 U17298 ( .C1(n16266), .C2(n16265), .A(n16264), .B(n16263), .ZN(
        n16267) );
  AOI211_X1 U17299 ( .C1(n16270), .C2(n16269), .A(n16268), .B(n16267), .ZN(
        n16277) );
  AOI211_X1 U17300 ( .C1(n16274), .C2(n16273), .A(n16272), .B(n16271), .ZN(
        n16275) );
  INV_X1 U17301 ( .A(n16275), .ZN(n16276) );
  OAI211_X1 U17302 ( .C1(n16278), .C2(n16386), .A(n16277), .B(n16276), .ZN(
        P2_U3224) );
  OAI21_X1 U17303 ( .B1(n16280), .B2(P1_REG1_REG_0__SCAN_IN), .A(n16279), .ZN(
        n16282) );
  XNOR2_X1 U17304 ( .A(n16282), .B(n16281), .ZN(n16286) );
  AOI22_X1 U17305 ( .A1(n16283), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n16284) );
  OAI21_X1 U17306 ( .B1(n16286), .B2(n16285), .A(n16284), .ZN(P1_U3243) );
  AOI21_X1 U17307 ( .B1(n16288), .B2(P1_REG1_REG_15__SCAN_IN), .A(n16287), 
        .ZN(n16298) );
  AOI21_X1 U17308 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n16290), .A(n16289), 
        .ZN(n16292) );
  OR2_X1 U17309 ( .A1(n16292), .A2(n16291), .ZN(n16296) );
  NAND2_X1 U17310 ( .A1(n16294), .A2(n16293), .ZN(n16295) );
  OAI211_X1 U17311 ( .C1(n16298), .C2(n16297), .A(n16296), .B(n16295), .ZN(
        n16299) );
  INV_X1 U17312 ( .A(n16299), .ZN(n16300) );
  NAND2_X1 U17313 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n16720)
         );
  OAI211_X1 U17314 ( .C1(n16429), .C2(n16301), .A(n16300), .B(n16720), .ZN(
        P1_U3258) );
  NOR2_X1 U17315 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n16310), .ZN(n16304) );
  AOI21_X1 U17316 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n16310), .A(n16304), .ZN(
        n16303) );
  INV_X1 U17317 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n16302) );
  NOR2_X1 U17318 ( .A1(n16303), .A2(n16302), .ZN(n16469) );
  AOI21_X1 U17319 ( .B1(n16303), .B2(n16302), .A(n16469), .ZN(SUB_1596_U53) );
  XOR2_X1 U17320 ( .A(n16304), .B(n16309), .Z(n16470) );
  NOR2_X1 U17321 ( .A1(n16469), .A2(n16470), .ZN(n16306) );
  NAND2_X1 U17322 ( .A1(n16469), .A2(n16470), .ZN(n16468) );
  OAI21_X1 U17323 ( .B1(n16306), .B2(n16305), .A(n16468), .ZN(n16307) );
  INV_X1 U17324 ( .A(n16307), .ZN(n16312) );
  XOR2_X1 U17325 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n16319), .Z(n16311) );
  AND2_X1 U17326 ( .A1(n16312), .A2(n16311), .ZN(n16316) );
  NOR2_X1 U17327 ( .A1(n16312), .A2(n16311), .ZN(n16314) );
  NOR2_X1 U17328 ( .A1(n16316), .A2(n16314), .ZN(n16313) );
  XOR2_X1 U17329 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n16313), .Z(SUB_1596_U61) );
  NOR2_X1 U17330 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n16314), .ZN(n16315) );
  NOR2_X1 U17331 ( .A1(n16316), .A2(n16315), .ZN(n16326) );
  NOR2_X1 U17332 ( .A1(n16318), .A2(n16317), .ZN(n16321) );
  NOR2_X1 U17333 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n16319), .ZN(n16320) );
  XNOR2_X1 U17334 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n16324), .ZN(n16325) );
  XNOR2_X1 U17335 ( .A(n16326), .B(n16325), .ZN(n16327) );
  XNOR2_X1 U17336 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n16327), .ZN(SUB_1596_U60)
         );
  NOR2_X1 U17337 ( .A1(n16326), .A2(n16325), .ZN(n16329) );
  NOR2_X1 U17338 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n16327), .ZN(n16328) );
  NOR2_X1 U17339 ( .A1(n16329), .A2(n16328), .ZN(n16331) );
  XOR2_X1 U17340 ( .A(n16332), .B(n16331), .Z(SUB_1596_U59) );
  NAND2_X1 U17341 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n16330), .ZN(n16334) );
  NAND2_X1 U17342 ( .A1(n16332), .A2(n16331), .ZN(n16333) );
  NOR2_X1 U17343 ( .A1(n16336), .A2(n16335), .ZN(n16339) );
  NOR2_X1 U17344 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n16337), .ZN(n16338) );
  AOI22_X1 U17345 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .B1(n16340), .B2(n16341), .ZN(n16342) );
  XNOR2_X1 U17346 ( .A(n16343), .B(n16342), .ZN(n16347) );
  XNOR2_X1 U17347 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n16349), .ZN(SUB_1596_U58)
         );
  XNOR2_X1 U17348 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n16346) );
  NOR2_X1 U17349 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n16341), .ZN(n16345) );
  NOR2_X1 U17350 ( .A1(n16343), .A2(n16342), .ZN(n16344) );
  XOR2_X1 U17351 ( .A(n16346), .B(n16351), .Z(n16466) );
  XOR2_X1 U17352 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n16357), .Z(n16359) );
  XNOR2_X1 U17353 ( .A(n16358), .B(n16359), .ZN(n16353) );
  XOR2_X1 U17354 ( .A(n16354), .B(n16353), .Z(SUB_1596_U56) );
  NAND2_X1 U17355 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n16352), .ZN(n16356) );
  NAND2_X1 U17356 ( .A1(n16354), .A2(n16353), .ZN(n16355) );
  NAND2_X1 U17357 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n16357), .ZN(n16361) );
  NAND2_X1 U17358 ( .A1(n16359), .A2(n16358), .ZN(n16360) );
  NAND2_X1 U17359 ( .A1(n16361), .A2(n16360), .ZN(n16363) );
  NAND2_X1 U17360 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n16366), .ZN(n16362) );
  OAI21_X1 U17361 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n16366), .A(n16362), .ZN(
        n16364) );
  XOR2_X1 U17362 ( .A(n16363), .B(n16364), .Z(n16369) );
  XOR2_X1 U17363 ( .A(n16370), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  NOR2_X1 U17364 ( .A1(n16364), .A2(n16363), .ZN(n16365) );
  NAND2_X1 U17365 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16376), .ZN(n16367) );
  OAI21_X1 U17366 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16376), .A(n16367), .ZN(
        n16373) );
  XOR2_X1 U17367 ( .A(n16374), .B(n16373), .Z(n16378) );
  NAND2_X1 U17368 ( .A1(n16369), .A2(n16368), .ZN(n16371) );
  NOR2_X1 U17369 ( .A1(n16378), .A2(n16377), .ZN(n16379) );
  AOI21_X1 U17370 ( .B1(n16378), .B2(n16377), .A(n16379), .ZN(n16372) );
  INV_X1 U17371 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n16381) );
  XNOR2_X1 U17372 ( .A(n16372), .B(n16381), .ZN(SUB_1596_U54) );
  NOR2_X1 U17373 ( .A1(n16374), .A2(n16373), .ZN(n16375) );
  XNOR2_X1 U17374 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n16387) );
  XNOR2_X1 U17375 ( .A(n16388), .B(n16387), .ZN(n16383) );
  NAND2_X1 U17376 ( .A1(n16378), .A2(n16377), .ZN(n16380) );
  OAI21_X1 U17377 ( .B1(n16383), .B2(n16384), .A(n16385), .ZN(n16382) );
  XNOR2_X1 U17378 ( .A(n16382), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  XNOR2_X1 U17379 ( .A(n16397), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n16395) );
  INV_X1 U17380 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n16390) );
  NAND2_X1 U17381 ( .A1(n16388), .A2(n16387), .ZN(n16389) );
  XOR2_X1 U17382 ( .A(n16395), .B(n16394), .Z(n16392) );
  XNOR2_X1 U17383 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n16393), .ZN(SUB_1596_U69)
         );
  NOR2_X1 U17384 ( .A1(n16395), .A2(n16394), .ZN(n16396) );
  XNOR2_X1 U17385 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n16401) );
  XNOR2_X1 U17386 ( .A(n16402), .B(n16401), .ZN(n16398) );
  XNOR2_X1 U17387 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n16400), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U17388 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n16405) );
  INV_X1 U17389 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n16404) );
  NAND2_X1 U17390 ( .A1(n16402), .A2(n16401), .ZN(n16403) );
  XNOR2_X1 U17391 ( .A(n16405), .B(n16412), .ZN(n16407) );
  OAI21_X1 U17392 ( .B1(n16408), .B2(n16407), .A(n16409), .ZN(n16406) );
  XNOR2_X1 U17393 ( .A(n16406), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  NAND2_X1 U17394 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n16410), .ZN(n16411) );
  AOI22_X1 U17395 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n16413), .B1(n16412), 
        .B2(n16411), .ZN(n16419) );
  XOR2_X1 U17396 ( .A(n16414), .B(n16421), .Z(n16418) );
  XNOR2_X1 U17397 ( .A(n16419), .B(n16418), .ZN(n16417) );
  AOI21_X1 U17398 ( .B1(n16416), .B2(n16417), .A(n7573), .ZN(n16415) );
  XNOR2_X1 U17399 ( .A(n16415), .B(n13113), .ZN(SUB_1596_U66) );
  NOR2_X1 U17400 ( .A1(n16419), .A2(n16418), .ZN(n16420) );
  AOI21_X1 U17401 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n16421), .A(n16420), 
        .ZN(n16427) );
  XNOR2_X1 U17402 ( .A(n16422), .B(n16429), .ZN(n16426) );
  XOR2_X1 U17403 ( .A(n16427), .B(n16426), .Z(n16423) );
  NOR2_X1 U17404 ( .A1(n16431), .A2(n16430), .ZN(n16425) );
  XOR2_X1 U17405 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n16425), .Z(SUB_1596_U65)
         );
  NAND2_X1 U17406 ( .A1(n16427), .A2(n16426), .ZN(n16428) );
  XOR2_X1 U17407 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n16433), .Z(n16434) );
  XNOR2_X1 U17408 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n16434), .ZN(n16438) );
  NAND2_X1 U17409 ( .A1(n16439), .A2(n16438), .ZN(n16440) );
  OAI21_X1 U17410 ( .B1(n16438), .B2(n16439), .A(n16440), .ZN(n16432) );
  XNOR2_X1 U17411 ( .A(n16432), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U17412 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n16433), .ZN(n16436) );
  XNOR2_X1 U17413 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n16447), .ZN(n16448) );
  XOR2_X1 U17414 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n16448), .Z(n16443) );
  XNOR2_X1 U17415 ( .A(n16443), .B(n16437), .ZN(n16445) );
  NOR2_X1 U17416 ( .A1(n16439), .A2(n16438), .ZN(n16442) );
  XOR2_X1 U17417 ( .A(n16445), .B(n16444), .Z(SUB_1596_U63) );
  NAND2_X1 U17418 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n16443), .ZN(n16446) );
  NOR2_X1 U17419 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n16447), .ZN(n16451) );
  NOR2_X1 U17420 ( .A1(n16449), .A2(n16448), .ZN(n16450) );
  NAND2_X1 U17421 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n16460), .ZN(n16452) );
  OAI21_X1 U17422 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n16460), .A(n16452), 
        .ZN(n16458) );
  XOR2_X1 U17423 ( .A(n16457), .B(n16458), .Z(n16455) );
  XOR2_X1 U17424 ( .A(n16453), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  NAND2_X1 U17425 ( .A1(n16455), .A2(n16454), .ZN(n16456) );
  NOR2_X1 U17426 ( .A1(n16458), .A2(n16457), .ZN(n16459) );
  AOI21_X1 U17427 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n16460), .A(n16459), 
        .ZN(n16462) );
  XNOR2_X1 U17428 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n16461) );
  XNOR2_X1 U17429 ( .A(n16462), .B(n16461), .ZN(n16463) );
  OAI21_X1 U17430 ( .B1(n16466), .B2(n16465), .A(n16464), .ZN(n16467) );
  XNOR2_X1 U17431 ( .A(n16467), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(SUB_1596_U57)
         );
  OAI21_X1 U17432 ( .B1(n16470), .B2(n16469), .A(n16468), .ZN(n16471) );
  XNOR2_X1 U17433 ( .A(n16471), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(SUB_1596_U5)
         );
  AOI21_X1 U17434 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n16472) );
  OAI21_X1 U17435 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n16472), 
        .ZN(U29) );
  AOI22_X1 U17436 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n16642), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n16631), .ZN(n16479) );
  INV_X1 U17437 ( .A(n16473), .ZN(n16477) );
  AOI21_X1 U17438 ( .B1(n16475), .B2(n16587), .A(n16474), .ZN(n16476) );
  AOI21_X1 U17439 ( .B1(n16637), .B2(n16477), .A(n16476), .ZN(n16478) );
  OAI211_X1 U17440 ( .C1(n16642), .C2(n16480), .A(n16479), .B(n16478), .ZN(
        P1_U3293) );
  NAND2_X1 U17441 ( .A1(n16481), .A2(n16666), .ZN(n16482) );
  AND3_X1 U17442 ( .A1(n16484), .A2(n16483), .A3(n16482), .ZN(n16487) );
  AOI22_X1 U17443 ( .A1(n16724), .A2(n16487), .B1(n16485), .B2(n7821), .ZN(
        P3_U3460) );
  INV_X1 U17444 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U17445 ( .A1(n16727), .A2(n16487), .B1(n16486), .B2(n16733), .ZN(
        P3_U3393) );
  AOI22_X1 U17446 ( .A1(n16694), .A2(n16488), .B1(n10668), .B2(n16709), .ZN(
        P1_U3462) );
  XNOR2_X1 U17447 ( .A(n16490), .B(n16489), .ZN(n16513) );
  INV_X1 U17448 ( .A(n16513), .ZN(n16504) );
  NOR2_X1 U17449 ( .A1(n16491), .A2(n16663), .ZN(n16510) );
  OAI21_X1 U17450 ( .B1(n16494), .B2(n16493), .A(n16492), .ZN(n16501) );
  OAI22_X1 U17451 ( .A1(n16498), .A2(n16497), .B1(n16496), .B2(n16495), .ZN(
        n16499) );
  AOI21_X1 U17452 ( .B1(n16501), .B2(n16500), .A(n16499), .ZN(n16502) );
  OAI21_X1 U17453 ( .B1(n16503), .B2(n16513), .A(n16502), .ZN(n16515) );
  AOI211_X1 U17454 ( .C1(n16643), .C2(n16504), .A(n16510), .B(n16515), .ZN(
        n16507) );
  AOI22_X1 U17455 ( .A1(n16724), .A2(n16507), .B1(n16505), .B2(n7821), .ZN(
        P3_U3461) );
  INV_X1 U17456 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16506) );
  AOI22_X1 U17457 ( .A1(n16727), .A2(n16507), .B1(n16506), .B2(n16733), .ZN(
        P3_U3396) );
  AOI22_X1 U17458 ( .A1(n16510), .A2(n16509), .B1(P3_REG3_REG_2__SCAN_IN), 
        .B2(n16508), .ZN(n16511) );
  OAI21_X1 U17459 ( .B1(n16513), .B2(n16512), .A(n16511), .ZN(n16514) );
  NOR2_X1 U17460 ( .A1(n16515), .A2(n16514), .ZN(n16516) );
  AOI22_X1 U17461 ( .A1(n16517), .A2(n8944), .B1(n16516), .B2(n14819), .ZN(
        P3_U3231) );
  OAI211_X1 U17462 ( .C1(n16521), .C2(n16520), .A(n16519), .B(n16518), .ZN(
        n16522) );
  AOI21_X1 U17463 ( .B1(n16524), .B2(n16523), .A(n16522), .ZN(n16528) );
  AOI22_X1 U17464 ( .A1(n16526), .A2(n16528), .B1(n11462), .B2(n16525), .ZN(
        P2_U3501) );
  AOI22_X1 U17465 ( .A1(n16529), .A2(n16528), .B1(n9798), .B2(n16527), .ZN(
        P2_U3436) );
  NOR2_X1 U17466 ( .A1(n16530), .A2(n16663), .ZN(n16532) );
  AOI211_X1 U17467 ( .C1(n16643), .C2(n16533), .A(n16532), .B(n16531), .ZN(
        n16536) );
  AOI22_X1 U17468 ( .A1(n16724), .A2(n16536), .B1(n16534), .B2(n7821), .ZN(
        P3_U3462) );
  INV_X1 U17469 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n16535) );
  AOI22_X1 U17470 ( .A1(n16727), .A2(n16536), .B1(n16535), .B2(n16733), .ZN(
        P3_U3399) );
  NOR2_X1 U17471 ( .A1(n16537), .A2(n16663), .ZN(n16539) );
  AOI211_X1 U17472 ( .C1(n16643), .C2(n16540), .A(n16539), .B(n16538), .ZN(
        n16543) );
  AOI22_X1 U17473 ( .A1(n16724), .A2(n16543), .B1(n16541), .B2(n7821), .ZN(
        P3_U3463) );
  INV_X1 U17474 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n16542) );
  AOI22_X1 U17475 ( .A1(n16727), .A2(n16543), .B1(n16542), .B2(n16733), .ZN(
        P3_U3402) );
  OAI211_X1 U17476 ( .C1(n16546), .C2(n16684), .A(n16545), .B(n16544), .ZN(
        n16549) );
  NOR2_X1 U17477 ( .A1(n16547), .A2(n16702), .ZN(n16548) );
  AOI211_X1 U17478 ( .C1(n16705), .C2(n16550), .A(n16549), .B(n16548), .ZN(
        n16552) );
  AOI22_X1 U17479 ( .A1(n16708), .A2(n16552), .B1(n11359), .B2(n16707), .ZN(
        P1_U3532) );
  INV_X1 U17480 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16551) );
  AOI22_X1 U17481 ( .A1(n16694), .A2(n16552), .B1(n16551), .B2(n16709), .ZN(
        P1_U3471) );
  INV_X1 U17482 ( .A(n16553), .ZN(n16559) );
  INV_X1 U17483 ( .A(n16554), .ZN(n16556) );
  OAI22_X1 U17484 ( .A1(n16556), .A2(n16686), .B1(n16555), .B2(n16684), .ZN(
        n16558) );
  AOI211_X1 U17485 ( .C1(n16691), .C2(n16559), .A(n16558), .B(n16557), .ZN(
        n16561) );
  AOI22_X1 U17486 ( .A1(n16708), .A2(n16561), .B1(n16560), .B2(n16707), .ZN(
        P1_U3534) );
  AOI22_X1 U17487 ( .A1(n16694), .A2(n16561), .B1(n10732), .B2(n16709), .ZN(
        P1_U3477) );
  NOR2_X1 U17488 ( .A1(n16562), .A2(n16663), .ZN(n16564) );
  AOI211_X1 U17489 ( .C1(n16643), .C2(n16565), .A(n16564), .B(n16563), .ZN(
        n16568) );
  AOI22_X1 U17490 ( .A1(n16724), .A2(n16568), .B1(n16566), .B2(n7821), .ZN(
        P3_U3466) );
  INV_X1 U17491 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U17492 ( .A1(n16727), .A2(n16568), .B1(n16567), .B2(n16733), .ZN(
        P3_U3411) );
  XNOR2_X1 U17493 ( .A(n16570), .B(n16569), .ZN(n16591) );
  INV_X1 U17494 ( .A(n16571), .ZN(n16572) );
  OAI211_X1 U17495 ( .C1(n16586), .C2(n16573), .A(n16572), .B(n16698), .ZN(
        n16589) );
  OAI21_X1 U17496 ( .B1(n16586), .B2(n16684), .A(n16589), .ZN(n16581) );
  XNOR2_X1 U17497 ( .A(n16575), .B(n16574), .ZN(n16576) );
  NOR2_X1 U17498 ( .A1(n16576), .A2(n16702), .ZN(n16577) );
  AOI211_X1 U17499 ( .C1(n16579), .C2(n16591), .A(n16578), .B(n16577), .ZN(
        n16594) );
  INV_X1 U17500 ( .A(n16594), .ZN(n16580) );
  AOI211_X1 U17501 ( .C1(n16691), .C2(n16591), .A(n16581), .B(n16580), .ZN(
        n16582) );
  AOI22_X1 U17502 ( .A1(n16708), .A2(n16582), .B1(n11365), .B2(n16707), .ZN(
        P1_U3535) );
  AOI22_X1 U17503 ( .A1(n16694), .A2(n16582), .B1(n10748), .B2(n16709), .ZN(
        P1_U3480) );
  INV_X1 U17504 ( .A(n16583), .ZN(n16584) );
  AOI22_X1 U17505 ( .A1(n16642), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n16584), 
        .B2(n16631), .ZN(n16585) );
  OAI21_X1 U17506 ( .B1(n16587), .B2(n16586), .A(n16585), .ZN(n16588) );
  INV_X1 U17507 ( .A(n16588), .ZN(n16593) );
  INV_X1 U17508 ( .A(n16589), .ZN(n16590) );
  AOI22_X1 U17509 ( .A1(n16591), .A2(n16637), .B1(n16636), .B2(n16590), .ZN(
        n16592) );
  OAI211_X1 U17510 ( .C1(n16642), .C2(n16594), .A(n16593), .B(n16592), .ZN(
        P1_U3286) );
  NOR2_X1 U17511 ( .A1(n16595), .A2(n16663), .ZN(n16597) );
  AOI211_X1 U17512 ( .C1(n16643), .C2(n16598), .A(n16597), .B(n16596), .ZN(
        n16601) );
  AOI22_X1 U17513 ( .A1(n16724), .A2(n16601), .B1(n16599), .B2(n7821), .ZN(
        P3_U3467) );
  INV_X1 U17514 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16600) );
  AOI22_X1 U17515 ( .A1(n16727), .A2(n16601), .B1(n16600), .B2(n16733), .ZN(
        P3_U3414) );
  NOR2_X1 U17516 ( .A1(n16603), .A2(n16602), .ZN(n16606) );
  OAI21_X1 U17517 ( .B1(n8041), .B2(n16684), .A(n16604), .ZN(n16605) );
  NOR3_X1 U17518 ( .A1(n16607), .A2(n16606), .A3(n16605), .ZN(n16609) );
  AOI22_X1 U17519 ( .A1(n16708), .A2(n16609), .B1(n10759), .B2(n16707), .ZN(
        P1_U3536) );
  INV_X1 U17520 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n16608) );
  AOI22_X1 U17521 ( .A1(n16694), .A2(n16609), .B1(n16608), .B2(n16709), .ZN(
        P1_U3483) );
  INV_X1 U17522 ( .A(n16610), .ZN(n16611) );
  AOI21_X1 U17523 ( .B1(n16618), .B2(n16612), .A(n16611), .ZN(n16620) );
  INV_X1 U17524 ( .A(n16620), .ZN(n16638) );
  INV_X1 U17525 ( .A(n16613), .ZN(n16615) );
  OAI211_X1 U17526 ( .C1(n16616), .C2(n16615), .A(n16698), .B(n16614), .ZN(
        n16634) );
  OAI21_X1 U17527 ( .B1(n16616), .B2(n16684), .A(n16634), .ZN(n16626) );
  XOR2_X1 U17528 ( .A(n16618), .B(n16617), .Z(n16624) );
  NOR2_X1 U17529 ( .A1(n16620), .A2(n16619), .ZN(n16621) );
  AOI211_X1 U17530 ( .C1(n16624), .C2(n16623), .A(n16622), .B(n16621), .ZN(
        n16641) );
  INV_X1 U17531 ( .A(n16641), .ZN(n16625) );
  AOI211_X1 U17532 ( .C1(n16691), .C2(n16638), .A(n16626), .B(n16625), .ZN(
        n16628) );
  AOI22_X1 U17533 ( .A1(n16708), .A2(n16628), .B1(n10785), .B2(n16707), .ZN(
        P1_U3537) );
  INV_X1 U17534 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16627) );
  AOI22_X1 U17535 ( .A1(n16694), .A2(n16628), .B1(n16627), .B2(n16709), .ZN(
        P1_U3486) );
  INV_X1 U17536 ( .A(n16629), .ZN(n16630) );
  AOI222_X1 U17537 ( .A1(n16633), .A2(n16632), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n16642), .C1(n16631), .C2(n16630), .ZN(n16640) );
  INV_X1 U17538 ( .A(n16634), .ZN(n16635) );
  AOI22_X1 U17539 ( .A1(n16638), .A2(n16637), .B1(n16636), .B2(n16635), .ZN(
        n16639) );
  OAI211_X1 U17540 ( .C1(n16642), .C2(n16641), .A(n16640), .B(n16639), .ZN(
        P1_U3284) );
  NAND2_X1 U17541 ( .A1(n16648), .A2(n16643), .ZN(n16644) );
  OAI211_X1 U17542 ( .C1(n16663), .C2(n16646), .A(n16645), .B(n16644), .ZN(
        n16647) );
  AOI21_X1 U17543 ( .B1(n16678), .B2(n16648), .A(n16647), .ZN(n16651) );
  INV_X1 U17544 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n16649) );
  AOI22_X1 U17545 ( .A1(n16724), .A2(n16651), .B1(n16649), .B2(n7821), .ZN(
        P3_U3469) );
  INV_X1 U17546 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16650) );
  AOI22_X1 U17547 ( .A1(n16727), .A2(n16651), .B1(n16650), .B2(n16733), .ZN(
        P3_U3420) );
  INV_X1 U17548 ( .A(n16652), .ZN(n16659) );
  INV_X1 U17549 ( .A(n16653), .ZN(n16655) );
  OAI211_X1 U17550 ( .C1(n12994), .C2(n16684), .A(n16655), .B(n16654), .ZN(
        n16658) );
  INV_X1 U17551 ( .A(n16656), .ZN(n16657) );
  AOI211_X1 U17552 ( .C1(n16659), .C2(n16705), .A(n16658), .B(n16657), .ZN(
        n16661) );
  AOI22_X1 U17553 ( .A1(n16708), .A2(n16661), .B1(n16660), .B2(n16707), .ZN(
        P1_U3538) );
  AOI22_X1 U17554 ( .A1(n16694), .A2(n16661), .B1(n11066), .B2(n16709), .ZN(
        P1_U3489) );
  OAI21_X1 U17555 ( .B1(n16664), .B2(n16663), .A(n16662), .ZN(n16665) );
  AOI21_X1 U17556 ( .B1(n16667), .B2(n16666), .A(n16665), .ZN(n16670) );
  AOI22_X1 U17557 ( .A1(n16724), .A2(n16670), .B1(n16668), .B2(n7821), .ZN(
        P3_U3470) );
  INV_X1 U17558 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16669) );
  AOI22_X1 U17559 ( .A1(n16727), .A2(n16670), .B1(n16669), .B2(n16733), .ZN(
        P3_U3423) );
  AOI21_X1 U17560 ( .B1(n16673), .B2(n16672), .A(n16671), .ZN(n16674) );
  OAI21_X1 U17561 ( .B1(n16676), .B2(n16675), .A(n16674), .ZN(n16677) );
  AOI21_X1 U17562 ( .B1(n16679), .B2(n16678), .A(n16677), .ZN(n16682) );
  AOI22_X1 U17563 ( .A1(n16724), .A2(n16682), .B1(n16680), .B2(n7821), .ZN(
        P3_U3471) );
  INV_X1 U17564 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16681) );
  AOI22_X1 U17565 ( .A1(n16727), .A2(n16682), .B1(n16681), .B2(n16733), .ZN(
        P3_U3426) );
  INV_X1 U17566 ( .A(n16683), .ZN(n16690) );
  OAI22_X1 U17567 ( .A1(n16687), .A2(n16686), .B1(n16685), .B2(n16684), .ZN(
        n16689) );
  AOI211_X1 U17568 ( .C1(n16691), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        n16693) );
  AOI22_X1 U17569 ( .A1(n16708), .A2(n16693), .B1(n10985), .B2(n16707), .ZN(
        P1_U3540) );
  INV_X1 U17570 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U17571 ( .A1(n16694), .A2(n16693), .B1(n16692), .B2(n16709), .ZN(
        P1_U3495) );
  AOI21_X1 U17572 ( .B1(n16697), .B2(n16696), .A(n16695), .ZN(n16701) );
  NAND2_X1 U17573 ( .A1(n16699), .A2(n16698), .ZN(n16700) );
  OAI211_X1 U17574 ( .C1(n16703), .C2(n16702), .A(n16701), .B(n16700), .ZN(
        n16704) );
  AOI21_X1 U17575 ( .B1(n16706), .B2(n16705), .A(n16704), .ZN(n16710) );
  AOI22_X1 U17576 ( .A1(n16708), .A2(n16710), .B1(n15805), .B2(n16707), .ZN(
        P1_U3541) );
  AOI22_X1 U17577 ( .A1(n16694), .A2(n16710), .B1(n10975), .B2(n16709), .ZN(
        P1_U3498) );
  OAI21_X1 U17578 ( .B1(n16713), .B2(n16712), .A(n16711), .ZN(n16715) );
  AOI222_X1 U17579 ( .A1(n16719), .A2(n16718), .B1(n16717), .B2(n16716), .C1(
        n16715), .C2(n16714), .ZN(n16721) );
  OAI211_X1 U17580 ( .C1(n16723), .C2(n16722), .A(n16721), .B(n16720), .ZN(
        P1_U3241) );
  AOI22_X1 U17581 ( .A1(n16726), .A2(n16730), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n7821), .ZN(n16725) );
  NAND2_X1 U17582 ( .A1(n16728), .A2(n16724), .ZN(n16731) );
  NAND2_X1 U17583 ( .A1(n16725), .A2(n16731), .ZN(P3_U3489) );
  AOI22_X1 U17584 ( .A1(n16726), .A2(n16734), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16733), .ZN(n16729) );
  NAND2_X1 U17585 ( .A1(n16728), .A2(n16727), .ZN(n16736) );
  NAND2_X1 U17586 ( .A1(n16729), .A2(n16736), .ZN(P3_U3457) );
  AOI22_X1 U17587 ( .A1(n16735), .A2(n16730), .B1(P3_REG1_REG_31__SCAN_IN), 
        .B2(n7821), .ZN(n16732) );
  NAND2_X1 U17588 ( .A1(n16732), .A2(n16731), .ZN(P3_U3490) );
  AOI22_X1 U17589 ( .A1(n16735), .A2(n16734), .B1(P3_REG0_REG_31__SCAN_IN), 
        .B2(n16733), .ZN(n16737) );
  NAND2_X1 U17590 ( .A1(n16737), .A2(n16736), .ZN(P3_U3458) );
  AOI21_X1 U17591 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16738) );
  OAI21_X1 U17592 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16738), 
        .ZN(U28) );
  CLKBUF_X1 U7810 ( .A(n8994), .Z(n9345) );
  XNOR2_X1 U11591 ( .A(n9860), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9797) );
endmodule

